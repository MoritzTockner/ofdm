-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
JusLw4TzrVK0BV0N1s/ARQ/ca4bbIexoIPbB+aH0x8e9BqxYzFRzx7t9e5TcMsmUhF5alohsXNGC
RO+7vDq7/PnOCVRmYlnXE8vQPQJbu2w20sQEQxbD5ishFGXydst1KqlcHOI3RM6kOVrRskbSdMdj
etZA4K87oY5aiN5Il6VupTYxRGbE6DwDpHTYkR/er+zPo9UsuElRwg7Ex8MaZagt5Hx2G5zOn2WY
B58L93qQ/muBM/Ii7ieMB2qwg+dQHf+Ts3eMUiuVI7vlwSvvqToZd7Um09+h8xdDyo23hUKVyB+a
RcfAAnQwjqxzlnq6HADEI0/CpEN8KGjXOYpIJA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
kIWwcvSgyunKjovrohDtPcU1+SsBz7I38fq9R64E514zU33xSYHEoT/tp6vIszGasDToQjub9cLy
lNUrhY6wA1ueMQooEXvjaje+bTAwhK4ej2MOeTRbdCxzxHm56xaDCOtQ0qOVKOTfL7ncUXLfK9ZQ
FaXRZyxQ1yRChce+kSEngp8Pf1Al+AzD4fjRk282qvFZedIES3iC7l+KLiaD8CeoBgrBodInJXAH
MYc5Mc4k0oWzLFl7go2xO6wPieDZd5zJL/GsTMobSGMztTwAy83ua8QEKfM4GtAMx8fSsO1/Ti9m
ZB4Dq2KZOG0fezlgakMCgFNaA8aa37TvnvZ2PhvhI502oEHXu3X90pBiZDzGirTkc8UHnEZoayBe
d8Ef0FVNUKec48Rgy5BrkkEYAATKOeAHDAsIIImfFghsSXoJUoG9d7zFPv7MFKGRnS4OJMJWwOrE
nsjNN4aaEhAau6Cqdvq8OqHAgWyMp62zhjIA63gTvFwCGLk9yw2NS0p8MHTGpUBZeVsn4V9rAPBB
lAy5JMgCeMc2xI7hpkSPHGfmTrEMR6XTJ71zhBOZ2Jaufoxo7qTPtGHDUhL0HFAgedr5KTvjcXjH
uQnZmkrNoVsXHgAzQYkzMr5ouZJLV5bQ51sxsnODYweN3/4ErR+QRDucpb2WnMb9oI0ywZ9bcGIQ
T3UomWUZzKL3t3MkldKApgGbqXgmgI5EY8z6wKtavaFGgIqXXnRAUqtrxQD3x4eZ7jd1SbeJ5bu/
WTwcmje3xHEPYMqv0cj46kbdt8LQu7FK37B0TYO5PSR1Qt4ENM0+LGo9cCgc8+PYA/6kYSDpQKId
5gRFR8CQ6rG764YEwHCH25HlBjcv8uY+jobYX2EBeGTBrkmC20wmxTYrp2tde0Rvs+uWfaLUoMmu
Bi3TKNszfMBt2/2BDZ7tibJQI3KI5l0d1Lzrtanv5EH8lLjSDAQNKMtyq4pUwwosPEwqdZelZHD7
y1N1fBWLpy8chcIvQFajQ9aZi8Vqs45XnGLED8sEF0c17FjFyNzk6iconHd+7tW7KXRjj/+aX3e/
YOiIbUe1hU4ub6JUHTLw0iDp24+UX22GEtVwe6OPBXPQw+j2MJwP7YBB9DgFQeq7+JW3nJikg/Vn
9x4cp/YDpLwMU7XQMEM2CDeAtsV96mrFsb1pJKrZoAb8uK6wrPAZpjuNva7h+GaEK8+3g9kXEEGA
Pyl2uL0EHoLUAv57KAhqnd/jSV9gPqqLyOuZ2wWJy1X8V/pr0e17kYEPSRFR1VcfFLblG95zAPXa
HX3UwTSm6bsm65ebW9zih881xhuxk3O781yaK7ehYcBHw67NgK05Fy7+fMKF23ifWa5cSX1Rlpzt
/74MJJxFr7rj7j015Lpa/33/K+ZCRaiL1SVbJtJpl8+zgMopfDJFbcejMCMG6IkxpLwZbcsrBuj+
xTdgjoHYM8F3QLn8aXxqBDEea38Sjmlsx8ZvTNWk6jyy65YxOctIMqBb1rHWEF8+BOOj9OyUoTYN
3eJX3y9hufl4IG/UNCXvc/YCm1coQdm8i6BOf9S7uzsu/1XCaD3RUk30EgDysBUpHTAovg7UnUex
X/1qMq7ojZlAef70Ezn+sDMAJEQmJFv+fjA8enB01r8LcjxIyYuCJxqS2OZcFxREqBM5F2Spp7AS
gEAwc0ShQd/+ELC0bCpNbds2TiG0BdjDub9suSd06WpqtHjB2ZJkXPIcKc4uIO9G9NuTFgKeQ/sf
NWRqbj8s6xscuIR0VF+RVfPQ/DNYd7H9FNlmw7LC/fpEU8dsbABdTTdiOaWhswsEdqTYomQprNUh
OduyUJ86fg8Ex4v/1b3nADXmcBuqcS4a6akFG4HXj7LFis2SyTPkZwqBxyv17seuaqLtE1FaciUt
mClMYl0A5nSq37r3aAxYlDzYkL89w/j96C0WGJkUn/f+JYGnw2SaDSGLyru1PKvkNR2y7tNapo4K
5+w8bcrvvk7+kFIz876WGHkn5gt+t8vgKeRJGehcoObQ8xYZgVZPWxYcc4hzJ/bI2MnZzTiXvXaB
SpPik0GGmGJWvWcN4sg5oOaRAiHe9hzIvjVYuOEaY/k1OpvkzahMBIocLxctDRT32UOL1rEK0XIx
F8GPTzEmrRySvzIZiGfAz3Bu+5vA2PEdHagCQ9RuQFu+6UxbT+9RcfuPNEfRnHFBGVCwwwlraEuL
TX4PqYjFMG55qHymnKByd9h3pFbRBYNswoSGJazoHdi4q/3006TWD7Bm8zYHM6B194s/chHxxOj2
GcuVgY2cvV6ZnquAm3hNnDb6kbc/Jr2HvOzHVceyrnokQIN7IWEgThYr2Ga8YrRreYvEgV7VCq6f
tNMiXj9u+Ix/Lkz/0IaWHnZcKlmWeafG6JZxYsZuqVPOWbVnVf+VUWyt97ie5cO9SxFf1pNCqZXs
r/44xsvHGDFl2vHXQaY45LIqMZYwgd5k+xWjN9Ra9d9PG2D3Uz4TjAWdD4GR+31C5D7mPAKj6NJQ
S7zNr2HmUFlBtMBQScVEzN4GXloJpHulmDH6BkqC0JvHrSkAwSvpfUfe/kqjQDG92OtYa1jw6QwP
OmcAAgYvMrD4DWmR7EAQiIA73vZEXN7NXMENiSQN66i7KqXKke7M2witBd2qQaUk8gvtr2pGKZiG
uyKGFfv7Vl/f9Hcbn/O7ZnnDmHqOOSC1LifLLEUSzaTXLCNxDdUKRLcy9pc8FhfSic71eSAQvUOO
xLSMYixr7nluO6YLLVKQk5pwDpiq1HDzHREeiela0Q3MiRo5bril1Uy+jwCeQl4n4dVNvO6BkTtp
Q6Hzpk4Dwf5WNXXqTRP/Rd+vUwxFmPy90yE/2+5MjagRG9QKUC5MFfUUy+gS8txFoPM48Hl4caIN
QugLcnFW92lQV7B9IHN7FiSlXbDQb+dE6ojOJuYjnDTwjWlBIDiLQVSgdNRYCO8pDkAjtImHbOeL
+rsVGsb2jGzstgmji/xyplIvWR+CYQP2ULq7Oxc4pGG8Bj0/mZmptWHn5D/hnsb9c94rrUfAD3WA
90tYySpaIpixnuYTed6GqD2Vru6H11U/+G7DZ6wP69I9c4WQgZcfTKQzS3px5Y1byScRZA5mH2Pt
Ru0T+sxDDUGx7WOM5Ad24KnX0mG9EzdZZdeFq8Fu2F9IORvqSlYd2/QJHNkD93fLqIP2TqSePbvj
Bv0XzMaLGrWkk/TOvh2cuDXZeiDAk/7zUELFUGIfxx6uldPDqWH1ploZe5BOVtskQ/3qnbO42cnU
hRP1vWZp6vvtTQACmOQMTrKImRRN1uidiyZqvZAsEt3sBNjvjwfwAGBAZd8gS2HTXV5ITNM7nZOu
SyabzILWCbwzfQBErvmbBiWdx/2UDAK7HMRne9Vmx+N/08Xi11TcH+sSCgFyg71Dutw4RRAolriw
tgdJVC5bGVHQuUG6edDF03u77bOGfU1dCoOsrFpPAftn0M6FWwXjEXJQpFjbqpM8Y9GEwSdLWuPs
6k0PmuSdi9NL5IR9eUSYaJecD4icVIOyZfxsn3rKFGlKbGsj/SGihZM3sIKqzax4bGUlyRaQHTJ1
eNsd8CBD0K4wpthmhodEBdxgHJQrJytzVHVuBCovSgZZPwiE6E6PS/5uK9jDUym3pTC+KmMVu6G/
mTOgaAfpSc+dQSItN8goS4JSMypGQ2bapo5DrdY8kLYweQ7J4clRrfzSEOsD1vd2VXxrr26SV/us
Naa8lh3KKC7hr/yHiUsAkuvSnMwaIyBItb8uEG0ba8qXk7udp2oGkm+iM41T6CnuVl2oNNzZE+nk
VTV95Z7DfVEhG6J1uHuX0vZpBNoob+kUOfwo7xbtq3Fnk8PICwzxaUthpNqT9mAXx2dFuYRQ751T
nngd8skUcqCcjc4SmiWlUq7fIATg+ITAzVIE3JP4EPzznsub1LeIrK91OZZ3As4BfUM3WrNC9mMd
2UYFCBxkpxXfkWeXsSSrQvuWoyo5YwzT9mlEZGUjY7fSkvaIv08VTit+4Z0Z5nH1ReHm0rbkqp0/
hjh2Op2ENvK3QNmAbnm40RS6VJbMwNUhd4GRLY9w8scGT5pgbLL3M3r3ZPkRLdzPrwofFWMFs+E1
aG9UULefBCI3At24PcmiYJ0nKiMC7LEZ/niLchLAgQTPgtrIYKYyF736N9+OtgEP40s0pGJuR05A
2mOnoI6eePnxJ3jkVYBoOGc84RNAn8mAG2Dl8CyJu8Scuv4e7CifjCDVd2boXlUDKPf3AqeMaZyp
mt212dfrLBai6MArKFbB9D7d7bVEXcRhlXahrsMI6wIPx3UW5QtnHiUHwpoKXqxmWG/ZRhsnuSFH
Wsfu9/eBj4l+qq23lYjdowCpZFYYAwk32PjIb9kWhE4/f9+vDPLtS9KlnEGcx8Vp8XUHb0Nvqp+q
1gC7hrb9FvpH7nN0z7XhvMxMBkQa1R9tWSSUqUysJLK+y/dMb6pUA+aPMeasM0sGXtAwAjYDJqB5
0CO3UQtxVtpKi/m1yGWN8egHLBPist9l3GKPDPHFIgjCNO7oPBD3tXrUIyFBbA3uzwhpvZK6CIC6
x2FgfSP/Zy5/qj3Y3S4Fy9UQZ516tNnnc/6qgDmmGeVtqdFjqaAtvmZZQ6fOQ3uJ+6VmDmMG6+ZT
7FNkUNHoBm7TXWFYypCLaWFNJTAphhAOZHdPBDSLLNNmYprp1f7nhrkeKz7qByZrBL0aiynymhkC
e1oUbbMPQ2IZh+8OYL2rN570edWjosWSTZI3otT2LWf8nxYnGDVBjIraCSE69GrCz5Vz3e4dDV9G
fVuRgNkY6yC2nugp0hohXkfdclPfCXpcfnpIXbaUWmLed3ZZcr44l6Nau2aXwy/uu5IBWt3R/g9b
ykuif6DVVmQ141yMpFC1Cx2lngtY0UAv8Pdf0OAnM3i93ycWQ7k3ONFFdIfhgrFi0ELDXmWPbTAq
66wUUPAKUkZxU//Jk9YPGg8Gx7OvB/yISNDM9WGb+b6liaa6Er9ned1/DSVtXKbxcojxpVZqCtRe
4BUUrQv1Ui2HFCtznsJRzjTsBDjY0ARRsuXHEXYBn5pMB+bqgYFyiGWlwqKg2JXgzFcd4ZjbXv8k
hOoy3Vg740VSVdCBCQPVXfAifH3yHk4/ExT/rCw2nVloAbgOYBjwTk716WgVW0GZ1yX2en4eNtkL
uxSUl0a+DDK7mNE1LAZKXYI3JTpUrExI0tXzq2jMLKJuHh27t73QrajeCHI/figN+hGztge7Cz0Z
cggx666LE4lBX4INyAf6TpIB5rqFSw0WCmWJ1c7m4eX0jdZS9lAynVCgf/u6NpTOFftCjunm4BFP
k71Y1l3wuZf7xo37RpdZg/A64b0pyXwlu9UcvOiY4oEOtYp7i2KnpDxCyJ8zMxGil0x8Sm49d+rm
Jr9RpOwejp3ai6/UwlX1OHF9Yn8m+Yx86XZf5XB+r822DO8TIFfP3utJz6yhRc1AAjNq3cQEyytZ
26N2eo/RwsU2iP5FZkEjHtcb7VTnzK/fXQ0JEqUb4PlKKk4WtDaeXnYvIcIZjVSv2r/J0aWAM7+B
D9Vx4C1lL7KHu6zRBHUOKURVz6pLUGHt92Fj9TmuGgBNOGxmX7L+9AZ0LHg3JHzNMLbMr2Qg1Fji
YgzJ1Tgv5DS4/JEwceFGGGG7/kQo6dFwhn3rfgdjA+upoV4Gcgpxs5qYhdRUBktw1xDbGbMq8Hik
OHDVOLRjt1CSaUrLCqxYuseml8MF2nkVqeMoNvDUp5xOgZQ9FqX3OxjuqRbEfFFisT4CarBtgIYv
dLGZBeWDyKEU9MCR5RafjCdOA8TeIUEDxRHKQyJlN3+aBUMaqhc2DePwOxY2ih64p26rgmgRX5F4
1B+7Zq6mI6q9n658k91Ovq4PyAJrSiaVdQazJe8wkgBrxGVTD/y6/7r7yDkcKnsi16wghTAnKWTW
gXU5gaU7PMlJShzcKbeb04XxoTXTvJdv7qc5IFZFhNVbuqoz9TTbEo7Qry3icAJLp06QEdXyFAfI
LKltPTHEwSY6z5XHCrYm33lwPBlvl/+CU9+g/xBYE5RTOUOlNYLYU2ylI3wbN+GEt9VHL2fgPRap
5cdf3wONo9weAon0yWUAODPgOjdxr+SvjUtvjRhesIpV3Uf28S3yGqq92RD+fXoXMfRyPAku10NC
9kCPDxH/xWEUNfP3NPvH41WHQGI1ou/TMFQqhKFx6HK7yapOltXgQyhn3vGXdX/N3N2tUwNPLm9n
tIR4ue4KAGKR1Elw0pJfk1iph/Y+NAFbMkE3Sbae33i4UTqXUCazhxfFAgLdAueQVHaZKuAyVOjj
w0n68XgXfWGwLwoGrtaoWigsM/Itjww8/pa8YDadN1sIw0n2PdHH9awSGg5vZwRlxHWhvHmKmbSO
5Za7GbMQiRWRJ4A2CmZm4TnlI6RxITHyKAGMkVp3CT0yGqEzWdmxa1MJLPt65orgQLsd5yjUQeuj
JHMXiBI3AW3piy3wEMkfvrKTBHWsaFVXcbjELGLodn5asv3uC03ckDAbCjKUoYO8yGExJcvraszO
tul50LG0vNQ7S+62tXxferCwKnMWOc4d26nzjd9e8niHgLrLZG+cBdpBCX+hfIXad/ubK3wUScPa
TWm3k8YAQo6odRNIoWmtLUDQTbAq/coerAiK8NBv5hKakws8YGsINECSGFM9tR9EVmQn5s76vkm2
uGsT7zCGTYN42CMkZS74G9NwiwU6XJxyfK31YCrWXBGP3/ptax9CBSka4zuK3FjJqCisaB4hmFmX
WX6YUscRx5ohXDb8PkJcb196Es2wjYJNnZlqRwdMhiBlSdcorzlHEqJ8w4CAuKP+KUA7arZnV3he
pWh9E+8zhOfnNxHKV9UnAX+iEJjX3ZwPb942qDxKOT1ifOjfhl0ioOoq9jI5FHuNhwZv2gjnEsNG
RPwtRsSTwYbJwWa1K9f0xQIMUc8RfJ2DGK7h02AjxPbbc1gWaeRap7qbGcEliZZG0IPThjDWo+S5
G5i3GyD4PLYxHGUGPVzpUTPdw/l+LsNofoZFCp3bjbF7Ruz7yfoGkvLutnX4I0eNy+ftm639Naeq
HLcY1dk4YJE3/9ACv7S3q4VDDchemEVMO/gl/YGQwzkt9z5Op8ZYYZ7K7+TLJqwJDAqWX8CUPIWd
lmdq4HQ3RYHEhUD0nNJjm4GCCFUj4rPNxjllxv3bg6n9spHhIJsA6XqLlnp+RnJb47olPmyEk2/Q
uyIuLB2JaYgyQeEsel3ux31jJsNgr7ZCj+YQptWzt8afcAmwze10Ae3dZXRHQks721aBWSE3I0CJ
hJqCxBvyrdzaYwK7GkdHpywUQjF+rulsN2RfGVq5K9hmN0TdUHxiYHn343cnUt1zmxJlptHdOpZW
yVDCG8dLnAJmL/lECwBttHPKpk644hHoJrQ4Fc2rWGt5bR5VpKKvdq4VDiidkwV6OxzF9516LyjJ
dPhJIlO7gQD/dIvmW0jnUm1/Us2QXadHwpecKIgjNJaluwaLPp4Z4gH8Tfncj+y93W94KDQAsib0
TajnGRlRxhk7sqlSVePG7sbDg97UUsFiA9jHFM1uI+sgd7nd8vjiAfmXROI/jssFe+i0z0bIq/LQ
Wsg9s6SZe0W25z2VgV0+Xcxj1U/1kofdhUKPy+edmUhkHs5SW1smVG0Bbz/I8d3wDGmrIGvhrVBn
0p9ZzcehastmO2Ca8akzs+2WyjYOJU736hs1XwxIxUNBndO0zuwSXaP2pKnVkpb3zXT01wypF5EJ
LGDlDZ3a04WZYF0p47CRGTuTDQARdBIwOf/lwFbAIjWZfkREwTtiFMoTueKbxzooxfC748Iyu7mj
eDcdKGKyPZp2uuRNwMCB4HMjMlryNQxjVrc9vUbwjDPy4xIFUKqXoFGChBGAQQQltagcIQ2IwE1v
JfwS1oNrOCwmUynaJv73oP6LZ8PKTbDOPhkVXND/0abzKVOFu9bRs8SwsNVlMgGqyR+nQkmQlCgv
guQuyvN35C+jVQUaz4JRtyf+n7H7u8SVpWugCr5jM9oTtIGWWOheyS8EmkibT9vXuDLAXlmgQtk1
dA9nN/4EqbwJaX+smXBxrHmNJ5admj7yTxWmaxMl6YdPE+xBD6qEFdc6jRZbqr6Eru93lBbwGFmw
CNDfsJcDqzN80fdBZ5+rFhq6MrzOt3x8+JQ24amsj3arUe3FPuDWupf9jpdj3Hd8iY6puQRhzVgJ
FMqKc6rHRFu9l78gnjvw8nOCCKlKQpChHNZXWFN14942kRJF8mgBNOVeSiDqpB6tMof36Q==
`protect end_protected
