-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
t1TpGzP74+zWKqWoOqyZOkPSUvL8P8mlajEKNv7lo4hN+oeG6Jdy3ifulDT+//WjbFvL3QGR7lDi
ntwCa4kheIIoNRCGg6e8f6M/40V33FIKkgwQeDrfUscnjKxzVKYZcpewRS4w7rhAmxaiLoCxCFs9
QykZZtI1EOWCvJSIJA/ghTQ+Nf3D0wrlCg7vlSPiQmwopbohxCaIUNsExpxt0q9hqtdASNXBA8Hy
Q/kTD7/LhtW1HFv4yQwKU3DxvaY+xJw2QiVmGFhXdGUoJjOFbSp79EtG430oQppEDwnBbIGYUWgS
jyMekfLj6uNgl/R3u5fXF/dJfbu1NoKyjT/XUA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
a4FNxD54QcK8S8+58eyV/al48peN9vKfD6NkPeUiW1jcs4pnzHVhz7fonahMILtxzmoeEvfecz5W
ZL57KST6rPSZ/+uVdko0o6AOML256C6mO8MIyupDO27gA7duhB54RySfw87/m8LoAwf3A92MWrtd
wIfZAxjgbj3joy+rLla3sMksPPB0O03ohu6faf6YSSnsuN4b9wgD5JpS9346s0My9o+LD5zonCkf
cLPbi2d2nlWCNRizhVbG7uyU3BvXTFkUt5lkm4L0r/iqfydCW/lzBcMLoe5WQwUjgNB3cMlmADpa
t8PcZr+ROF8vZ0Lq5oKydjT28npK4Oe9vE/692OUI4/j43sD9x2TnEYAPyiW3Icq6+wZls9T6LkZ
eljoc785FaLgkLg1QTRustJcWrpcrXVRT0MvPQcv/HVZVlFv65pKjDoB42OVWtQLY2XzXh4GdHg+
tnYKKnrKb8eV03x+sQpTFramgTsMqv5CArVOzMnCqG90MHUgLQLUDpeaqwHtaTWxRz6cOvutA8Q2
42RDmK2ASGLSOzRFAvPnlvtyq/jht1XJDkZmwrRx5GsFnqMMjRFXT8J1aYdZqqaxH1NdD6ax5TP6
dp+Q6oLw00pQB8PbUvpKsANbvn6jPJdawjnMIqCCVC2JrXU1DxIczAPNxd99k7F/5nbgOc1o/S6V
Ohw9lsK9sx0BsQSfo3l+qG1j+KhvH3nNIvQmVHBJVQHFgx7sjZJeJXRJJ1hELuv9J/Z66pdvzStD
MUVc7ttR6OXQER/kCWRBe/3t37Pb7NXaDryrqX2j2agCj1zPQvGaHQCrFCLVIkNCCgUnfWks0AMs
+U7iAWUBJ+us7wCvPZAObG27miWclG6iGEakFPhKpr+UtTdQoSTNb4wJk3OxbCMEd3fx4G+YnEe0
/4y9yIli99oR/jHIIMYJ56MCVBbQ7chPazHVxig31Pn09NQzdZIuNQLmHNnSpTOp936hyj13kSbh
4gf71b+i9Fw5WkfAE9nHTsBte+82Z1rBbBSAExkRu5U3cW8x2VZXlpln5/B9jDe5uVKaqTwW6AjD
3YN+pSM8bqXVkXIFAqBQS+OqqiuPYYO91VFloXmN4UHdoCKYvxzlRIsx//Sc09XC0Nts6sMAgMWQ
uU+jEv9yFRew8LHlmzJoVkDLo2dZVVYixkqjqPctigGxvVLuyuAPEI6nmZ/g05kvf7T/adDfj3HQ
KR2P3ypntSR9siOavi1S28GDN0gDPAAPJz4I0/qC7XtN7Pcmz5TYxCPXbwmvxlAU0ChWeT9PdJ7U
BxLLS5nwRFAC0s6j4ruVBg2Ha/hyZmtBOXJql17j7/DORcko8jH4WRMtvShr5sXxl3rW0/019Fy6
LmWUKmmiu0qUlfDQEI5jcy0bvOxlG04JoVAUNxlUPiJGRIARi0tp00/pwZJoOm4OdxiDS2xYXzXm
0HCBQ2RWu6Dig6lxxbx+ChplN7tNQD1HUYsR1uqWPUBOvscD4pCuoyu85kQiqL9oYqGQ8fh9LXVR
/myxo15JDg6FrJAQflzWKYsPkbuTP+wlOeWmmAU9x2ebfh2YFw5Yef0moCJF4My6VwuIcv+iY5XW
F3OWcy236e/ldqbITGwfB4iVxZeojcoThWoDSbdhYKome/ALBh7s+ZLQneSTb2jb0nnlfEdiKMxk
5w+EJxUFx5iN6nGDq6tDQbBRe3rbnCHoYu935FEJ6HuwMzcbW3ODunn8K/ftsFrHu+PbGFCmNI6u
sFCVG43+iaQSMBmXD9vJesQprwgHTVvav6KylGm9WH9IrMnUXFk27F2x6CZO18zzszdkgHD7o1D+
1cOE2EPXiRAcBzu8eZbOATTk7FxpbWUYeD0ZCsK760b7bREQxCQQmdYxp7ZrNot6DQVYuW4565nt
ndkCByY0kyoJGHp/9pCVZiRVmBg+RCEJieTh6aVjbebrogMdIlq37ZqWZXM5nmkCDPCDrK4vFVYc
ULmLxynRpJ6DZkx9e64hwP7xFUKmFU+z9jh1Bhr9H25i/MpjD3/2icBUPuAIDX1Ex9WwzrIWpPWl
Tonu7hcwnkiF/YHKBLi0FFcgDeLa6Q4GERy4m8YttL+QQ3IiWCuIrCmskpRAeFBx820cKFZkeVUO
TuzhyQ6jgdN6rzc8D1bmiWsn3p+t5u8mkqy7YluNtl4VO6SgM/ELDbfcigPl7io/PzFwOLVSzM5P
mQJaiRMXe7OKLzgCiOhaDD9/R5mcugt7RpdwF6nnt0P9+GvBy8GRfVR2tjx0SHEGqifpoc1GE754
o4NIdJ+4WweEcKSRlH9HmMs18C8hGApBmMPC+dE655vqi/2Xi+apXlAhFFUB+P+xJGoMB9Z1VKwZ
SQNMuf7xOsoSJNimy50dhg+DX+uB8hfXv6ISPZIl+5Oy9gsFpfe2yKIqFtrm9SDrJW6xKjQy8Hc7
JlqSKBQdC9apkNtmQTss4bRqCcgVZHa8YAlLtwshksYUA5NBP5iMrJjFHM9HJJktK6jxGfid7sGJ
jDwzScppHOj44+Ew3Kc3dEhrD56DnGanq+DqpHoiqxBTblMH9iBYc9FBrBuJiEl3ErEd9f101vdC
08MCpJWY5rkya5V53Kr8sK9EexZe3VPgAcHGcWMFat9Z5g+mvlql/yG0WOYQbR6Mo5NyTfDRhY3s
zv3N56VDAaU2w0smF0aviQ/Q6Wt1m3wFSOlh6lKx5B6RPNDfCh0S7npdDXjvIUHe28fxpQHRwtRj
zHWlMHRvU1WL+AQzkyrMMDjsqDVQzlBlgTosCCCTlTBtYluDzFnFVJvbEH//ddseL8z8ZfJPelku
8g9oD2GRIsYcv8C8qKRt94k3pAybD12K6XItJSPJeh4ZyPyBzjauoESIkuHt1/Udq15kR5EWG4g8
aOoXqfo0rW7jQgohAvFl6mVM6jA7xoa5ljgdhMVD4qoFW3pnu7PeoS8be79/6FC1KuVGEsTnK8Fi
4jaOVXEC2WQwEet8Tz48zdJWe39AD6HaQj4UneoS9as/Bm9vs3usvGIZnJ8ZMVDpZt6kIEc5J+06
ozKle3/bHIxN8bEs1lzdJfPd5Mj6dDLBwjJ4jEsBqWLJtCH902phZphgSm+NBcpIFKU8KOfgKnZN
jcdreGjguEmqX41TbzeA7LIEdAhTnrTabe6RVD4EQtChe0vMAB7YQW77uLluh/b5Kjcfs1yjC2k4
n3jdqJZ6+p+mZzf2SyWpZFVPHQxJLRlm5175zKU7yD7BcPH7gxT+iojwEk7iD4X0jWsyIyHklbdt
ec7eCUa3zpAPkVn66t2NUdHBBrXoQPfAklVXAfBN8lcTDCgd7/yL2l75/7d4/GFwgfQjbbNs2UI9
Txg2vlds2Oibrr+khxTm/AvY/sSFN9xCZwyYscHQDFdrRLHCNu3wOretnZy+IpcuQ06Q3HADaZwV
/IFdhCZV0NpY7zhjugrrjLDO5piaGA89lERQbO517pG9DzKYOa/tSIyL+4kVT+4fcAe8pj4ukPdA
3eW6zK5nhL1IeBa54Sirdv0NPRz5a9r5Ff+7wWVIuNJyNljkmTdVvDtTdOJH6+5de92k57+iu6xa
UO6/fyuhwiYAy1QFTKKrkjXqXBTBst1nWk8HPZPnh7HJPGn/s2vKBfu4hhWT8kXrz51eTsJx8O9s
cmt4THkriRIQdUkJko25jmeacz7YizfljixXJtXoNi+b8nPr5dJKhJ7CNOY3+nBp+Z7OlYu7YrTA
x/fzElkyVplcj9KrWVfJwcOzQP9qecNOitBgJ5i7ljhQ6VPFDtX5j9FL7ChbusIximhIp85MJJHQ
Ey/o680wAbpL9JV/j3xnyJycRx+VN7MVZq3uHwajbWjJ41kNldiaONX5cbfliDFg97WAzgaKhYrh
p4duwSjqFEyZz8/BcmItYtO+q3agh7lj8C1JMaLo5KXKncGYViJwTTVCzff6b5y1w4HrPYZprW8r
6RaYnfBX2g/5AGp6kY6WrMczndGrc3XSDV++uMCGl8IPaTlWea5/0GPjo3da29KhXHmwNieBaUL+
b/3QJOFTqfbJhvJ4+Lkl9Gdaatpdpd1B3cn6YWVHppR9sIRReoxhUgN7Sjoq/m9UGbUWooV3rx74
JGwHBxSbYW4Y4siM6ZPN0vXOvzaI3m7sGO1uKYGc0J4eNm99Preel/B/2IPlEEF2fTqJQpsbvrk8
REAwrLerSqnEu//wIneUTPIZGod2uPJVN+RybDHQzsC+XdFwzuIQr/kncUdoX4vhyeWp10QL+3P/
OGJ9+akSwgCuZ2I7YjZhNAQrVuWNPykvuVfuNGlWYcE2Z+O1AI/uZqgJ7vD6ZxF3Ad2LUOZgcyks
MWQ88iWtDZvr+/lO4bVrlgfhRIec+YesyybQyUE7/CO7dUmNk/05PvSk/0NDqI9JeHKTwb+3HbQh
+GZlIYUhse+0uQljMwYwl9/xanEe43PhCEgMl9doBinQ6ns2dvHVLo0o6tefzzwJ3HHzZmSJEDF9
wTKD7CYNn6Th+oyGb8Eralernu0acqUPuGmZmMnjVuDBRDwl1Dj5Ze4U+uNhRvEhUOAX+1IWEzcq
eK3SzQ4RgzWP+wG+afTJj42R7or9Z3hy2W1XwgixVbt4kJit9rKjULwT/dMjyvS0aUkmKTS2x6d5
h4ULSKORJR1bwwWG+xtbyLjF2+GcjWz26v76wZwNEEa/Gei+djk/OmJ/8TQ5+eCFcLR18XFxAkJk
9huMDv/n+zbu7oM68BwxqE2a4rzDd5lLETWJmQ0TOGsdC+mi6bQ3LUguUR22Nfryu1dolHGTMHl2
XfFp+R8x9mzYQ2sMdVpe0eOOc4qMv9FCdmNqPVhzCmNYN4XbG25XuYQQEBn4QwEnfTS8L82Iwa1z
2UFOHM4zLS/H2xYgrcsImoVwAlRaPq6YMInuSc+OLAYp44DzhTC1BT4QAJ/hM+ZD5ANQnuar6VqQ
eRrxFjzMJURYgWNobX7oVGNxftqJ5n+/SBn3nhJQ2t8eR9BE78GHB3TH4C6j8gv49mZh8z7kR0Ne
zb5Me4+CutX0O1r3UqkQZiuIG/54ZAEpEQNZnsKtv9DtiZ5jiwQbqr9WPB6S7I7/X2U79Qzz+sDq
1kOTzM0YJgNd3eX165yHpHEbu3GB5ZTLPst33nWvGXtcfUCo0CYCIzV5rsOx4WAJaaZ/my4ffkzn
xdUXauZHyNjIUlTGmon37zCqAuqu6Zd9y0ixHuSQw1iMoxzrmToRDfHz48ibfWhCCoRsgOM4qC5J
+NjBi3aEcd6hIZG483K2aLvfEcWkrkBF84bfiRHKJCXDDIcxs8RyqwAOXoiRK4Ne2C4h2OhnUSCs
Mec6B4bjViCpZajWc6v9A633cVBt+K0hceh3hprhA3yUenlUDNLp/+reHHzAGXWDY8vy8oMnYXuA
23FiaB/2NFh1xvsyjjtzVIQmMHeugjtxXZAqpCGYLowGNb6Qer9Hdnzw2WzehJQGl+ul3ffp6IMo
C6tJMBRz8ZUX8RfiKdW8lkfF4S00JeZYX42349UNr1JGHspTLmorXrOCUCOfMnwbdUkxrd2yV/2p
Ue+jrZcTN1zrERH2S1w65jPIqCdGC1MTsJDn3TlsnRM2tLvquIV1TT0lXyK0ieEOGcNAU/vjAD4m
FGuOcLbd+Fpb99XrHKbGhKG12ovXKNiaH39bcDfYJHgSN6uLu0RKOeTreKC0oh3kzVNe/WF4/MRF
HCfeDUu075F+5wBES4svE1uTxYYolmFtL4FBWpqx/SIK/P8H7Y7iBu3hLCRGMbrdvBD09Q8OOLdJ
Kkj4Lgr91fhf1c/SOKojf6xm6WpSSNaCr54lOOtcMy3vbFrf22+BSgguNWmINWkFsrqTe1KO9B3/
lGZg6Q4cupnRXEydnbS28XPgRmb/CUp/+YWrJ+i6eLVeRyjdL8xjcTF9OqbT2mebzKINpIWayz9y
houuCTLuXu271JaLiaPRK5ZdmPB2CaR6w6qr7QUbyUESF6rOezrFLqQfEhZZcvjx8m1zs74BU0Wc
Y5gxZLTDYXegd7ha18iN9L9zIJh/YcQVSaEMO7fHtkhYe8xPLMeem0eFuuNjLX/3HF575wd7Eo0w
OqzKwg8OFjrPyups+/fX9u985bBukxf9WLAPlwwIWzTlhDtKvbJZR4SKf86czLVIZvJUlZfNyql/
/hJnQwsyIvUuDQfIK6Z+kCvQu9CkVF0AJZD67fT819NNuyFjUzrOOcn8efjg3RuYpKtR+Ujvyfbx
EiWH91YKAMZkXoMbNExuk+oxd7Asnc6FdUttPyB29fg0yMNJtEU1HKBqyeTceeIjCCZzF2v97pUj
7hKuiBl8+KuvUWixiy+gUSAwHgmVXvRQf/rl7G3l7cIGEKPAmq0IDYYj3GGZu7/RL+afhXFyJjRt
ynGbDyPFlgp1+NPkVSJ60gffkYs3pOO0c9aU88Cqf+iObyuBMRVzu3bfWyCnytlW0QyoHInljnM1
5ELi1yQsAtxJlGyON/SpKhp8O2AYZCE9ok8qwgx9ddNvOmsplycsS0x3AUFbsCSh+kK+/RTelLuu
vRU1U5YeEXr9WCsHD5oVQdDgo05lX6yBRo9EqdsdPQmbaSqFA0v9AufCI12WBNX4/BL4vni0Kc00
/sTy7BccRNoHfQwR3rK5TmqFYoMK7QqDXIvwZjEM4jfolw4ur3rQi1zxMRGkmSR5kydR60r+TaCG
Xeg9nVL0t2cHfBkm1kI73w8pZjEsx0hWbixpS2XWhzFs4iFDyX+czP1FMhc+2eFS8uTubTQ9huM5
8/WnaopqFTUud9nrp8IgT1N7Vi/yLZg3z76VkuoKQDCp7JohQnc8lL/qp4NPnUQAevtIGASk5FZN
E0N+AycCBiXo5JagnjOxu2MGIGDw1W/2yhMB5IkkUOu2J83w5qdvoDkAI1DxR4zoc2GhKNZGje0x
nvhsz8Ant72mEgQsOXam7pTow0SVchsAAtsXHrrrR9kIdBpik9RTlKeYQz4lKgkYoIXJNLxC1fW6
3Sku3nUw3Bxgauyqq8m+yHJcvMRK5VAVNhqwnX2Sbk8uKRxlDy5zIMGqxppYT2gFVRJE0jj8YJer
f0awk63Dkr48v29Pa9b11RwWv8xfv8hVBDD3+m6D4ZOH5krH7zbgSFzvUWfUvQs/Di9rkCtYzLd1
DUg8dXhKVeq12qd2r1DsQUgA+h++0tyouvLC919zXssydBeakCrAv63vk0puwBiCDSuKvi1aMK7r
KGTbySH9n0WzzcHnyEfh6cHuPYCU8GrRbPRM6c68VKOps5cpZuF8vgnO64UcoKM/3xZVG5HArPKK
4FQtL32Z6onWhQMbjcTMiLN9txYYjgEClAAjCiDck1gFEemH2ihnHELMu3/tBc9GMjq2hmyuMn4W
PHiXu1cw/Jx6WozNltFbMrvTny9b3NDN+ko7tgcRmrdBIcGPSQOjv1GRxdMWr8L3zMvc+kKEEASP
RwM3K9m/oXanEad+sogjQSFke+/ea2MvJsokmInkwv6EzhuwYHig5k5ABB6E+aq1KllYMna7HjYH
/7iBnjMOqq6b7Otwy26otbU3R58yrUT+PnLuH0lpvW2GIcEmH05EJffTUF+GrrFjB7IDC3OoIJWL
UrX/ikJ80E4DoiAvseVgM/y7igMZ0lSfy4e+jY1aw93zpeVYc0EV4tnKP4i2AW+xW3WIfkKZmhxp
uwq2PMqqANBgPJzVQnVxLISQ9v1w29Fzj5h+Kiu0wjctAqhXTjCnB5yNQhvwUOck4z97JRWUd33H
04+tgvCX8AviGLGjWEJYnb+/+CT9yfRgPiTqLq3GrvgYMPj6/WUeZHTyOIY2ambgwkrbts7ID+W+
DI7zMy63iQrestbC0LGu+tf0XtEktpzmOBqXSMGCYL8T+uWu4jOqUPmYyCGsyCqqzOBkr9Y3C+Qx
/s/81RA9sy3TM6w+qOc4TV1qfmGj3kEY1KDYbZ/67jWdc0efDFPEJhhD6SykeHsuZ3/Qz9OPuDBE
5k1OSuDFJUTj/GVjWuFbv5pMVgonO5wFmsE4AtKv37ZctgvJJdPMtpDeRUuqpFD7VmwjN66A1JWK
2GXYuOlSppLlsY/bcUYZSnltvXeYCCd8Ma6YPqaWjsTOP3wnxXHC+ogZjxSNAJ2D7VM3gWV59o8n
L+F8j29vek48Ibive21PrxtquHJVuYt3GVuprMQU/J/aQd2bOAqH/PE3Yi+bPpRbtIQLUENhTnR5
WPmFoEUHagyCpRvd/fJbVyH5eJgb9OcKoAO8mY5Uu8Q6NSJM9jiPVyFBQQvxOxLG6agmCzgSmgHN
Ssdx8b40La+EGjEBUjDH1DjYbv/K1liMIDf3LPFnTD8BQxSii5XQqnGB520kKfT73szKGBLr/kD9
yVYpiuq1y2IsQWlbFnu7mtms/xU1U8eXS1ZlkZO1omeHrqvJN/qS5kyYpCuYccJSUVoe9yPAaKux
H0Vb77NSFrbeASkFVteWaUdPK//mbU5noU3uYXQT0m+U6F6IiyHn0sox7kKGdrxDK7duzltfqeH2
KCr+4wUgZ6KJOfFVN+G9Z514TtUDp+qh8EhTg3l2mcWL1rSYzRANkw53s0O0ynHAtWEJGDOOyj1Y
HNsBNqkh4nsOfo6O5a0g//u3AOuVKy8Vj9kI3zdrQGcT8HJLb5lGle7N6QUTUW1DR2//ubztrzDT
IsSHBCR7LlxxovPGVa8AoDK+dOdyZFadDSNh0P13aPTR6xc0pXdfthkz/WsqP2vx8lco1nIp+kN6
126uM8LRm284QSxXaemWqkkLyQzM0nbasvf+Mw8lLMj7zK2hyDdy38M6nuxhkXukcxcsPobxV6rT
MnDQVHWVmUTXnGaYo8tM7grtGDLhfKfK3RqXWvPneH7m4dpNCBnSgLXWa7be08+qyLI/OJso7jkw
6jhn+cTN1QYs+FRYEy355AZfKd0rS9HS/zkkHYLFl8OPGJntYoaP1FdqXuLnvlHJaZYcWLk0zcgq
N/PpkilhyfiegIp6O3MLXx2kERD8pIHFtJ3XdYHEDylIAqXHctZf/4TpLUC8wSUywt+4+Hu9Rell
f5qds9YJ6VbEcXhlvEj2j2g5UgEIJ+e81akuInpjcyf7Q+QK8fnFwbb/utquzb+JqzFHQgfqallZ
Xj02+WfyECXYvZWbFMARkrQy7lHI/XgxN3RR2vzZs+9DGvpisWYKJbnX8hB/WlGGbW20O3tQqg68
N1bJhZ/yrmfNguXfOpqVtN6zxSnFOUkE4hL57K0DejxJ+hosTnoQ0caQG3ypn2peCZjVjvXkEXTs
jFK2xrjuADUkOEC3TPXWNoV27lPgbhoeAAMrpzvajxuVxNbRqM2vymYAKvg+wQe4c3URE1g+XYXf
9RCYCsvnLaQk39LQW8o5fkEtqszvRIRezjpZw2jPVCqSApXcwTv7Yd+DcdWtEOXXflgoEgACfmh0
AVtT4W2V5fP9bpUtyS0xwg9QpTf3SeSxBUV4QsLHe1zZXvVcMfUfq3eYPK2W7qZgBejSzEj6U0Me
CoHv89tnJu8/NSFQ+lm+d4p6mJA0nGhHycHYW33MgLlJA1ZpFZUIrmaCyMj1w8RV9l+gztPIwgIp
HSnrzjOsUyl6vmX/IeE7YIikbfjE9XoX/8b+IUThOxxm9BpW7k7I0rg4TjzWduSzlPRs9UOShut3
vtXOlLC1LUi58qxzEk7cJruYhlwEbYFyMRflxgWntQ0T9sYB0gnDWl9iyOulDCFlJa6TjGUtR8MA
42DdMaEHe0MRrzFVw2F9sL/kPAfTwPY08kLXDG9LliI+2DEau/appK04zBTNKbat6Fwhc4Cx/W3b
G0hKCAgKEi+8b5Vtlx24E+APBEWKBlE9fevc+8aTRE2VN6e494fb6zCEEJN6w66/tTDLu/KG883T
iOtTqvsfzvkCxWAtmJ9AB68d2G3mm9+41fQxJal3lMn8t6LIF0buUznTUacaKOdLM251EgtUZXfW
J5JWCtpG9C+R5n61/M3/qas5nsQo0MjL8Gcf07N1+Xea81MBE80dFJuv1M51r6KcF6rWUueHP+qo
ocpxSLdbdhYxOyNrtQIJ0LQeHLaYmFpM+je0K0RdSlBPpRGYfMk5vL9FeaXNvl5F++bsKpvVFKBZ
Z5XSuhWkkHURGOmUJcdQgOlPq7wRzIxL2DMadEeZE05XRnd4cPhUFOtyJi3JS+4jA4+FW2fSpz2k
rP7lsnbPGqB/GSwItzwAwlYntQMLSpvEojExCWBIP/gegLe8DWzAYmoYi2VPzB5OR55R4I9YQUUZ
PVprSovQ7TGSdSdDAiGXQZisMCJRC0QKEPgF8LeBhp3ClWgrJ5V9hu9yAcMUMyEv4GPySZplGu7a
LgpSux94Rr3vX7ex4ZzjSSTFrtVNKnxyC0R7BSZfWoYaSZXU/0s++ifhYPCJurlAlhYx9TiAg/wd
HGIQtD17r6r5qXcAqGblnTnIv6mVwl7XvEzZL82ODaprFbyvWRzX8FzPU3PwhQC574n/O7XN+7x5
4mD+jqv64wMeVVkDI90c1gm+RnWsSit3XcudZ8E1Gz1xetvTAVSJcIXo+d67qyxVT+wa5vu3OLUw
rItte8nZOxwIBkbOGgwD5k9ZCjzkO1tPTGAsQjG1DTarOVSwqcX5w0KIFwGzGBYrMoxo7nniXMTZ
jmklFPE7pq7KLRcEDaIowUyxOYU8swqCZraOE3+c11KQstn9SsmFJLnUa1tjKNKovkUDZh4meZOW
jWKGwN0JwiDPqIvYgDwjip683yoF5z6dM3hHCod90xNFWoc8U7gN0d5aUhksdlFCcwsPM/WnMAxE
o+vfPr8cSYOCw4eBmLub23aekHdgqR6q/69Hv8q9c1/RtnvUdrYTZ/+TnV5Y+8wOd/XS3yln72//
gXcm+k+1RnHCcpzXgcDmj1WZ5Q5ZND56xH6J9+QbNpzd3Pk5nZIA5aDBNrgJ13qWgR/ICU6HbFGk
StQP/WArTQbbEGQei1+uYFn727/4wm8feQLTEkLTfue8iJnVRadxqlL/EzYrOx0eaMO6lCq5X4g7
2tY2vOlcHdlwWp4cyyPo0hBAnD8RG8eQBHm9061b0Y9VJuSUpbt6yRS18Ba/PVObDy/caLpng64x
MimOi3g/bnAA2PK4k03/C5KSa4qMZi5vZI06J/O6xjrYvnJJtD/Mfxe6xkQy2XUdLRBb8f/xEb1S
kYTr4HJJskuIjxxllPd0hcKSi4ET/d3fdede/EGwmtzGCzP4eHZAcwmVApxsdnW3mzErpDnTFGCJ
k5LkZ4cepfwP+5iCnmY4aNXMvSLle4JJSkaJFaEF6AP9eoQdHxbwhlreWUng8SDXejUMAicdadqH
alt3KMe6dSrKyGDs2TrWRYivABNEEFbFvTYw51cc6L5aXdkmjY70io7jhQ/Y0ZXoZIdNknFncIkm
9A3vvUhNDsUOp+gZcXPy01oacrq/ibMPlNX4427t5IdXYRqEXiI5Dyifo3WsPf/rbidzMKXrbmjw
NtG0TD4Wl5Ofx/mN0UfEym3F5DYkK4iAs3eqBrs2dTCox+nVrX2sBy3bZUM1eaReR6lLcyX+sPnJ
E3FUYAY/3BKawxGM26CC1tcgAH6YOtxnrkFJzn6UFOlG/tDXyJzcmj/Lmxqxxe3AcxNwYrUV0vZe
UY3E93YIOhCsOIV4fq+z1SxNm+txokasCxwcOGkpivQV1Z4KcfsGzzeBtvc9S1qU9UGGIxSLE0o6
YYkwrtRn/Zi/qAZNsZbeewv5OurEJx3epDRqESrf1IHYwVSPa1nZrJRRxxQCF6r+NPmiZ0TOY5Cn
nyVUvDASmtF2qdiTMBFx8mzO1AQAxPo0vGNG+ErS1uKNmI24bSD4U0qA6ienbdeWNbTY48f/nMdT
YX1f3TY9Ynxzqq+Jc1PHzZSFK3EX8ENYM/zL223GifI00UA/wIXb2Nbx/OLAWXzP9PCv96FbwBsB
S9KnSttE1oKyYyVjZWIm6u7uMxdyayezdxAGG7RmYrey/oopbQwq5OsDQPLQqJ6+h3gly2ps2IZx
AcrA01X2bGL1Xorj0ruSolgvPpYqcylx7oyKo+5Ga9212SJ+xp1Mp6xA670YZKfi41zJ0oFGGMUI
eWI6U9x061BQ+ijbQPx4uxyqi50nMP2DlLnpbpqZICyrBsAS1MiCJLRq4hfb9Lz9vqsHEZ+TmHBu
PxisTzZd7y9kYR+H0viG+0dVeBN9r6CViXKQkcTDtNzOIYb5lSGUpTd4XWo7iq3UVYVmPwc5wVCQ
iKM35z/khfBWOTzJ3zJvogaU2Fv/Lsb9AkZQNQFK9GVRwt6qguJGwq9NXU2maR1Y9sgmbTcycaNb
0krM86Oq5xjqsZpjVvWP+Vs8DZuyng0TBC0tD+lz+tphMH7M9sXF17/Vc4+AezWtL4gYBx3Pvqtm
ZJHQyPiIOJb9euDVafZ1UxGt6lh1Hxy/6fHt4Dl3/wIcUEU2rrRtnT1qifApyG96iGwo7C5Vyhrq
iop4to+UFkqRMxkywT+hlHozxR2btGvpS0sGLL03Jb6D11hh+X7M++KaZgMZWB8H+kgeNVH11JLw
EW97Cg//BYN9nT09waftcIHkr1V2vD3yjNbVoJop+w/0EoRJa14DIgyQna9KFoRPK25Pa+AWMB9t
Kk6SqaXs5rG7SesySq+5uRBgvkDZGJ1d29cr8p6V5JyCwjN+5upWk40g/XgjFwngwIKu49ASTLy7
4pGUNsyDifUS0zIYETNDpBHPAntD62Pw3IFMbt3tGZFQRFu2L1OQFQswH4aiGu8yjZlytgHRNYek
ehcSEPaogbOzLaYxWy2ILjn7jebQKki9yZb2JWKjfdoHTFEEmzpLNKL77S7kefxIvpcjXlbQvszY
kcH3D932HR8JvrBNyDHKCHbJjrAEg3a8VI1gMQxEmHIDocVgj7y574Xupn6FPlknb4qXYAom6xXP
zUbWKB57p9deTGDutjayBWVxfRg2O4C/phRbJhH2J0mDtz0+uNofBXdasoC7vXxUUr6CSgVKHmgo
6lB/obPea3yMwVaZUItLTb3CjrUJtrsanQc4Kc8403MOqQgbnU3M6cxTOHlh65JBUIu6Lztmm2wJ
6I6my1J4TJorXzr22kQlLmy9miRDcGFoZb+CtU02Z78ykWMGbGkjHIxSkv8nhmJ27RT1AuBPJtdC
S3oHoJZ1kX4qEgh3gVvdixtqo6Tu25pxARLUOVP+jLE1M4YFT4NvlobJQmlfHd05Tp/vNFoeEmDm
dLr4DmmmP2NKZZ3qwANZyiKPofTysczTE0p8Tfqh0zNzIoXRbpnqECse0XwxT7/oQI0PwqxanzsC
mmbPAUIA5xU1PxgQHUIJm8+/6H0EswElpysqrAtMzlT08BTuKAyPd6aCWyUNhEm6cjrSuJwme11G
L8GLNga5YLTMht6nNHhzVTGTGKyw7kZJuC3fr2F6UQTtLoXzdxuG8zJRlwvtpJ2XlgckCnKGUDZF
9EzV18rsRstaasuc+iFib3K5PE3r3V/xM82FUTRgzVfY3qApiJIOqqFbJZr9Jo7d9UMZR5hqi3Wx
Wu0+NhcEfN9PzRa6uBErgj+0Nj47TmBl/CJSWaDFm+VbXLvs0hfg6cS+347EjKXMd6kvZf4yqkOv
Ag8JZCm6gLQYDg4aHd3Fry5OA7MwfL4lhTt9dGT/4Rlem6L+ZkWcKaBUG2LQcViOmfKBv7PrJYUb
+u0CdlVUJSXX3z0fVcxOzoSCrC15VBD/4GjEfb3XEAFZna6tqesaCVFITm6nvLZ5TsE26TdsgLrx
6swEXRzJ6AdORShPklfRR5g6RPJbO2EEU2BhbKf51Y5m/uo4aWC7YM84haRSeE2gI3+JAo0Q03vL
3exysavbqKMr5AbS30b1BXTR64eDtyucIU+9V4B1iRGafkS5hBIcbU+rCjAfu+Hx/fTyh+pxxqXk
tAVoSZ+gprQRsWRzAMyBahrL69nXPTWHmraBtSLXtfOnEagbbfVfkX05uCuNEDvXoaUYn91TnNEu
7TGZFLzZEuSp6xEAeqA6iRx6yI4yfnWC0V+48nvOHM7i4R0LcXA4CpybMxhzDR0QIRdfC1WElnC8
5Q46jChZ8eaRYq0r7K44xagAea5zFeHDbIE0EPIZAHEAehnxD/4WtWZ0r6bg0m3X5ZlmdmeCHqY0
1lXWR79yVchrRSEoc8YZtcvAfWCc7tDqpFIWfWaPLq3f7uLFsAE1gldx2sEs6+IzzGCTl1yt8G2z
LLxJvA2LUenmkGsASkEvgSIAyj9P3hLEs/ZJrDnxRz6LLW42nnz1b4XjzEvy+nOO7ROYxOY5aNVm
V5zihQZ4UAZ8xfjLPapurpZOFPXKJzrt2nDAPkPNqZQFXPv4LV3gE67DEFdDFQozJjQx8XUDMFTC
KQ3aRWz6uZBFhrBlIAEEiG7lLoNloLQQS06ft4Gnq6qbLLLvdxAcd+NaZ1xk3Ya8RlOheFNP5U0e
1bEf3vmdznimwHyJJToggDRtaqfTBt1d+us54g5mGOCMXKCPLwRgIqxcIudB1lDb39UBI/FJdTIy
64EtZ+WF1sSXc3EJasQgiGKNEnUXxlYjlQ1WcFhMguI5gB/cRaJio0/AYuvMs6HguP5V4fhvYFRm
rcm7t/sC+jCblqcnzd1KZ+1u94DVXPPIT0qnzAbe/iqd+ExVXJ5xXIhihDF6Cun3Y8nvIt4v/cMu
llwp96iUtXHZsJaATbLoMYkHinIKErSbiAM2xgnj3/8TuqzBbi+G1IN6aTdOg6SvS5Bfce0gHa8T
k+i7IN4rEWB9zLlxFiQzWmGPWTDTIKNLc/3ZfPyjg806pXxyyPw5xtR9zbLCax2eaKfOTfyvUwZN
6R81Oow2d5QsDXqTufpbk4PpsPr2tuOpLrptRebtxtN/r1P25GWJNyu28NRMrAlDTICXyv3DME/h
B2TV24ukVZlzSJXOy4QtAW11m1ywwFsuMFZ0rZZyzbB5rJVrFMdA9PVxdQnteYT5Q2Tf1y1OxVdG
Swp4VcO3fC88RY0ShNsljA0PkDkiX/BmzRZOr+UE20XAoMzriM4qvJbO5276CVRZYXIOj719IV0z
FciV/nHmu3sAL+++xzq7mKWgkxoypLDDyqlaTlVfqh3F21GhIsWoQkMwkz9Ym1xCUvOsOoqzOsDE
Xnd2bVka1On/4iclsr7Ph3gMhytrubOAKA3KGXppsMFKKWw1h5FofTnT5sBYfjfuCa0CcfRSgoGz
lMO4QHfpeTYm5ECgamG6j4or907cKXKBkmyL0Nona/L2fKbCLepyeKvkcrjaqm+ON6ptYB51zJ/5
mCNuPIGZLBGujZprihPEoc9prFRAjRCaGEulBMBIbgA9KHPi/xqkQFjeJBooNdk1rR4VmECZA7x+
OayPIIz5GkizGGTT+gkpH7Eou+M8AhbeqlMXHIT0rocaWL8OPMXtbRA2xb0ag/9GNJ5Pj5dREZQD
rxWM+kwOcgG5xHaGtkJQs3YydXfqmemtzYLda/TVB57vTB39PTIEyPH6Urf5sMGfE0dFghvRLVzy
SvkD4JO0HFaItKtNh3Y5rB9Lj4z+RLQqLlfBJvhsWddJPjYzWRGxJPIosWhByUXHWQS1eF0putsh
oR5sIbZhZNw/HEqxS5FVo3fcOUxmwgkBkqXitkKTvFiv2KDJ+QrFBYp3Lg4DaLOkMRf6f2tHoQJD
2wYaGIeCm/vtgK4tp7JFlzCzWrb40e0xyHbE8fEC1XHpLOq6TMTabXYu79p63wCvYk/Fdf8dy34e
Y9GYjqt7vgBUXS8/sFZnZ/z/WfhQROQvtH0AaIh34kXurVBGaNN4TdXEZNOuh7ZeZFinwCHaEIz+
c6nIP5gMkZR1svdmwfKfp8/GTA/krzlgPaLco+MDirbv9neM/NLhXw3FM/+yyaNxBROQxdFfNog0
LtB2T1rYutSjzHqR3WwudgkKaT13y1qsCUNpHw616tWXiqMa9OaR8cP27X/DJNNaFDxgOeNVAeBl
b+K9z1bxrWMAPU0qlAdNhyj+3fR+v3nTA6XAVoPW+z0jmQn4q9PKf1c2IxKBnnkk14nLWP7uKERx
t2r5enl7iaB6cjdadGBqJrkd/mbapYZlPP8xUcE3ch7BLnX3etsBR/nOnKV51uxPmo3JCzHnf+pW
yrjxC4hT9oay/c6HWB7JUNb2OpRVE+4EcMoc/dKp8k8P8u2c7hXv4gy8gMwDanYuPJr0EmUswchF
aghZGmBp2lr66AM/iZvxosj2n+FVaH9jecQJyri2gWezIUJ9pr1yZC3T7fWnbJo2Qs6X1WESTjxT
x0aiZAr0UJl1ZWV8jw5DHALA10XPsx7FNsCGD8zA/4LQJgWB4wWJsGxerYQrx+JLSiQbKeRjcdaX
jonAdnx5kCrpcVOkojNGVttBEc1DyN4iY50MWD8DqQAI/eI9MM7yyMjwH7Eb8K103QeTvIjKfIU6
rONJJwXnzGirb+yqZ4MYDc2HWIGNUlGhBeY2X7xIj6r/Kyclzsmx9nOA7P0hBrgWRgiPFogvEDV/
4YVf9Z2UjzoPuFEOWt5/uiE/CZf11A9F21hEqhZP2VMlSzheC3jQvavqiRHdWO477Y8kSUqcsRDL
hdcXHgZF8J8efVBc3tlGa5QmL/3APsvCzsCfHti9hRBANz4OQcmNFqEDcjDZEf9Np481u/EyLZps
Wm0a/m1HDwNg2gkLikgsDYz8NBedQJelRbsKWpycwM025fRsDGvMsmxNrG47SF8XZF9ofEg5LMj3
/zXXzioVi7567Z5sJ+91nDODnwNXfiiUkh4UXdfRH8p+DM1xICV1FSOy3b5Eig25j5UW4uaUD0+5
HLM6fR1ILmP+7WyFKhgFDqtNDzzaeAkEmdWk7zn4Z5izp8javXC//v2OHLu21FkF+QYWtBllsPLa
PCx/AelE7/D+hHBPVfdjDbeHsb9J+6gpn8Xj5iZ8IJW7ywqhLcn9mMbFl9JaT3/Lp3JlvK8VEExI
c73165Z04LNmVegaFNoMy8HoGGHM1zzDbXfaftZ7z2cUmhyIvjfLh63Bw9xVFjgHvnIA4izdVJ3Y
moR4yPxRyDhF9VyEg+n/Vrqt1+XpXTFWNjL9kJroAt4fbXR/7S63fZZz77nXXcF1zIr1X4fzlU2L
RQoDh0P/o8yE4IPnnGhzioXP6/5CL0Xs/HYeQ2kkePkYBSP2xjkG+05VUO73Zhi/UnPJWObRIPjp
Eaf3b5eIqYBKETGkZDatpOxJfF/Zztzf4ihyhW45j+nojQd/kBYFF+iPSBPN2h0UKEp5PIYKNhBa
b39g3htS6KrUV8skp64FonMuD9rm65oXCSvG6QY7Fb5NMuhGCjkBj8P9RGBxHm6f0k36tifb8rsJ
lUW5A0vKn1h9Fo1uxoh2rTpEbtb+gSH3CRbJzF9BaXVX8A4sUd4oUav9WJ4EirfCu8mDERC5hzqC
Y50IZH9dqiVb0xYyNcuyjYKK2mWqQ/bAas2EWQMKOiC0SSeqKeaRiokF3w/fVJGRKQtVRPmHIOeV
QYN5MpBAQ4iCOXT4Phr7mmFw4VqMPnLhb/pj5bK1QQaE3TNBnTlb8Bkm3sUU3b0TSz/0ug+IovtD
zwK9WrMOflFcYsGBeGPE9chOCGgBXsskn4KjJ+VJ49x64fF/LWcjvLE8VYgfajE8awiqfhy/bbCQ
S/uoK42bvih9YZRFaAn76xbSiUAM1KOWop3q9oJ0B+M3OmJ/utmiMAIZUu7uUDaKQrdkGYqmHxBe
59GULclgFzJJSjdKufdulx9A2HGubU/SfdMF6rBdc8hEH+bKU/TUxVp3IXgRCQPusARl+kbByT9u
cIIvLkPW8iWass1Kkhw6w5Ez0kCYFruY+87z5c8X+TeOM5elcU7F1YlL7lrcdB2wPuqUYvJg/54g
gA4SSvC2MGWcBKkCwxu5CeQQEX6CV39wX3hnC2ndLuFCNP2HA20BbkVHHssdhaDm8Vd3m0jrpndf
2+xRhwtsnXypjUcM9xzSHPRh9P4paIzQTg5/VEBHieX4J3cFxfFZJ76/bnktjTS5aRSQ9HswHngb
/FmTWen7zMRC7A0tn5JeuBCFbk5gzp1JM+SdcyQNfaQrMJY2XzoxNEJRuX7QFk+wfpCwNw/aA3o4
AAWYZzxwiq9ppdm0BJ3WwBGhUAU16d517BhlqDYZRpRNYxSEoLjznlr4zfhag8J1UbMLuJKcT9UA
Khx9Ohe7RB0TMxRi6H3EjWxPcha95cIjRvKSwdRLje1h8QsvGPqm55aBFEAno4Bfe3aFbaw9Dglg
tbned0akWyWkVY60pz83lqkUhz+uE9BTmMP1FiQGsWp+rsqU6JQLZs/CuJ8Ue4Ex8ba6Qo6AfS5R
z1NfadHY50mjYU0phk1yvOox0PvHZFkvW7T4q/CYIrDSLN9iIQc+7CwXbBtTcJhq5EF14YV444Ab
WT+nVs29bmpcE/TJPW9PoLyAmVe9EklmSnAxLD2XP8oEY4XvEbDeru+WAM6KFDPBQPm4sWAydL8R
Gv7xb7u3Psy36jiX7ca3U9Wz90UXi19zl+1kwedCFrTJBWyZ0wSyAtwd0Ewvq+5SQFEuFdh6vM6Q
V/KGLDRBUKSqtnG9zSlXBu1BwE2styR0k1TlZ626fwQK8FlFQbY6pDIaAo1cF6a22iQmwEEUgn7s
OEs8IKL7Jl6QFW7GYIjTrW6dcdAGj54iQS92QyoOWmbrVyqEYWXo3jFm3Pcqw/xs4YhUHlyxQfFO
6UcJ/dT9Hi0gFagMUyIKgoS+w/bFp8ucHs/+oUjBSuHWqcA7NlplS9FQOzjxBew7JaAcVmEUb1ju
/tHSfdz32wRvcOEgCYxem80SM9NXiUKvsisEIwwslnD4hquXzr1r2WiUvKXKV9Rs70NRRZZZReF3
3zTS5snDlQqih9LsRGoySdnMnK9d4xWjqI6LtGQ7QIaZWF/1VqzBXYidETycdGxFj9ltZK/2uTRK
pK/cmGmVcomLT0Au2lo+absWOq2brpdSLD17am4g1pqQL05eIFF1riQhYdVzAbkdxyZN32fYVx7y
xYqCzA6Hsn4cRT32vtJXB7oYvD0mrVkTLljYY6teUiBnVTIDkbFnefbVCJDQdDyrsEodRhkWkATk
8ACMVEfKD2pI2cNaYrCgBJ6zZrz+UIlRulEUGPrr31XT83iseWtL2blPlxDeHn8/9Vy813Y4Far8
wD0M2NbJXaiLB+Va0wjQQe3r6nI5QLtlc0q3C81Rf2AB82Als2rhRY+zq9N/IcsnkjaOdFReifRv
jXSqyIRGho+QJFBeEIYBVjUoMkYPS5xbnwg6GUgWY0erjsvroU3wRSlCjskFwmOT6+XBoROk+67z
meQ7uXdx3vGhdbJhrZY1S0/pszizBceBMbbEppZvP5jFR2X2uSOIGxAkzewQHml/wezsknkyPZV7
bWDK+HOu2D9dedH9LMk8wGQUr020e5TakmVt9utszHSlo7efYH3gRQ5EYER1x6ik7LMsMahB4HcJ
zqbYmaRUtnNzlsaYfbJt0qr0tdKXKWJ9pfxflCLXWbnnRuRPEFxP2CTEYVFj/S2WIRc7Gx/spmAr
/lgQeMBS33GL7vw34hxZFmtZFnKIPcpy4ww585NOVRe9j9tXxwPFoIOGReflbZuXp8GHgH73H5dN
KRqqpvONCS0lVLXrrqtT7JgHEafpLaopyn2JWq+W8BPKCcxWLM2H8x4g7A2sOmgJ8Wm+vHOYQ0zp
PEwhMST0eKY5qFysDu/WmyxhPGzrAIwJgP9i+sSLcFbgY5ZTlnSCNQAvQqivTH3/XQYz1JZgBMh+
okx777f2okS6JMPp2j6gXpDIhzb+koU2S29eXTrFJoVnHo8LI/YmbNggd6xtKry5wzKpc2I4xHUV
WfEEFIAvQOPlCK/EmcTLNF31XgLCt8FZO5dpvWQOSmEvRjG2AtqFtE/4G4nRUxa1PmOVxKPZ9vA1
w1pC6+w3ILJazfxgfS1qNsay8yOi4RSrq2LOSWRMFHR45aAaXP/DyOlaTIaXvdzmwdbIEsftObNg
0HGVeXCZh+Cgh41KLkd7kuBtNy7xTKLwBXsA5a3jtqZegMCjI7+NCfZNDhfbMCe2x1XAecC4ncnR
rrqJFskaxFRy+APTk2ClGA96SQUa/3XNGob2InbuRNnw81w6gvCCbC54LrF9ckBsavM739Fjm0SX
1bnv6BAlLXHvauwDaHiR8s1Op8whiWZdsE7/h85cS0JWs5wR8uDN5omlcVqAY/9AermC1xXZn03m
xk+WkXhT4rxszPwqaO6qwM34bha/vySmKUSPw1qKiFD1CFSJ7VfvtBBqAFBFUZuOAgxe0RioxM20
sUSaVjxxYG8vakTAIXfHzdLTevgnx2OT7wUbDaPvEJJE8qZd9g8oyIhM9np772yH68v3OCqWFayu
7NOEUhTMMwifzE7x42TROpcpztRw+gatJXryJci4wsUjLp5MDxCN60jWx77e6SeCpcU7N4SLhXdl
vrqGbU9a8czheK4VVY37jwNveT93k0vF3Lop/VAkbEBGeTAWzLz/jAEW7j+yUu+6DVbCkMEGjNzl
OD7STYbbzPGeN9pGE6Qh6m1LJVZ8CRU3hjkcJoZeMQNUYxFJT9Msx7QxRcOD3wGyemmm1xoasx2k
gsqefRIvaPGhHzGUg9Dkpar5rOdTwy9Kc7wvyz8i39L2glhBuDaNmmabW9wIXO5vRE9zy9p3x0yb
41hFlAEA4os5xZBej02Y1uVJCIXUMoW0OHUp+8PmlWlqixVtakPVfuN5fPLMbQCMRZUx7PXhcLXp
zvx32HRbIW+GJcTLoZjrcvmG3I6SWZMZQJLk4GVMk6ltXTbBcB5O9Z8SVzmI0XR8s00nCi2MtjXq
7GnqwtrpYUbNfHKmrTM/0qO6I5yX17w/des3RxlgiTaniZcPajo60dEzA865XinBTnAaPO//V0Ds
cSzLnhkyIPZ65TLX+SihO5/qN+gt2SMutdzl3f51UVAk37eZCrm6t6KyYSj4gSLe3+KjVJxl9hCp
pCxC5ZpGeEDlv+lpYNCL8+QOrfCJFZhRbVBn51BdVNa/7AM3+FnrBsKQxDgZYivqPcLMJhPLd4AS
ogpdR9Fn2/jBKxYXC1KZp0byi3bt4svf3XajDiAKllpDMTXRNSjfuhdqhKGhpAv79ON8rmNDEc9I
ACY7KrFTY2c6Ja9p0T7oAx0zIpO9DLKYqaW0lR/lAOZ+KD9T1PkbgYhahm69JS4E/GnWgiaGlANv
QGeWCaQlEaDn6bvTJ1blMkVvJMUW7kW4b1GHcC7wkmFEbPYE/ST9nD+lVvGCcpWhcZOLZQJQUrKo
QRbyG+DT5xnbyZ8Qis0wZXZ7P2hJG7vEaIIpTYmFnvfY0GqV+sePh5a9wGFVj9TZq21/WbYM3AxU
Q63vPVhtq6mpxggD8uE5eTDsQfCL7Zy3d+56qqjDHOXOySj3WywcZaqsoeAwMukp1YockAoBWSo7
DGgQBFyMt9t9rd2giQ10LIqUelmeccFIZceJ2aI0HmgpM0h8wVB//E2F2+7FcVjaeROSlyHKZTib
gaw+HmiO5ZW1yYRvtqXvlrHhMujqsN4pDOUIimxRKT2RFvcqZAKl0cbDzx7+vvqSCKyq1E2sD4WP
eXVKMXqO0tJynbdsV2V7BhMutmbfjOxO101Q/Jtiial2wINmcb2bFnyMkUIyovW2hvwxvbXfh/cU
Nyf/X8+VAnzl9JYZ0nDR1FoQpv4YjlracPdpm9zeuHt7AFJPM5vbublo2bGEvnu+lJgYlCYshhKY
/ioY0gbFwI0wgjvLQjJ078X7t0VVtY1itJqqAFvKtcCt5K6EJmdOoEl7bR/A94a2oJrQZcT1g2lU
mHlQXxXDos8i7adetr8OzgvWW5JgqWxo9QijKRYNzQ7tF8+v6YsA83shsPK2/KdFx6jpbOQUVf7I
ZrW43Vl/PawUPmWYXvhTOTge8lg4STKvRjvUrN8VZMMviANQcwYoajriNdi0YAoyuU0vu5MlI024
LG2YZvJdUT7evT6/ruNdxE2tQwMXP9peiE2NP9zHzdttZt3qApGoW+TCsuq3xI0rT6h9+O71rQu4
ocHT4jxAsjoc8PMWEMiGrdxsKROKkX+FPv/m2kqK0Ze0+BDCcrceDBt7vLItRjZ3wRJx05qLWiWP
B6LTCZm/jGbeKjcx2QLMC/odmomvblM/oVjDkA5MRAZm3mynfq02FBPSXBCasW77ayrLHuRb3GPV
48Lg26cIeU2Cwa3EnBWk5Wm5U4hHI+Xe6vr0nxD/LK+K6VmpH3xJAo4/nI9WkBn37/3UJgYUJnG3
pdxrJkidkefwqXeepdt52i45SAMOpbqo1pGK52zBJovZQZ8GHM6R4JohDJa3ZQrRlSsz5yrzdhp1
QoL8tb7VxBH0XfZBGthAFE0jKR8dsw59R0TpJ5SmmjAay5stvaQelELmKzfWmrohCv+hUquqosxl
aRtbMJquzin0kkmlb0ZfJWWwssHwvzS3UvB2OXkKlVoOogaW7wuT0pH5E8/4Ji/sOmslN8SDrSYc
0+Uj58+HpUTPsjslTaqpEqIGtNWygsavipLIWob4Nrtq7XUg30gGj0JX9wdaWWnvgOGO6r6O0VJv
F3HWenIEPrbV8ntvnTW8Ir0FyzfIWEynUNlVavoP9VXMWnj2WSho+eEmbXgZF+oRIQJcMdcHWuaQ
ijucfoTuGdBi8Ekf4v8CvN9j2wi+f1xAqwie3SYt7LB48VA8cuywWyhFU9qciDjVXa44rC49HoB4
4TC7Xid+KstNIAIFuGoj+n4lXAQ7pVYdgyHwmEbsp3NvoO9Br11HHAA1xjtFsb8iAGgS0rdiRNx6
su8Vt2uah7h0JCaPpEBfWfORT7AvPCCfHj9AgyzmYFojH9RXSe2cM57V8nN3fpvsVNxegCAElHeZ
p2glE40AKqK1QXw7CIxIZV7O/tYzroZ9s6sxSVbZ4ahDorXNO/LUZw48qG8bPK0beZ4GTB7ddQE2
MBb15hBR4RqSwWsd5frhlRdOCLYJDOlh3hdAriB2PXifXHlRIjMhFaCwyrDSBUY/kSeg93XJB+tu
zdUsQLG09xYJ5W9fqxUaNoz86osEh92FTLlBY4Grhl6oXSReZrMOx5cXPx80WUVbKigObZtoFy3l
EPUl0WTrniGgdk94icZuOib7Gxw66PXPM8My3xghRMvPhrDwOU8SGEdpoPHetaoTxLBVhFDuFt3o
gl68aY6l20XVcicO3NMyuPbGoGtY6h1ZuEI9J1oPolDrBf8jJ91MeQ+MMpROXhuZuhP6qikxx8sk
PeQUFrHmmX2SYOs/hmMWOgE5CAngpcChpqZB04aj9z4MfzFsGfHgE5uENOuWbJant/JAdqQxw88l
z/19Mse1y698norY0WBinjvEuXQS5l3IdAXa9/k97qrC/SsLb1fxUOoYRZ+JeDk7ZhvTqn4VW4x/
rD9bj5oeCNA4VfnUzltta6dSMBsZZgRd+N6J6TknsiHi6RXRgIUasYzTQdnVLch9aghJ0dopdT5s
chEd0HKwFsqdlPWNkW/EtRPUEdJ3h7Vmjm7aKrsDkrruMA4+nEDS8iGgRihR9xe3Q7X5pUynVCBa
n5i6ueQuC+49rlu97iTNoelVNnNc2HF/+w97W15uaHNjBwfnAvPYsmj4GYckEJuHObT/g4vXAunc
/kAfXKJTaJ4DDUnVFaoX0A7AWcaBftBMUYpCik8Oad2ymOWD2bcgCj6MR95Elis2BHfRTyPizGMJ
i4fIA/VhdC50STJ9897n/6NEcwVlLAoSjKxYQzbm+2WlMIHu/4HjrT58RPcNPIg4tAckiVkrlANa
/A3s0qbO34a4eTgYYsQkKeIlf3IJ0wtfZuYijK+6lzF0/jrvXGfXCG8w1XTxFoUrrnLE/YnjbnqT
R/n1mFr9JuyYbo3Avz3Sfka19P4E1oSFmDV+5GswcsBm8P6DPJPZGq1rQZWG6fdkx72MncOQ8x+d
Nk965KyqkoqHliOu8ryxjnnxbtTc4YmBIMlVZfpIRGsLXuDlRqpfJ2yD5lYJ/HqvXS+r+X3qf2JY
Hj2BUljxtDkP7iK6FparSS1TaeYWObdslR9froPJYIqTdsITQ/H5OeBMnKy1Y1Ajm4WFd/mAmbXK
hyAvEJJvMIbkfbAtjizrmGWUdj0mXWD9+FgX9Sl3MNS2JG05+JkYeiKz2nXTp7qim437upsAQtnI
mmP018TGNgy54dK/9sZQUBDlTdozD/3b9qOSp3eGIjP6IaDlNJvGytsrqlqxskHHZEPpJpu+aSyk
a8c/9HtMCYo6uwW2eiAUsu/6LjD83Ov/mFK+CmAwa62fYCOCqgOrKAriRWhKKCWxwn2mfdOzLJWt
2WDyspOTQtBhN2v6ND9AqjYZCnPrGOfjEVsC2B6yXXMZfkgezTVELXncaKRigfqYy2TCSYeechC/
CLw5x899/j1j45ql8TZxZBLW0YPNM38Smc0kbuYKDWVIUbqQ+fUNZM1hUGFmeMAmgpwZ0Fg7WBEb
NVljV1u8b3ChH4ZI4JmNAsS0oh8wRl+FNSlgGS+GH89BIWb6WQouFgqmAPWGgcC2P8tEpyoC6wHb
uDs901LZTngHW3bCeehAfKp/yFOjlzHi7u13WOvnTgvGGTrXAlEgjVs2QEwLpaTn3v0ApV5ldQkx
r1xg45tEgKnl0ZXtKkyYAmIrcqYuPGtmALs6qGwuqiXP2IaFymEzckF6dpCQ4WtElmOFSV+LY0na
Y+9xmHqpkcBW+xbHD1XL9eOVshyVRoouJyf8iENSIGvA7bLlmVLLfrjoMzUF12rvZGiMLyMBqEMN
fNuuEK2KIuiSw/Nm4fVItwpF2IEqQ0o9yAL6VDGduCX2fvEaTHA2IKvXw83zhHM2FHgfpP5Vwup0
H8idmdQlWGJWHs8e9xOQe7JAqW7+GXgdJyd6rnC/YQBRxdSYcf6rrQTU2Fqy9WB+npBlGn6FR2Er
iMKpzd+q742dWhKo9D44vv5Sq/QtGJ/iQHOCUWG5WS8Ej14vKCN3ajnBc6qVaHXTQLGY0Da+7ZrU
jc9TyjWB4W161c/5214cj5gFB6KaVkT4Upo/bvYQyHAv3rUDVq3ON7u0m+kjbfyTVD1sWf/TghZo
OjI9GcVKlojllL2kcKCvkhzjTcymovrA7OYVltZb9nH7CLSrMBNAhF3kQzqd6hh9EGrPP90Eu3pf
/Jov9nPAwKzO+2Ew5jhgG6nvujRS0zEGx+kZIOLx3rFwwSphY57y0gSFkQ7EvBlizCmTtvIPJJ0i
yaUdOMWv18p0Fq10SIkVMbiy46Af01eqhJaNnwTUIQihNF/Mv6siLgFANhqku7EopJcR42WlrvcG
nEpNyZJUSCe63koJiSuLXkiU4OTXl9Z4U8gBNryfahc6DtpeN28Pz0mQmEmovU85bkp48KXrzX1m
CFCn68osEUjPLYdS7xPvhhCrmwxTwQBucT7NHU3AkiPAhmbtpb22RlHRH2Fw7NYDbbOx7zCVCn80
/j0+AIsiG+WWlGkGar/E1L83MQyqPoudEieoArJzDtDuFDjv+ZN0iJu1KTPOnjp8rHzQc/a/d1u4
+pA2PQl9BO0FH7Kb9cAMT2zUHewNtWZ9BDHtDbsnYakiLJU7ZojtnOYoJC7x76mUpsHXK23jz4o1
6YWRFTShPVmYRQ70tfZID+oEojU+QMO+0KN3rEFBMEXvK0lEA3xB5PirEkmonpwVbEbd4jb5lZNH
i9IzR76UIK2KgFlsHIvg82By6Dv/CfkLthrQfzJfVFdw3EJ3eEMAvzTmLxVP4lcVaz5x3lH6qJ1P
WpfVOQZoq89zEY8akd8WV48u/DiV6Pba4X5UXqMXoGihZprSyjxzOy1olyQi6zxWLjkSm3Xy/Hqr
8WVJztYjcXupSN+2eLilu72k601eiM15dG7ljiPQLvgnZuGZ2S50sSX1MxkiOO/FgFtyvtp211GF
R9hIZR0DukD0VY2aiPU4ONm8l+79ocTvxeQfMKEX9YfyZEpePvfJiThaSzCCJ1ntBraBeloqV/CJ
apdrFRYgnP3mU6Uud2WueV4zq/sLSmBRKNTJMJKamcqRTDH1nlFGM4fe/Cl1BkKkuGwvixBGcDD0
0WfWPhCRz9gGKuudOtsfGk0YWMpYP3p0/rbTt7uqPorcQt9P/r7SU8Xyai6rLHX4/OuAkr8/Qi1M
19zYSBGQIz5Wh+K7qsOpGVoL8FBw1z+o4pAIVa/SLlvfrwmMQJpA2WasVcdJzKEwA4NXnu/u5Jsz
nXPYd5lMgo/OWXzez4A45HgU34pjS5qmDVMv/UpSYxFa7uJ/EctC9NwnvXH72Vm/wyinvftRmWae
H3sUC7Va6HEhuMG+oZ0SZ6TIj45xfcuZpyh1Gu3vFQbI799N3vkIjL6TJ84BrUL42+LodREp2h5H
JRIJYo0Dzek38xA/kPrXJiEmWl+l/85yjh59swlinm9FHalKRa/021s2HHua5raNbfurHKUJwTGY
ConfU+UwJF5LR4d+Am3GJpsFbAirK4Smw3h60HGPrjNouOpgMFMBBfP4YyoI7J+cx4j7oWZ6QzLs
hfZZKe59HRxGQDd3Edky+Zt/6vjFc6nkiWgkzX0tMGrRfVAkzBWWGJbASWfr3NVrJ25CErOxoSHu
Dun/eJ24fN8BzepDH+td+zaxMV2lck00SVLfdDXHZb/DFelnscx9IB39nq5Q8dakj/hkV3vh8VYT
LwRPn7wPuF4YJtBU84Ozwn52B1SuNbFu4BMGsNONkbCSECf6yUeONgPa8HWhO1UMG4UykBIOff4S
8KdbQaaZuzQTrM/aBq5nlBeaDM/XQPRY8Ez4/gowZUREaArsIqy8zxtSHtcOFMC22SLr+oqAnnL7
Qo4GXs6P+0H5aj20QmsgAzNLDX/MgV+6YgMHocb3tVuFErm2IvYtKOZYZhqY8vSpv1wWre6r36dG
2XdqnycoOadYu825cmJFMtoHP918YtRbAeIIjs9nyAk8MV9sjlKl25iZVyejAxRp1PjJmgm2Ppp6
46tZwQYIoC6ktL3/UkcdAbjEQSFQRFgBymwHMeljQ0RWOIkHTW4mQR36shKvjCVm9X/C05Ta/YTJ
QxSb+/6EuBUbH8Ia3qaQs88BzrqZURh2kuvkuk0CwnRVCSWpuX3E76oDO1Pre6czfosXY43d/ks/
Q8njpSGj+kfW3yi4PbolFgrdCL1nCDoel3CMVlhqj+4WF5r7D1CgwWFCmXrChdjO3/xpO2I9rVsE
aG1joRfxneNlj5oOZ9YyfrRDtROeOgTIXDiwGSrkZo3ZVjpkmQsVXSOA8euPMX02H7YC+65ib7gE
rFqxD/1b8s5Qxu7gwrtBh+hiketkJ9k09J8CeF+AZQpir4yBfgrl0bghYeOdhSRrGMwAlxTIfAPV
+fXyPctGCKkY3rDrH8zxXY2DU7FlJL/BSZqXiY/FB8bOn714cQ2VZWN+k8Ps/MKs6rcrveRleaIS
QjHUIWmGLDwkuqwu96dQVWASVNJ+DxrMv4cqZnkstFqm6Ain0Sy/bC3n9wUogye8wJ3ZQ16iXhmD
yv+4d5i1GCiTLbWOzvUU/MaFp+mOFbs3aeXLmY+4q3rYaSu/SD8jOy5Yg8z7DhdcaMeCgNXebfEh
objqQ0SDyxRgK4e3L73jQwxC0/g+6G2U77jnMCfWTwQKxgXMMckD4N3rovZIN67+Ef7UHoLa/Ibr
JkmPwGiqhGO+xOn+FNaDgEpDGzo/zB+jusC5sUlIogc974KWohus/TMgYgvzl+FWDw0KcmXH2cY3
9F4MyCTglBLUxVZ5DQB3zYxVygiTkScgJxU0MXj1x6Xb0rFrmIN46QV8/7XZAjcgzRxqzXdyjmKj
YGSInlEt8LZAVcX2SJHjKqoqHJLAkUy4m57Q3RpZoQqoc2nTWnRSjH4kfn0PWyOGHZeHNkuJ27kG
VZ4qtW+vO/fNYLhcB1p8DXSQnykmadQ7UmG7KeiDCKy5DOWEo7cQomkmVH7A1clD1GRz9tguhJyt
GoYW7PdSY4xd7SJoF4nYg8TvxrcCgWkhvz4IEwoFfGbBscTdYpTcfZbr+E+frg6Xh+SFqHAluUI5
1N+d4jo6WwBSM8hhDBrhN46/C0CMtXx7dYRkyq1QVXZMwullEDkfe54wgKrADa3biyvU3d5hGcH4
4VIf13S50dR4xKQZZfvZBQb/nW53vn8T5K9FbSrLtcbDgyxDbobKczItn/zr9lPRO6TtFazNS21l
BBFCXKoz15+SG1gbMn9QNMLXBK0PkrXzEXIrhHsZ9gktHlsrQUsMTwLaqsY3Lr/cEHs2yzIPSLHd
a64spKBGgLndC8a/GNVlLBHJeheWy9/WCpv/4xooqt3gU09sML5fOf/IgwrsBMVLEPL9k/Zvmtpo
edfE8xumSS/zx+YLLiI3s0KpXFtzUiGc05rDFcQFS/5+IldEIB1aSHZMudkowPp+9fbAElTAQkHQ
/m0eSzjY6rUeg9rALIxdTzDne07qGCdb/lnQj4vyHoLovzRw1k+l/DkpVxN2Nfue6WSKUUY5RfYB
3jfpgq0ieVt6pzKutwkm327ZMoYVDz8LEarCaxqS9A++4XOWo+9htPo44itW+zHiOUHTm9kPYQ97
5YYetSyH7jAN6sKV9s5uezlJc4vKuMOuCa18TT9UK+W2qqmKZB9y76Ra3mBNr0BRruazspJiXRC2
Y5y7MYW8zHNrfkdDxnT8rJ+ylv+SOgf4H6UdiFkmoexp6qMpbxOY2/SXkaBFcVhFqqU2vKY1s+PU
jiusgxnVmA+Ve05QKBr1oSfX5xy950x+wGPCaYhdDvWA29TAZFzbEh+yhsTBSSrIMeuaoMDtFMsV
lkYFITvksIhHQVnM2CptnYdqnZS67Bq1x7ZRn8dEgWOlII2PB9919x+sJtZ8q/bSphX5ufw2oM24
zBW8imZPr6+NpG2YQfUOJAJotXXmRSNNJQnlc4xd82mkxGfKUUoCB5SyjfNinxVY33NluuR7ldvn
JTaRyJ28cUm9vEFqqyU2Qpqvz/oFFyNKNRSE+kkE/1Y/w5NpBFww4HBMbNE/Y5Ti9/Wxo2lnBWZo
tAa9oii84KxX/y69ZUFQkrVTYu0iI7TphXNhdzF7kL0BZobvJdB2Expxjfc3IVlNfRU6c9kgLfUE
7o/Uqfb4xPyhN4EhR8VtCk0DzFU+eKFj04niqd7VdSE3JtF5UeRz3SdnS91QZaFkYeMKMC+h8Z7X
wGIkx1T50+EHuIymPfJl1jkAcwDc2Z3HIlCsAssYoVbLyseZVOJj5JoWLzRUiLkxqu5hr7yNP7Yb
bCy3Hj0GlIzlTPNfm6kQ2qzNGykS83St7aewePmgObeheqmqxqJIkNcdY0WINE4lyKQ+Dk9PK26T
+oHn/PyzRfQKWaQ9qvHTM34D4UIdPS4s1GbQBqQfpxE4VNG2foTSQMplwBVWQeOhIUKdV7DdnpwQ
5o2dxmwjSH+pxdT9G+yV23hQuwx1jQvYD0Dgt8OEjt8p3fkXbqo7eVbIOr56eBzLyRr8GzuRn9EY
dLnC1yq5WoXsUtuXMD9i8Vm2lbNLHbX9ZLZ7A1IO70DaNljka91znHgUKwjabuiQzTyJNjqjAU93
I3HjjaEcHaXVPzrPYkW09sXstSQ0ZISeLixrOLVsTFDdMuabh4SB2Ob9Lk+q9Fal2Q1MSVrZrogZ
uP0RQfzM4IsBxFU/qx4Y6KrPuShIBRMqZSqYCgZt8xYwDV54Y8arr4sBu0onq9uRcdO6jhYlRCTe
bgJfiJQPhP8R/xeIno5Y8WvNk6ZcpIHaQeO1IHzH4zouurfS/W4f5twDzVWmj1l4xinM9FU+25Da
CrLiQqjKe9uaI2TrNZdfvPI2z/03VnpJUryo8XLGwL4lmvN/Aaz+KU2ZpqOGQA+5WGOLTIPrK+zp
KiO0TdeX8tbO9aORtWy3Osa+t1bKQdY3LIv3nYFTAO1CIdouFKegQHrhLRGjXFyDPjZHYD5Q5nZN
d7sHy9GYFDWI4XbF8wvokvAbnGFI4/OqSNCnQKJ7ar5MfpNVF9jIp6mrM1/PDbspnewu/aebzhVp
D6ih2zYQsIqhecQu1BY7ajq8eMnnfkD9yTmrnPq0iDYuScFjkxatccmh0brRnCEsvKKXCimva13u
hAV3vBN2jH2OAHMloyeh4SxUB3KGAfndEoz0w5LAjuLlPJbldt2iSXtOWif/Hl9GJfOP+aonaoRg
ezz7hzpIKQQTM4NhQ/V34GWib59GOvBz00OgoCXiW50F9lm2v1qbe5EYegg2hS3mrVHAyJngK1Aj
VRCe2NGj3/PSuq0G7PIUohgqnnc4tzT070CDutggtV51+DOX4dxeiZISSuQ6pr0IpthN9T/mhhQC
af31ep4HTk4uWEa8NeBZkR+pLSgFlB3uGD8kfERKWY42Lxnqy3XmHeJgago28ziqQTGchSpN3un0
alx5WzmPoCv5XTUchvdxIBi+JENrGCxP9Z71g0Us+I7ErcZ4f1LpcFtxY8sSY80Xgs7dvecLqfbS
erEporMLFAFtjIAs4aQMEAm8QJnglcwQ7wV9iDDsq5E+GpknLqp7T6vW4Aq8pn/LDAZOR22wnnMn
04TJ6pVlrrRsGhgYyKbSbYxkulFo7GQuhqLvasmaMDn6jseBsBWjGnMK1FFivQdkkyVKIEhz7XFv
GHgyw0vbdo5vmfC/uRlCDpPCsF0UaYpIGvv7eLGFAdv0mTTWuKL/8lRSPVtdXo7Gg9oqtnxSXTZ8
pL/m8YiMyjw3ahk4UtB1noIhHqE+5gVE5wgXslfXpWb5zwG5w8jXTH4tNqXARr2swWAE3dhL/ql0
7W9gw0kBzJPhdjo5QmFipdvpXhGLnDMZ1oDy56+hk7fnycBu/PmalTmbFlTKp2DBnsgS2WMkA3r9
BYO/vH18Lk7vg1ylPfWtCTwgnL90EfW4pHrwW6MaNSGsdiLGXuBybS+ZUz/lnMK+ivDDkH30hVif
C4kZ4tI/Z6XyMf6CJXU2oNMJkXHb3DS8M7JGOdQmscX3Tp2hhRYVhMNI/Q63CBdJjRmJK/cC2wVV
kuMt2L5g8J7mteapZgIJSjAk0sxsfQ4nNL3M8RJ/e1TU4HVVHXNZOzsd6gWwNcWiUWv3eZ/YtKgD
t3DNU1EX1zSuDCl8fVQHblvkkf7e5CFFYBM+oDSJvTN+HUalvtLsjVX5nkqzUuv5RpqVfy7j7QhE
IfT5fSyyWDWd0fCV7XvOuhu1bcKXH8OBygReFXVhRSYr+HEWwnw14XpcostwiQYtN74hZ4gwuaCu
IGz7MFojgYvb4EW3/dHhVRRlO5wfBYIf1LibXVOR7VXlXlyaxiJDh2/ZfopFrLa5Q9OIq2r0+NNZ
be065QOgoa8Q6IF7O4YBoUwg1XPSZfrUtdPZZzcLxgdry/BBgUMY92B6EY1WL66i5UHsfQnqXIdD
PqfBtQKkAKrMbPU6Wu701kfro3f38Uwy/HT86ztNJ+GZ57O9GxdhE+jrcrrCoe0TYLkgLJ3MnvrS
XoD11bWRplJ9N7c8EfKPZSJY3Rh7OFABTONi7rZg5HQKHHF9aiER6lldLuMetq9N8oMrjyJVx7xW
pLc9vVAxr4rRft7PGPuMvNoSM6LAuTpg1RUcSPBNtoys8FnSkWmb67eIr0Y6RCVXPXihqjGbVNmc
8kZyhnDp+iEYyvFSJKkF4w7A7G5weVY73HDCkV9uIaMy85Lv/huzFS+SR0dBe8eRDhmSjCe6H3LF
3MCvaHsDfpXBFDpJ4x9iM6qIkh3erKEoJVbHUq9mujsk+Jfi8w/H8+yScb1+piP0mSnTL4ML9kXr
9TolVxsatNRw/mx0T/KXxjtYqj1p76BRvBINdjo5WXfDTchhe7zT6oVBzAa/3NUs1BMOrHHikhrC
HLF82xZLC0EGlaqhRPcO+yKEDjP3ipE8UWUCD0DstSSim4v3LDknj0UXZtfqFTBAnH1CVFqkCO4P
r8/OLmboLVqcC4udG5p9CMS45fzdVZM2CZvQBZcGwuOlTLVV2L5ZJ6Yw9Hqhvd1m9DeZg27xQqfb
30FEw9HFODjWIw7ImPqMfUOo2t0HKfK5YfNvA3Z+V3GWpJGZ1Q75aop8w2/MIHhmvEzX4HRMHTEv
n9ZCCThvuWld8+CYY+OY8g6Af1M+WG7tQBFV371uqs1MpghXHdQY3Lel3ohydlVoEG/rBNoL6Bz4
U4ukPsX8TmahR6f9gpKDMgA3phfef8xm00i5IHwOIBcu9f0efQyIbZKrXZbT+ybHWS3f02ww/Qad
Mf2y2/kWpLwaeMzR67n3mdl2kiX1yXZdpY4cj3jW+goLB9P5AddjHjQ9C3CKcERRJZPfmjV9QB9O
MZ9Vm5P2tHcX1TZ1WZbi10pNqCQVmKaPSWS0U6sqi2/7LPNaLbv+Bso8Phx+cZ6aUvtzaOJELgOW
MlN3eNOBTu2R/gPZX+KCzgg81qdnAdYy5EaSgxCy+yoavIKDHvPA7zHJB4ikDfd4pdnXvyCepjVn
W5jtsFreklqutsIn8ilVow8OtwcJvr0XayLirKbuna06w9zQcDOdHx1UwTWb/ssg9xBg/Zi7ka3y
aVhjpLFzKmfv1s9ZYpHcCpzt2hrBw+IsuI+nV2A9gDk1RIulv+X8xdKjlu/CytIYS/MYFupXg/+A
/WMtQJ1FFzJUBqZ9mO2w1nhwGPIqJFnA7mNTc58aISOGtrBAz++qD5R8VSfWTGI3VFdmzIx+NHEg
Yr+jWL5KRLuvxzyEcH4CAqYLErEI4ocw7vuRvomkvq47VhP67n9tcpI68EvC5ukKA2kcLwH7LHup
x2xsCKdHhwWBSGzn+5N49KMtC4U3OigJR/9xwy+dMOWDkGf6GbVk7OOmTOVghSxdTJkfNls5zgKO
kw0nHvnntb9Ccjyk9B7CH6hsVBFUyCySoL88LJn8TELn714Vupai9TOsPOMlnzDC2BSNh5Wf88xm
jGiUdnAPCTC+9LZrxxs19fb2fWNFfg4adG7qxudwlL8ljyssStbHOeIrHWELuypVF50lOu/RPjaI
KELvczAceXhnmS0DDN0OKzAAw7bLJVkLjuaWAj/OSwltlCYG0BxoPKSjSm5HUe0GS5nQKcOxWgMF
w0Tr33NtZr09bB1ywJnoDW2SHYczVhVIOn65RHl1+1NbXgOVWG/lG1qb8asKS3fiDN3JFtLf9iq/
VzhFEtkImGvHrMVND08U9Co4j70ka0mWovvFG099AO+KEDrMN2Kkv6nFcjEyVq2WRBFbEDslFIkY
rpmNOSVS9xiW+aKgKNEq8ER8/0VNT4ahN6a5QpJ/fyuxHB4vb9wOIX/p425f5lILbguc9l56gTPi
bfgt13oygDH8DFzf/uzywJEwJhquYyy4FF4H9P9JP3cMQxaYObqho03zYeFYxiEAO7xAoAJbFfLH
jSEjZL/GACPIidPBxkm7673GRH84Y6ExxxLJah6LaDEjYqbZPjN7brQp7U1NmgeQfWNfnwEgKugQ
BIeEY4RHSFvXPCdFafKclulZv0XPKNScV49GFEux5evPtErKjKuib1V5nSW21N1vpSdZYDE6dOIc
GD4G0Tf7YJzpJ/j9vEGpAitG9gArWWB8C+4BHv8j4gL7Mt29oKrMPSC4dM//krN0GSec7lhXLTSo
Hf9SkTuyhnNZFw3LALTVl7A9rUWLMVmwG66z8Cz/zxbQKPvIGLsWivDx4qUeH+32sCDoQtcYq0Dr
3WHxb0sMVZyqueKKHe33eFL+sG9cuQZMa/4NKisOqvk1wbxFMwOCD76wXQhXN2j/EB9OvCgU0u43
O+3OEuf//DecjYCCXFpy164j8c41TDUtvi0noiQkoT4SCMVOlob8QdrGlwePlTMTECDSkhQoZLeL
fOLmLeXalE+3pP3mpsEOu9jgQ5fnW8Qiu+4hFaC5JNQYQBcWbYZjPuDbKRdsmENzbLnrXTaZBlR1
bSeBqw+WyBEgS7GabxEmQMXZxqLbooZRd+JrDym5K/48/cbPReVqrumqV2P1Fa9vWsICZ1CljKmO
YfjhD13LSmcd2wfH0tr+VM17HJs2wizkxNFz46KEW613rC6E7miV61qota44dpezt7bTIbLRWYRu
FtNT09frxhn0MEATO07aCTImDVAQeLHqHOx0hxQGQiK82GEfNbse3JhZGga2w1Alw0aGkRNmSJ4d
5by9Qc2Tl76PadgR+7s7W8oQYu2U0FSJ4nLWOG0WrkVuWZBzAiX+GUR17zTKDxXbniHLGNOhlPXv
ImZJAnhgOdnzmsb/w9RUG0qH2QlcO8dcBOzs/bsdhnjqd/+R7cAt3Q1gKg6VQNHcrRs02eIFQd6G
K+rSeX3xT+wu6SBP8nXptneE02dBNi8texmSyfAEXY9VnEZBNwHdYUCpz9TNCu8ujYKi2UvDezDB
99FRo83kA3xwCn9v4/DcvJ1ceik0bH7FE418haiLeAbVP5eBR1wpYM1FeCNFMq2wf8zVZZ2zXQDR
xXlu5VGNY6QJ+n/3ruXxIpzKZ5iJaLZ4HcZLv+Ijr4YhTHVvfRtNDHRtgCyzwiECOT2R9pRQvD3J
7NfSc6XTxuyKE5hgDXA4/rB2YazCOiQX4msaWayYjjDJ6/uajkNIVnKbEgB/DhcofmhuOOG38Q4a
lXLK+ZFxZ4A8i7YDdYFKKTjkEnmzqw1w2IiD5EK9Z1rPhqc/lxUmJYh5Pg1SHa4wlQEP7mwvDGeh
FQZ29A3bEiqTTuTZma1ziDNNqxlkj7ObbHzhFCiczf+apjlTG81sf8EHvb+AwI2cjDqnm9YmvsHl
FWwDmzGFvE6Kmk6GplPMYawUlNwzUBbWW9PSnSGGwJC2apZNPfpz206kLZ04dTFrPfGYrnAdDhqE
xMNcvmOyqdB5+DLY55iwU7MSBgUQsVz5lTp40/gBHY2iBWqZ1gJnsK4xOnclb376A8tNyKBsaWZ7
8RG47IAAR7DB2cIFRbEk373TnU74fsS3pHeZaAbLxdGXud9jIBbBZP3/B1GbTWHdAo+Zxsyr2ceo
VJGUwXg5/I3RYDZhQ1jYXbiHI/0eodA7kGlGCQ7vQgMnGKsmMZ5oAm6Tz+/QI/xdPGz2Xjh28Cln
Krh1CR3326Z1xD/WCCuly3EVPb+Zft1UrLNI5Gn5MfqAnoxaH1iJ6uj/VMMlqfuMYTnpntWsvEKG
f0w2b8DZ3fH2RlJeEV4PFjwo9ZIennu7f0CdXvfvldC6RJf3xF+j0faBGyENiL1o1eLjDg0Uu2fZ
QnyAvXoD8LGgLkTL+88uRggOgXUGCgVSBuCKsUOx34122x68T5jX4kuOeB3CltpFJGG7rL7T7V+M
hFEDcxgEzu9G7dP84iGEOIjzEQN9FDjVzX0GMbbNc727YLpLB7TRKQ+lH/lBxwiN0viG6z7Qozpw
WP7jnvKm3wC5+ds/DrW+Vp63hE7weZ7cea+SFGzO/CMlX34t8xifne3mGX96KVeLRK+UFdwlT2sb
Tu1O9aIatulBSG9fjcvP281vr/6OjmKYuz7My8LHuuFcNF8+6unX1Un1JDrYsjmLo98fpq4MPVXF
+eTS9MPMg7ZmUCjH1FV5naAWlMAft8rbZb8o3iQxzwAuN5eQscRuhJR+i2XEHGG6GBEuWu2pyzBP
KR4cynKcd6z6iTGcw3or6VPLkJF7QtOV3Ha4lwJz80bqhGN4BhBFgCZh4SMzWKhBoYwUg84feaIx
3ruxekXu/TJ12JUo/KG0d0kfetB/1dLKp4Tai+2GH1Yr8USPWoCiKkhCUglUxGwzs4cKLDDRZd0M
oXw1kj2wnR8cJf52vyHtI50HN02T+Vu5U9hxHycsTPJ4okDRR0kQqeUUlfhpomzpZhXxzYnhQ5DF
dIU1s5QKVfLLYuaHSxl4HZCkk81fp5nySV5A9NqI91fxcfm+sEokHXXY1CJI61uF/2Am40eQoz3y
2XSA2pH4a3XiMKK+Y9zIQplOQXY1AKT0lAsXZ4d4pdKzpNAkYUXBLinBGS4/+/suKYUj41JTTvOM
HVejPLspqhI68CqRnh9N4ngk38160NKfMpFRrj+nLE3bM+Nn4P0GK+tZXz7U1kYcRwblxLog+MJ1
PSMhGKK52omRFxlWChzAHMsJPbzldGRq+7hsS2Q1lKToDrmGkbPdl3kMOk4t8rXzKONBYhyFONdG
AWQxbBapSBZBrBiFVhUIrG20Z4/17erzsY09CYkL/yi29zrPTKsUgaOhfQhJPjRaXP5fzSItjIVh
wcrIpTteDPV+O4r/ne13MLcuEttpUjRlE2vm5JWKeRvUHLmpft/kgfPbDiOpSEuzJ0ubcQcsm/u1
A/gwKBBbOgK1y0bFKE8XDRY+IxkAFiCtR7wEn8dfu8P9z88QjtJ14bXzg2+GtPVzm3HJm+t5fIzu
G4I1hqMI3y61UgfYGLf0fCC3sTPcpITDGrYc5mt/JJ4lOZmyTfjzUUXGbKKpVDPPpbN8f8A1a9Jk
0eFPHib4r1lxZ//ZMMXN4zNhtJ96MQkzgSfVF1p/i3B5ZZXcIhQ6mJZCQWSEQQRbrf70qvPD/4Ci
QjOCKr0HoRqhvyWznWxJ7LqZAHIkvxjpNMMmND9H/epxB3F5gfH93kNwc2cYrdd1je1k6KwCXzhc
m3G72DC0C+uBVJtPsauYlo77oJhNN/DMb0lTfD7hxfLDDKOeUVErjPVYHBxIXbKic7J0A78ZpNxw
jriYF3gMB0kFUlhb2rVEE7eGX/RTMV5IJbBWGP4HxX0uKpJ/vbfafcFRv/Z/ULeycgZ1QAYqkQR9
EVgW3KgSi5NKLPfB954t95jyDiuxxOWnlvVej9I3tRCfIBWLHo6K5qMIWOYkjky+bjpr8O62tLol
mQYtPhKyZXtNc5XBeKd4N8YcBoVpZGpMoekERoC8/PKn0atD9u6EU0A+E49/qnhdUCPULTcj69d7
eOcgnegaLYiV19ItSindPpsJTVzck0wvwokzMJzDuS0IfTmpai/LO5vRvy0JGNyn+XujJGJOd96q
lXYuPS86LMXN07MckIiP3ANm/m5L4yVlgW4vWhaUk9SXSqS7BGSnYTy55rJFanDy36K31/dC7D27
X+xULsnmw1Q3gDT6L6nsCofZ5oh1N5Kr2ggHVHLHSIVMQuCi7iC1wCilvX8uJGCZkCflhWEiypfs
1Giq5ZmQaOJYyopR6s5Lm9CbOJ2HTbP4PtlCRsHnl+Hd8Za2KQRb5wRrZao3bU+h8R4yQWbeSxBf
dVBNnz5GgiMtEIGpc8tvELAq7QhGUpkyzcYVm9EsDgAkLclyAVEFohqK5DFuEchfe3QlcptiQA2V
44rhJJODb6kRuXMCOa8c/DbBhnDLcuVGcch4QAcIqaKIB0V94P7nDW3Pp5U3ncxjrAX23FGfFuAc
EpUi0L1IEVGrJcfn7b9AEtPw1UgcLGhJYT2dldBDAiPn9634v4elGAEwgSU2EK7kHbRghnqxCBDT
CNB6+9NUpS8GQtMaHhICbsRKk1cf+vtBrvUjQZ/64ns80FqeGsinLpRAhDdwM/FoYUd8tsQiyzyC
3loOi4qPGs76CYg6YrIb3dj4EJ5s3wYWuBkjg2sQ/z4KOonAPNgAftBLwI846RZLIZuscwYv2Tzv
FsBSwmiHU/miCf6labgPkqg+VrmZFKjljNiy/q2I9xY20WVlRkip/arAtg1UB8yrKR6zKfz2iy5q
YICYJtqY0PlsKfF2OZ40C3Qf/ik5t1UYbEpAPfkIFZOgQ1P8dRa8W/Dvt+E1l2EFON8FosCxAtwj
l3UlPz3Laf+yrGv1/3UMaRM5HRkZcW6CnWXcG04/pKa+Y7ECAb/DNWrftSc8qd6flTZYz0ZibxT+
E3QoNiJ4WFewtzdwNbrDnI3yep0HpNqr4ujke7oVZuJGwc7Lq4s/ZNVf5TSyt+FM2UmHx56sQwDK
LcF+k4i5LjgSo8DDNX4qeM9Z+dvwpXcwfA8qNPwCMR/4snArUJbNHgpVSgKdY66DVwKOVV4rIr+X
HFBccvqUEUgW38+3kMBU+cZm6KLCpwxX/1VjsPZATQtSXATgtAMpSZAe3IdcYpA85WtsqKbNzu/t
touf3SNlWQLYA4NdcVHMIj5JCOdqQIAIN+m4plevdvGdgApZHaDZ5aqsvChXiKpC2AZusHL1KkwY
0dLKVqIcVfF9RoxrdEy3uGKTYVhvQFV+3L/k5lsY9A/6EwI7MLIWIuI0TRcwU+B1eLq2X6R+Gf9e
DtnrZdNrjrXsaqaO7zjY9ZNgCUbol/bfgSSfF4ICMKjXhFZIlI1KxsWFUbGMIudAm532HuvnCUYx
aXoJRNRNbu5B1kc8Ayq/lYgwolf688jVlP8fc7EYIwsRMumfzYR27Gn+p7XS2DzuhA0qKvszv7zH
Q38mu0jJXfP3i5BlI9XD312yZSTVUE4i7flSqyeQFyJp1yBsr4Pm/UZ9QtrYP+P0hW6VuIabHfYP
S0odcFiEeF89ibcsoDv9zkzcvQbwKDMD/VhXzoyv+eNR26B4CLTBrmS+v9u4sWCeKt45/LRmR0Jb
0z9aFJqwQEfI2jyArdUvcK5o2iJDxf8ZKVPJOWcOsV/3giycYCAfrN3U5TxiySuPeszvbn7spW6a
DnckXqITwCJfmmRE0oEgehEbVGKgBJ3ZHw/Df6cDauOwXKgIDVXwunNhW3vNS0UhA9iO321dfyQi
6+dkYM4bHT0Qj07UZwfXcXWBG7fJ4C/T8y1vBIF21vMgzudEBa1XuKnpzS0T4btd0n2gPu25gtAK
0xOXcTq9PobPith9vLF8XKrBXg2xCikiL7N3xghgVP0CHapCZvy5yI2+5ANrHYmLn0z1vC30rnnb
BpCynFec4uswpzqwPHJ1R7+EqB3NZyS7/PhdTRLA9Un6FV7X8frxHFCEQHpKz9JSk9kH6L1CTdVI
BpXkP3KaONLMfZBPj6o1SKwBdRJjokVa0y3Pmcjzbtm8SkhjxSQoWMsoY2aoHwxvcLWmvAmEYX6e
Z+wxXgmbX1s0+CTreu9HFSgtJmh59NNhJAMoiX6x9oO8lOpAaidFK70uoi1A6GJsVaVIfl64I2Ak
huayDVP+KAMI6ZXcX6L5LQoxb5Y0r0xwFXkidjJXr74Rh2jFJGGc+IU1DF6oxV3ZMtQxrkrVmR+H
d2Mxs9Wn0C4TVh8UY2qa9l6sFDxcbjYzoYYcQ1U6R4skbTGhaYs4AKZT/nuBd+7OgRwYmY3gvo0x
00bs+WhsPGsrKRiFIYAMLjImSs/yNb3UuAUm2AvTtQOXSwUTdYFGlV+lZXx960Mv/OFaSgObuD8r
70p8ISAW9654R95EWNT2vvMjSc+Re5oiYYVIHPO/sN0Ang0k8vJpulvVqe0efH6MsnZPdgh3H7pd
oxinTpu5GwsnTq75RMrzO9uZp79U6nKuPahT3LB4VCJoAKSLiDY5WVEnqrPskNcFkxcmB+wDxv7T
SGVkSN2EYPcBUiH/pamQjL1MBD5Vp7ULQ9+EQY4QCLtFDMZogp2gV6lXc52EnbjG7tpjbD/Admqh
+QX3Q43zHtw2E7TUeOevUEWs8SwU4k2BA6xL/65eFs8QyEngHvoNdtImdoRqNCuRoG7qYyP2FXqm
GQPfm2/UIlZvK7rMy6X+4XNENUcZb5rLbxQLwVydj2iScvTzQFnIvaLcjQuQTfTy+0PjIzFg2NQ3
3waG1ZVzARQvNlFHjNWz2lc/yvPuXFuVEwSxYKpOPQms8MCODxwoyC7gsVPujVEAOyz10Y9Q1nMb
t9cSCbHVoL99rOd2XETjkRGjIiQj3n49VnZnFhMZkF6tuG34zFETKo9HpGk/ljRwinLbfD+th1gH
dtn54ZwUXc8oM3cH3H/oczzd5k0utm99zmTpj37cVvzEFqvyCJ8qxCPB7vzEgSFnNDG4Nqt5bTpS
u67E/MFV0mhD1UKbQMbygP4Eyn8RJGPqso9gGNyxUAKV/Dt2Zln5KeQi/wCKxqvCIfLggMmryuvb
tixebRL972fvGooNhUkN8alFpN1ynHI+AjGN4ZzZ3BrJBlWrhvuhLgm+V06/dZOvxpMMvRC1l6NY
noLqe5F8pOlCEwJnMWA/bT1FJG0DACtCbN70oD/4EmKsHGBd7mOsZwzLsPOdo+ND9/WPy5tRoqGK
8/+qC9aoLsl7gKpkzxnmQvoCC1mW0gEUE0Bawo2J8X8JRAC7RAgLNIvyhWEZX9PIh/TVGjxSSc8D
ioHOJ60rXR86fMM1qRgUBAaslS93+vRMxJI+wJ8S9BkjLAeZJ140yP2f4gDlZPe9s/qHddr5VApm
xYhPsKiO0jTgtpZGklvjB9sm9Z3cViN7DxqKCIZ3iCfiF0+J6/ehSRQhRRM5thv/ztoQ+/wRhhGW
3Z51oXtPZRuJE4lFQFRZnhJ8bo6+U+ZfNM0WOMOHzRNTB6EzwYUy6AR4aPhrXeipIqczGuB/E4lL
/fNgMGCNrZcxQsmoc3soiL+IjUYxNBmEG0oQlEeeQ/it+Y1EFPJV2q/n7IQsMDwlvLspMKv5GRj7
fek1mOdRT+ElaXJDGdVGDknzB5K6lHqAiVmqh8wPT2rd+o/UdhOH5LkvN3i4HkPyMuMfhAO/C87e
ADWb9CvA6tF1OCyCiQGCSfpKgI8axmTG1WKhEGxVLi/kznRpj829+Z2R9muh7XVDD241S3Dxcv5l
wehe/m1AukXjLduLKFxaFxXoUmQXICeIHGJTd2+YiOhslBibuDAuplq8WXsUW57F65mD6VLJBQ1C
YCfefAz6jQza/IzzycSHjDzCtui3yzuyd0fiVqnDyJn+e0XCCnpsjrpWPlqPSi1ryJyBBzHppm6u
u2v6cWHNez9KW/HMeQZVU4TgIoG/jOGG6WqmAHqRphyJc0k3m9j6sYwOH2wGVwBr50nRZG9Sj3y5
vZXarw/Tx8orl6AtnVq6fQ61hgdvsUaNtdvVkt8FBwkoe/HOlguGJCuYkBhrVEJ7TC5pnyOL1sk7
DgRXDjuNy0n28c4v1/6YVg+Cr6M+QXxzVanL35O+t7hDiYFFW79gL2HcQkZ4JGZQ9Ht7+Zi3a/Dn
FNlUNxHArs2M8/Yg4SgJHn6iVhiwUy8ICqYu/GCFpJ5niVnqBG3c+qUKW5foUsIiaOuSOl1obMko
juXsiIYdwYMfxSULpAMYhgjjRCYldAnFp1mH8JYAkxj9h0JOiRdRz3PStdnczhT0cXaLqA9zY6fp
l8fxducSdgBS+upIIUKJiq62D1F4ovU1J8zGrSM+z64haLuDxQIwgFboJwrnwjWZtVaYLSpOZgDV
StZi1WZ5drsuq6JatbmuBhOInAoSCxkRlwxDitMmaW2nB4Kx/kJe4NQzVH9DC4TeGUM8Adu0FI6I
+Rd9K+dwVQvW+K4STiJV/zxsPgja83w9LtDGgzONiv48wO38cM85AT3y29zpqNZWoFMaRQQqWIP0
Rl3NIPN66/m21TIVF+LcLKTyJf/GMkVaSMHSlnml2wr1Sux5Aw0GZuzFOs7Q/6bk276EJyGj7KAs
M8tGnv9iq03m5QTTjQH+NDlYnospe+1zpDV3WhAC6q4ka17UjltCSWDfwp+0F7Y/wROuRtZrddde
EAPvTY8gspLktjBfe+Pi7dzMVnIxb3ZlDbtf85CfjQRuQ0rESk0U+WoVN23TGdXMRiTguRcMoAcy
xDrPrP7lnuxEs1sTV9vKLE7y1vKdDw+MyQ4/sI62zNQKWy7/JrqX+jGUhCr88R0pIMPIRHzQREJl
ITymbEjqh25MOLldFbDvtE4jVJOjOOFNs4SQkmvtnqWPv3dkEF4rjpHg8ItgYxf69DntO9GOAPJZ
87zDZR4HjqQjIDxXzpQt+5BByookSrUxT8ahcUichE+oSpKrFGNwkBgxmQk7bWFiLC8Ln+/REQvF
Y5KbRZKoFsrNVGCW0B7x9gDUIL1b2k/BuN/iCker2Qy6lSNAAAp5k6Md3EUxpcfnT15fmKO9XQRd
CWiA3r8HefzSX3dyN6j/5vL5XoMctZ5sc7A9LFA4klOBJTkvlTwhSBjfwSAAXQOZoJfrakpSw2Mg
3w53pyEWF87FYhS9kMUcpSRlUtE/UMkGwQQH3hoVdhYP/QPsSa/T7+Z8GTy8ttbqJk045+0eX/4n
DV82t7rVJ2by9MyI/2YiMR7Z4YM+ez6LAr3XutkLDCkwfnVoOs5IazmiZHBDJiUiyXGmGpZEQCSh
yb9C7eEc+BzId34eb2Cr8J1NDPc2xzHkUxqu1darWHahQMHkNo6kWmZpwHwmSlBpVbARxYLb4gH4
ROK5WGR5+wrh1eMTSFT57YOYT6QoRY3YJ5ULv5IqCkI5jiwg5s1KF5u2JCQaxY9vRvNkn0htdlGS
gL16pWxmqQjO1SnQ3K5wjiCoSoiDIVIbTWbXc7KpYymAIL5xxs0V2sXOsB1Ng/9GiOGv9TRDIGHH
nDaR59ZwCqm58nGFEdu7W2UT3OxaBVRA2rY5iz1RreDTX1FaVzmq3oSrrNNear6k/UvUVLx1gEiw
kNON8KJWvpCtY3tFKw40xiE59JEam4NP5U2mUUe5gufd07+lA2Jxt1ERVa63yx4cKq0htnhgmln2
TyadihKwaUoUyDmmaoVcI9NHagl45NVdHi7BHt+89gov9uQYlBYaTBKAnMPbOwqTjaIVdkXXng6R
KTlTcshefCXB4eHAbIjxLHw9QhANkdyLvkzqm9s72enOgtgYbPR5Ul1qHRAsOYQ0ZUNvfAqn9Qal
pr1X1KGDxqR2N8q4xzAuoIJWzrvaApexWVpGfbsD15bxaM6zNcVK/0pIOfrISdYKJ4h2JMwcMLFe
O0GFvbq4nVzy/WwcIpxMfzZzkSVGSx/40mm3P21AarkeG7ckeyKax20zf88VE3B8YBHN+Egfa4zD
vSd9+rlOxDX9J8W67UhQ1T8ZfrA4+GiINgZgo+XHzPEfQGXK/qKQsBD6JEuTI4BNKUjmG0kza0uf
2B2iSxyvThJp0IOLkkYxiMHrUs9ykeBdUc0jTdaF82SyiBqA9CZ8dh3hO6/mqHxyxaI3rIQXBKSu
enzwU3602pzEmdVJjtj0iVT2BSJyxTEvq72uZUh2xzUmQbZYFHKBY18dRFKFY7yscchHJWtL+DNj
gUlDvnIoP6HrOHtwbaHxUItr3WLSXa/FfIQMQOpTnsKM3idA65dvYBCjuFwGk1WJDMwVarTopSh7
xYchL7tBPFG/w9tSY+WfH8xMnGqZ9JQj21wuhmaikFz/wcBytV87/kNakOHEdeshPw+A9DcvmT/O
cyb9uVzZMnGWs6m1gaEzFdRUdXeuyfNINDqMq0QJ6al7fA20G+EMYwx6TCwtEJgguQvQ0Yew8e3f
H8DpjoNw108u8sHuF2WrLNb/Js2tqk/loQ17aGr1KXhZsMtKu6YHYCnMrxQ/4fyBqwXnm/8yJkoZ
ucyBqTeFm7zPztE3RoiWSvYvC1XfIdu4cx+n7wyieAhV1CEyX82Ndp5avoNxJ9H0hhJ/CdiCOEmI
7krLVP0yUEHJUPztOa/vRjazqcCzIqf1m+tnkHF+FMSxyJQeyEIBaT9rYXCJzUp8kQYcI8Wu+3m3
0fbN/8lFr5gw2V/BfSnylwfgbs8e9ypYPETYIxefPG5iPFkFEYB+W2/2SFMFoiXrN+7LdWhTmV9U
2c0ntcKHHZh6Sy86klxivKfAvhQV+EX7yA3pI8W/bJnBo1W5yvju/JfViGOoSsxC9VGyhWMN1xEl
rpwAOi3bh9XGxg5Gg0g8Wa5Y07sN2XmpobPt/XzALACgrYdMK1DLfB6/cLpGY9mVbgbbZt2aiopw
PLA+352Jsodsj3aWjeGrJJXWFvLMWz6PdzB97HDyAtMMRRtpMWWWaAf4Ju6bHgPC5zBQUzVdJjFq
z6vvTdNiyrxTDMRp7HqOga68hKiC3cgA+OzHiUp99Xgr9csR14VnaFmlDDSFmZcGhr19WAvEPzQK
Hn2r5O2vWDxnFJH4I2/nGwRoif3/zFrYBE8yQyq9jrp62opVP77h2swdxU9BNcufDEYJpf6nBKVD
nmfvCj62ZN5rXt602nlyf3LqKuGFhJY1dDrHZnUEt+gsS0CFzRtXEaKxOjWrEgKlqE9Erwc0gEN7
4cU4TOkhNDB1lOnCNP475BLvTYLR1YZtR/7a2BG6QBZj8LEuvbTNCcvwM8ZkVb9bPm+3vra+dwjH
MARYbry0CwHtxn259H/xEqK9eiHPYHjjudtn7+G42BLOKE9qTObQF9AxJbuXZ5amiFGv1QSgF+9Y
NCnUgtT8bXoB+A3yd7AgnAr9FQiaE+HMSwjcM+hvEg9AWMo0lLpX9adwGYXYp+MJlypZccr+4VIf
F+hEy7jAIynqRdAHYrMKMcV+sOYHIyd0raJzEi2LaPL+tJ4ODgWUtn6M6IMO2Ll5lA8YgfXnrZSW
QwufdCqBMUxazF7O4ISSGOKKHrbEv5RFKXU8uNdGhjuW9+vVQ7dKA27UosSpkS7WKtG4x5wPQKqw
fgA3qlA+tDojBimeMWHcI7kLLYtZ+x6apAjU/EOjCM9bX+Zik4oXXetpHBHR2d+tp66UXCxicx5H
qVCP5GtJwKSpQWgcvsJRKIirQ1eSxaRSJ/v/rMx3r1/R8OLvQ/w5lDY9Xa9O5Gs+PVw/G/0dmK95
7LLS18waWwp3CeJVF1J9JPptdTG8oB4BWWAcL9MSLzNpQ0wHNnayzIjuC9kYS2ebX57NWh/3LYax
NT9Keh/7YtbHtNazABBl2yBizzdXAWta39gL/+LQICUDQt1ixe2ZlEXH5NPrmCEEUlzWB5qKE6b5
iB4eYq2azni4fsPNH82eAkibOnSUUoBkJDq4p4anC6M9snoPVnYuqfEUaS3ElYIiG5TpBQ6nKxuk
tuET24OQ0gYBn6ia0XOe8N6pww1KdjJkeX6xX3/C6GlRFFKp3XOpoH9mXmY3LtkWOpJVV5k6iOog
71KCnixTKKx1DWG2Hsgm1CaJkDCgSfrli1WzHfEpBsto5HwJuMHYvnhdAoPJC894HFC98YcYMu9w
lWU4sLB4RtgkC+UB7UPg2hmJ7Op1a9fIJ9O7eX1i5P+1luCPeokTrKDDQWYPD3N5aEROxzFNd0rl
LT/ziBztLUufNteK7RNiB/DX7RioCmCkOLwoZe7BKDYHa4JG7FVlErxXzBO447K4ZxSD+B2loZBq
+SoAwrVsUpr8IAVrpz0vdKa6TKdGGaHIoESS9qfXVmFFD597YBqA5kuJZ985kObipJHH271sm48/
JDGeKZu72p6/3eYu00YYMNR+mkWEeWBOK1dVRqNCt7RvoqpdHCa0zqHuILGifegCk7RA1YXV3raa
0QJbK0K8YfXfiSQb5/mECfh6+DbUgbnJUHL28SQg8Ti27RkVDODuuI11qld0NmTUXrObKckbpMV6
1F0WEpC3Rrf/c/S707oqWqlBSw/crjWM7X56c0cMneAArYZmkKGtUMKot4lHL7fDiYlN+04SQmbN
GaqCulDwhAwqZS/+CvWJHuWcYfDjcwTXZCLNceqbWY/7GDcIpaHjmqYjHZMyXEE7UllvzweGfg8L
HoAjhdOltdkIPTEvoNf9D4vTstXVH4OyuonFf3968Vc+Fa/b4Ma1x0icz5I7udVvgqdB9FKNyyOH
JJGXuYBvdb+UOD4fuOxy9dx4PROuM05L3vy4D6AgyUAJWzTnx6OIgSVpplKm3l4WQwNu9i6J84nC
DIIwX033bvf4YewMZeV6NGe5kMSR+vo4f3IrGCK02xCnEPxyFMs00ENyU3U42VruyCLZpl2W7R6a
2hnAnLxrX1ucJv36MVTDMdaBYYc4nSdmAsdxWLRldRA9hTxiw9kLrZNFEuc6VFJXbzj5IzpRioD8
6L7n/KG2t+skU8s5gUdcX/YEaxWIFHll6t3px70mjXjrpfxnrEdg0bl5aLgNN8UFQ5lPx0D01XJg
KPXY7oXInFuDSHfp9ExHsRxPpYx0rW5XqjBAdxBlBVrAbMF3wcfoR98ZB0l23SeKMJc4y+MTN9wj
/raS5fmYl8akP00ctXp0N2LfkdijhZOcfZd2ovjCgFl0hwKbO/iQv124yzAfZOulSsH1IJGMoRE/
NgQJC1Ue6iRqoCeGfwcnuE6NFcHQX6VyVshrihEfI16+mD2In71ZwNCsPw5W9m+Fg0u3112uqnXM
Ypl4TL3eO2BAGQZoSJtgBBbmn3bGhKqJY+hsaCjZm4ROZdUhWHi31WKZNl6hXrTtTy43u/bKd2b/
ORhyokx+IXuV9t4bEjwwvkY3fEN9Ml79WVF0Yl89/pFjA50yd+v1CQjVvT7eIoKPiAwdrqAEjpdx
B8ONM+cH8pLXbkShk+iFA1MOwPNd9KjSh2gYVL8RhgB88HN4OVmif+Gu4AricWJqZiuwUfpGGg7v
Y/ztkBwcGZ/O1RHH7dHoPCi6K6yyxGY2gcq4LfvXfVFtDBn3ztYqIuzAI1Qqu4vcy2SNcha+XkeA
nQRBYPdZeyjdV5ausWBkbDsAa+0A50FQNqEY+xECxP5VnaWZXus7f1PsAZsTfjB9Y+CSeGzYGeNi
kMJyQQMXDj7TeBPLuR+ifH65uPtgoSfewfQgZynHfT1kQCEitatl+Cb8WYbFsTYepYFivgJ5Ce6f
O0b/m0xCI3MLxp7NP67rvuk5nHgWqg4nxde516weXBIhuDBwZ4qxbF3aMXwvjXr2JwTkJA89GzEl
kBuMckA+R/HfQKsf9/ZThKVJqFwxW+0Ykht0joIhkytYlJz2pZ5qUw/8Vnm+m9SbukZ9+x1AYwL7
ABVXoVXuiou5lN37Vn1oqKz+EjLhrwGACAOWB8AUtZaQFNc+N7e7s8BJOz1kglYbvBJfFtYTVV8J
km9ZL/6kAH4bHE4iB8kIe3vhclPWsT9XQbmkBb98osR7R5JmU5/uHK9FUUQbN7v/v+WkRdSA+yRe
FzLTZOO0Ws71w4CTuqUhc9P3zus9lABb8JzOFdaV95xAb9hZhHcQceGTvmBNqoYbgwdVSFSOtjBL
QKjXalXi2VWddf+iWz2SGuQ6S6o04jyuHBBH4l4Jw8dEcuMqIt1glbqLl8lLbFOPNMST+yKaXFSv
9BtbB4sn2GdKHRv+skn1E77K53OATwQz3ny/GT5q+RbS1727dtrtCZYOLk2OWY2YX4AcPocVv6rr
MVrvXC0/qPaSfGpDc9foUEFZf8IiZVnxabUmG9/dGNYaZjaiQfwlZsCFG3yMp+iE/DVPlLxvLKv0
oH3vQaYI9KZ0G80Dzpn6pDYK9GUnKPmKqyIZwnsALwmRItIqXshWGw0q1xnoaTD2Q7SbND7AFqYv
SY/Vz+zMy5KaUjh/09Ls2pXa6fk8o2DuoT4vAULmMn255//eJb2bkuAoeI51VeWhfAbuTYLgFO8Q
9um5+pAZI3AbEBoVEY+cHn9xua3bsGZkPGaiQ6oNcoKbTOF95e1ZMhuIY1Q3YPnw39IWMpmA3wKO
YBIrYcIu18ThTM37yBUUZtzs5n16P47FJkpZO0/CNQNo/4AEf//9MsOkr9d44iwY2HZR0I2d540d
qqKTK6EjZ8yOnIILN3pXJkzCm6oOKtA34NlGzPEaT/I93ZNsOvcIpU+C+9/ZCtn2HhhGaTgn2rsO
iSplZ3XNtuvxQ6FH/jNdKbgSKr8nfV8XkI/0/luQcFDqypMEI80aiVXBXquIT2PtUNx0ZHx3xp65
s7/tHiOz9D4eEujnmIogruOD681dcO7MTXTFm7Ie1zhlOG2U9HFNnLluX2lmpbBpG4aoSUB9AZ/o
k3hocmx4DLpi0tG2WTVTYs3rxKA0cmFX4fWb+8YuNTyOcq0ioj2/QPu4QGSAzp0WSYWOLepTyuBf
oWB0n2DODI5TJvNPF/8MzpeBr41l5ImUxY15U18nnxMttAy2/Ry7FWOOpivw7PzE3Qs8i8w1LM+p
bK6grk85X4REZqpUfCLCCe/KsrHT1l35LVudG1JowtuAezKTKvRZ9gkBGpGyTebnDMRc/m3TYsKl
03/q9ZQ1vt1g+YyCU0NUtT1G7EhBT702o4EfuouJe0SkWZ/tSGpgLIUO03Pmn8Mv2yB62jWOcCne
PrnNSasWRGEjpYOf2/8dU8sjiYytHoZWAZLE3aH7/HvpW9WC+KXHRpfWPJ7ykWegPZQyDZHlnc+T
jWGtkO9+ebuBtJpOQIYTl565UCP8Xmghj9+SNoLwuTDWsQG362LuhxzapS+M2XRsYtfz2Po0z3AC
ei7vPmqSzUoSJbhzcrwL0tuZ2d7pWG7nZhtvnmL0L4sJOqExir2LF8sIiEBfFZq+sHEJtJV4XYzN
uvHpeWkHhq7RNKio64oiSne+ELeZACjozTLE/eUB38dGlEBa4UC6IHRC3x7ELhAvlMeMMp1sXfNS
Vza+bKw8aunTGbarinShjwbuerFxL5ONOBq1V/j6GcNsUnWhdeIMohy99YvCOUv3sFE7OC3tewlg
RRLAn/nqJrdTYcaYhFS3ykYs6Pjy8G4sQi/YFlQUn8lsetHVqutHSy7McT2e/kvMBkez5fdBlsyE
Pm6pDhrnD5Tu2yPTIo958wDmr6H95zkBSo0qWzurQGaDX6QUPxhJsa9hIcqBFqDSZp8fgiZP8Mbz
8y65bcDR0UPulxbtOBtUwgLOoWTvVHUXgHTvU0cOq43mSjMVYlKZ/H4SzrQcHXgJCkkA3cK7oPwY
00APBog1CcS6pjFWbCDei9qy55wRvxQJN3K3DxjdndVjp5Pju1/l4neGNqIHJ0u6zRF9Qx4W9PK3
muOVGSfp4EvykxHoW1ABcaNY8Vdmlz17WThYEX9+EwqrciVpiqwRFB+GXbSgjBMqrJ/rEIzREh3E
BNew6H4Aq+wVBKJEKbXH5gZnStapMcchX6F/5ZS3uVn5KXMT9yAgNgzqyaT89WSOYozEobpYtZ3a
R3m4IYkNQBMsekfrOk9JxmVkZ+qBVWSyTnv/EUXoCHFynrXvX9LIszU5rc7a3qjWXVNLWb5TEdPR
Vj4ZVOmO7BVbLmr9349jrpL2toyKUx7bApD7iddY9sPlNrq71HTMJbVYBtZmYt5ERndS62Js6LG+
yrabkg7eV2hV2J12WOEW00JiRCDEK8UjgBSfWZAOmYHYqiRDHJsfTV26mG4GZJ/Q/vsHNMQIRSau
NeN3m+qjGSHIPkbg7Eki1dsSjIzfALYjzPdQB9lFZoYblBrZdaFKBe5XAtrD23JDv+iG266/JJzH
Yqi09y3SJHIolvSvtq6YQ8oYPt0OxFxFgqcee7dazHOYmooMD6Z23BYeJ/3uchzzJpZdtiuIkc8f
55tD1BZzdBUTQ0mwFeS+pwv9VLTuGpInv9eW67RSE41E+PWQfbQlWRk4coMiy+U4rpre14hSxNFK
MNQc67HP48+xL56WbCdaMFkBK9G2SIyqxRB0XQx7/9t/GhetMag0b/UOAHMHUiR5paCC32qzvnI3
nJaN4nqNnnN1ifXEGLnoOXqYTR64tR4bPvoqDQow2Wm5MdbFFzyq6mQGAFHksOq5hPSomhMQ7bZ0
zoxVl5FSVOxVVvfR0v9L+UimqEyXD8bKOcig+I8bk/sI7uGtW8ftnir3F/Ht981AcIUFuimmVBct
Ks8ZJy2ZRmutHxsVmFWFOmWzXAOr4Ijgs8Twxz5grWZX106NyprdzYtOrIUFxhzd4Z1nAryk4xG/
7pjYhA03WJoC/XPOqjwYr61cXbXIg7JCL3kRPIGr1FwUPzQPB7XP66exFlS4CJXOy3zGABK3qwdn
i//mVe58P/UpDa/A7RTt4QufiqNPM5lOV0BYGdyQMOzoi5tBffhQ9W9+cdxxBvLs0i9B7N+0CP9O
OnBEiPm8020Hevnl9v29taOxQzL//jkMH2UMh6TCRUasgHO2jMMWg+fC4qBqxReR0aiZExpY+g4g
p5xMpj5Kc6FR+N0up+EPwxWVNRZK99NaFR/QHJ3xSD++D+/d+ub8ZwiBMIGyDp1s2z/J3tkXmjx+
ab1UQBYf5JqxTqr2k0LbWBXckCW84h84H7bCTO5fVO9S7Futapznzubgwsm4gtj2Zk2sSyI/7KIP
Cc7L+P0xzsAzozy5dvSM4YTgSD1p8hjyKR4hjGTAnzQYa+kYVbLOqlW2Avujjoq9OZkQDLwe37bB
ULVKKra9KJ2sPc4i9JZ03kclBuaxF431RivvX8D4f12uYWbM+matJo3UARmr39QHn10/eBHDfbKb
ZtUv21wymAudazCJ9d6QBpBJvPCw7TLobS3u5sO40V38YBMKpWzSTZV18GiIc38gsmhlhzt3FlxY
acMsSEBH5muKUSDQCYFLWm1qdUDPbJsISEhr++C++TEaZz2EnsxSKv92yyAiLYPkh3Zyk5NUJWhV
lVl02OcaUxE3MIEQnz2WwLsAA5n6E9VFW/eCqncCDXwC+UyUeFixyowvWDtUmrE8SS2BKiCPLANn
7a3+SJxcJRZP+4pYUHwWF7TDt7sS1nvQiQpvC0PcaY0Vi3zpMhwmEGLWUGznvtAl+VXgYo1iCOYx
RIqGKKL8aCySkgtJEdu+9hNwSpD0bqQsT5GpUheP308GOIo5FJ6naSF6iki1Ye7vnzVO3zDBa5EP
ktCXFaZ3B8kSMYFohQUgC4GCWjClR/1NIy4HXAsj1QuZJn5LcvQXBMF593X+35SUCfUa80qV8LAf
sdfNyqRmV1+Sr+jwjEVQY1ONYIHsO49TL8pt/Bm5eh6c4uoW5eZClaHvOgeh5NHyKijOchVk/2nD
JQ0P/2iECurzXMPInQjZVq83aB7uQbyOavPBAck8oeP2J1P90rinkYbVR+n3DD8darORHZPT09qU
7LHNc+GcINWZy5T9Kc07g7VN1bSvYyUtEeWrMyp+gGxe8ZjGtC2X5vEq1lb0toXdwMaJx6eflULJ
vQp5GznsEKT7WT7cYa+Vtiq6rnbCbkGdHyOYqHOHQzJ6wj//3sk2mcCLOR6oJsFX5kaRh7wPa3rk
+8SpBxnwxkdZ3QfjCZbnI5nm8CJuyFibq0EuU6xXpBfXUILe9NYbxFiyc+YwTVZ5UsN6mXzR+crR
BSLOvz5+wrWIvbyiLFnFOvhiYZ/PnasZ/MYlhjqK5hGR2l0L1gsf8YjleQqGz58sp7Y/GjajC1vk
9y6mY4WGyu8gC6L+RmEquV/ohjfQXpJnivqzFkjsU1ECu60XuwvlaAgkGZopyrk9079psqKK2Xqn
fvXlteuhCjYVy7ummVI4mD4Qcr7af8DH1NcFNo3t5P8VfXwiFgZOZfIJoR1sNow+WEVYzT7tWLzE
eCmACySEH7vRZ8xERFOVkj1P1QL5qgAnsMNbFz3quZXDDKFYZZ4MykaqsazTuUX32A8fN68RG3Ur
LguuMJIet/+3HxPxM+MVt7zFBWY8g8XOBdyvNLt7+saKRqs/IZyhDlr4eYJ2G9xB4zaDcHYpSLrR
tmIE7wMxTKrEZQiZrg4zGMTF4yd0KLddXgq72FIn/TBnBoaM+7dtq9rhL8zCV2rQvfvQsjoOWeh5
b7Z9voI2jI+njLN0bH0ryJJtECW2kOADs6bdXuteqzYelPXcsQfFnBjGSa/kyvfHrJQ4KAyMeQsO
d+Ym3MH9gbZPGFWZFfH4YVczzQEbhfDcilkTVrE5xvgfwVpbRGll3UVecRf0dQDT0R/gK3qRbiCb
eZYed2bbpG9HVUP6bsS0adZEJfxQMG8Nqq+tJ3EuT8RK+k6Uic25N/rQJLsyM5eAvsLxM+dxUitp
47fFooFoZsUY8xhOBZ9L1odbueo9KhrLpUtZswKE0JemdE+NqZMZI2YztMl92r2C/5ufdxerUp+i
XMJLx/htDqpYiavRbo8XzSxmqJS7cj0VmzdWCT+R/Oso0WR86YwetJzuf3b44Mg2x7DxBBbMAYw9
eTpAQ9nzRCprB+PUH6TEClM6UjwKzJfgPHgYfXc2YIUa5NhV27IA0oo7JmPHnQ0beHKTHvaOcUl8
y5aiN6CYj83qvU33bTq7mFgKpY8UjUbqM/SrGDLIAobhxiKmGTHt0oPyxPkKz50bJdr+V2fc233k
H/ltx6zi+LSGxbjZphXQ+i3C575C4NAjv3+MQevRy/Jpa0Pu8bOCofq684YkSEqayBy5DkEtLx3K
T76sHhsGRu8farqIh9TROCjhFgJmyR9ZUQUofXmzjON5lXacwUJDuztUQRk03OobJhsX0SLxEy1R
O+amIfyoT5USFiUniBpFu894IwFrKzMhYBVcv8m1sPgEkN7Mto2aDK9exT+zvWb1WVWg/66fALpl
NHXbTy/Yx5eyCbSiS5Nr/v3wqL7UqMLPwOoclx1AJMx1Yj4eQaHLJr1Zu67NBr9SXiPz/HNNpGpW
vq1cNai3jUtyKytrrd6RlVqJXJ9H2gplkhn3GsUVgWVe47a8/TO7k45Rw8OgrtX/ZibkaC/dDBXG
2vuvfEbMaLRfIK947zOI0ii8xMKnPh88JIs5w3qDEt76t0F9es4HhB/aFZstbO3Est+7q2gp99Mp
WyswzWH40oDhGv0i3l/9bXmxi1FKEE4xXuoX6awRfcRFhJ+KsnuB24yqXk+0cQuMd72g6S0fO75q
o/lHrylO3PFhAkgJM+c3g3vrzds9WsRlHOngyD1N5MzgUYkSIPSS48S0V4U+N1Il1gnC2W+vpyOi
I1Hfq0CB+uxE7nLnkGWveGod2+75gOceEukKtele7vaUS8UImYIxM3LTNszsWuY3Ovq+k1caxqTW
MmirP5iSGmSfTnxzoihCaZ7fWbAP6b/m9unx5Wy6SYiiWeufd1dCEvTTsUsuQFr9t8KwtVYef6+D
OMkwHYnMyCA74cs0KeXjq2cbMr1cmmY1mu3uBC98LpMprzwygbV36vi95TxHKrCApw0OV10KmehJ
LRl2B3bUx9xZfvpNFSnDS6T7c80Sg4RXpLTyvbR8OVjNNNm/slugT46N8eCJnWUrO3j5U24y/Ajd
OemUH4tDBNSf1swIFbWotvVCKMKsPKI5i2iOLqKgDrc8zD0kwrQRREV8mzEOsWC+yh4Xra8md1u8
qJgggYkdGsj7j18pbEh8fUpJflOvTPd3IWx9zXOtg14ar4UumAUBJ7NnIUO9ii/gpqMSfY2jNLVT
ji5YNJjYFAWbDl4cX5jPfoPHGR80DlMa57u+KOmTKCY0RVDjigBz5eyC6xPIgPgNRRWRIwFqSLHf
N2Pe+jiULrw/Kw5ho0K8G6u3VRkwd5+oUkNIYq4SHHNnLRDRL0IhZUyb+A+ZhDDdYH1mClGcyoGo
QF0eqNQfXgzp1+zZHEhuCYee85V4MChyc5r4bbEKhh141+D9CC2otG0MBciCCO/GoislprOh6awC
ETPDTWRrKFssvLn3WpTTrQ3CaTWSkCKprQk1t0GH1GCyue/w3Se3keirssj9IXE5W0ImvxJZG+4h
4WXBdm4umiVM5tU1qre/qdo/iZB+Sj/6fGLslQnQATbBsPfBPfB1bQrboOWp243DPevhOvHBr/Lp
9mHgnCtEaMfDSy+Gn9TYPOMqeGqb/L1oAplyAz0N3/dHv+EVVPTsoEkd0NYR2cnvRVm24zBcvhPz
Ylf8q3DuQc+w5EC5XuM9e1qRtJa+x3LUXg8iaH0ilWMCBT+d3gUYLC1BTvmEoCb+Sy0QdTWzCgJM
cBnKRi92PiYgQFt2V80CEkatVhUYI8Q75biy3ZN9zkKDn89PoaXMp8KvrQVpojlUgw7wQoS53MFF
6r/nnYj2eq6ljKeQG2CJDoa/tD2vF+bwyUtQGa5rJEraJb25eIAEGly2TnT+1kDChFSJc8nBv95b
9WAImcRrVY4fnJW4MibSeRjB7sW08Ftsz7pZwbQ7a7EWhsP0cxpHXVeLTZVoxkiC9IRoJhUqppju
YPj57Udb5Xv8EsSf9KcuDH5hDNUXqAZFWhVDJ6jJtQX7uNy2VOHV4jMT2kZScBCeRoKBSOvgBdCH
nwCmDmorqgmuSxEHrBltmKr1ih6D+ZJh6H3kM53JLrdmVAMf4+iDZ6jPgu+NqULYi5Lc3Cj/RkeB
OEBacqOc5pHzOwBrZi7JnqDVesPAAABLtDtwVIza9RjBM+4/B7CCFGQtEOWsFTwcyLjQf13GwNJm
FeLCtXdYOiVIt6BfD1QrYGBDBMGrLxunLJLlA4MtjJHjFSyTx7EGUNq3v6Ud4714LInwLKRDr5XS
AJWOqMRF7FnMG+EFDEVUrV8L1sTGQXN4G9iZgpQA5oDhm/JdvqiluD8Hk0CuqPFdl2m9hXFeuvCO
xSJeEQ4fMtBR/HBE3lIen5auXZDfx0UvwT95ZK6LyZYobiZCVpkNidfZ2fqUitxixkmAHhNJCl71
PtAdFBudZbOOmLr4HYb16YlaeUA94hmxCqKA6jIaU2aH+PkpU2cxkfaP21/eHXdXhA5RyKSpy+cm
KpDWjBBTpgVJZOzR3+CHTZd9vS5gz6tRmXcQOpoGIS1v0wt46D1W02TO+fT4DlGV1PJRitaNnsXV
vbJbZhKaYsplknX3ey4ndZf96fvmDk2rWOQdX4OBZIGMLC/YJDiFDkTkWYyGq0vL7aNy4DBIk1QY
7t52y6Z/60wzj/85qobhH29rBfQVc8/w50b0jIq6uyX/CVGFMVJCdFOTGXN76w5dO/imywqpX04W
Vc2e/DBV2dop95c8m74Fz/OJcla65i0c5KQEH3C0TML6rTDZnTU9s89zlgqvb7dqdPFcQNz2AfMK
p0mnDnezhwLiEfUjzCD/IquAdCtSV9ommuAptvOopR7i+0Diwlo2SOtRo/H4LHIdAbusH+ZCbMGr
0hB165U2qwlKHZvt16tk5UEQCmeCitB50yCozdb6krl6QLuvGz5sY1+LPs/YUkW5XtrLVVHeFCHQ
uE9n87pbUhZ7cX2XcNYqdKsCd1ip+v9P65uy9CVLxvaNiD/92plOjWt9NrfVreS6QzOL+iXTGgRy
A22HiuIwd0r/fG2vgsMOklsNi8NgCu7oIFyk5R/h49kuZXnebmsu9ZCsOXmIdAz1e0Xv3y0OaFKy
P1RNH384aMRoUEyk1nMyRwwiUwcWZ6gpbytHl/99XFSApgS7Z1Z8bJ4bDEP2e2aZETl4DZkaNUW+
RCXTfN+flEHrD35b4Y077A1lp9PadrEninqPZ6d7YlTV0kbxHQMQWzMlVC5/dcy6A12deQgeTazf
OfHGdEPAg4GCyKJkqvnkZw3vXcOR1JN4N1ai0DqVwr4xiIIo6E6fesTpfPPYJxzDNNDq3jorhY+x
MEKB2RApuuvoMeebOpd5/w4aOEVVDBSFwxt17ecI4D2/IcDnu0u3JMQaQrIf1swHG7In63N8xoNR
b+0yh+8Qe0M9tN6N+ki5+prRqkaIcJyQp3Fe0duKUdkj3wxJFWLIWFpE2mzUKkg7E7Uv/or7YYOm
KjTX0Nwnj1Be0fvE5jy7PUV183bj7kTw7lelNxE9BR+Wc/z7LI75DwyuTZddpnY9L54hQW4VjK6g
FFbJZjudAoG0dDatAe4J+Uw2hIS0MgPGZKvzeePfcPA9RF5vbU7cAxldJqVSpAIYNamAfj0xt2Kj
1uP4rxfutdO6Lcz2tgN8Bgd2gDwBwvEpd8mF+MjSnVCO3xtxsc4iS7unLl+v8MoOP/EJgaELl5df
IevW2UNCMKh1D7+qaDcAJbXE3NQmY9fRWxcRx0QXfgrtyDv9Ucxcz7DBVu0sd4ooOLehQAA3oa/+
CA4AAJSYvX8Fr/oTMomc53G/i1+o/ys0KwCa/h8JDecGY7d4IDFrjjO6stHAY7sXg8ksaJtNFCrw
2yIJWX9QGLrnG/EHgI0AZS4oj5irVlybvy/USxpyETyuxJ4e0KVvpoJ0A4ywBeHr3uFOE/8yK+Eu
t+wpNhwV463nLfE/ydfEc7ySD+NUO17FXEcFwqLITU3tqy49gQoyH+R422ek4rsAqcvt7Hd4sNFX
2rZxpGzYqU+0GyMGe4ZCua+yLrys2cc2IjIDLr3eRJpJQzJkqgN/ItS/zFwVzgt3hZdEiAzEsdxe
uwv3lTG1l+20iss9IZY/OtyxUMdmsWFYNXObqJYPzh+V2F++czgl3POP6V/py2X6QHbMSrHKqg/j
MN5zXsMUs6hhCAmaf+FxzsLzaSyy6IipOC1Sx+u8h/I0JUb6Lvy+Ay76Vod3hxjF9lIRG0StkzCm
eM+IY/YS3j8d5/q1XxUpityjV3jJW2UYkCa+y3BykSaOGd0BtyQMACZSDp4uobTzFU5RA5lhKhKQ
3dXSwt1VlzPSZlIlGXE2E88sZ2qFRBA0eqtenzbm7Zc8aga8vUrUsJoaCjVf8Mxg/ilFDSmNVZvu
hE91R7W2fME+B5ZSs300VRmdcN9BEgIOIm8HJeMgXcnMKcddORHZ3yQMjc2tABbYP5cihZvAysOr
+YP1xvVyyOTd/lVhWsIKb6BBS3KZjSef6ZwKL01g2bBLVONEGkIrjNINsZCWmn20reSMsvD9ciwK
Zffly8DuPnMsfDm5L09mG1/i/SAnuQLxE4g9ynPfYUuqi0uEi+1dLTy/LnD8xWO9awskMxA5PW5d
lDNa7Ui/F593V2MTQJMJmY323GWvEhRY3kdplEFtcvuhA6x98nSeV/0W6SjGlmREAWZ55E++OzYh
ZbwO9GBdGWbySqEnQCFWEOR2qcSGPP3Ecbit/oogl+3kPcUpRF+RVT3Orwi5eLndDQ8RHxvEvFP6
ay5Aas9X/tLI5ahDTA3lB2sCuU9/RcKhErT+tRDUqDRTkkJHpqGACBlZj2YXv1VBFQaqKosFLnZ/
EYFb4/aVaaAmBWRXw2OxPJvUQ/Z+++9cAl8Wcs+1bogxlBbVkVJnvXMHYBfy3HW3ArxGEWArItmZ
aqFlf80sVFHw1BDIWm6v9mqxReauvMKISvRHYdbzS3H9MdNuuBHOFUQK9X7y4/Bar6dfGHDJrDg4
fv/8uSzEPemJUUTVArvRJOwOEP57IvElvHRtiJlm1bvbD0DEYyDI7lkzFDtHZkfBfxzdDHJXvyd8
lxZezh7jo5HdxFsXiMn90WTIIY5ZEacEWlvZyvOKzTNElhHNIbJPZZgdpWTmybHNY8HRYsp9Vsf9
K9lPIv/GlKd9HBzOXEZgwlkRSymgOzjgByvOYBtmCByKYCqpazVzKfWJJe58vSxlM8UZKcaXD8t7
uCS07Oyg2nfgi09j4PexM39D9p5QNIsRc7QNktjqMi0WzRVWvJLgEsdRuw8d45ksLNA1s0Lo/FxT
/4Kn0P8RQa9Kkk+QU6C/tFSxQJZCKIL2+HewCk6FEXxUN0cOwzj7TuNOTed4KIc00M9FjP0XRnmL
T6BM5um6D4AZgESWvjsfWFn77jjNO1ZsqSHbT/NsIvus1ZmLJ7wpLp9z0msIqiiNoCd/w+ECGnT/
ynAbHNGC/ip5xEUiDsxeL7ZMttPam8AKqoLDlAwQioPW5dGaShiak6YS6ej72aVZRpTlRCMWkEh0
gV4MMNvFDSsxdcoIY6aeyrPXRNheCGC8NdbY4kZXV4nq0BgjxWr2VOPq7nG2+zBBiR6VGBfK5N72
ml9BvxS+KUYTLTbJB4CnQJFSzI9zVwGo9VnXA9sdgzZVJgbOuws6fM+D75pkCZIah6t35SlCI40m
S/bUFP+PytwkEWBErFw+oBsoOPaGJy8d/pIbZ30DMDG5IQfI/wFfzKzFCLjqAWfDq3F3K36CcwhU
SqiC5XVbNWj1W87u4C4thC8m/g0qcAgA3LOPS6w/P/3/jFBvpqkx/F135tOjkn/TFvGBx5qkuvjg
/QAGAInMCAaYTX2HGwbLBjgrcsmH0d6HFmXCpdWqZKEwgEXOlJj96CxUVLYGRKSEkkOYb3bE74Hh
M1q+nxZDk/0nmsfjy3wMNRJNLCTexybzEmUO0zHCrGrM6JtkyzUslOmUKlGxai20oY+nB1S65lHx
w56C5CAAjl/LrGZjCgyvuS1yalQvvUlXSbBWpJAxNpPtR1ykrrdn1HBwDqK2h42W1JPREmHUcsud
N5WQta/KMelshIXjPFtna7hmcIi/8Gfgdbsu/zZ99JmFVPOmPrm9TXf9+nUVwXrulnvycK21dASh
w5cYYZTUw9NOgD1ERVzHR1xdknx2Cb4fYLgGUPBD0LFPf3p6CNI21BruLcjQqUOlq8sC0V3Hb0Sy
bNWZ4lQZ+8cuQcfSTrrgUgIF7uozgQ4rdBG2OdkMzX71VyXhh3ad93tse45nsZKqXN42AlLRSE2V
vgtWUqIb+HZjpY3V5DFSFP+Klr1pwZtErL4TMlMSUoQESUxfB+4bq9ea0vkdlpGlekaDngLfL2su
eqojYzn4TfvPJBCooq8I0mmk4yQ6Xzl+1HtsOnq1so4x31pPIWr6t8MtmKwsQ0R30rIE1C4V5puh
Y4QSIKJIEx2dmJKUuQX/Mcz53+JEcPNhhfEoy5dGxeM5DpSNSbAYDKGT1bU87FCWtA6Jo6CwCpn2
CdVxR0kSlAwTzUOyd63jdB8GHo30eY1pcEnFjSqsC1dK7sj8LO550RrHujydf04mP/gj0371BgpU
mn9B07hVqRga1gakWXPUIw3pU354A5Hu9M2PPc4k5S0sXgfovpz7BX5rW13qiMNFvDXaHGBBMtCw
ESI1sOprONwS2HT8592UFSfy9kmLrN64VCc62E2D8U8/lRwkbGmaYqJE7UmXnxRuBIxIuPGsgBaG
1K8o+IOokwOeivjb4ALFnS9qYF1Pak5Oow6QAxwwIIIzaHH/lXSd7qZa9Jo0MCqTahjflwy3dg3b
vUhV2DItCqfmuPGxokfkorz9nQO0HYR9YHFBqVANYMLidTbEitDS3aQIc+IphQt5PUwjxHBXzM7k
4KI7+/qSDwLbDVRjBl8BifCtuK6Ub6bT0hKSmVvJxq6rHfV4C1Lol/GEFWjATloAwryY1Baq4H1O
w4PG8xIQAA+KnRl6ZhNGwUyHm/wKxK+wstSIVfSdX59jcAycSramfBbqaGfgBm1lR1WUGbXr8xJF
hefjh5/Ox6KTtQ0jp1e+2p7V0vIIQmHtefPHpJWQeStXTyTcRo9gAkBAtWJbcXdwQltgHEFdn5OZ
i6uGpSHGSVDVPop+rxk7aG7QFgzQPqzAi6BDRSfSVr+RZfC4cyuwJTTo4N0cfndwU0DC63o2lZjd
Fp9dMtHhT5jIcHO5Qt/sT6VRr4SEbyW+YGYHky4O5yRo+j7Ik2dcrRN9+tlx7YKcL34uwqLut1wn
RyHiKpZbpKKyCUcCgl25mlW8TSs9Te2qCIFGF1XjCAxBRGsuIi/NESjLUzoS52nM5lzWXzaG2dvI
HK6V3TtC5ybRpMO2H7d9XdXErjCHxd5eH4NB0fcmmqMTxOQCUnOUcVe+TWJAAvou9L+0+r0pAMVe
DBHZdL87Qd68WPq1E9wEi9xidf4cfjPXs2uLk3eLC5/3070X76HflDG9vFx7DDojB2hLQzm5/X4v
KU0WLR+pZ1GY+rTIDiyVMulXiJNdv1ywsnreMQOxoDi1Cw/d2RjhewS/VmpNGDo5EozZa+4wP5ty
ulYn4Sn6/EysRmU+jZb7pIsN570JgL/8kxjC+7qiqSvsaISgd7ZlIaFd1K4O5VVwHVF4AYPO1wra
LwLWEgqH2LR/59Xpt/BQZqmeRLtPWTpjhEmtVUmZiyTgoz4qC6hXbcgAj97rK+xNhUxjh4K8PFxV
DmMdqszz3iuJzRcpRuvJhvehJJubnDeiBm8cIZNYICRxe2PrsxVx2HhGMKFzFp9EwUuhDCWmS8qI
eNfL0ob5+24FgtSnqizVH6c2OVvJnGDLnFwPMF9phvQnRfwg9MNhXiAdpdgSU2sE+2arZeqGP7pi
2QoSycMjZQJXgqvSj55NeOZYmwBP/ex0kZgfp6Ecz9Vkn/2rskzq2LejJleFzQ0BirWDkSOs9OIE
FPsLDRqPJwX7iDoiw5uoHdlmHXabZKKhe5K2h20MzhBfacTc09jIFNBzQcyjmznTcKzkIqlzeRPv
nQJeKIWqoN/NLdTLLVYtTEms7Omtru8pFvqznMx1/67tlPaATByoPsQcAVaHoC/zm8+Qia/8aw/d
SFqXHjVj+GqVfUcen4yoIoYqXW7hHGB/WPTWn/luXMcbQceafFGomdLTLrKVpXkSXmUPLl7BGuGR
t/EzmnL6DKXr4epsrCk4S4d+XjzyCzJOzd7sfEVK5792P9OHLG8Qm0VF6GBSs3LPZKiEguS1QLDH
M/AivY+ywfKMpAO2J5DbXnCwKj5yPEyz4R2X6Ve8ofDDY+EMeA8bRAZBkn4wvLGVVi1HebfJm2qo
EBLGyvkMD2WPBsg2eIdEoi24uwtfWwRZ4rv/ZYVQe/fdjaRfd52jBZyWTfJrZPnW2+9ox66pXEPp
MmUWfloran8vajx6ZJyauqhkF9WO61kQPaoYRtFZucbBbed6xiDHGHHUDjfgDcyccVDrVW31uLcW
dfIcvarbQeWGgz5MJ28rvy5ZZtN7zKMgwpKAZryGH34k45KHXlOmr/UdlUXbxwRpHfnMO4axid8A
nAH7WLbfcF60arO1gnwPLbsESe5d3IA0jSetDvWm9wNw9YzC1rG2W2+DGnB4nIOcMkmGUip3SSe0
InBzf/KHWDzHKjUR6+xrRWernPZI+wtFkpTSd/FjQMans/K82sFt5urbd0PVDG2ZzzQQT8lK/A0i
+lmtgcTcw2vAFOq+Ee/bXmsHY1yG/rPqKIIpgrgNtP9Iwav5CmQd7rT0oYbL41xrfksZ0uEDRsLh
UwP4hYmhGQdkPeMsypvPLjIXvzJkRr+POuhy5jog5fTeBWoR/Rmmhke5QfoEsXp2pEO4KCFFbRAx
B/NtzYkKgXFAOMAe6DO+4kP77wjyDKR5BhddKKituk6BOrUW5fxmX87nNaoioszB/Ihc2MJsIfGh
Jqe/UydtqLoOBprrNB95EZw2sL8kTY/Y22ulocv33jNna9/U8xECh1msdYfESxhCl2KmsNCP6d3y
EdWexTbFA298totfXc3ro6rfmj820Y1qFbpKQvUipKlBdfZ5p/W1iOCsZ4IQDXmUr5At4OOKYWiY
bLlVt6ycGeWVefbkRGU2NqZ6nXGRjDiUrNf2WnSZFq308H8S/0XwkcVx5yqSLxoo3EL7qKEs+wll
7dIblWP2MC0Lw4ZFc1qxUH97UCnDYfeS75MPKH6pR8hQbhl8upHOxzCINhEDVrfc+FNWKN77sIni
6NJokWnTG4RfalNXS1hAu91dkBzTrUmGO6/Wjzg5LZGHpIxoFndbb2Twut3U8mDJOiHk1a9a+Vmn
JBSdEUj/T5aoQLBgMci4TIT8MYhJDf5wcd4ndQ6Srx/ZnE2kFSZ//WYfGDAXleO0F/juL2HLPeeC
XoId5rZMFjybHd7wHGc//iiYJm4s44tcxVbEro85NWn0KOSsnRuQwEERyQh4fuFnKd5UEswmTbP/
/R+g/jxIqGm2sZrzZxEqtrZzA+NL5llBAPPXn2CqVJJx4MhnKIsxGtUiJCHLhpscSvUTf5l+l8uV
T37uVa+nvBO56Bowq1qY4n8UHPQynGtXJWq+GGJoMQOPW6mH2jLz9VzOt3Ypyre7fkFsxCRzHtuE
cLXzTSXEwMzh9lqPbNr1gA88PBvsLhP55e4UyGFe+eXXJOJvIjgg2RjxX8zERq3o9pvelcjgxIOP
kIoYu7K0pL/HUMXfF/juaM3f0bfe6YlVZnyk6mttsK5N8UGyGnO/tNqXrfhSlFP4jDNLY0Pkmn0c
dNHjkiazBN5H0mWLO6LrDEcQecxwUNTeVtOPNLMTSDyxa9p5sfnILOh2RZxnZVibG9Be9+AP8yFR
ZQI94lGnhBJGRJpEYqFdDST3gcv1WsP0BTqy0KTHLKF0b1K7eK83mbKuDx6H6uSgmZXc2nChwpCo
qSywbPUwNIOlF0n2/xB9mJ13cMdQcZLds3nr5pWXgZKxiphJcyQroJmICwE9E7WSZ1csp1wZYyuA
XhtP9fabHchDKsdcCy/O5Co4BcETOEfwwg3X8db6VsrEhE5Ol24iXisaZXRj0KnbcwOkrFDiGmvt
f8W1J+hcVpx77V3c5WhFJHDhPVgfLrYhShiXXPLBbVaYR+1msYPShkZ7wQOcaHkRpadu/rNKw8bR
+53yokbKZOE8dD0dv+asuDf0j7XyiYx4DRpQiRlggds4i6YpnEUJNcTDNjM70tt12yTPYAtmGxx1
FE0ZvU8QHuwp88umIAqW1IVm6tsWaz2lc5h7WJdFYRwWrYPxYFNGWhDxeiWoPsFpHyTGqmHchS1R
NSiCIno/jwyJTGzk2VhKOXB6213hTJ9VU9Itll7bcUUcl6/qo4pbdFOSs6pUKRjkQlY1aP/QmP7G
6YqLpbopjBAfLFYeLHdprLqW9VSjZG1CRH2kNwyTOLLhG3fdL95UVQIQRpJg7YLGt2nMb5fEs353
HZxT2VSbZEbs9gnFeiTExMUFI2SpZdZNN56GXMDTWISWND6mYrOSslAgok0xcxoRftAmvrlOibE3
xv9tXDfOacqJu0YweDSb7DJxmi0y6K+/J8X/7Qgi+iBiZXVNtg7l0SaBRnCqZDGzO6MQIR1izD4R
IIuCHBbucl23FB53fX92Jj3WIhisW/lAW5DPyTZK3zqubJPx9BBVbm7f4OLioLQmwUnzx3eB13/l
lYnAOKqvIQI1tbLCcFYbYmXiYbm8K+Fwhu6OfEbL21Pa4ijk1J59/Pw2odhL6fD65yLnr+BQwL+I
oaiYtn7XmvUoj6tbVvVzJJCbJA8ovNTBc5H5NrsOishdz75C9s0c/3xBVEvvIzHcA6dItJBhCqRM
rDDkWFNu5D1HQsKRDXqSIqAVE/QASfVDELaG9Qn67/7OMFbFcVopZSivL+SMBgqPJoCZSSdYhrDP
p5WQN0FvpU4dCbwJQ35pJ90tj8PkIjIZKb5FjfwtqCcfFtLUUl2EkCR6JNi3A/+BdwuvXl2NQL78
woXQWKkmZB10c4wlA/t5i72iIND1cgkME8IdYujErQfIuRXSXTJiETFkBmxhiEPkmpNZDUcTKXsj
jFsiiZI3iOVnCQRoZqE9D6VSiG/uTfhotPOuxXaD+rUDHNWGggNJFTWKYKB1s8UtHmlADxn583s9
mxgOCndDBCEU+LdJm9kJBhNWYI7OnEnkBTu5MBSIaeifq55wbjZcfg8WMoJYmlNNc8h9vtoFDhUb
ZXhG/PaE9rf7jE2xM+D8zeKzqvdweSoOgEBF6QsD65k4M0BkQBgD74CniZLYGklDF6p2SZcB2L5z
eMC4LnWy0bI1+KzPJ8HxL5xw3tp/E04RV+J+fmEh0HA0PMjimiGyPbmm7A/4Y2f7QlQXgZABE3xQ
Vq9SkhaEMKcv6+8S4v4OcCE8t9p83hLtvpgHvy9eed92yp1xneJIEUL1Aj/RzZ5dkdPE4cspw0sl
Xtq14QRVoaN5H8J9vCvVGSBMbYXPOlms5ajJMrtafu6/uapaRFwRuSa28ei/C4Ek9fncrAmVyeBK
ryg8mZdyL7+h9QjfYQ388CeDvg4Rr1phe/JgES+HUxM7lAo0CnGoPJRtjCCCu4QiO6kvPXOfZFYZ
ry1efADjLY7Ae1Ndnpi0i2IDJPY0JRAmXgA9QYS1C8O3hf3mUgZcrEBMzGWC71C/sGLtVMhgijUT
9Nu3Qg0M+WB/5hwMl7sVJfg4yPSYrG8mpeVJHAn+/nWkzlvzOA/9sw+U6EchJX7Rarb2xbD4kOUv
WCw9+AkspXGcv/l9IbQN2pOEIpBXFodUUGr+V6aQZQYPWjV7SI1A5dB6rK3ouh3LdO3fOKzQANgp
r+tPLqs+VgY5Zhqf8DY2j03EFUgdSiaQIOfsKk6syTKgJBntITczg6Ft22Re0LWhvbbE3A+utUQf
+hGWH+2bqA2iOLQYL+OZO6S7b0W48ssxiFLEcghDYGInTHFyuTSt/5VBp3sCfcyI1B+vrV0TKt2j
MW5TbJmDzPZmpeWJnOs3a41Z4+ytqFYtuozFh+kQRoGDDVzKLslig0cR/irweVUJsmFN8/EnnG6U
D9rNTleCC9n7hKR/pA1D1cEgLg8oi3P279Xsx09MyJ1u4ROU5D2vSWgUu3MU0iwfETxH7BWPSL5K
jKeUjqqxstaWgrAr0cP5RGTJEGYRYajFv5TjYSKA4tWyjeXmt5ziv0AxWWr2IE+aJ73uhpdp5ija
dJUiU88TLL9o9c2xPAmvEsHubeP/bXsE7jGXJLkP2b0cG0skcj9aI2cU3hFm3IZhPuGyIM3SoAE2
x0GZuGjnNOFClIud0lWw6dIpPLzK8ufcSsBPBoDNbW5JE66kaAEU9v3u9hxs2XbxdhHmpL6eG2DU
KhJdgRsgryc1GtuFOK08SPVFA4cTbw5Mb+emuigKHzRuN0FXz6iOvHjV/4sXdMNSR6iVPsU85PRH
RD4oGJAkwQwS2/pFLH0cW9b1AQq9ZVLVt8UQzWpICaZHpw16wDRzVFiue1JMmMF+MhBMonTKMBm+
aaqSzPNo1oTP4SuILgUhXxsAEKodW7yhIPGKUfUuRRvH9Y2kqxMoy85h5gGXtQZ5IAven62CyJEw
bCvZnf2CrsjZhSDU5zgCcG/FzEdoMm0REa4gfKaSkOT8EaXgIIJwuGc+8M5LTccddeLoSkowhV5H
cy9vbCXLXibCBhCZ+yKfZ6Jgtw4VeDQsPVYQJTIuqadccw2Tg6UZwU1/iUqvWSlwe/cu37DBR+p/
p65o/9JLH2eP/1wErfWjEHl2EeF0leCgwC/E8qFpmMpzQ5TCc77mMBTuGFxATO8ddxewaUa9v7ll
+QUu6jKRv3ejnhX0HLT/lLAbnQqdCZ09V0bW/TXZEgbjG9nWBh3yT71aez/uROnNqR+j3/4std/P
x4pMFMlHagguwYNPTNNdm3is7KHVz4X2um94wjVfyfsYvjqEZVnqbyw2FNDTFoJeIu+B9fK+ksSq
If0SwV7ghFnhlG3IZ7CA6knMB2sDNZxuXSvZZZhP/0HD7XNCDB7qzMz0FGba0EKZzD6Ft/+VuuOu
GBLuuxAtZWDOijU2tnZSEZTajLeL3jx/B5QF+eGuJ9Y1wm7+zVd1Xn8hYS8rcYy2w2X7KSCmM7mJ
k52oWE899vr1/PtqHWOIWVbwlg3gm5xZdvkxUHi9HbIB+WEOFznvpMEuza74nDQpAOKcyCAYQZH4
WfSXbqupaLsOpTyEm2//aQ52PNtSm4Np/VtLDO/AzjVbsRW6X8nXZjdSNA2aOfurAkYZbB5Wmr/e
i5PNTRuu0jzWZ9GXU7DsH38GZuCbIUSH9p4WW8q0QrrYM7O/Savfy7ymWdaBReDo7PYawBsH9L2H
buTGi7jW8YawrqBEF1ucDVjhi9CgDklbHwFnOucw5drnQ1L/csHHYeX/2qoYrDZFvpgJeBNpK6g1
yzGRI/t9mohk1eoZ5VBNke63jXPArldzUqgwOdCZVNPROqhW5rQ6BKqPHKB5VyDuoln/RbCeiARe
OTtyOkhKbLPhdA4moo7uqk9abQD/1JWRIR78cAbdB3cv5gSKHjR13qp8lz59k1I2SB3mVlDQ336m
FESXV0nSpgUysl9batboeqDGplZIO5imQPtpcjZ3E4/wE/qgS/g2wVSQIwxWSbrrAfh4VpRe7BMe
sIZLZTNTC91bAwSluwvToEQaginhIFUvNZMc0dG9Xnxk51Jcbp+AeDG6ge1run1qmQS1r6Kt1t0s
IjpvkT6Ffss9mjPOKO/9DTqs8qeskniE+mqFzwFADz2W74+qpiOQk7am8R30YWV0yjFgLVprJjYr
ZGlHfEw99W3D7puuQ3EI4RtSMRv9GXU5kOMY04GHPcBZlZc8ex+m+tsmaowVKuD1QlDxiUOx6NEw
Dzl+0l92Vv/3WGEakCy3mHn0vDrLEOa225oBaX0jZvKDAVYGueh+G0Tp9/U0b7xBdhboyw4eQo3A
2mde7D/C4ktktPao8Ez5wS08MBvhE7qi+RUEF33752qfSdgDDEUoN0uXqzDLKNk1SIY65TDQh+sA
yFCuGzhR+KUKfPPM21ANuKFzodCbUDFgGZ8j9QvrfAYk9Y77G0ItPKhDvUj86T8AlSIDhLq+Wul5
6cFLUdD3xq0or7ec13X6W/AGXqKxKSGGl/hFlqGDl0k0e3zgVycnQ0T0gllklLk0ilOdQsQDaaeZ
lmnzjtLAiH93WAh8zHuRVZY9qSBeZ7RAzrnffYgPZmNddL1b4+B+/Tnui2CnKcQJM6OzCvnsttUU
AVkpc/dZsvjJhq4YbyHUpNJosuXF2y0MmT9i1rz8BTX/PdzRRay3/zT9Kw/iokYqDurpr0P6Gqpc
AKrja48ThU20uSZJraUk8/HwHNpmJtnF4hpOBCMTmksAWc/Bmips5BYoCppsaAYOGj5x5WjRMpQS
uKvo6OFLOEcmW9j5+naUuQh/K0u2ZerAWYuzqAvGmmznX3F9rKwT98/jZKDoaBmeI5znrb4/Xbg3
8ETd+7Q3ALwGDHSuqHwFasQ0L97BRuYi76tKhAK1RwBj7COfoqfEr57ThnZmdWyW/o+wPeQzpel6
3BXEts2D139LYv5MlQp4iezXrOsNTgNPhxpqguUj7vX5R6XDPnG7YyXo8a8GvckE3BIKqQorv00T
sL+YulSkh7RZxws/AtI+g5pDf+xesY4oOXWsTnCKizkNqC96jE9sCVVTaI/1KrrVAp2MW0n4wf7P
D1QkjOF1X+zvSbkiVQDErXZxwurwgWgPd0haITHqYFmkeoT6AtRyA1bip8K+XfCh3uqmRkVdVjIa
RtfsO5iybYoDllKXrexWSWtWhPC9q9KP3awlrTZlSVfnu+Fpc0xflBei5yGuCitrFvFX82LHyawN
H+VUwGxh0Mv3ZrHl6lY03itL0XKpagqR3U/68PzpP7J+gzZNl15iIvtgk1Em7wjPxapsAGi+fwqi
V7gVFmID7lfUuszZE9ExmyBChDG+g5+JOzUfTkE3h6ed9vphTv2PjpPBoda48bTWpmqxnbooQe4N
Mkxi9bAZTc1vo2gw+R+V22ksRkj33k4AhXwMWcwJIkH2vkcBvF+EaBD0+wQp4X0rFY9mvcPRkoF9
rA4F3DaI96Edn82eyoNW26iTaLxRnL8/sLDtvL3VMAmMXJ3sl0qpfM2WTc2LFA81bxFKOdwuU6SI
Kckd18FT1nrSYTReRy/45tK9WF/hrsZGjoGrgOrKnJ54CaBmns3JmTCal22WWRuqOI7F4x8Wrn0x
POhpGRLAQhdL3g9F9WjXy+fGG6wIGoaHEz5tfyWQeLRfxD5Y7X5rynjabI39ehx2r6AY3x9/wS4r
XQpWIc6en0mUp8V+UeOQsh5spO7cRppytxJRHVHed5cJUjvF0aGlBHrHnqUcLngO6M7tUB95spvq
O/fwXxn1ki/2lAU1/SnqNXoCGJ6DXE93fK2t26iBZ6HPlHMyNxttYGzknf6r+Z8K0ZJO12cbJCRt
xn8WEOaVcmMRD33uo9dw154mUBAuMR5Y9TZjhq/VZYKdfrR3biNhv6/f0plz6XFGITO9g76A4/Sr
SegYm1lb+S91UaHCSoJWbeZQzN03UMoZDmH2FMyq1DCJYGdofCb68/kxitZDDeHgvSbDhNlxHlDn
mqXfHOyFNUMKYGcvaXQxOMi8blcxpOBVED9IiQ+ifsEp
`protect end_protected
