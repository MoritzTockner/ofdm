-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dna4yTRcJpQwcEdCVakZrl4WCHVudsWo82EvWmwKO5FvAMEfLsvdQbD3NHna2eZNjfXBkxQVIPG4
OmkLWsbPJJA17UeeL7GWMp3QE2bCJrD8FvpciW9Yz7s8RLCfuLVqD3Z/WeGVwNfyM5UPEyjOhe7u
cAMIYBW0pxx3FegzmSpUPuFujjX2FXIcktZ4PbiNeCL3Vq9pGW7rGvFwHK/XZYbNgpkqr+sXDp5x
9Z5yuQBIEmqbti+ZTj/JWsmdxQhYoL8i2aNW1fwnbmykStaw2wDMeAA0rQNnkbp1NjnXneqWGvpq
x4ZphLvmK/L7qov+LVm/6wdYghJz7M2ELlw5DA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
SN7biTlsJUk6rvMpqBbYazSH8w9WHymBJZnrSbrkdJAKXF7/tJ+aDlEJXM8JKYMUs3VeL2he/Cqw
iZs3t0c95kfpAK0nVEACDO+ITgVm2PveqCAwsAniz+pC84W2UOc5TQHkKmGgftS3ShMBuU37ZQND
DPzXU/aK+1lHHsdUayFXbnT98ar0vRjXYKxnWYC9BgGtk2Br0Zo5OV4ZNPL954Ned+BASzjiGbPm
cUS34oXjAf5mJBXItnaWnDEATAswltijcEjJquLeKOMQ2+WvI3X4i+AcXhhDJTxUhKqd3tM34YzT
r+e5T/b1ZyAVgNjmbhj8aXVm+SjGECod9KZEDVSS6o9m/gNeE5HdDoYng8lQpcwHH8eFwerDmc9N
EZCYkd5GCfNoQI8B6P5gtKNZfC7QJfZ40wthzZZLP17nKugwVZQG5o2oSWNDPT1GSAhTekZbsXMV
U1iiVF7HxxdwdDWglQRGYXX4LQARzpkfMfXFJuWgbY8QhjuMdWJSbZkFuZPyCvtI1gL342HqYizs
N7RvvUobAeQSGNG+ms3UAIkC3zdjWG06Ks433qkKwWJts9MkjbIod2odCKeVNsV+/zcmfnMG4WzU
hdCFDxOiRow3OaMZxQeqbh0oDeR+A9G68QSizOjzRBZ64K8hHQ5ujec34qSBrdIDRwHUXCshJDXj
0OYdmGUQ31ssVk4WVrSAiiQm5LSncOUAIoDnTqDii/UpA90ti1eo6ImBW23Cgz79AWWmEfcpjBmN
q8krg+PluqgHjCi4Iq+glLdCxKTKY+6SGR1Uc0/siOLMeakNyNwDA71PNniHAdxHwLmt/7uvXnf/
Fkw1JG7gcaFzjWWlXu0qYilRaxY/K56OUGT4neQ0tIEhJACEsXCwJFWiTuP9KA4mcL56mEocKyeU
NatfLvgwpaH3b1LcQ13vsZ0JLWfztmmHdgbXKPLa/18HUetKKdlB/aOLhoXcZmEPTeVNK9DQIZxj
W46BWhB0sEkXIaNhm/B69TXlehZjBT1DkA1RQfMU4CzBjEy9gZ2Kg+wyxehXOCT48/0mJXnVMTKM
eLx8M9uUFl8X8EADLpTB/48A9Anfnf2tQ8aQL54q7bkO0uAkl2SA35VfhSDISGNfx85mcVBgupzx
ISDOd0H8ChF2t0m2mwkqNAcSsaKzx1sHkLBJy0Heyd6/GyiPl9aQX/XS8G+ZQWrKK7mA81CFZAf7
uB7sjycb42SE+q7ZhCwwiz5541MhyglqpApDK91lhNBKCszi2c2i61m3X0u2c7QOLiA+drzgZxKN
3tKNBnSzOhzA3mWCXo4FbL59Y/afv1d7q5DZtEeMLj9SfF6tYb54wv2mmALcfa6XxB8Me/sC0C0P
HcBKO3JyDsgub/0CNfB3KRcak5NVRhW2t0loNc31QWv9IBSc64owTBAVjz9vFikI3F44qZDR7DgN
ReJc4+nJbitiwKj3hcCVw6YcTX6M8ydtxwxUdNemRbtSEaEoEcaooSjplfxcN6W0qRML+A9VG1HM
xjKJdJJQhcERpFG2GKQIkP5NCkKUcOamuCV8BHKatSpj1V0hXl3BomstAsaoj4t2pVc9QvIM47Yq
BjaO74Ndi8zHT4QUNdYUA4mw5/U+pgDYVdo5ppO/75TzXpYQGWWa7XLermac9QuU5sWPF3su7uSK
KB8AaYm2ivEpbLbqN2lD1e3UG23DE+6eGMulSnDMPdYsIZQiYdhkvllrB3AGvYs+QulHHWnAjHZP
dmKmYrzFrSs5ZvwBI/VpzgOFGEtYg7Me4Dgjty4eFIGFgjfEGLWfk4XL0P6Yf1PQ+xPrLhv4bYbK
WXgF3KQsDym/wINj+GP1n6Qo3WXTkXsaUqfc1sRwGC1+nv2u21fuSNy6hCiSvhQf6DoFcQDaoVp5
uuoBfjOrv9CcVh+6IeWli0VwfvJyaPzpawDYABAsHeCx4GsU+ADxkL5RaoM3OgnsN6gwgBVIzMdh
volKuMAJVNTV4H/Aw5NQAXFdn6E0JhIYg/3Nl3DldBkMDJNGW6ktsxg6y+hba0qVurLmapHY3NKF
1rwnJ6E3ApVR13MqhJf0IK/J+NfO5GAs7Ag0TSi9c4lZJSPhMKJTP+bpcMwGEu53yKWYxP2C29wk
NH2z6fqPInaKG2tXe8sknsjxiUeYRkIC3B4KocKATaJ1w7nipKA6/TYbJHYkH13xySIntx8aslXP
8QiOyOhHmj+EhNvPUFvzO1WnTDfT/9rTrw6x1/zKDoPIAsA0NBzuDt/duSbgNhCZCW3eTvU0nYTn
6EF4cmXQG8q8qKiUCEdrpsUo
`protect end_protected
