-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FP8vOgyVHfI90yPL1J01FbYrOzUilsHlmzky/DG5o0Se2qqzCLdO+N6KjaRdyefWZdWevyakGxyj
EFD+omJ1J9w4NJf5IfLIe9g4H9oLUWkIURjHDJM1LsfYkuhbYS83nAUB/FE8ZzWsei3r/5lL2NCJ
6p/UzM1WdEptFgGr/NotacD+D8sAAEpa5wCrDYC+L9ZJvghTLhnKxLZ126DiJ/EHx5H8Ba2cL1IO
Y+qqCc1QDOgSjrzmcE71+tIr1dDXrZnpWCNhpq95Vc738mFEaA0uA5nrz+0j9URXB4hgNoKWTfb8
pPoNXvVStYib4UqRByd9ZYvq4V+YKAVju4EkSQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
w9xoN72Ca3DDdhfYo2qMev66a6Qry0qS/vxgchN5U+lKFAgDKZW8YRA/yGpgltMYBFgDfZDc/c+w
n4dAdn9f/c9yyaWbQgzCHFJUsrbqTmiCkHWFhxrPz04dYw2K1G3a+i1xuTkbVyPnF6x2nN8qWcm3
jCyCHKmHzzRoqCVzC4xY27H2iucPlhLv4uXvfecS39zVbpaaq7WEQ7o1DSV1AppaGM6KrvDpP+IH
SF0BcGsStSMFx/if1yvr5DhcfKY+6XzCFTv9tARitvD+SmwRvfrLpDslFwSFDVW95lRauEbbQEN6
MeOtkR5qczOKYKnaXCKENE6vXFZi9xowy5gSvFh2pwfJ5pw8VghhU4Tv3KGLyDLCYIT5UuvejCgq
SIGQUT1ZmcSwbq4foj7f2hHJmQcO9gO/u2q6Q7sf2nvKPz7uXE9shPhnQ6DIVHVCg/pLQSgWUTW9
WvseP7Hi4N9uXn5Qh+8w7cIYqqLzOjf43wMfsQIjKMC4OsFQXNh+XFdjqYBQsdEetIYIfWRR8uCB
Toh6mNuLxQirWEbUempN0vvPYJhjBSvU39esK/D43MWEs7eqIuJ6C413ZIGET6AokFcp8jX7rbKE
OIYW4YX22hXbTJc3FswzI8S2THHui7qmAlP1/ZRSTqcp7N6yzgZ9q6TQyZhlbb38fl9aHr4oC3Su
GCkXPfYrwuUAJfGIdSvPe6bufvUChNaU4McqZAktBpKYA37+J+zu6ZZvdu3XI1PgJazkLHrOEbaE
lQrbOEeP5l2HEmlv3Bu2ZkE0VI/YFlS5bEWv2JyHy7Hud/0/utZl371TjBe5/I1oM8pYyiuDTkhV
2dBVsglH43o0xCZc6NInP9U/HL1SpmVqCKAILrrZao6dy1x0codPsB68Xv5DvEx7l2EbmyAN7rHv
P6YOJwSxfB6lzIoCa1vlDllpA6geSQNGYQejejXvFWBTdXf3IFPbQ7rWMqnm0eO2EiARYlkUEu1p
MOwtKggp6NPo1MKZnJeRj7zaffRjWQOH81aLD5j77lPaa7tNT50h4ITDkXJYOqJqM6WYlxN/V0Pb
GAhEiHrQOaO2DVEOfVal6xro+rLuev4EKH428SAfcpguXXkBWOgjOdis37iZKGX1+HjNlMocJa+i
FLOVfFq8oefyHq7x0C+ACxFK0E+EG1HaCgCH+GJIfbWGHGeHv60vy2ML4OQ89TPaosKRnmjPHDCb
hK/MROM4xHBebAKsf3rHIjjWxBBxs2BAi83KzVsUp+x1tdy11OOF7xOjT8pyHubhJtoc63Ac5ymv
/k+ppiaGGMltkxkVxlIl/okz/NoJK3t0g0k6P1/BZcemCxMNJQ8rtG9UDM6DLEIV/TwrBKGXryD7
RlXdFPUpQXTXf0uY6Jp02kSSFFeljHvaibIKdOudhp3fOubPWUFOQVMew48Li0JEp/lwpuPhaj/E
RQhDjUqPqktikGmB6aeOawAWdQ6H7znAnE+SUSOx+XnHdbk77a9dZ2d5llhOvZqGUxz1fFQWS8dh
nJHKT274IxE57L3WK1M1SWMWV6tvQDGUS+zrm2XciHBHL0SX8Up+0HxSSZ6Ac8OUW1qBJ6sUDjV0
Ofy5EoVfeA3XToOBCSWOvbDGTSxs8LBX465Btgj12N9ptr3JUJYQKVkYK9Y851ePPDSbcdamdst5
OHW7NwId3HMLBpnM2npjPyWaSvL5VNpRIo+2Pn2ErzJVz5GZR9tDdzgxhf4tx+xiD0y69ajA39FG
1an1O/hcOIgbpA3BeuJ6Li3F3/705ay1EbbVfFab467kPCXmruViS6GyeObJ6S4ylVLAcdXH2Rl6
qFrDGG/YJG0xXHOS/ZtVqCubtOcFBFh71VsB0SVmYQqKFzAAM1lRPmyHVZoaXfyje7bL2BfH2KeR
3j8eVD3MP9Ncek+YBG2oY4Jeyy1zoNT1EI0iI4NFllvbmfKXJDtJZCgIW0mt5xhqU/YB6Mg3jKqp
uDUi/ROAdAxjihST89+3SAG803h0o+J/ktYr9siYQfCyRkmDiAx61euIHBoYDdnESA9RA8pr/rIz
WOsiioqfOvhhQMBQEt5H+uuCxLUodejAlLb4qt4fnMNI6ELF4JY4lOiMUZ6ilqvcLSFiveYb68k3
Yk06M45DheRDXjVjRbAe220gNeIf9p1DWANL95TSlW2fh3Qm5Gk3ITSOSdueO9HKc1SSSgLzDTcG
aBC9RqMN9gSzQbMdDfTtI3QM64c7GytCeBzcuIk7BuT/Y0jDQ8OuPw+QiT9+pO9Vc6ctD/VoLnw8
CiSACwc5fs4JJdmZLhehT55YkHVf2XGkW4LpMC4HYQJ3tYUteGULB38idDitmFVTx+bhPUK7QHUH
QtAqG6C2Wy2VGBEWbd4Az4wnwrA6kivXZ6B2lkJNAzowcR2vMQ3FXtVRrmxtiCTahAZm+EujFL+M
xU4sOEc22cbLLZ4TCsLtiWZQTFFL2MDDl8AbDwjfWNwLL5rM3JwQVnsfC01V8pqB4hHV2TPCkXtK
ASd9xj8bXn8Vl4zxkat3GZ5pL7nhsIcnQ1GLs81mLSB3qCIY9mH8U5IC5AvvL++Cb9wvBeso/raH
NLwB6nC1gwdrOxelR/SzLbYBpDTL4//BlSa3j9fWsth3/LND+c+NDKniY0Bo8LgcM6yiwBF2xWbn
27lXWH9Dgtv4TP9gYpL/UhPaxeGknX1RxaQ5a+zjJCIC2Ernw4lUMoicS1XlmS0GbbmuTSXHwdbi
l7R89su6h0Xe3NtfLUkYYNko7Q6S0IvDwafok1Pv553AHGO6OFGWI15imzD5lwB78kzJFxodLCzd
0u3miwf64ixHQ6OMsJMUkMDxCxa2WwJysfoLP6ipmWbmWCjAyanI7TRkqcHH5+ugQfP4rJ/aT0B0
5aTd+FbdtejlVFXWGpiGfYzMGb26QjsG1N1FPlC5GM+hv0/WZq9Bp1QBEdiFeNo7itxewFuuzbY+
XC6sldYdGBDH3dGmSUiz8EpRNFpnsC6Ls30QEJn88O5kd3vVHbnk5VmW5vDCc44p0gmj1JIDPNns
cigFUGakR+ogutrH8cP2v/xIMI80SXH1RFbdaO5jHV9Y6eiNFAqXW+nn5QVWmJn1rZrH6k9Krnp7
CrHZaEH4v2P9JpUISbBb2iqvFTr3o9kPYWzD/EMbVe/529fNpaXv7rKlo0bZRngpM+R1WjHcdLgk
Ub7BfAsYk4RQkhp0V9thv4kra7aqZcvyNr120/w7nadHF5SPpaeREVJ7y1JUM9P1Jk0PbcoRXOt/
uZF6YIaWTAcOeSIcVjTHcPNSJ9IJLmionKZDOosb1N7cLIkGsgQFiZ8g9R+j3JGb446WXLmZnf1l
mIYHJNDDZTX9eXMEVPtBORTYYiGN4KcD75wFpy26VkjV7d7jyUoXeuO49DW0DO99LUJWgfPvNg6r
M0HH5dE4xckxsiErdwbvzROkwRx/OnMVXd+InqBO/3GpfH/S57Z/yEqxTSORayTrBOBoTbfeyxpN
+JcP7cK1ApZ7eszC1WsZkBQd2ssOzBvBJwfOm6iA+MoVPOwpG86uyfFZQXXw8oasR3rf46oWe+73
b0zAyQWCVnTHOJJecwFInYKVDN4CoB/+GlEqyfcpS+XjGVlQXnM09t8SGn+aOXOCrBYQhFpWZk7M
Y5aD2DUsv7HuUD+1XLqKsToS8PU544SpZSedVH1LNn73DGb7Zq4uHLk250K5V/9uHbdBuSKiU2h/
3bPMeFsMA50xKfNvj7UT2CNlQDKaHndSNo446eMfTYmUrk+jwq70PHkBdUEo/CEU5M8D7OO12om7
EKrdeQUuoYf4iJA2iaeugScpO3LjAw+xlI23B47WHXKiOUvyn0aF4tYNJv92KKjWbkAV8+cxng4A
T4rVGstBfzsxNcL46lpOmQP7i9bPZNEQJ12Bw71QSbFfRz/kN5WMj43RPqVvgeGqbpZDLd2sCHWs
SnfVqYIuVXbjOj4p1pXVW0esjXk/eobvntJuK6ZwCjNRnkHtnXAbKpY5AV6zBbk3SZhkn3qCF4sS
LboLO/FleyljMNygcaRYn7w/q3wk+QKW6b981y5/ARa0MDzz/Bz9NrII5tSmnLf2Ac6QgUMrbcxu
uUCoR28h6yX0GA5uuSc0+geZsxbMLADpMaiiRCSoo8CKhOtCCvl6QaFSvgqAcy6Bz28IQDP9LW4x
4GJDcnyxKuzCY5VZ2psor+gckMsIQYgjiEFZJpL5jfDSuDpK0d+UH4KhRXxPpNOtfrjhnkx0baTS
zDZ1Hsl7nWFd22L3/yBpgX/LfOnsoJtNurqRMdMVtByDPcWrtzwoTG2SRzcuk9EAII11bDOzbJbm
39M3GNS4E2G4eNUA+S1qobRJNT90VPrPHNrjnPqcWx4+mC+krC36q9Tq4hJto1XxueiI7B9k4v0w
gGsDnHecZMYRDOR9wgbEaBxxYyeysn5/sXEvIS/w6sWg/d2qYHX1jKU1m/q0uWlbypWmFhLKsOvA
ir56iZoa+cuq6OZFyrcV0eA65T0mC/WqZbxs4sY5ICoTWrNKNcjYwUO9vc/vET8C6vGdUtc3LdQM
ohUChsBWBGadpi7BWSWuh98W+pYVNYN2GA78ciCRRaDpTuExOSjSKQiMbRaCq2f+3xp4ON6hlsUe
RaLUQAQVwPclMvY0w5cgWPgUdPsTGp8DsB5v+xhU5RBQupxp7bqLy2QsFh2Z4ZtISlNA2CJVkV31
wkupf74SwOiVESVsSMw3CTk9DPDNliHDvmc8f2z3cxtBSkWBJbZSnzmerbZQ6hOA/LReyZvnbnW0
p8y8C1hReqfAa7JVccZpbM/d5Hm4VLCwQz0mDiMZfP6Lj4RRVcahyKZO5d4Rl2QU7MUYtVkwOt0A
J818OYbbnlDimb7nIpTSr1lC3n7+CcOqShWx3cvSc2Lf36UN9OPSw+e9MjLt34lA2VlZa64Fqp70
X7/KQj2JpeaeAfMeS0dznYm4IJ7wz0Cr9wdQfT+zMwv5qri8JGKgQeHurn/Yrx6u8gVsTa7Xu5WP
Q4ytBJylsXHj3n/pl+p3uLrwqftAEs2OG1Ah/oN54yAazFgufLnt2lVOYjlnPJqUocZ1RbbqT5Yz
zWF5H+m6pU6Z4heBQs8+MFjyFN3eBiH8AChgllzOrvOMUPwzMnW4zKz2U+ioVdTOnat0Qk05HJAQ
xxNXSDy4Ty56KkGQ8MXHdOOpN06NKYpi0YH//3g2B8F6uOu8gRiAGqRc4Rv+C4B6SppjFvoBUSaf
aAUgNRS69ktjNCWe7TgtDHxknik80FtLuT2djqOLcA2+6vl9q+IE3gaXuREdsaxPQ9E8My02mPeD
NP1b8hV2aZUJe5nHZfkkh5QUJcG6XbPiuObkyhAMH/Gl3mFuDb00Kp8lw1LM8obQ15iwbWxlAc4B
20Qk2elnsFFdJpLnL1EHXWFqOD0Do78wgJivP+OSZNCf3H1iZdmwM+3CJMwtFtlr0lpB/I7wTFio
6x3L7OJR1bZbr39CtUkzp86K/TKNySQoUQBbG2zYV1mbSN4wNBlPh2ExXqg7ILXw3t7dUBYCM3lb
Jw9FpdmmFMgo6LQX6Wple89FIFPa2Llqkem97iU1aGoAIowhqEFny0xzIyJbDmZ1hWc+RGv76BjH
B2/O8qry3ldLOTVa+qQLAI/oZFU9wzHXwHjT8SI8F9tjFXSH3AorkXZJPCP29eJ1Oq9ZMaL84Bup
SbSf4WALRQDeii9oI4Up2pRYTt6HZ1NaNhVtF5O6vwDMLq885LjYjJcql6pOT/sECTCTJ6Xx40ih
gdeDfOvzeMwer4o6wHagkgWeUyJVRZ//4oeuUziQ5aNL9p0+B7XP6sr52UoEFL+OuQOB1izLMnPp
4jfjhQYrOE4Bqxh5rE6Xrq76VYAAvGSJNb/Lo1FpjagJ/QvD70pqkfCzIvJwJbImgmGPlRCbogrb
PoGQkqPPAK5rLOem6tntMwBHw9LYqLRJa9stVJn35eMnSDvywiuIk+P4c3B52v2tIpw2hq99i8wz
W6wYrGTggL3OA1wKp9GOvsiuPx/whIT39OV9nEjjbbehpR0c710PrtXEeZe1gYKGxcQtL1z3hJgR
k4vSoZBce8Vw0tVGsIkc5OJv3arfST+20UjsnDZwTpcOJ93BQEuwEUp03DeTW9wNLD3lecTgdF6B
NA6XvSKzPW5148lb6c8xZV6EDxHJ0obsum+70PPQ8eHn0p2uflLcSqFeEpUkXmyRnZMAqu/kNi19
8P/+OZGExin2PAzQFz9wQfuGzWWFSNyqUFlZEZAiDy+UXQXKptuk/5ipy6BhImOpj56erWfVZWCf
d86tMbbZr9ARHyDWiH9ZbQmgkpciuMNuGNH6C9qNW6/ZOFqKbalbt91XH5HnQZ8jad2aJo40681H
kali5a9Pf7YML1OFD88RkllAZbUEWyOUTEJuJ9qYOlhaOzehPhiGzD0BEgaurU75EAGLC/9zsccN
HGOtrD+38r7lBIXjOfZW8tPk9U/ixWJ5Fwkrut0MA4XRt+tesN24jf2YtxLgXLlAYeWIhTTT1BlH
zC9No59hgHlNfs13LG/vwxPSIg1Lz/NaRvtKt0mwV9/F+sHuMPbKMibKThO62qGc4uXqczWfw+eL
bXkLYMgk2CLkIrmN9TKcxt/vHlL6hAnAku700lvifGs4vpH+Yzch+QG83pCNqPArXAM6X9AeMbuU
+rP3EpW8zOonSerC1sWQTnQqbGae+hKyhsG3Vgqb8GE+CgKEi9XUFtNApVUVbJLKHgru9S7trHmV
3nWMKBfWnRKrP6k+9sQyBPtQGdb5mpPdbiZAKHBTTzohFHHAAbBHbi/RXfvgpOfsS1PXJEr93CLb
+cQ1b3z/CAly10ztVrVH3faZNWs5EOXG03k5zqln6xvj/VDrFG3EefjgOT0e9sDigCn5lwXD7orQ
s3DxEmXlrdb56HaJHySmmH+/SavcKMO1o4AVaWe//w2/2pMAyRzbsIqGXJq8n3Z9FF0rB3hb6ltC
uDqWCI39I1iLjy0VnFRpgxsGqzJuYItSOaTTTz+ObSAKCIS1mnNn+wBX1Hiw8GwPDFFEqpxO+vjP
XWEmmXrce5aI4+FFkPojTtu4snytWbcmVW2a4UXVKTISGcGVTp/BB2EeCXemdt6BdqwM0cPCm93f
75l2Hy/T8Yc//xlRO0TNitMcD6ES9yMCtVWtzpGh/FaJZiHmRBBYx4tbHQrlbzmkXgrYspS7sb+7
V5HSeTm6KHNDxJaEO1NyYdIVvQsVdmBz2GDt+/HotJMv7JvfwizK19NOaXY4YC9APyByJKtSVx4A
xEciGjCgjULCBpYkkmTESwwETBHpSV8L9x736gRm94fNFY9ks1l7IkmEPfixfff2Bwb5R5g+mFVQ
FL7KdySu7LHUFnwPwNGlK7yiPliEZuHSclKEgy5owXv23mAb6LCF9t7rXu/wxyPi0wk3YzrhwIZC
pKMH4LijTOkoTbabsqXiQ7rX+9BchFN8frbDq3SnDxXA2D4pJzkek48TVbBkp4uCxNQjuEqQ5+IR
76sHLKNirHdACBvcOM3prG0qsUlCnkonh7WIHbGjRFzEIgSa2hBCyhq5hDwxkVkhuGzFttriKxuU
uYaNnHg4wZuUoiL1DK1gHfKsJhe/K5ngT9DecyTscU7tJT/b7q1ETOjccSIe5L9v6bl7r+rKmzRH
AZqGc0MwwtYIjd4vY7AX3VZxlS5zRDqSxGSgextZxGbBJkfB4N0+F3Uw1a1A0TsnjX7DWzuvtvf4
RsN1tgEZCV/TPTex7c/Wr8qY2XMGXZE1AkbnBYtx3LOBOBi1jismA18uJb3XB+khIwfjI3h5KO7C
dGeZCtohdI0gwfMdncFlTAPMinB1PfGfK3vRAgs2JLNrJ/9+o6CtOTnMJGVeJk0hf0V7G9wsdAtL
zzNEWtaRgdGLyyC7egQ//qMpqHApdjyx0Wfduc6c9LZzDLLY3reV1lxoAYVf/WUTo9WFKRSzlico
XMDHi/ixGv7HTVqr8ZPR5RWZvPHg7OUbr6iFVVcp6E9f7Xp4K2QYq86fzR7oEeWO+TFBvkW7bKoe
wdpkjfnXGhiM+GrQPa8o2O1G6uzKZ9ZpTCOKlwwY/kSPDREk1B6hlWwe0keNtRFApxLzZxpr0/0j
3TCbKEkWS7bMGmy2hR36xQOKmwO/khu5n4sSwYHIwpMF1T/4HO8MOuWlWnhRlDF0HwkAHQPyvDD6
38ceKSj9w+4H80OOU73hmVYRS34eltMS4k8h0V1Ml/4zA/0sH93Y8+GAhlJUM/SxfV4x4oo+ea0r
BkhBS3Uq6OtaE0H2ZdkHlExS3HvzN1vZuFZK5Yupn5EZ0NUrFbjvjuDBAFp/zYdRV5lAcEKJs3hw
/dOEfx9NP39fsnYIR9ndaQCmnIydjDUnOZ3Lx1NglNe8N6E1Db1boQSB7oeQTUdv8eGAmfBKoBKI
RagdBDqD3GONfnhErniQC3r1p6yzxx8B4HpqcspJY246g7OIDzjT8KYR76Dllgq7595JVVsiH40M
cR9b7IjY/npwb2KeobMo+TkLd91bQuzZ+t8mPBJcKkyyU+q7hEtRUETJns214DIGXLDzNfDD3l6I
Yi7hR7bxbZwv5aNe0FGNoLOHUSgXBSLXp8SjJ3KvGfGKLNkmtoeIri8s21+RoC8QfMQkLEfP++FB
yEFe97eDqrLhjaSCKzlepoi22cGs08KQ5E8VEDi6k33Hx9UwuRKrDYLBQp/VeK64HqUBXpSQrhYI
Qc/n1X1kRssb4MvrEDyTMp2dIt4NpdYgkB05tBL1H8caNCPIbDGfj4gQ5ObKM63Z0p0SmVVnU5Ml
xRQAF+v5GVEgTVZr2xho0aOwDmilzPlfaL3pje6y5JiQsYUZ3rPfzwY91e9+4u/qiMwiaNnVrCiX
sPjxiY8YrOKgNepqAxIoU4XT+TPzeQyR12Oaxmex561MLStfT5bXJMb7yXgsqKWNQZ+dINC2TYdP
j2E38FeNiFwIfKnDwROxz0N3gnecM56n+7mD8Iq4AH8N8TjHIGzidFcuX9Kkz45RpdV5upcuiTYt
mQgiK2LI/aU9gynTuUkdDVTdS4cY8VnrGqaXHka2Mvg8nyiIsNGPetHhUnzrP5j7x11dI8BbKCy5
FPecgirBQhkWf5nhWphFIM7STsyI/pVX9UW8WPvk3z/U9cEAm47lYDzHF3tvXvb9CQWctu61Y4ML
JZ4xRxBSiNTwrELqTSA0n0fwpjsomW3KwEx3UDdk51Yan/DrIJAnjgpLbKUWqTd0whaxI9lw0Dl0
TjDeX4IW7+CGxrNr1PXyTmWXmkcYwefnfTASKq5168wvt2tM+cXXGOvDDl/O2PiMJUQ2nQLhQeK9
/nFKQyB9b7BUsMRJHnZZGzpCdTqQMtbHkRumVHCgXltFuGW69orLXuA21Dj36tyjAx7mAh6HyExV
FN7upROqebCn57343mOb1Bv2G7D3Qg3Rd5MSBtKoKlDPsJj5223z2DvYUm7SwPMHntDeenB2vRzZ
7zoEf+qzkOZ5LJJhM1QMxB2xjPwtz6FidtyWUkgutSyO6i1Sx39VBH2L4H8snMswtoDcTTbCWEaq
FbYH+pIHzx1qFzmHlVQLUFpveYiwxrrLFjJopPcp2Ex7varlZGH8xQ68Z9QMhHeFPTqTqmU4o5gM
9iptKvZjWQDNPMFUzx9jiS/1T2VtqZW1/6aowKgfSReaDRsx/71dMLq5gB2kzLjqjBIfIQ0M1G9v
c0WIeKon3hbPqNb6rWHTqpXfKdSxuSO6cGZjRlP0a3urG6KqlG3Y70dVLZo5aeZ0hjnq8JIT8ISq
BXZCa8OJItJj008zK56A19O7In4Yhk5zGTbuEcODgCoeWYU+OJ5PAP8f1CbXbIGyE0rg2iGuYmvh
KdOzWhfhc2BvlfTCpgBul/ooJ4lt5qWada/HoNpoIVJU1LAQicbbBjvIFP+wJ9sjMyzQUjROiuUc
+arQVRHmkaKdxDP9PAWejlurB9s+KGHVb2E139qw8uvwmL/9fx8uAN0MPbCuvcCp9z+PORmmms7u
7DVL3N8hfCY8uAJ/l6z1Q6g/6sb53QDtScBgunVMT1IWT5YuMX2yMmVKIC9xWpDas+1ZzHW1Q6UF
byaFlhn0l2mHZ6J3OffiHT6Ay+Zy+c94ZSn1NhQn3Ot5rb/KZ5fL3+IKDT1q8591aJJzC5sZvPPo
lqqixnKtdSW8fvsxylZoQCxCIRtlRRv24Ls=
`protect end_protected
