-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dImWB9VwERj9JsYyDm1GIaV5Z/wE0PL/7u2hvI8NBPMtAMA+uDQGlOe6WgIydoTxEdcMAPURvcKs
VY6XoK+HgPh6rYnyMvdDv+RTgGoLdap5dsOnvZw012LDD2c7Rra7IPGi2dxNpL4sSQ3zFcAWc2W+
xWzf9Tj8DNOUXwCTMHHeVRKfsXEgxsStM5nfg6y5lY7HPwkl/u9VVdG7uDb1xSpF0QqZ2uYAUjmV
rlqvQm0JokmP7ubnBsrIQ4Uf5zTCyStJWW27w9FKeps4W0Ngbjh3XS34MUMOynL5Y8YwDm1K+CFp
N4n4RzBIi87SIOyxte/1rOkCmArw4+bz7/70MA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6224)
`protect data_block
5xAiYB0gbrHK91ZWKcMRH4hwQSQZVAQXQgS3uK1Xny7IxgQc5OklWr/PxRZGf+u5iJzWNCKF9eyO
pRyJZBshKJe7nLMQps5ZUIeHjJ0V62zueXDPldIOa/BqTDYmORxXkPWPYs6JLhXf9Jy9PlxwIj9H
ZvG65dKKv7QaZh99DuawfBDmHQaupjLE8SSB74l3u1FtSj1UCV1414BIo7RAq+xTWxj2OU4KGsj+
vWnH2Mol4Rf6zz6dJm8JznMNLbubU7ycJOO8vDDZlC+b3AuzrccOLieHhAg2Z3Xp7A35rox+weCM
IdDLv9j9PwmbWKmE1FPf2s1qrEE7N88XAcjoOH0D4Hc3O6kHeg/TZhdbpxfoIoLVPK7BAceq0J4D
tK1muhEjMnKjq9FTz3srlNmAE7Dj9xx2+vY4LsV+zvisuQUOzbjtA3Zd53WWLH1aXWo/ltkvNThC
B3eCGZWc3T29rZYsFkCzE/beklg5lRvTBnbTHewGAU5Q2O9Vx5srrVy5Hdn7tT+UZ521p1lki7sD
BiwSkUegJJ5NMYg/0nkmVRpDdlBXckxGmWp3hpaz9UUqBlZXg3hh1kAhT8GT/xbzsce5qBz+HtDu
dhmzWwsJcGQYInhQhk/DjnUwPoCIn+1B7qeqXWPaY71MBcSBOqV5K2RDUuQTx39FrIzkp9pd5Li9
0r9Ix/nZMdBvNCewa41/uAnFlL7K8X8mxc4VcpnUhY8c4C9JuctBBLJmBxlJh3blCzyQqJqtQGB5
uUT20kV+8WItfgSU3Eu1sSAgVhvow2GY2XUk8kTxFII8uM5Ge4S8l4iL946ONPviWYLnACguN0hb
mNTuLAsF1gBsVlN1GxipdzNCTeS8hkf6aJJ8kpcNXr6IKZ/FGhuQiOPrTVJecFUQ6Wk0P6XximcN
qfh2zMOaa70pDeyVFKvpMYicicl2DhLuqKTsI1hqYa71z9wfTQ2+KePtsWTHL54CJDwE5Tc4Zpm0
wWb/N8zh+OA/jPHBKxYVkcAs7xHXynjDM/QsqGJAQ8juIxfnsLusbAPpByJqfRORh1f3guWvp4pU
dRoTv1sveGuxkDlF/KLqz6v6W9gkctjmUfhSwo8r1HDVcnuGJReFX9PnMguBL6aOxVMvWWWjtKq/
r1/DDkYXvBloyBJDMgN7jSHqspJnvsOFIKRxoOkTvEb+3XzR2RxwVz4wSuevGhk364idiOxiSqyI
JnTxmcTudt0pw99OAiTMHM6WWHFlT1qgHit3t9ogCfS+kqmfpw8KvCSG1hDIGUPmY8X0hFDXR70c
JjQZcHpj2Rneq6HSd4pHAVNJiHY+qLQC54rBzamqn0k6G5cI4e0SacZxe+P5J7PGVrwOzYq7bfbF
lLdtGWOqom4PTnge3o1TvsK6ipJRuA68fYTgRzOKQXy6zrRZTM4p1romrCkGCypPoXpGRmZGxSQi
A8FmawbT3FK7jxo0kzEEOPc9HBxZsJ2vbX9477CHIu/wug3zYpLDHWV7+5XeEevTPi2fUVN23JyN
8qDeFZKIohX/2kwcTuFdWd/c5cOlJLk6sWdbtRjAByW37c2sx0skJi/a5Zeg5HApSvmmJ+FQAjfi
nypPywbJWbcvQmuo8cr8+fZUg1gMgdHHy/3gHKuvr5AZMss8lng4M02l3ByWzr6go4FZRdLfNKdA
NanOOuVTnk7r4e6NNwBWpk5+P3RCmquyIcorMFsTjid5Pf8QAX/uVlj7NhbqX//onFoeTXhzx4sf
VZByzSdTvOqaLa4KWdlCpWWZwL4IFFfOMlzSgvnt49BzX7E7l9Z5pSz/F9b+bMyVyWGQq3cBMEuW
5Smo6ltd/QMra5JGLbw7ZAanSwjD4QCbW7QL3tp8Mx041+7p2PQepHZME7Cbk4Bia3mwKRK7vfp7
TlASbYJ7fGLz4OIQ2i7B42h0cCRUfuyNPmLaK+HW9w3u0ZhG30kquYxG9O1zWNQ5IureaAX1njF8
4xaQaiQmOO/rE5xmwva1ZtIS+xonvBHORVrxHjwycOLSkZyHG412sV0Hndb8UZ+H2SJAj5YQfIq8
lgIbfPwkTTIkrU9c2+dphcV/IMr398/Wcple4eD8h5Fpn384mq9w1tfgwRehGAxnBta7rkGuY4oy
wmkq1bMudxX0/hJIRBT7qpby3ingFE9ACXMqpCygA98AL/iwonBiN+Vq6VOJgSGoyi93Q0+ny6iL
V3wNQUNHR3guKkc0jpmELt+KIgeiAUbBRLMxSDCgP9jKOxNbEJTsRMJvQ339q5UY8OB9vlRLM1MZ
fBe+6AzBDmTJA3FrpRBHtJz8Y933Df827fYtSpWlIiLfI5Y9QUhY3xHNaNfXSIbKhwRBREt3LpX2
nGZKuoILg/V7tBxFIwM1Cs1CEXRJfaq9fSCGmig2PCJFA7VPG46WtSDdT9L7FLE0BwZJIsGDKKsC
5s7AlAHeC5BmHv1/FkFhsoQWWbfgt6m0796C7WX/wsIqFWPl8vCCoge0TztohdKuktAoRiAIQRpI
oU5NXCC1aZiDPxs4PCypKKimF/O1xwKEFkPyYgl20Nm3Wr81/RC6pFX6u3JVh0OKiAJa//zfZfC1
2yfb9J5OjAqmZ0SvOT/8pdwBTc+UKAE8JWjXICJ0G36RPA+JAHT/VKTg6XPf0ePXvFLUO3HYvUMW
8153NIXZBOvB2KzGDVemHmJF24bZfhmf2cv76KGBwpt1cBB7ndQ0SxarRITtCjPU8XnsbQDkXAW0
EBfYgRxGeFsr05owIdBxsFiI32IDpNIGjh5UiqHimC91D7eNX1iSDuzKRDlAb0+hePZP2mEp2HpQ
YMMnJHn5VqfuZYru4eNHPBTn1YCv3w2cutS71TLnnVx2kAWyFXvg4ovh9ltjrxqRZJwgHisS94KA
bIHiCy/Ho6Md9A3u/CPnAy2fhdJVtH5Jspk2g8t262mDamPer0rwITgp/SdtmaoVNRTDkNl2N5Wn
UsSlMvOaXZxk2AkZVKgImd+2hkJ7xZgxRCPJIKEtItIdMAL7z8+fjqByNYgMCsII1H+Cmc/7jFko
ZVr4lcMmrsE3Q0bjeHk/zfYW9bO9rao/MLEvB4JDtnAlrZyZPEypjFbFFxqqndWugSR6o2Ki10me
i8ZfqOOrnIIlLwZgOT59BQNE0qjSLm7bts8HfDl803EEE1Zdi+0l13G+sAATxDnxRcrPA+su3CP2
x3BzTUDYCel2UyULEZ4IZTSaiUCfRjEUs/2Wc32FBybFCdwOE/3Cvf/bs+3/Jud8wDnqre+Hguze
bnTh0vcHhwyakoki/gm2QJ5S+/hpF2+Ffmt50iQxFoRko8pLaNuUxnm/ctMDsJpKiRML4mLChRBh
fgNIbh03eN01RXx47NvDXyEqEwNZRpkgGXxMxzAP6j4dClJdBpla8QzazMUYrY1lIJNfuT1a0K32
JLccD/c/rjjZdxF68pD3YyfxgnHRgOpGZlVjNmZ9LLFWQ9pQi+ncktZI+EG9AHKUXsMOLvYyUYKR
J0xJOt67x5rHIxa8QkfJ/0Lf9Rt+Fs1WBXgGUFtBPUk+YhbwpsS83Oe8V2HFYMrjaqfoZap1w8Vg
CY/b3Deo0MGMs3BQXOaBoGk3hvx1TQpfM0nWpB8s4fYYZ9LQ+1lfzQ2Ht/QYn67GcfS91FeidhVN
A8CFbzwd7Vb0zJph0MmJZCwGpg4dD6UYKgqbXUW88J4FRnyHXWGj9Foa7OgXLOdw5pVPlMOP7u5f
7xkUAVlkHRUXcWfcUmfwKsnDm3Xdow3EFgKwYOtnkeyzh2KAHQA+BJQj9VNPcrD1YuvgwoHM0+b8
9tpJi34ZxVoVhCQSCNsYdLA7uQWK/olEAYWznXJwtHG2SIgeWD1l1tRxUV/zpBsCBEctb/8DFsOz
RbwKICyKnwfi2UgZlB4GL0pakDHsXR/eb2rhuxffobmb+q4Oe8udjSb4ETjI6FqqYNjdDPwQqG/J
uV/hpcVeSft+hkcroyQfnVM/yhv3wWrDr2Z71sD1iLFtGQMrtZaKjNh+3VwrfP+1Gj1+/G2ytBzw
9QW/7nNPBhr+D2osDsJl2HETYxC0UVhMzUb7IJmUlnmF95KGUOHzWBl1YlvpYTtpiI4cG8M1x96+
YLC5rX7cvJ6sE0+Lpy0cjWS3aQ8/HOatgcmxziOGTAJ6GpjVIqBENDfX1LGJygyFVhl/h1h6Hp6j
4MqmHDAHz1DSvCtsuuLfuM6mbYR88ywX54emzdLbzapb8k7rLRzWUzNNDBvTB3ZSptwV2EDhcFWH
MXBLnfBZetJcqeDF8iHr2GeQ7M75EYF3Wg6SXDt3kumItRe6Iy2/5VZ+Vs4PrQqeuTdp52pzLKQh
nBuS/9VRKvY5oZ+7W8b9rCSIGmzW+Mqg8vniaUUGE20PeUhxNZ0IUj/E1LY3ttAAA7pQ1z+08rRg
ehOxjAnAEWeYkq8jjpCbrvHV5mK7CA6xT6FPBfHK9298axT5rTDy+cnpGlQc09wmX8YdZSKzxSNv
vjz78z21yMyZFzyQxewMt0Va3zEupqhNdn/xAbSydHvf4n9/TTO3NsPEugAeHBGYis6jPRH2+ZBQ
L8UDKlnabIv7LmWxZkCknBqWb+Hf3CcMdwThjiX9aKQ3CqqPHvKkwkQynsGA3cHRnCl5YCNi5v63
BiZHxpyPgqqTa1dtnY5v2paDSfCQLuT9l3/OmiGmqKkblXzQ9Km+2zlNelLPMcTLsUrxcaxzd4uZ
Ftgn+jwxMWBHIaaqHgq1zK2Gdqsrof12aLsTN9rq8yJTBsFHr9PAPQG3T7PR4Kl4HW6pww4iRFWj
ohKP/B8Vxioi/C3TnXjLwW/T3DsVuKXvtc9u9N7cZ6HCX1LOfvUZLm+upcVmzZ//2hs8Nu2Qep0o
JV8xJ5XFKvcWQM+ZtBkhDFpStiVSyrtsyLw1Vz6Ho0VssfCwrNkCNk82ljLWZy7x3xVjHDZ65NCE
G4v7bu3wprDgiLAZmleIYBXP/PaxOv94jYusQsNCQFadvfeWC0tNFiRQHIqTkRL5H8dlp2meQd+N
VBO6vzBPE4ZYM09yBIQGYeE99ZMLPy0e5I9MX4DbzoAtEmlbvlpxWy2L4udwvS3U9oCaDygvQeSS
cJ79PcbjAhKJo4PXSCjOCtYV7D16nuAKoaV7LPja/2ABoiN+QYLywc78G8R2PJ6Ht/fnrYA9q8jd
BD+b6d6XYuuDrpS3zvThMTmLtGzJqtqWwhFUfgjL4eEKAT7m1KIXiSdtRETaKKKGeOPPBGIwof8O
tVSnXdmouKcddPhWsexnBdkWngwZ9ZmTvg/RhjUz3VfRJ8UidOmLTeMEIuVn0dja5RMp2jDfpK1E
S6zG8niOe4gSQ6hjwIoNtndfdeJU8JhqPbtE5cWFQLoXt6+gmjpUCQAKMjkYK6mnjNczux0J4UiZ
H1/Y5XiP27A96as8+Nuj3iu6iAwgTcUJRIGQMZQczBSJwBN7ESf0eA3vEko1aZfwxRQNj8hpwE5I
gY7tVe3zzvsDnj/XSEBAJDOuGupCWeAzlVTgYjFR/GgXqS/TY6TmFRBtGoCAMU9B+8RCEFWGemDd
8uw7HR5f8hv9kdN9pYITPg4IDKij2o9xraEgKkY7aGpWdaNYf/I3sh/vy1EovbSMA3zK97dS0WyO
ia9A8yQ1m1la0Se9o8gVfV/ggMU9MZUKNZPTtChN12v+ebPerR3JG1p7bajHhz4t7/PXeSWOEppx
6sBExYodwLdoIvvreGOk2KEdegwTWw27WmXLG3kzd7vPEQBvvyWlsz/bERSYoR1YfR6EXLS1iBWg
RfzxgXSMzkTQAarn31alC2ndGRzsCfIOIyWRV7bD8wGrMdtoAQbhfcmr88JgDzVZqEClhLAcyvxb
dAdbeHI7PG2ecGFmY7wSaJqYUc8tEuZB6W4ClRupZHb+vYjJa+E4kKQhaDZV0Z9frf4NmKf24IH7
ezv08aV8mZijYz5Iqu8//WiZ4vJyt+NT3oMvbvzIyQGMNKynvb0Nw5r2b3BKcevU0b7zTyuDGS2/
oT7kHj4CRtOJZgD9lvHVXORRgaJ8+f/CPZJLz19KfrDiFtStlWJUwibExFrlk9scay3gbp9EB4Rf
T+2Axn23nrTqB5REqtb+ZeJ/c1tLJQ4nVEEUkO7THjQ4Krd1MyoM9nJe/+8GnHPHKxeI16vRGTla
MghfwWTPa/5bMZoGZcsvRz6Z3+qArOyEl/+I6lAdkaHbQHd9lgsDPPivUNxLDLkjiYD0OAnzfKfF
ma7Z6TBJRgvlU5HcHWKMkM/oCRXGn9wyq3kyeQWkXl709OKBFh02ZwpWay61Ih3s0rrAUDsyS1W0
Q03UKrWUURvzTsIEWP0Can9aoDfbkyJaOatcAkQwZkSAg5eT3eGVY6/P0MfSSd0WU/FIu+vkUet2
oJaEX4ANWyL7fl2iaZI5YNKoaSY2E/ueTw9VQoz3ALSxoFDoJK2UOpcE4nbvSde2PIdjl0i83azq
i2qeueHYPcxxtpkPNdQMDPPlcwN4VDlUJMhRaTAIc1jrGV7nDkbpA2pqHXBDhEB9xXRBtnNjWRmG
70TosFoKR2a3V9VFrcYSkhWPiJ83PHtXwELioxTHVGoRWXY6z+aC1I+xLJF9QIF72B14L/y6+r5e
gYNMKwRBIcGKu8Vu5IqIKFDBI3Gn7OhRxnS+pVFnHKnZtBilKk2geJMqB0S4gNU6XPC8iBmJoCzw
gVr9D5sSoKaz7SBMZZ8qPl8b5mdvnzIDPnZP99wI+Xo6EwZKwrDoN1VkXxdIfLupXj+NTCj12LaY
+qHxVFkzE7FPXUUpVjCupoqc66OEkhhIVSCZTKwhuX8JpuGFi82LUWsM5koW7VE75P/TKceMZ9kp
mOqr5z4AQKlVLcLowKPHnMIzHC4sz+DU+2qwBLCIKR1nDgN8c/Tt4ZM3xOAFq3ektVxFzWOn6K5y
QIWehEGJkd9q6/sJ6QRg0JZ8PX27FP15EfPFl8Au8iAxpNWKFcg2bcUZ/z3hFyvlu/QAzAdwl1Ei
z5GkPjRujBtYBn8O2F0vfofTEXW9kwRXTFCKuZSDz2vtCID53jV4k8I+/1hM38QwprFoPFxy+f3x
GHOl/bxCjnyYGuTWapBXBbQeT3vg/VgFS3ACV/B1GDgthgNKC/VS2HqEfjaQmrk/IDdk4OHe9Hkk
0WqFUxNx+6fD/21NHvH1ZYAqDRXxO51+gbYNwlUcicWpFIbpuU0dPeY3tXS1K3H5kBohZqI0ODnH
nEw4TM/lKBwY2CW2pHx+12maFMUysjfzJt+0n4MQ74jTPMyBJcwMT94iBmh5gU/5ZwJj5AQ1IF9L
ujPkTHPJukcOqBr68tcrmA5fiIMC7bPZH/eydui+NMEFTl/Bn+mq5pg382+9c4FgCkFgNCHdDl2E
rftYa3KPvCcis3180g9vXAdlMWXkeIqu+hQYWsPwn3pBFpFfTxP0gfHsMqhQbK/3ib7TGDCXCkg+
rdRK0gW4oEkWDO3J3X3MQ/rWXLrEm9B+g0Eg4w0ulPSuy5feLB+pLWgUkf7h8LO2etLh6wkKoV8X
gJSvcGEm4Sq3S75S+Im/XepdoYNwIkGn7D1UZK5LaPIs7VNu2ScTfTmp787JfwA1+9zyUZJ6NyFg
+zFPwpzIOwVUSBalnSHh8UMlLNpTQR2bswPpXFtnD1PMhG11lCm94gN6hwqeMhuppbXT18sUp8NY
jzmxQy9WvasqMRgzvzTTXtBz3DOfNR/JGIABCmryQc0vPHs9C1s3s5LljB6Rpb7C1l2XvkfZuovD
iVEnPn6yntXF58qrE1eccUZcFA0+674REZew3p5d71FbX8ygcrguPsXp5Ak9YumFVkr4tTBnnYSh
3GSQMvB7+e0OBz0uz0HSwQ/WXG6gfoSlEt6nI2yJHq4h5+vUIifJ2vLiu5RfqmbVFxP6/hIz8wav
8HAqdy7Zqbf5U6RGT2XrZGLspKQ8+axqqyuidg80+jss1JPr0KKEtQKVdZAmS9NlRYnx1rQ2jr1h
9zyPkbPTcYcfGl+Kax8SMM4E2Cof+1qM/uZLVkDoiu467V8jMQNzdv/DxGBqYkX3ldJ+dAVnAnxS
xeGf87Q6Au/rdYtj61VViAHZyTuKccoPFAHxB9R6PW5vgRcIYMBu8iOlo8EiYBQDOACmaoy1Ro8D
myCdxbJ0gRd0JUxEk1K7Wr1wy3E7T/czATd59wLDmjDOghmaGBadm7jWh/3AamCZknQOIyBrqN/o
poY+wgozFmULUd7eJBXE7zsdReKKcaoRJBQ8uYbwLLBdrItbDrD01F4YSQoqLI/lqWOW1X7l/ZU2
OUrXlk7BBNGgUts=
`protect end_protected
