-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ba/NSltYPbGBOEoUT50CoP/KJaA6228Re9Eipwfd76KPBdus40ayONIR8hxIDHO7kPSfhsr5tJq6
zJKmD7cqnlKhKCqaQQHwb/RTclLPz6VZI2EpUcCO2/jIZXRJUw8QMgUgwsMpl8aiZ0Ta4bOdniP3
k2xGAitvKDMkLvo81byEy8Y+pDAAboZ1QvrjbwlmamIxvJUYeJmWPUbDWwo2vN1f3jkfCpdjq4jL
XeuJLTz1Z8ReRV2FbIFYIxM9kH/47tV5Dqgk0V++VnIUCLBgNVDkId5QPiO+pY5VdvmNCIczrMH9
T1lfwigYlp4zEuWp8cZC6EA7VcH2DISMCp2w5A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
ZCjfzd0b9bzLPsd27qcuI/6HTaq0r8TTaWfoF81qD0oE5vuh4dYWv/Uf3X8rRxXPh1EWDuIFWbI1
+UR0pBD18tKCmsr0xwDRkNFA8K22696VED1/2fNAqN7EcVWXSbKEZeJyUnHlCBn6CsBLqdvy98SZ
mLXbOkh+0XmCUfXdP7Yfiv8kdaB01aM/lApv+RQMjKtHwCgnVN7v2jGF792DMbxgVMaPDcwe7vu+
HJg9wsuhtwoaOtR3ETz+yaQ6rdOvHE6HOfxJ8V4zQCgdfQcE18IaRLu/uZLhHL6ZCqfaSNrDlN9m
jaRCut4VnIZPuHYWRIuvOF5VF1A0KBCSMxfP/lsCmYPd495cPObyCk78CTYf70GrmNRUZRj28crc
CGd8xtYUwVttAhCzgGKsqEgmhZRL92DzrUm9Eys/UQddMhKY9qm0+1AjbAbTkFmRAFsU0tmTWK6o
Tx9dsF1lO70A+m74/cQ3PV04xRndKTYivhmj7jCk2vQUIadf5HYmj1RFRlMf0enLN/l/hS32kD1x
eKOCqsUdODdvxQwaQX+CbwG3z5jsY21p2lM0wdoOr8Ol5wiG4eHkw9WODY4ceNd9gNy5ogToq9ZD
jCOwRdwEa3JVlAZo84tpRqK5ZlHgQTAo8RcUK9/r3KAMngSFJfefRch5jS3V2bI39Y7JgZrXb+fI
k9mj87/ZKaqVrXgb/5sNsN1w83ZKAQjilC4VMuRFhZI8FmSV3vqQCkPK4WXuoC7GE4LQ0oCXqabi
+p9KM+RL7VT9sGWs2wZWV0w0/RC7JTlzkR+kGPSA3iyG+SMVMWoWcbg3bR8M893kF81IMCIy4PaF
dfg7MpHxEPEaZl5ebdV9bj8TynMRt5cJotz42aKiljo/xNi1zJZxkMCQr3lft/7mpVAkK5vlcA1+
i2d83tCD+HMf4ibGZTIH3kMQVoDTAZmzuIl2j00Z9OX192M0cDbY7CA0lra4uRO17MEJ6rJvXpGy
o5ukm58Kn0VcmmR6HEumfH4Reqt1F05TrhePRn5g83WF8dT72g544G3apXs5D3XwUwBrPvHNiTzb
YZmkskq8U2sFHtoPQtoKugc/+Dk/sbrc0ujNy9mrymRyehHblqnvXFqL8paj+OsdKDUNqEOeZUPa
vBbGC7LiCZOdI3MVUMrX6gRJ0ZEe+1WILpiawkI0byYWNj/gEx2tPlhWMXgyeRW/TQg9V9ShDYo2
H313lB5D0ew2+bWcpAq8LU8U0EMvUI2QzTSCLp1IjiDqDDxZhcqXCIFz0Eh+xnwsCK2HgACKzGUb
0/qYZyAFbQBB16CmsWkD6FhqsfBePuNj5s7tul6FRRGuHz2rOQMmV04tRO37UjNuY9yfyTDE1Q0P
fgP8+xxJOOPnSCUd9j2vvDGjSnVYvxhwK9gBC3IBoX8PWDHlNACcFg+wYYNPzGmPBLidMvoxtgNm
0MecB3GRU9egyS/jgU7ORYrWwiNzG8p8dE/F+yM1KGMDERb7Tp4F6uKRZvemvUwaCfUznJQT70a/
dOABqjsz2p3zpvK5cCQmxtbDeknOUKT/UN5rJicQ3X0Ns2whW/RGnay9SVneNDOPIx+y9EzDjolh
N1wMZzMTLucimulthRYCVS+KgkZUaakSGr3VrNZQIKWDi2ZkMYQNQw12/RZtXvvStUcGAB9VYINc
AktNpE3TyyOk1wQXtFLN6p7olmoKlkd69b3SYld1I0oE7Cgxb/3Fs2ny2p06lVmKyuC46dNHN9DY
WF9x4J3nJqWMWvPr7oxUWarHHjgqV8ILYJ2bStWF33XCfqu/sT3B1a8f5abnFaeHycQoXNs4Mm5T
VcAeshOY3woSC6nYhnp+F27H+IAXIrxznIAPXY6p4LP0thStoPCa1lUPOJkhgZmvm6DDSfzqQJkZ
6LaK94ofnqI7oLb/FXEsxLtNtvnrB1Ws+WyUfU0WSZu8SHH+iUeO52Q2XNfy5uA++S3zUjJKC5lQ
8PDgX6YodaQNfFtNJOPnIWdzl8qbLAjvryfatCxfEJsZxSIJt/+XupD+GWqXrxaR6XYCyFwnayoI
6F5G0h0NzaYlJwq4qGcgWq84Vc9Nxl9s5/Cox/DegmiQeU6sojBEulDf9Y6JUw2Pf3mQ+hvL+aJP
3SqBzdMGtkFsRqJhKuxJ3r/ROtsBjZydazRl+4sVzoIQCr04WsbpQrI6aTFZE2KCmT7/n8qxljkG
HZTYByPPI47luBe0LNY9uwvow83Kt9++1N0+U3lFA6pT6xHTHZFyV3r8cv1Gmz18StO099kOcTgB
jgiYsdb32sXDPX6unTIw8e6YYhCI0/ULGp40eucthO0O53BKSsDyy0ZQTok4GQVD6D4axdYSnPP/
Q2cXVs0pjrP+b5L/Z8vFOgtCXoBn2KHQAV3LMAEla6oYRNKT+lAApTBzw3ocletaDHACXiOW75+J
XPIKTXy7C0LJ61pGYVfy/RxMlLK+a3O91zQ2sUsWUJX5XNdfaxBFkWlVjLUh9rVcrrKFWjZ5g871
47NtDEduwH2fKarrOwDSMEr5kPWqzavZJyFWDyCWsUCaEGqgHtIe51rSH7tzu7EaJqJP2hf55zn1
cv6anc7zRhdswwDhKKv6qUBiC/Z766V1K7M4wIM827xsWdhPsBedgBSB6B4GtPCYATEW44EQPFZI
1Q21565HD21cuZsH8DKcSLgZ0KzxkCdWgwbmgTWG1Lk/gy6GI0EmTdrPy2B4MtZkRHqWxQLlA4Js
HuSxxTKmhfV9+PXxjx67WqxYChJHSNwUI6CfgTw2b+C7vmyjkF6PSx++vfjpGzJRlMf6nX6hkwFA
FJXaQXqgcPNz1DvltttsiHEOTKfcka7lGXskZp3Xt/JmY0dIS7xpcp0MPGxqSe75qQCm2YigzAZ2
GkIxZWyt9RHJ9KLcJIO9BAWYu9HQCMHi0aB1JqD+2spev5sSqhtcmOjiATaWjPHbthQaCkExlCIF
j0Li8ExbN4chGTfvnicVC1ZxWY4vAD62NtmeMcf6AkImYUG9Tmn9l9TkBMCEfYvU/AbvyRJnxLqg
7SNSiz3CkR7rC23+SW3PK5yUB+Z+DA2lqkdqySyPM55kDOTZOlKLKWuwgJnro0DMdzUR79znFiU/
3FLles2GgDtEX8JiQZ1OQ2ps1rbZA0XpVfqIJN7X9t4qIJ/TjmzX2pLKaEd96G2ikuL57eO2ts38
t7R1bqoBoU+etemqyvmjcbK5R4GcfKoL9TiY6ovZuWbNgeBxJyYZGp8z1467S2R7cRPhgUQ2YQh5
Sm4WlMpICF8xxuuMPef/6Dg6K+sKN8Ugq+B+d2YsOfFpHSL6uvrLbDhhl+Lab+fvipsQ7n/vB/ar
+ghCT03qgl3w8JydWUnl1uT/8nWep9a0tNarawbh6W4zDPYwd9oK7hMgQxLTGjCqG6VxENcSF3zh
i9O/zBkbZ8uOO+iXO1JP8Q1Z3odtvMVoJ+dfPNzR3pvS1XvUrzpjLAt5VgPlkXzn5/RwSU0E9Vfa
heN/ZUyYJTUNTenB2ylmiHcWyEsPnOY8v/e+/0TfbCQCSMsFOORsN3dT1ncaNaZ0VilQAjiFBTIC
g8yIYy1QInFV4Hoxm0etv9bm3z5yV45DJJIvcUQx3Y7vI9s1HDinIg2vbw2NkK4wzNVUI8lzYwPv
T9ZlC+w2Oso6guQf7a1Tj0JGu+wsLruDu1Vjybd1ukJLy/kh//ld2f9aRbs6yGmKiniAMdVmQK/A
559aqtej1SvQbgC5oVfVRekuHFhFDI3YWP/ULH14a9NOYJo6nWFis922TUp5C47Q5xecwTH5z/kh
5HR8d71kh6v4am90GHmndFIcY0v1PGE0umfGWKI1aOyM47mkIffqe2t6JAXJcUXJd3Dn8SPm3C5s
Adxep+X0MWSSO1WBwzTzrkJEe4aWTqXo4xiSo/ZkENscrVn1NgsSNVnRxJbhu9JOZo9v26lQx822
Ke6zqUQZve+ktMXtEmJkpcbGtv/CSSZC8Cz1t2dS8+VGDlIthaz+cv5CxwNbsoCEQEPSliJGmcfs
HYFzTPFe+ZmVY3uaCxLaNF+yxgPCrPrAgladApU8N7Xgw3lU9FVHBOMafv55an0WuckP+huwOAEc
Sp62bdcUqCcTwDuUkcWJ2wWoofCiHcYm//VXiOrTDZeGwk9W7nW1IBtWlBPZdCpgbupT5W+WbYl9
ibv+Uedp6ZCX5wPXKxoLV+gzimLWZXYBmt9RaIopgOe76KKgVkGlhqK5vZ2W1lgmMvMCyodNUG6i
4UnVAdjnWcBcsy4wC7vFNTmuZklHUkV15lr9NZrmV2urmOZbqC3n3U6hvkhHAAupMG1tbvIdKEge
t3SafSSuAUZm0Upk5j0HhARt0mHilZGcoMZ+kenr0XguU3f+Atdf1Ee1f6xoROvtdH/fxK+vkPWu
9r9hv2qNhyetE6wg4CwdqYrdI59IBvARf30RuJBCvm1HWSQL7BMHRIzMb7N1Vj/wXNbxiWw77fm3
VXbuDulswgLE+/WtOH5Rv78RFt2ajougk/GNLIqgoUbiabzoHCPeCv1pV7KpV43ICyeIWTHXV2iF
nQoBLMCSgjsuADR1ZFrUaA1cTbk6Wo8Pbvfe/R7F5f02gUqBls4Ba6Es/tZ0n9Gd4sqTwFEaHmeo
UzCE1S4W7tiRM+zhiIt3BmAtkPFuaXEejMOgIPWaHZIbQK1lzxv4X9FcTlqhFxcR1qnbjzvNIFEL
+HmLaiEkOQMBMgBl8jilgPL3hdoiW1XEGiLRHMNa488NsMgVgwdRUVVIPSXSRGS+R+7zlZOnVZoS
W4cSr+iR2dfUQNegWgIhaGeYTbdkQ6Yx9R10QXMNo50DOGGf+1YeQ9DEJJG3R0VzdeLhquM07GNh
IGDtd0jsCJTHLvhyG1+jpAxNfPaCU1FGqqM7yQVcW9AIlL/zxp4rzfRP59gNehKoFhpYEZO8KYFi
iox80tXO8YrH3UrW9unZpbxjWJDVBTL+ntMvOT68bunMt9p0hVFWhjtLy0ZeEwhet+6UpgENEOgZ
k+z8+hjIjGtWcOaq1qszPI9XU7R+Pgy9vHAz7yMJ5ICtl7h9jhc4DGXz3CqDcCabBydiOUyPHUVq
ctcNfJcgbvAU+XMkvZLfL/pZuXsYMUoIYgU0jAKSUYZQpIjbHHmchgMoXltYq41B1FRZGL7N8JqC
h/BKg2vWuRKdPSXWzS/v1rho320Cqf9aS8x2CSGmVIQXEWf6rCDxohrXWgiKogsW8xzGWW0UI02/
YwWtZTt00TQVBOagkBRVxiOUBOvBchUdScUKAeGVU7FS8jahUWjpBjYCt7Exi7hbHo+61ETI5j06
qUI3cBLpCNitmhlxLziCQnpF6kba/AiEMkeXuLmfB+9FJS8HUGPFkVGAKmqeyTE9LKyUF4Sx/txh
UldjglvrQNabZhjPzcpnhHIxTTbsEjKLttxs72yXSaZEXHyT8iiGc2Nvn/SY5ui/h1+npirdFbdV
jfMBWbmG6XQNeshoQvsTdmnqcZ0DQSpQOPuPRb8bZ/5mLSmkeudoqeMDRdC5F+jT6zDbAPW/lcvc
BPGlToz1oR/FXFO41nqNIM7K6GwAv9ZM5MHhSILapEEO9gUI/UuzgRS1Ql2ikF14C+o3KZbppHa/
t93tqEQbMBxYWUh1gxx5jiQCddLG1mFbBXr+Tvkx0KbH0QwcITXZnNq6AmrWshrpsX+a2G1xBFFo
Ck/Rgam/3UcC4IuBghFIBhs072+U4LUT2LyNKj7bTVrse4S7sJYMXq20FLLICyfnAIJp9yPX0dxb
nJmLoApqEt8LbDukIQA2zxJTmCugybVe/vOBpALgHMAQ0PBCDVLHTYKWWE6o8tgcMqPDguKzI1wZ
BtAheJpZmR76Fiq1VIs+PzTeutHqszp+ywu3VeaiXWVDR6LDqZ+tyRuLuyJc+KJ9Q1QBuolaOINu
x/bKF3r9szudLE88Sl9n93ee2Ncq2oXtEG6tJTdXDuRxow7zMM7NiEFBoh8qC+HamqMu3kb9CnXA
/l14SfNNve2tgCa+go8253B5UC1/rLu7ORL+FF5Fb38wqsRtHvtDXWHHqjG33qgldQ7ZwB79QXHP
rjlcSArPoN84NmQ/GD0Pk+0x0lGv4VT26ij99HMJ5Qns2scOlffhnAYETEaux8nKzqSQAtS2U0eO
QRkMOr1KrmdZwwe1h5YrWSkhmtYv7YtwavsRKwbrHM2GR61H5YAtNnJBm+jag59pcgVB83SA1Lae
SkIYv5y6TxQllaakfaxWXyp2n7xTyJaFrk3h8AgbW6WO6/1PR1qdfb6tRehCQ6I68rx2pHxv+M3l
9Y+JYZVmY4IjWIjhjFLHJzVSkzYJ2IYD7p04hL5+OYOUBcE5mXL0N9DtlCEEqddYPkQfXuqfa8iy
/IrfUoZvSvkNjqwCBGC9eotZKm90/24FZ7t3Zy4FI/hVSBZB4u8KSnWGRRvM+adTj2neoq+e+pVM
IJM7hvCH2cQ9BAsxUdXew/VXl/IJyKDOug5NmFFuCdP30Gtq6pWDtjBZgh0iV06KZCscxEKSXBNI
EUIyenRtlm1kmEvhDOgXpx6iHVQ1PI/6VmVGzLSQMZjpFJOa4Idz2KHLYY9MPrLTHcUeERnvxReh
bNRA/gFF8y6V5Yz/UDYKZ1V/PvtuEF8lkt2cQzU/7Xd5L9X+fTE816z3ObhcFI6B3UYFm7Lv5cIy
Hl5+XOI5LgzJsSa7Z4xpwyim79Kja/dVYEcGfXCE0n/OxnGVGeAgBTjroyqneK/WV/Tz/wHuXTQR
d1tsUjnJqnTJbVY67n8HoTmED6HKChNvCS1C6kLagnyeOfUX5dtHXoXzwSvc5PyYCzd7Dns84nBj
kpNGEX7hCW8gUrQ6wlYH5ElDkLVUn6vaN6vJ48tRCVShng86Xd1UGpsTPe7cGM7k9jZ11AR3rPBi
nXX9RnuQBqT/c6Mjr7P1/9fRwwH1CckGdmSqaL9yyn9hfSsWl/d0UuMtJAzVBAxZCJC6XdkDoyqO
ElUJ1koHJs161nzLQdAXFqJ1hilxCgFSSDflrHchuuBlTMHmOdvXyftJlbwK81sZsb3Axd8lLwnh
PP/4e2fg9Ad1o2OceqwIUd15pnefdI1uyG/+lPW+HnWhJirhUfPMEt5CIrNYXwVKLjkRlZLHXqbw
nWHxcf+x4+MqotU6hMyj6tTdO1qVbn87wOptRxrFbFkeZQiO5iNJxYp51cHriLlUQkmQ5JmPLML0
uSGfLnaUeQKG5Iqs7xf8vJilhI02IjAeNCvaoFwTagB/7vsrRF2DZrdnQT8Chswo1iMg5fnsDSc0
gc9nQhQ2T7QLIDYIaqiqvWz0bX0yPYwJuvp83wrSgJDYagWGHvPr7YtnRYaRY1GiECIWl7xUUxUN
hzKAxIJESt8JJVkCJ9Ex917tBvg0gbuHDSCb6WAjjOot/TDQFZg8EsFxTqvWYxlla8VaWtRo3hDW
w8w7Md+SdClZKoSsTecwgQrUEGVggLS0aKgmOw0TvALjaX1R8szEgfsiH1NHuQuvVsIOtejsu7S1
oe+9H+FEmx8aqFFUysrVkvrRoALTKuSgL66zd2ws+aewhT5Zile9aE1II+cOTSVJP/wWBBKX5b7v
CUqA8z2vJSbBXWzpBQjFhCZFizupAieIR9x9OwF9Dnj0D3t0pEY5OwJ8mT+Plk5IKMiU1aTBo6XL
2QVuPQ0p/BrAPstuDEBLYXxqWgrY7xLmWRA9kF//dRzho+TTGICzFr344MLUuKnxi3j8lwg0ici/
uzIRHNdf5+WXyu6SeTiQNLUcMFDEPodqVnCOoUXKjvEdpCG6Tr6gK3T9MvQnRcBJ1fGmD0ZCeDeL
x4sqtl5KRLdoXAwEQmb6ezkZTXVckxmNZwaLCx0/tAXX6yGa64rTZro7Qs45vTFf+19/EkkhKLND
RGhzJwbvkzvpXpHOS9X4pjrAyIEG1MQzNZoR3Nwv6zbPbVETSMWDt5zz1XzVtrWpAotCcpKkd7CM
jTKrjP1Gh79fznY6at/nbbpTG48WB5P6WuE01GCJFVEA0v2E0NKmBYjNEUp95lVfkC31omenonb1
D1w+mjr6b3nEAjZqDaovBgswHsg9cSzBOIt+TlsaUzaZAFA/vHn/GwN4Pnlxj60uy181OW9blI9u
e1pZoc6hQ9/h3t5eOZs9Qo+8HhCGmxu1D/LFzJI0szDndyfIk6Ppd20aznoU8NdLvxt0MUvlGJQ6
EHeRexlgAUuIjm73ZQTUccyidje80IeC7iq71PZHcBHc+mBBnqtD7EW2G3CnUKzxX1bCO1kTkBAM
hm65o0076gIpVAyYC32u/ShBrSqLB03w285vZJSOtRHHRC/Dsu1VQw7kDNz9jXAd6u+YGHZ1Xq3o
AdxGtnjAvT7jDqHhHq04H3kv4Od2rYEbRwLIOQP4tY3vFx+2AQO9LMleCmfzJY+vKbMR0K6iZ8td
SAwcWGSfEyycnRpgUV1aYVSNNy4RLw+rv8W3L8LaHWFRSf9VKcDw4CtxEk5CoKf+Q4XV+bNQ2S3g
tGwELB2J2zt6cGla/1rBSWRXRE6O6YcHXsUPrQ0QUBR0Rt0cuCFo1P7Fyy1Mggq8tnVIi5LYoUe0
i0yOk3GcFLcutyEDrYztSTKxPTvB3yMTjpxjnLtZFWYCJuSS/8M2Wo4noQ7qpq3s0XKVcKVORnF0
+rqFoedJ1BkcJmD8COnLh3WFJRzTtyP9cPP0toKEfQVnGhnc1cWZYv0LM32w7bInNU1i98fdttj/
sBGaH7CIYmmPlLJWWuB0VMe3bo+SaGacwbS38YpFWHs3kqr9k/2MZLqshunNxB3WPYcCgKB3kFD1
3YvPAjo0sQUC97bpVoHmbw+X+Ow8fztfztUNizse9RiH/yVVxYFNO4bHyi21CcP7AfbxVqpq7e+C
r/zJA2jQbRrEtRc0veBPhOwLAT93dVhcasJIIWjDVqpb6qCb9DLjG8kI80Ri+cupDG5K9vUcB1TQ
pFKoJ9Uc/7RItpgqMMqHnjos5VnmqyG/4iWrjbt3tjb3knx9Qx9c+lBzkx4uEKwDgzj7Iz/G2MGi
AGKyx0f4c0OIm2K5S6Hl3217VZV/lK5tQq4PHjIm72aoADnGD5XYCjmR/PRBCOuX13u92qaLGJNb
hkbbrtQkbn2yy4l7yjqF6BU5plwPAbNnyS63MqA4dXgcL6RaVglfKQlvgGpUjNmN2vLDvcdMuQfk
AnykhYXZOVumswFSVNQvJTOCXakdpinOefeJ7z2h1BK/HZPNh4zQ+Yv9v+GBYAehZop1O+y6LDAJ
2r0GTMAwvqwd1J9GENL7suXMbV4AgRh4V9s1754Fk25fOPM1MaoOLCT5bAHvhIBGROD1AQxliSCI
qFDKkbAfVhBlyMgBcrwmhMe9Wp8slO47+EK6xIhwsHzDKHjNbv9zWZOAEfdl6JZhv2FQztCWxVPe
7qdO5yIoccDZhHTQetnw1rqPzrqL6hJNlmkNu0+1lvPqAZgyipfBKuST8dLyWSzfIGOe6CNU4hvX
kbwDpAsNb6ZHzAr4Rft1Mek9U/wG757ehsbZA1mVm5ZV8z9BX2giXAX5I8yh1E/JiKwhfQcXgcy0
mSBStzYj05P8luCJEMTRjb/wlbkeQIuDrtAjTg8nrXX8ZrpXB2EhR/30Yh2zwjBTDEqREFJYWE0X
4CsTvM5toyyJeOZFEicidcSS95mzAnn/9sL6P4eoC73ezEvkIvV18yamu07erqayZFWwqeJ5jqBr
/3m68Q15eJxr49GerYI3s4yPpMqIa9n73nW8p5fytcwTcFxpCEs5y6JZgIdQAhL7o5kLyXvIzPTI
+qmFuSzEho6Ej74o4DqHIh3smhnmfugakzSVvKrRflsbJgU2jCIQiecEyu4tk8ERtw+GrEBpTYzg
YQ948D+b/H1liKXA1eYiWVOie+rj3i/5Fz2YFEX3/k8PdFnoSlZas3gV1moq9Z8Zww8DHRW4k7v2
WhF8JI9aj8QJMqF75gopqoGIFosFvtn4sz3z2z2Xc6H7TbEQnHXpdp8/U9ktKRJrBBV+T7jFOQv3
/gW5yuAqCcGhT5ankA3RD+603k+FqIeqErFG7OcLg4fr5T8zCAjZmDSr6eecVVD40RKuhfoyzxvj
V60tlxZCJRgmhZYD3i38Mog1/APQ1p4ph4rEfYWzDIxqczd6/5qgHIVqAhsC+DPQtcc1luYBI+Zu
Ibiuzmo4tv5EeA41FUYtjZt0DbC30AVlMIkgzJSpWlqYuPr5+cNvF2egIX4jZn1mw9G0hv4PX/NH
Z4WkiUXKlDPjj9O6rKZu5bMXVEHE4JtEOMf9ZsrNi/U+FGjhWlaifLyz+YM+1G+c+1/xTOJfGlxD
ntHF2xGA+eShkuZsoi+XpKXM6RjgWSXmAnOroL9rLDrgWOKi7lAcyRGIVdpYC7grWDBV2hsEaxQ2
vhRBJKJRhSM6cDRK+gHJfbm5lSM18KiKr/MpSPMF+Dma0zNH8bOehgXL2HIUsQPVWzo2hnVczpoq
gRpCopQoyxbXKMpIDG/F2KKK6ahR2ctrSxVA21hQHz2uwWyv1uCy1BgQI/29v3Zfty5l3AVSDpar
vql943oRX65/vFT6g4e+9+CWrgWB1V0Pvhc+XcoJ+7XbakKqxOaHxWzu7kjtmaQNrLDoimkRz0pz
lwr3p+95pXc9OXze2/GzeWVN3UEZIVIoIBFGrCKZ2yovlpZzsjOPohiGa7rbnicjeNZTCxm1pAc5
mwYUivZfu0pwfwXU3hW4RO1kzIgTD2Y11/jrDT90itRRJbfYZeFDEGjDdkymkYBx1t5PPYPBY0zz
qUT9IWHjeTNnjVwEkI9zrb+3H8GjXd+YzNqbtLBPmCF6HVmr3nc2sC63fMvOfOvgeYWHYuHYzqCN
uEhgx1ewmjHay2LdFe1mC7ypOtK6+RKvQferugcMYTjlN8w8uC0oU5n3Eo31iI7luf1LZbKEc0WR
FPTZZZkZVV4cfOA1s0HlwS4opbcDEK+TyjhcX+yr7YBdzdW2VynsgsfU3ySAOcHuNZ73I+AKsfqq
ya+w+zbn3e/v0xD04Cx5Q2v0ZByF9epwFhlh9k0epob9DHNq7kmETXhE87uLQQ0lMwW/GJTiHoMb
IpZAW1tXE+yjdE8hGeP8vn0DSvc8UCfmLHd1BrbO0tf3ARRyttt37vxxpwY/56hdw4LCOZuxsjdE
57vMx/pM6fm1QGW1i3D4E3R8ey6wTDCNJwDq1N/NPu+RE3VxmjYYUKc/sHCo7ujbjZ0Yy3aHN8lb
ZvSqPyW8jAMoIAL5u56CJTAP3056oF3p+oNJ8ECS19thhU9r+jWQwh/2kDJj1PnFRHy3yO8vpKKq
e/xli9F9BkvlkhjotH6w1YpKXQWIF1o1uXDzZEMfGM6CEv12hSst6doyEcsCTPHOS0OJ4yytqfAa
g+kbRFqYDrNWs0f9XUrBtCSb06JTY//mRz/Db83AaymYSQ7SXD9zgIC8OGLOQwAln9dGGQ5V/jtK
pwqRqCplXaet3XGpPgP2gszONH69QzVkPkw6Xfh37rWSyNhUuxnW7G0QPR2SHcyMhi+9ezeDXbVO
b9MOeqQ358sZFrpFh13Vo45WUUqZREFK6fOqGRSUhPhka731B9nRnW8o3+A67hV11mVLqaqrtCuQ
WvI0hJKLQa+oirwfOCNsOIQcymcwcKcSllB7zAwYynapD8Ww2tGL8sn6HDMI6LaT4Ob1qi3DvYIm
6oy2TXmQc9BBlqMYAjS2Yq7bAOJs7IooEFc/PzYTzDkI/HKmuvAETkEZMWC7rhQn7v08/y9UCHez
OGQwhSqRqSQkMDEsXY1S1YaquuozUzPQfHrg0v0Cf7KPg9jMJHAZGJieHLutqDK4LoAyj8lyLdbW
iAMrczxU/6XMFDHf3feDbakMKT0slJWyn4RwWGqm+QtNbMz1ESCy9jcnE7b+eMEqsraj7uDS3j4J
boGaAqm1ecQaPjPOywopI3WI+4Z1A/z7w5z9J4e3Oxo0Oy4w4G/FQ6Yun8xCZoxqBvs1yYiRYPL1
srwccZ+zrfTJpsTbzBO9NQsHyTVHDvPV8ZNsAbEQixG4WuAdt3n+gAI5IQbKrjnqfqgTydlPzTSd
/vdZ6ur7n6d6+vEB6Ln8bl9SCZNg81JxyM2ddfKQWUU3WLzXPndj9WjXwTXoAFQjytbEaIaStwlv
rzGdV2qbecyNBksevwRh5Fr1WSCmUuPBH6NuFtaPXCOf8IEGqQFyikAMs08SPk7RZE6MPWcvBGRf
HhFhSCEOVqCyA1AyzmBwtxGuzr92BL7DaHUIv43zvzTZxQToAiH8xxaJuCMXCTWX/zuNXvjfmiin
rzv1FSvRyBr50nEy265fWvs3+/rHE+BR8JxJH22janAUach4mI/sJZHT2fZ1LtoGsUYDQ7XzphCw
/3RxYXGok/DsW+ae+jMcu8gc2lQHSG7majva3ErjzmX5tHZCtFCIWkYTOPHFjq12akr7ltkuCRiC
MLZfyog6wLpXYtoBALLJb3sGkeSABjkpVTwmB68NBiXM4qaRjQOjS+pL1zj8WIVHW3X/q0059+NP
vaDwkpMxBnhGgaQSrQ/+VNALZupwX2J9OFVXBrRiDanjZrpacpk7l0POhGW3wwfM+XnwwEMy2/hj
c6GT2anEoj/vEnzyWOOA4MBvFrACsGXWkn32mrfaepDTOtuQQugECRwoPrNtIPvPZ+n2mAaUzgWS
6++SSL0z72/8hYlRC4LBq6GTYFy+QFsjutFLqmnK3t4h14C8uXNdVPDEKC2v6hoJwOU2ydJgiZdR
v4LpXbw6L0buxduLVM2VJiBh/eIvVbEELCLnRYDV/ivehwkTaR8q25sEmVnxIHtCjObkboZZLzgW
9WiqL5uZ4srHJX4cx0BFK/akXoot0Yb1XTlV92+Sl9ULr3N73XBMxh0mFc8O0qJv5f5tC/SEmUsg
AQQqmbmy3SMUS0e0Y+aa4wvb0XLFrKG6D8kUG4bh4OxJaEJ1mzcdfUUuS4jnbga+p9Ng0N7da7tU
G0yvWL7ZL4DkAWrfKi1Rt0QwudRsP0qbiHC2NH6aa8CFCTojAfPrp5au29d83EH/2aVltqweISel
h0zE33fVFlWnlW0WCxM4DKUYUFUHSKZWYsR9XaCCoSx83TEuio9faX7r+A5MZduCkRDy/jeaAcxw
+EYuqRc5qf8ZUn4F4FIMp7zDsaWh8OXdEzdngzjpswRI18B7SXefD50PSaWB/OdroQlH8ZvpOObI
xu2D4xgcQqmtQaEd9d2omLFVT7M95nOaBaW20KBVxUsyq1SraLqaYA7oWAaSTEOTV0ZWOS3YEIlf
ckXItVYpcYraKOAU9KbJQkzdf/6ipfXWUUff3ukvi2cZUJ7kG5eGiXl0W+C/U5SbDT7t8OyO+9Fe
2zPza3poErfB76QYXeXc81TFBu7XmFxEEnfxrq7LGQmY4J7Mvk+JqWX+ThNOqlclXlE74YOCqvHB
iBlIX4yEax0kvZnFNPuyNKgTzSU8cKE1C3M0qP2wi3NuEQnsUg2/qE/P7BM5isBEl3xW4n+hlN1a
L1O0fKc3ILDIrQXacnE0ROgxd6fwSWgRDjK0XwaWjCZg8gj1N45jhF9abLGXlkCeSzg0JXgNiS2P
QetqaLcJk4tc8YYbhcv7OunsIWznwT7cab3147t9yVp/pU2r0oGseEdf1RiF26UhbePwxgi8ERyY
vjkk6hooGizfP5diQ5UKZEgihXfHdHHDGBhRXHQbMOKVTrph4FeXVZhW2oZnfhqjP3rGpsai/niU
RV+A7yZxrdah4RuVr1yFx1cGdvuxmR2WCb21tTBsOO2+D66Go9fgHzs+7EfoGZWEqleqBchNcWni
p2qEKTMYbtkMq+M4JwhwqIb21732ZzFg7AkuEa1XkdRZZW/pcnc3SpRVfRcj8qCTq5ounpu6KywE
KDLP7pcBFhwZksi/jYsA+ilGCHGkI3R9qBFdWjpE3sr0ImOJODfXNtt5toPQXccH6zJjnpFlCjMS
kK4gZ3R/V2JLC1M/bldVssQtuk8mV7iAZpdp2U3ztTNrydVFn/11lAlTvAZXnERnJMAYXTfUL3il
GPggukxu/uyKEuaA5vWF8S0r8icO0sjKZ/0b4n4p7Un8lqs2P6BIoYoBUL58qI8kt3t0ZOWvmlIi
T6h4zwRHAUXYlJ7H9a0bIqB8mtsv8Fx9xillw6GUIorUVMAtKrDJ6DW8Cryj4zZRdtwaCsDwNShG
y0fCcSfWjOyz3t0aHWO1T1ieELXKBbYxCyhXiUOy2aFj3bME1uM1kRcZl/J9m6ZINJ/280/GEsr8
phZP9CvmTnD9EITGnAqoa7p+nWS2RtPcMju8l2pWmvdy0AnU
`protect end_protected
