-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
z5cfcHvHZTpbvXLza63zkdtQei3M96voX9NFLSRhFsQgT8bX05M8Qx+mu6s0OZng/DF5qfpWc6ar
ZwMqvyGHr88jEmxUgUrMye/usJY3l50+n0brKr7EcCS3DuXDOvCvPk8tPylzMPL3ekg22YWo2bTI
7o0AMZ0/+QIfVOkY5KKnxO4CYzdyQqeGs64gcFmO2P0VtBHIwkF+5oZWKrhn7HmWcvwy4y9Onumf
ci+bXgn3WT9Jv6bi49yNXTKiXGP33fhSR3gMg27zXA7V9Y3JsT6konjTe+6zrcC7TSh9Kq68M/Uq
C8Ai6dDn42nQ/3GKKM060ml4KSeTdmrA1szUiQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
w/qX9TRu8MTUPtvsDj047tAeEX6rHoriinh1cYYv3xIeckmqOwQ5S4VE5L/eIhdPBt2KSjlW/Ptw
U4I7X7LXafYtuSnChHOnq6c8FuTmLzveygubx0XtT1JmyhDyY6bePSjXEip0YDnYsXBJTdzHv5wy
H2yeZ9TNd3VA6gMfmHudZwHQXsBHXRmpt5PR68jQm6AUwnXzZPlHNAIe+zHSE+ZBRptEYFbv1tfN
QKM0xCMT0qdkqSYOWyNcxP//FfxDmWQn2iaLrCwvzJ5poqfi7nTv1SpGHJr5ztsMoIkfPlDHKHwM
92M1LV2TBrBrnal7elEv7Y1tQFoMM1zm+my8fj893YW066VN2VAbeJJmhurC3TJOqqdglInMYmMc
FSqxkBlj9JLnOFfIz6APHdr6ojyJtELm+9vXURnoae5qz321tCZtgD2dM0PEnb8XuF5H+zQ845uu
FFkOQbwY1Dh1g47gQOy9PDX7ePRqe0tszT3j4pob87oy4gt+5cyGMtChUVtSo0HHSjg1UVFG9J9M
MOkFvEev47PkELFqQlTIB1SbNz46t/ctQbiRjZNJjbTKUxMVxhmoujeypIZ7XPG5JkH0XvIMgdSp
UBeyOvWo05j9LPDKlU7OAQrhUyd+/uuun46ab9ABLuhew/WzIfM6CmdmupwMqKr+b6c4foD20eNw
NLhz/0hVEH/KfsJb5PBgk4FWBEqsEIJLKKmXPgjVTRY7q7aN85+dKukSurAYVx2d8bq0RLjNmHyP
4mPnwk7yJ8+YLMTOYu/05QJbjfy01nugDyg3qOddYl/yNUIJ26GnEUrwyuwwEmg7DOzGW5oZeynv
eCLzjQ7/W3LatY8Ebn7lafrC1XvnK2yFV6OMohlVKB9kw7q1MZVq8yu7BSKxmXYCacNBgNWcooN6
3yoye8Gr221hrrBuUnaEObB7T3WNYCMslzvDuPH4CZEeOz+NUuRaamnDXmIDqX64B6OzvJvhDcYI
WMLHmJwtzhi8E/nSpIHmj/1SLPMPUmQYDDvL8C40VlnYKFbB0aMOpTDoETYiO5dPKBxbfOBpNRRt
VdGzY9d/J/NsX+caiTRg+mLDyF87FZS4g88pfqg/ZUuHmIM+GN5mj7XwZ8RKmMT8eREU5y9bRFIB
/MjHTm/HigExP+IJs0Mdh+9Qr7PzUvRpzqgfK2TJ7tVtZ86fo6pzGjt6GvNUJJo8sHPJ2pzycx9c
LrQ3I1JvPChLmvLiWAGdqsxLxddRM+aLF2RbS38lLU1OIUB75QVa6YUIdoHPqXeAizQAuiWN+2zD
xAwe3/SbAi/WNQQ7yDVHszsDL34icl1rig5/nYg2a0w0WG15QqcI/8JviUrQT3FogBKgzpFReprF
eCQAl1F8T/ToFR1Kmu6VLks/1BdckyE++VKj+KVAh7+wHRSXcs6lPuzNdILT5Y8KkF0iXMv4z1Xb
bvQxM6M+xQz2yOfk8EsTdSpdUoKLEFPzK16Wy5TV2EAqWvQu0utEtYY3r747hXKkkBcu8tOWjZsF
g21KsV06WU55ZB6UC8IfscnTaeKLcEwWA6/Ehs1CzwO2xkG5QEalgDDEzdwnnT35QsByqR7gxKeJ
JoFZ4ZmLlxWMY7G0mjMRqNKDzHIjzQlVyKoms9w5MkW/HYGstkn6SQGq6++r9rlf+JNnfBEc1Ky1
/rJEGvYsebF+umX7Md5JW4kiE8LJYWpKMj5UWxDJ/XU1LBUH7D+2Im8SOhPDfLU0LDlRpFwp7ZXa
uV7YJ9dthGGRK2YaVYjfxDB3OFvJdPJj/QtsV27nnVWUPKixQFjCuxnBwjw2jMcKtEpaROnsuF5O
KdXF8R5hTqI1OwBb6rD+wY805qCPAzXHJe2Lv8EgXnvEbATDd8MGNxqero6qau2w/iUE3F7YEvWX
6UmDcHamqXojC9voI4adDqGm60/+h2HLqtr1nAUpDzo+YmfI9j0pOxx0QlvvNDB8zFXRCXpOdiYE
4+6uqK9REkHIOOkiiTa9VjmWX6GCRApQDLCBy51k1BcWPW8oSq/YqOeCR1dRXGkKCgM85LtXG8Po
E68DUhIlHNUFnFb/aA7O/3rwkcCLoI/HWOynZBBHw/JeUFsZycIgNWwkfTsPDhDAj/ifMXx3rgwL
BFqbssYGhUQ+/hjJW8Na/H6hBbqzUVn16N9mDKgbfz1EBKbYODX7yEl6lHuDbSMTSAvNiMtaZy6u
hA5hj8UTuCfRj7yFBaZA9aKO6yf51E45Gij3pXZL8C3kwrLEWyJtCk0ge5xui4/+ikN4wtXH3vEC
l3vivsAKPt2ay01kBQyML2ZQTM+OQMPtd/8HpFmYIb+MDmC2/A3pIhbCOPv4T8kXF9O5PbhKdyKg
0GJwNnwdnQ3DI37TMI8AlvrdscTvRt6JPk8JltS/YiO7VXJI2q3QK0f4LhEEDmb7EUF+tcYMmpBa
1WLx8KK/7Seg0EB1VlTP3LzhoxZ8WkUZuAylZi80343S4C9woTH0ZH1Z35Lh5v7PFyJovnVkh4qE
xpwQJWbO/OJQm3Mb7mk40Un1IwiQ6b/0F3uKF1KFclBPv+5T/Nt4le/9KxdNfM8Mg4Fih/cfCeiv
KEgDEqT3z1i5suQQFwI5FBmkkjfRtIpYV2OgFzrHiHhuwOxJvw7olsa9R8nB8e0POCgydGpCWZey
JJnVYgsHXID2a0CTGBaq37xiqhQI28FGOyOCxbymOOWNWNP50lRCKTjGfG54Jb3FLLhRRkZ29EZe
5/stf9Vykn+m69tTHE/r/2EFoUldyD0ssFzXyqcoYx/kvW6KPkdGMc+1Oiifx3svDC+1Ld8Odbc3
gI0LIytRIEZSOcqyIER/dGowuzAEQuAr0UmCxZ0+91s0Mm6L1fyRHa3BSPJEsCJYHuuzUR1oAxhP
Yf/B5dU4zzP0KxFpF3ejFP6GYLpxIfccCNFOV61rVtT/EAoa25Ybu4szL8shm+nwWrTxx9jba3mk
ubCJctxedoKQhR2nUhQEBqNU1XCu4iQfgRgZF932glzPS44N+RAU+AE+xyygbbehO8tRB7keewBM
3IEKS0AXxut4w2VjivHGgixb/trn+fdINv25yI7lcjWdWJocq1I/lE0AvYC7xJ4XKsXQdc4VCLrn
hqXXy93f2bgfP8/go/c7g19HoSugITTv0jnc0maA88HcrcwaBjV2FN+x/wNrC78or+jjrDg4Xbps
R1ayjPay2pkc7kZCLIjII40vgCeZXMeIql2mRkVx1hs41Se7ioauUu+iiZurKq5ShyHgv3sLuz3X
Oes2WvXmhjuUeI1vG/YjOmtDyyDKXECrcCW1jokC4C4HjvZQiJYt/5g1ay9d7i5n29gawG1IejI+
eaJIQYdf9ixpRhXBCZ1WSJFGt+TqPoRd43OdDNCqZJBViHN8MnkJs9oQT789SNCepei647ySmoRW
ToAVpbGWabuocLVSFvtzFUV6fzXdZW5zB5yukexzNH6aq/Y4NNDqdlBqe09iHv10iGlJv1RPL9Y2
8g5vYSo+PDi7yLmMkHUojl6BJ5+jyAOiA/GIO5bQq1Rlhezw16SxP0uUehYpr6iuJx7pEzOS44xo
YAMkdlzIaDziN92szoUwuyEvUB7t3a4WQKano5WuWglSAGdOGClBhPEBbnp+mSAgn8WMgTxYisl4
m3XhGFZxI2gexRIV7d/cFDSG2mWx6dtuYAS77R9EyLCS1MUQMFfnclabsnDPg3xEYoA3EPeLr7BO
xwq68u8vBkFjz/wUoojyHPnNsFhIK3dIhGS1U+Czm74efPtENEhoS0LItUtrapatQgpyF5hdIErm
SR6fVsg7feHODLKr/zXGMdJvdmXyFUcLdoCGYayWSpq1TWXAJzZEw/mPfz6NrFeJsogoCgvDxzvu
8FAUY0Dc7RAct5eKXvVTy30ptglgciRC/hkf23ZaU6pTy1fMYjOiH/tpbLCTTPpxxfNa7t8zJx4O
V5ODtG1BMD1SYfWAIPJWChvRvLnXuBFephX2QimJ2B/XjDrN2em1H3tWPgA+PRNpMUAkbZcj9W4t
Bw5exWRsjdjkrHv+dgQSKrZd9oliPd8RnpjV3YbVRipKZbHzeT6mHgK/HCaES9C+okV4J6PfQzjo
rgRS3NAzP7d/BE1CeQOcRtHKjG4YXmzIKc0QmWiYvyOMecHVYDcR0Ag5OAQScQ4ct3gzkpURAJfO
8lMaqJ42VOlmqDxm4kLGeTa3FSDcvk5Anj2jCRuJOPPTQbxd5laORy1UrjWjyBbI/crIwBrBlKBV
99cEEVlUjA70jpXGupzjhVUohC1w7s05tX1lbHMFHuxQrQs8XlOFt0yHGxGi2+iR+vyQXDHSiDn1
me+5rXjzBYmbOYwKqu3v1/K3nbaEWZVA0vOwfER315PRzYyCTZz4YWGslXY5kYUOGDb+g9b2WrMM
y//7D6IxL5cPfEqnKM38UzT56uqaGsEF4bxUbXy7XRRRqAZsLMdjsoVXKTEeS9yNAgb/cLXBI/Xp
OsSry6UonK9v/oqjVNeRIbSgrNPlJbSGd4EGQCqf6Ew5LM/X4IOjjNrN0fYl0WdCuiMDSE6zEFtS
HCVE0hYfEJkRqS8WQo5I+c4hlaAoioKq1kQCR++XUAqdX2QtMb4/p5NRq3Y0Pf+6RyOhTCIR9RRB
rCM1+PFbw8zUdeLz0fp6n1VKhGiGh+CMLNMG4GDEP6EkjS01XzxW1LbJbi296d8LyPLARbIQ/ndj
2M7CZmVoPF+QNeFDj6oq/r/MTxO0JP5ETPPJZ2EEjVkHj4sHc1MT0lFNqOEVKkdoqIkk0pn8Hb8n
OUMUyoFxS2HNlSjvaidIkMe034tasiYEhZ59SDxJfPWCTCuebIQcpe4KVFmz/2sttP2Uwv6Porxq
n4f9pWdOheo9vf0CiQEnP8sWr/pCURvYUze+Jh2W8E1rS/wK3SO4RFv4S3L8xnd2MWqOIu2Zsbp5
rxq5wim0r8loL5faJ4wkts85JFbLiE2S0nO9ZBo+q99m9+hFUaxgxn11T7ERm6KFl8BHgBF3/xwq
RGA1+kP6eoDYsPbEWlvk5I5whG7w1eSigt5VKPYFx8hFTkua8Gx0UoJ5aT1tXj5+V/K99DUq6Amj
hiKo6i9J0/L5by9m1CvvCeCtUtZfZ2FLV+KeVfuLkadFy4pHT4l4Yo1W0q4K84iJ/QxwRfaEJKjS
chgNqNEGhQFps98ygYgssJIkCDpOv/yXENHoLZBBeUw2ybmW7+oSSakKZ8LfAz4S8zFZCVurchGK
DyidtUwLYHb8SiAJbXUzUBt+BaofIEAInktXbnOrKJqj8DbJgWjT3NbTsilZw0kXXJH2Fw30jXBN
HP2Oi6Zg8KujEr0kL4B5DlxRJQI0WLA340j7rO7h1gVsUMw7D5zLIo+bVZNDrA8u+hm7QuwEOx5X
CoFWRN7QxaqMgc3LLpCn37vIJVErd4chhORDPMsmc/R3V8vRfcAtUAERZwp0nCZ4YUFslW4AXiZ8
xgeEnlLiuCo8ZnY27XshGUqPJ79nr+lDy150wK6r1yqBY5RuUxQ/CpycAWEtngHE3+iU+o52i10J
l6fRB19jLaz/B4zeqye+dgLc6wvIZjFY/5Ws03701tFGnKUChNIlA5XTaFQiNAhuYSuQv9tSsT+r
t8zq42uLJFVkV9pu84vY5UTte+xmIERxoj23RFlPMgWhIeeQ2rLOJ+cfZb27NtYTm0FJCwcnUUdB
jcnHHhKBz1M/9RbRdO/2LZXTIs1IXZZUMbZ16vaUw4Y1UndnOU/0Fj0k3AKfnDifojD8PsaehO2k
mw4vax2hIImEw+0Z/d4ApJBt1rOE2nYXm+J7Its3gTyYn96DAucg/UMo80s393AVQXArTJ0ajPLI
ArdqqAsII5E8IVJiM8sHPlPg5IwbrcF4yWYLyYWzxSXAFTrTdR3+dtigwKkxUJr8UAFqVR+2p4Wr
a3YqPpfNe7gne0dZ2rHM4N4zrUaVVf0JOtjoFjybBhydpjkWNdCO9UbVImBLvu8PIz96otI47UD4
XMDUuzDQKWB6y69Z/cOnwBJtThdtGLr7lRYkQKK+MtG/ShejbnJrHUL/AJKBNHEKbWr2xZ7XMKv+
uFTBvIRSDcx21oMFJgliKs8ZmtI0iWc0B4uh+oftGD6Krw5XvgLFrJAR5UmD0W+TvBlWifPRvRBu
F/6PmDfCP6kmHs811FCWbyAl1OnuRRp09o67snJKRy2PaYXUP077wXUZI1Nmq1y7PFOukv86Yc6U
c2JBw5PKG/v2kcfrUnZmAAXbPs5YTs8sYkMSCRtOlyhY6rQAlvtAAlDxLoyn+cxZdeMpSiZsyL2u
wTGtdcA4u73eyIRqODqo3wTi4LT9zpTsd2EwH8JWEM9f5c87a8/QKk4BzSUgoB9tX/PwRuOTBzvE
gyWzZ0X1trvuttk4AbIQVCaKPWbly0t3p2YQHajn2YxRBHnHz4WxXSkd8puFmKuyFWLl8TSXR9xS
1usXtX3Y+kSVPpWJqKIvHrk3D8P6TUW8e1JlTU48YQttaK1C9nyHeVKYR1Omlzpi0azu87WfA/cE
7GCEfge9Y2A8HwtJiBvZEkX63F9wu4czETbhoFOrz+sn1GM0naSMFHhb/hkjTBrCzg5/uT4Hneda
EeRKWleHyyqUwDLgzfO2CRP7g0bdHlbthp4PCFU40OtpxDAnYb35E54FdOqFFOzPaUP4VT9IpgeE
32uN3rG9d2JH34tM+fyK2aec3TlBGdmBmRyANHu9JsuMFQKdk/0eW8hsVzbqdVEQy3wIh/zS9Mdr
BzJU+E0IsMS4VNZmpsITJ4yrE1pwRXg644ZtoQJrCxivUppS0x98tSOQmYiBFcLw07JBPuQuaD6r
siqM2Pbc3w4tbEps4aesSyXtBmsjmeIvdfc2S6MuhRe6ZrCMFxA+FYgj+iVYyDWUS+Kr+xhkfjrE
H7ry2rqnkQIMZUVOsOZr/msE8e2yvzvY+bNgAtpBZ5KegOcxsHqizatZGfyiqygoic3deyzwVPl4
6gqKIQcTNjAPj9WlQX/tUwieYt1hkoPGXeoyt5qAC+xuBpUuwH4C+Q3RSpnxxHFFIy+6ArblyClQ
/K8V+afERPZJ0c0uWT/7nMnFGXylRYAMHT/zHCB9TOKnbjqrO7mOk3aFIrEAk8etnbp7to1JqgdU
KIrJweBB2EF4WWVi+5Qi3IUUIY96fV7WNyE7RGDTHK77gFvMzIjPd5dr/PtVdcUT5IQC8tb0l82P
4LXVhYADvdY4XQ6/CtutmkqPvmY4kpXuWmd4RkrrQUggzKT2M5f9eGW8CddEb+6vPqBvpQkg8qPb
PExZRvs5n8Baj+aqdeyvhsMAlCSVP3l3eB+7JIT0wUrrZzkW6cBtsmwPxaL/ftET4CDfd6NtiucK
v3ZNFtRxm3uQccvYwxTc6RwbAgqlP9KtowtKKAudd4CJqg1Xop+YPLYDkvAIOdUdbkRd/XWUF+9U
6NlDCUQrqSuOb1kr2Z4jCBxAP7MOf22HxihV1JA2DEEEHjCKbpGrN0P2YGtz02pNkGD9rHumSDbn
+EStYg7rr7lldnlH/cvLpvalFwiEtvgSzNQdGtzIlTGhCQML0Xjf+Y7klmjv6C5B51YGo7xu0SAU
lIfEOfxAIV/5DoTzK4niHr62ON3gOEom6Nn3lURk0MUwJkOXRQ0oAiPqBFsLpsHMPBs3fAwO21S0
wux0LzuRWib2wLh02TiNpRV0FKDdJJL2oYxlMg7GLDPA2BrGsVieXVlRY7JAK5TSCWriAAzhrrJV
IJCPcJYSLtdKkPjwBKmPk9thGarrWNCR0ie7EJB+1vcKDKvCp5xhd9tcbciUZ8bJ0brgQCWfVWeK
oUAj4Q3qfQ/Wbcjd/9Glf2UQ2Hlh33Lbg0Zt0yqG2CSEmPiDz+u9a9aZjIKNVhC6y9STN9NgHoq/
K8Y03KxgzkF6zbdttqS7bsiI7qI9iKHWwYO4dFhx/cFsmSRTGzPCX9EEDJ88AbMnmQ6HO9LApXfn
eR900csaHfVQAnFd8QRCg/Qbun2jMmCv6q9PB6cvIiPCu0uaE2UbaOcDMABO2nrxEuQbysPKbCQD
vEWfYLTx6f2ejglM4F+k3DS7EYHMOgyO7LVLvaUQMhg5yftUZKdKHv8K+FCYEahkCPQj1ISmRHuN
aah8QJXFCoVKsdATCiRlhUQQtTXkxPMsW8TG8VZhfiLy0WJwAZV1KoIR2drmkwkCrtp2FUf6fra+
+MQMkJFoO11Zobammx6HhMBBFNcexqk06l1rY+mBiaXoynSAtoihCxyAIazLJog5dwStnqZsibv/
quIYGrNzIdugMyktH49/HVBMoc+L/lH6gHY3wFC+b52e7qwHLoRXtMF/OzbthQxdg8AgOTNlNJZa
uo0lXZBpWu8vKt510rLvzZHdzaKs7oFgNufqlC7p+iZbOwYsYKJVja7WqLeTi1o3dHp3u0nV76y8
mUfnKjMWaLKkEcNLaqWKJU7yWtXZ9GwQh9FWyEPGKDd5xk5ApHx7eutJcqoksLJqRUQ5Aaahv8hr
gegrptGqVwiaBKCVGejBi5U7MQzQ+GMLov3rDuD+6ThLnUmwbRwHj2sADPLiF0cV/C33yuG3GUG4
rMr7pqtC3mISKZYUnp2W4kgUE2KMKYAgjO0trBHIX36Kl3VbORZiI9X0ML7tfqxI4HE1wCtRJAVa
HV7TThqWeBlKNV3izUycPsnY9M/JG4jD4Cucwx4+nCFIgftVQF/WOcWcuPC+nzONA/ZSkQ+0MNXn
d2aHOk1X/vonmsu4kE96XZa/CgEmxM1TojWNBNql0CV5/S7QqwtM/Z7+9CP5JF8o5KUur9hBaMCH
j8s34wgJ9GeMrxj2LNUnC+VymeUY879xOI3VW2zanko0YDjuUv75xs+SjlK3C86N18bTEh85zN/q
d/2+OTahEbb3fXQpAYJ7EjEpMActADdjbpalS9mJMQBrplUZ1qmBLXi0yzgdCBdWSgIpASOjFspq
Yx1051aQ+ATwYKxUoNcpNeRj4J6gAQTBrZ7u0ztEaIE7c04Ctof1VJSQmEraR0QKDKZx5dmwUNH9
LJBL3Nr+aGivBJCnK4k2OjrHgRrrJdlbHKv6EXtOw1auNjpECt7uQomHnIACmFNEgtHCIZ/m5dWc
MVEfnrTAYoFubkot/b7TIpOIFWT2RG65jWsoYl9iiz/0wsKHzQZCOoHX0iNTshm/V2OD8148CjHa
upxtAJ+0xTAZk8qQ7conLARr0j6aGFVmGcelE8JItyZFiSFGJ0TtBD/05K20nemgoXgoGHIzDrAh
GMD/Digr5Yjqzgc8tK4Kp9ns+kYtVTrmsrJfELlb0m3Evyng8p2V9G7QIBWyszvIdLUO4QAYXF00
6dEOWJsx822gvOQfH4taCzCZRXTm2TSIKUyFKlBEehITY3RQw/Jg4Uu15sq3Aosp3Oc1ooPxt4pn
okwI283Rk5OxqMILLhbUqJB0q4dn1ZZCOfoL1WcTEXS5rTWLs8QsvpK2c2wTEWY6gs/L7tpgLzbb
PnKRHBmGIQStaJIdMDPmmGTeTvbsGbPakYsId0MEQhaLmg2ajn0M0uT8Fb19pmBfcj2o9DQWwDH4
xBGHBugoHv+40Tw1oqOu16+r4xB+ofaginu0aULVwnre/xMMDPUqHyNZuF2olQmVnnouZCn5Vcqu
XawY7AyQhUF8N+lyapLsc3hTJPo0GSxYQe99zXMFg+1fIq2pCSMnD4T2KfuzuubEiD0xxEO0qxyn
9iPFTDbKGbGydXpMhagUzIk0FB9PtB84EtjYEpPUY76tUvdol5ToVtux3m2xNmqiurrcfDpGLC3J
DBsogqjBGRCdW8N1+P9EXqv3E39QKq4vnz1Bi+DWWzml5gMnjg2WGKTxKxBP6CMDj3prc1dysaZn
suCuVaX9eSaUs/HqO3q8R+CaN9SOCa0pW+4zpcrcaOD5iDF9cvJrTIanvIkBWRnwPLSu/5IdKsMl
3N6xfsDl/F7B8poiu/NSBy1IzlgNuiUkES767zTgG1JOF5UI6XFB/+k1Olj6We2e9mWh89NyMuoj
k1vtNwwq8DjsMj0/oiSuHtUKzLMu9tlG6YyVTxkzA85nbupABModqzAeEFw/BwLcwOpThCkikhLT
nUd0gX+1Ge0ULEcjiawIG5klHfIA+rPPHJS+pfzc0HfN2uTgkiZ7H/g5CryF8p+6Vpo7EUNlRUgZ
loVvSU0dg2eyawcJo2S/HD4NKfZEi714v3AXtiDF0rXylG1xIZmgQlbH2LBB5Isd9N3BmRNn1gb7
JBiIqZX4GObEn9Uo02DhgbN8Apxfdj86/dvurfer7rBSemLni1Xye1cK9FbyoHLnnW3OteNM4AqZ
rvBu9s5GRw/JHDUUYbBNGnNPqfL3ASXfUUQ8vHXC8RNGxQNvD8nuijZDFsKiK0CHsTgc2uJyNWO+
vz+6HfrIrsxpARwnw8hzSO4IT/x/lAv+ZCe7EGr63IjRl1WIzcVhvvwp4HNX101/KL/F8V6j8uTS
HmgyBERySZKwQHG9LKl7JjbDXoW3SIVYJFg3NQveqyBm3bHokt+8k1PeFVWWKctezX4kvr13rtvq
0iI5mbGhvnsvSggNvu2xT8gCesGF1r+CJkT47tszAS3eN4aF4Au5XB8Ml3skizjWmsxPbIeRbxdB
8OiDMFV+LCvNlli4uAY/caM7XEXYtYpl03yLtiT4aVh9HtqBcICcCRFu3YON6Xy6ADwrySmX7PLJ
ZH04j32pjB1xNivR2IbX8PTYdS/AYyyfns/C/us5nf+xCbz5uijuGh5FdP98GO+MsbGcHV5yl52f
+aoZCi5J0vTOO22jFVLTQMVHuWp8eZlF8wNhFOu6//Hk1jaN5K8GkeM9lmKMdMg7T1VS44K8ct1r
FPu1FMttCejlO4/ekf45Cho9bUEAcUkbMw+z8ENYGvTVp+rTJJTS2wuyr6D3iNszsskgx19fYmdt
WsWt1Xtlktf5eFnl6wdqrLKxx1/3DvNgc8OKAfxGlKb6qoHtm+YEmz6wcOrpAZVXOUrONC3czIQ2
VGeyRdtoReKB13VhK3Y2nfgPPWEz3dIRLV9mlDQNElCQIRiJ/UJHQ9wu9MQexDTJ05q6+u+VWPhP
tCSGmaBT/2aBcpnNjGA58p36xbAT6baJmXZ1y/9AJaOMw3g9HcxpsgGkJ8NxTe92Oi3gOOF/puxh
uzhkhjbn1BThabpLWnxObcJu+JgjPvIbPIZjJy/EehU0RlzWxXyMw5AosnT7zHh+vqd314Yd2XSl
ZxP2lu7JRDOhojETjXbiHtua85N5O2rHZdkBXlGOxvPhb4+x9RTWIxjKDSz/RetSCn3eIV+ieJwt
ncVFjRPKdpH3c38CHn87ysGutaqREaaopFW/0//7IweS2jsA0bMSVLMgZEv01KkjVg1dVkOELkRh
EnJ6y7W9pmW4j4fVbFNGaNqDHqIPqZWtiRY7wJFqtxsHuq459YrjC70tEhAMDeklXQ3C3AVkrT/z
3CRjpec5K2iGism9KNpLf1aMA/JDyQD9Z5zKczJ49lCpitV2nQXacenNM1OleguHoF2uaFYeYXF3
UhT13LSBJ/Q765XisflQAc49DwcISxMtgwEx9pw4oFKkV0Y3TUAmaPcsQFI3vugybNudEo53zT1S
XXqphrQEA7KCj2tkQYfF2XOCwgub/5vDGfAAzltuQG4inGlqt7fLdqDuVedw4FiFkdVS4Qchpk0Z
iB9A8dUnuEUkMZ3xv7e5oZs1bjuPjzXlBsbpU6QG0WA92XhLf4GxtjUk0Qy9YpVPEKvHQJ6WdXJ7
IoEaR4DzyLvFLWaJ+xkSoVLDczBPt9Y1ISCkkg0oo0zxJNN/nDzluZTJLJbqqImZQpKqLrQrb+mW
BB7S91pT99xTc2CWtFfpdKnncsSgNFWpRC2yk1Fyn9zAcVr4x/T8eLwjo5AZ1K2YtwAK6rcdHCEx
+Kpd+Wi3qnz3Oa0sxwYnt5E7nzyBTt/QiwmF3DH8ce1Y2gZ3pRm2MypgyOZwyVhvXAQVpRCzDtfC
qTYqxbs6eTB+PloBC0MU+bT/YR3c8pbzPbQwf+KDRaiRkQtEEnyqwIvRgJRNXzuxrLJNORJWNwvu
eZGPhlATuT+HRlp7kvgHKO185vE8D+I574Yeszqa8bpL36Nezr6CrOCPEiCm170D4EcHQdw4MGDK
yEdKpqfeaU2FLs0ZU334GznGg7Yi8HtxcGo7VBYC8uDOvpkRz6SWk5geCnpRvxCTwX3OocWSD676
CbnaxHBVPHcQFgxk2pt7fGuyU1+RifYtI4RfyOAkfMs+8Cj+n8cMNYPLMmcPqR/OCk2ddeqlxPW3
Ql9t6DqAKEXz4z2hhwcyxa9quZGlf+k+RjyC5fmG56yFJS7iPNmswfYHvJAAX+rTc/D0n0L5kN5Z
TKgDB6G0puTXTAkanG3b16r4aMJIX0t99lMUeYFUt6uNgwSzg6AB7mi2QYHVWQN0F/FloQVloNMm
uydJ4WBnp2PYnqVEaJjNd7BgnnDiSUUHaf2TRqrM32moiMAVr9rOUvSyIyIVJcU/wXrqaQXHYjkT
A1y4nO0rIThYewusOKkVMxJjRHVBH1BEglYC6ASU9eg0YZP6hyammUOsYS6d0p+xru7gtj++3wfW
v1C4OwyQuxsCmRiIHADeje+R+kQci4+LjevpfMkdYj10KbIFzE6WQoGUugJ1s5cBcbPOQQ8twvcF
U2CMUUP3K7SAZ8RBKmr2574XlSLJsqApQObmjYiLWRHUPB4NWwoumyjiJlZawvtZ5Thiiajdc0F/
Nm0U7Rsso0/qgbD/EtD20pRw1BaWdCDIOaszwsFhjx16xcC7FnrzuWdcAWvWe6xQcx9vGS+OPaIh
jpjYPzXtWtB1zMeqN6hP10J3ph45jXchwPw1fbwGohiUi8JKTddSTEdg40iGRnVcCf9khqZg7HgL
/h7TrmmivLNZ5er057nfnIw0G/kDZ0Qyi0i8csWapwH2kUeoHLgyqaeTJZHK+W/i7IyRpcFyNq/R
LFJqUv4Y7CPxXYBqCrRBNtYmMOJ29lBQZFup4kvjjKEnd8NgQZobDhQdsEIrlebmUxNCSkNDbW16
bTLC0BLPjp/0GWLCvMJAp7mabsszXnnNOAKma9NwXcuDhUdfyxrwak13KGalIjUCcHAD5KFUeeed
QNPYfFz+xPjfKXYAvGRdlvyePSu5MzS8Cai475WslJX9Lrgm+Hk+Op9PPLAuiIcprwoeVdd6mG07
b2YRDVpVJNV5FLSg9G0hXQuhnnazHUDVMO+/1LFLQqYK6xcVOLrGO9RWItNcGIz3SQ8ROzn9G2uS
Lt07WXbJ8QIj4Lct3Ya1OFpDjiXR//ZrEobehTSacq+QKm2yc4lL33zkNZWhM5TcQqPfqvdY4IhH
TZSd+HeZV3oADa0uaSHd9KS8f5KqhRBs+pxP+/cogudZb5lw58+t4eib68UCZ8ElzM7Gibg2PJgy
Rv8qa3LpasqczkPRuuGHWDSHyJOIdd/4LK53h30/Norw5gRmY00mlG2j30IQTDQZORvIjH21S88/
E3FfwoW0EooxEUfgx//Ujb+CZMyqPxzOSO7y/DscfdYp2PFWVok3a+AXFisc53pe5kqF7nhjDpYn
mWSIHWZi190fQcSa8wA8vb6Liz78Bjmk5M/tpBPVmcOAXE/3wojXA0D3aFnmJIHKJJz/3njr3V57
jFbBXm4j6y2HQ6bweyARNDmpUpeJN8AvlTNkuxNY3k/t+OIkqi+A7olFJgfnbtX7MCTZJNkJ39EE
H5vvCX+pscMcHd91ST6nDglgkZ2rqmte1xAmFKphCwfjTgeeWKaHfaovYcjDPirCYjheFNbKc/5T
3CBOzTxztQJPhnmhPoC6yWtjKTuxFA7PJmRt0rr8jmqhnDe0YOsqzAY49FMeen3gFc0R0zRMRzC3
Ka7beznxp+NSlAhpIL9dfRBOBzIrpqWH1qEA82Ic3keJpCt3PAWYHVMSQt3qOCqw92YrxnfWvNvA
t85nO0TWL5v+T0KoV1GDKfALRGGFKgSsyoyvPqQQ0iFF6GF1AJRWssxZ8LNG5UXctcqEPcHLRMiE
TKAb4lOYtMIW91mRV8Rva7LLnn35EuDMwmfwb/IRHUCOuPhSUMO2AMfRA5x9nIwhZSAPIHw/HKvm
cQQXfJMexcfFTx6cRWcQdD0d3zhm4zTDXkHA3fCT3tf2K/8X0TlAhCQFoWes7L4d17zYA3L9SvaX
80TRpUQDDXFsBRLTVE42MJ3sjUdslt8vZ2dfCQ/o/6sC7hzV7YelBxJ7o60CO3wvDDg7yXZu4te7
ut+xRbrWTshmIzbS0CyRAD/x9saNaviRKAGcgRZ/kdHcaDZ2aglDHqGtmHRwamON7QeVhueoPOi5
lwtSeIUM0cL9n0ZJIul4c8IvxkG0GRdxlzPsMJGsatlkQgCRXL3hTPIEAGH2DeP6nY0q5auVwzzI
d1Z5D3uEqgKjmpF6m5oLSPB49qeTPDfxaNolQHyi8QGgOBP4CH8QkJjDjczQoEG9lpjMgg5aE7Yt
FWxnQL2Yqh1EqYxv2fMdCP0AcslmXZR+/yUz1ap9k3vp4oKp7s7Q1nFamBufwMlEvT6yFpdhAn1u
UupImqxIzBL7cVxn0gkGCYYZ6qFMnkCAcKT9razav9LNezfgx1fuvxf8Z5dNMR4WT5yuNnNvj/wt
cLk/N8MOU7cw469U3kNvhbzaVgm0SQPkteeEhCiC690P1r6S6Xo/0vInshuvo87frHrDvc95XD3g
Q4V+dthLzU6UElScX2uR+aav0LWumNt0S4yjaBmUkNDw0Sq5okrGLwsW5a8lf3W9IZEMmLBBZllP
GEC6JReW7XPd3Igfwt9tmFXMZJu+jrGseGXH2CMALhq+VriD+m7yYw1VbbIpiH8QSC1K0Mngp4Gz
pbim5igkToidNeJyCsa2GhUovTbRtmsan784DGodviOWZAs83HworylvSOtcZw62UTb1l4mBini8
IFBz0CrNbDTb7Q023TcCMslHOlL9Lyy7Fy4E9M9hHEXETzd5dr7WHbk/KaI0I99Fi/rnrV1DHIen
ZKOqAK4guTpkdUbH2g3l6/t5dhJGuZdqMpPoEpZg+KlgCpkFt0HcAwIQfcNYZuXpqCHDJdues7w7
jz79nXtR4T8LaNXcen2qrU8B4gKl8SesFL6o2TW+ePZyuAnTLcM/dWG2IEpU/UPZk454Aesb4TWR
n9CQnK5z/ZZ3xq4YDm6B1p7szTnmIgewq7HLf0i1PO1hJPGskvVIA3N78x5szBmjGZ7XKsTfMNVi
r11WN3Zz6Gx64Vzzgyi4STUBfQqS3kW4ndelnQUoUw5UgEKU0VusZzBCuCDbfabmtq6alVigKC19
sJbICVzLw07oUhZ42iqazAunOZ/d3p6ahVYTQmr0lQMBCPV6fwhwweiFJJgchJ7+JUipJePLVlf4
De7x50LFeQK410STZd2LdrBdRCXL+TCu3cDFI+ZNEjvEg0aeLwZGuD8tqPgJJj4nor2PXtc+0875
ZqtL1b94FROUDAPbR1VjzrdsBUfDMc9N8VB9Hfn2+L+8jFgmj7Pw8PowCGGg9xtqSZRVBDmUmWKR
08kGj34QWP8Ew4jCDKWuJK2Bvw5xMDm7IxrZUlA0h/rCWG1s1yC5etikja1/GpbaiLoiCq1mnrGF
6G7L9KUPoiTS38Ft2WlMxDjUXAyTIWbm33eITqPBFFsMLxA2+5djW2KcC19o69PxobbmL7qbi8x0
wYurrKFcr1sbkkTePRxi1oWLPvBxENkOIUoyV2VqsG6nToDFuPWhsJHTxQoCPIEu7NbzMal1gjbK
B5EIQ9H934rZxqv7Y7wYYmp/FUgPp0gVFgp4xnTaCtQqK742sCL6gKHTiAzZrUVz5mc7rwTZZk+L
EcpepzoM04VnkwW5jpBktVB39zfBUOjN6h+kOy4anpEvQX5omdhwfuahSh52RmxUu6C79Mw6PjzY
XyzAC8ekocTw+q9GImi4mycwlhhQ0g043C9dJJ+N25hmhZV8wBdr1LGvY1SCH/OmMimxAFrKgCnH
Ipdw3Ms6TxCecRlbEj6d9NzeH8UKbaIz8Dmo4gXoS1/UfW+v6yafzUbUdFJy6AmeO9CvP0ewD8Ts
ncyj4amNFwpTUQhTiEILWoClF5Lf2hS+FknDjkug+nWiLZX64zSlT7q2I9vAXzTqivweYFRZ7fkr
kICJs/bIuPIhW4rJZVz725SDxY37jeVDe7ZaCtfiJQU4IrEe6H0kJEubXHDPXhzi2c/b8PDDz/4R
BIEULXSJWDz7+DkUEMq5GulDN2aShGZGgAdNhEZpzAuGytp5IKuqQq2xNGeAvOKANwswJr9c4wvc
Ah4ryh5Tv8Fw4v3JuX/7/g5jQDvtiIDYKNGr25nZMhX5RHD7RcAZsuKWZ9MfpjFd5MgmQVJzahL2
WqgvJ6D3kb9RS8BWS5hgvY7C+Kh03uoxS305f2olC4BHDqRjAip+UzlrAt5hCTrWacJAKrLgSGLm
vqf2DjbTQzRXRst25ewbgEFmS4cPEtUyj+G/eUuZ1VzcdXsNuO2v5gb2A9NHukWWPF8DLVQFWNcm
rlwZ9ZrHUBHxMQ2Jf92gBhT/Q4mkDhi8sngfmKIn/Yo47OzH7wnNyee0i/usOkbhs2DD7Za7b6xU
0w5Xme6yTk+2jeLA55dZP8CYG6l15Qo8v1RW8aJLJVCaveOIxNtYgfm9PkQPH+9F6ZBUSumU8Xhn
+tq1CbpLbFzhqbf52EmdkteB4on17R105/aa7ESUqyWwjhGODBvJUGpu598mDL29zGpUaKjmIjc9
W+zML/0M5CI1z3/FFwlJa1c7CuUlmpacjwgRzobj36Owv/jT8/mcypZNba790F1Qc96HX8/u7piT
hUZ9BP3giJdgXQLgro9bO8BzOZTSBSq6p+BvaZlLwOr350vJxAe7bPlIV10//L9a7bOcwa0usEe4
0LyBnKFzBwGP5cfdKMugucGl41Jg6geQPhwYY632b/eE44gpHua/9/w07zUPPengiV56wjGIfyZG
n9xhmgSP7yIOQGWe2npx7VgNyLMnpRb2L5ACwJwiYAQ2G6n2lVqbcxxKXf8Vy7zwM1zUOTiyBc5o
3gY8nBvg6S5OKClAqz/ryQZgMnYhFdPBPIkdR5Wk4tnlhbvZiS0rz7xzFNhhugOBxQjB4BIJC1Qt
5gJJDeJyclTXnfRZ+kESrbxG/1pq4qvIwy1fTwoC9Ijd+PmbxR041zQGN6giaqmnq1GqjJPHu/dD
lD3B8W2kjTUfbWgTDx7j/auIp7z3zyCgkl01r9xIeJ6WnGrCdXnhMFQBa2DhhmH2z9kHF/TGqINq
U7jCFQhcmDE5jJF+Gw+KPeFVE+uuguewHfbnSwK8PG8AUpRkizBSp4cVEgcWpTcWinnrgjriM7RN
Nc3+6WEUgL6OeOIs9SoRW8yafY9EgXihD2ncKEZKo9XlWh2F9RcNAm3vXPpH6aKhYH/9LuhZQBux
LLTEbu3GgrZIJjTl3lyJh4M2JdHEocwCT4Y1r/l6yIsflMYwqbPYjIpEVStM9RUEw7eRmz32P4aN
yhGeustneMk874H/4wL6VZipXnHMN2uZLnOFfG3t0Rghn3hFWxGylfXn3GgSBHpqiWAA/OUNkyjL
UEpl4PYad+1h8ZKBfT8WkIz7dVUC+Z1l35ch18RtLAc2LnB/TcUKpMjEyin0AIqnNDgS626ws7yS
ihiwmlTHiBoWIQZmSO8JMOgAAHGpm82nGyiPsaW8P5fGpHqc5QvKwPiXiBF0Aln/5fRwqK7H3ZA1
4WUQvxQmo/hylz5qv7WBpuGK1zdMY8qIp9InwtkFi7sgeKUg/XqepoNSTPGDg2AcZrMd+HPqGn95
Azuh4Ei39aD1A+ggUpi8d1RBnpNPK+Y0I/xzjvCB4j12VJtuQJm5Me6P6HyiAoW/gsXAkicSmDDC
Wp9rNx45B0mcYERXfMEwnhWgoresYCPQc4FtqsH6iLDHBbDlMrUFjUn9vYoJru+dnrrmrqyudkAj
C1xK46OtUdq8SFwLSfpaVgcIpNIfiE8kzaCjLDqoCpAu/ftd/mnrhP70sDyGerSjnHVYDrrscP0U
XV67Ef5NJ/H/r5swsMRO5KUguFWnA8OL7+ihufhU3zCNtZcf95ip7+S9CQPpIowsXRmrnw0hva8m
kEmHnOzeorh9flGGbOH8bRTP73FUTeHSjaNOCufY80hzzmYk6E0MWCMT7BLvzT1m1JrCsOHkEHYA
JbQ8bL62d3SWs4r1+GfvkaOnb0fIggZgfE3NTsbigwrVgV+KNDhCuAShfEcbjdWqCVSVX7Eh4UsY
HuYjU4Xas+edrHbh15DcqOuC44HwP6qVqsNhYvYcGlNCzjqxkfg9322M3k2YolBak5jLMF/Py0Vw
WfliJxboqQ+bsRvAVsvffNyzzHpjXa3i6tovUXRvv/rjzkX5J3ApVJonc5aEmhSYYAhRnPfpHr1z
lfFL++lJqL/88o+gTjWsHpb46uN1/w5ol7yWQ4dlCopNyMteoUbs1DC5AC77lAwjOf12k9lfWHOC
bA+vj+aMaSbbG7TpAMsboV3poSLAMjy79WVTLd9DAs3/T/YiCdaXBd631bYW85fyHElggpMZhxxk
F2JwxwDdOMAqiHa0In9PPQPUHD9le+s4lVIT0qZi3AxULFIzqy0m22xFuw0iW1snSXaRsqWZgSsL
qY6R0Wph+vWjd415X+4dAv/3H41kwQ08Q8VfvfgK7bBf4vJafAmG4vVwaPRgHcg3oay12bU+KBrY
b9cTkZZW3LJlHTybbJg2n9arrVy0sZe5wnUYJXSxr/NRcV1D9UaeRtyNA8ppJR6zbODrJjrp5PPO
6vEJ7ky4syaCUt/DxfA4Onea2cfDZfIT0Zglm30ZJrX0z/jqRHkOxIbh/JW4tKnRsVyOIgl1muUp
twIq0YplngBjc+Ho/e2HUQYYPONR/qfg2fd12uSwuKWEs+REUn326iOaCBrWJsHteprcPzitXD8N
W4X82dAo6FneolVhFDBjI5wKoJcA83T7JINUif015YU2FkO35ljTw+Qv2qErDFbAHH3vB4yBI6dX
0clFf9/9YijFahqFwot8yKrHYfoClqfaTTFD5CeYSumtYLbHQpKKOBHn/407VWDVgCJPKkhIqTFC
0IcQh3QwUEY9PGluNdMj/vruP75FlBgS+eOlnlt7N0c0V+MM2UtSaZ6b75eSBr39qmM72Bh+PYvm
JXFO5ZYzL9FY2k8KdQFSbxfLT9L7g1Vd6pkfu1IHIgVdGTwo5Fs4PMTWYWDs+NaP8wuBZITdn/Tl
XtmxiPc+Xwf52ByyYBCd0mJuO5corBlFgx4KHyMtLEMG86ZV8eBcUf2cusN8zxXE1S1zOSJi7zL8
bql/sKWyd4vgf/lBBvjyN+RSxll1sZP499UxNvonydvU2eKTMtWMt9KofbWYD7pqb8+55LzujvQ2
W4r2VK8s1WFKK5c2PZD5BRed2Nx2rtM42mbOffN40wg108MKVBippXxurSoQ1wTpqTUkGT5RTq5v
EKjglR3KNpFspX3yAGuaxIIX2iua4ploC/kLVN7iOstSUai6tWuGWSPKU+K+ZktBOJ8l5a3OMkzg
kV/Cb4rioM4PDWBbhrIpyL3ljczmQMPoc2j11oTqTYrkfcGlQZ4tRSDKMQgzg5jLD2IOODP40c1l
+ZSp4LCtq/l4LWFa+YOdCyKPyhkVSOJAYS1/aNr7qwb7V3VFMoqVTuMIhHthcnbryoQAT6PRK+lq
N8KCaU1v7GFZHBTl+wv3khlCVwMF7V8A8/ttCBQaImr3XKix/7tKTwhxcS9+LyJE2FFZ3JfzXWWV
gy+z3MQFoIS33LTrET92k2ZbIJWTfosmS54i1kAOq79kYS4yoq4i1OFNt4tQT6yH+A6KhUpsUZae
hL1/2qtveE6cLheh+S1PVMDXaXpy0JzN+d181d/b5NdLVQ68eOv76r+XSAcgyx8/91uX4yKLfTXI
M0ZY2a+3WDPF7FFVZ/Z7nhHeD4+mGjEOMVwjcFGM2pZ+xtbOqWqAoUK/1s9Bu/5AGL1B0lCEMOxl
Pkrh+Rof8lWmlWjbfasTE7Hcihcd8LUj02zsmbp6mFg1nti8KtPKtQMKxS9BOagiEp6SzpEtasIU
O5QeW8nRyIoIJ7E8Zqmy3mxR55c91OMV3+ya0/K2ykeJ3EHC7pjl2AM3G1nATZoKlXfKBSdjwDYf
mFSVKufpjwm70KJ8s8lsXYVZ/Zkw68KA1QapVd2ucDfhekVzEfdORUpJ2p3T3+d4yT25qOycJje1
Ovh7lYJEfjK/Aiu9dhW2w/xJBPhtUVQUhjQzJ0o/y5+eVhGBem9KPjyDSt9bbT9IpljzBCYYfdAB
Hk4bz0B/qE8uHQrLu4SmGMQAMfvri3F88cqsQPLwnt2Hg80iTAZdmPX1AtIVyFIJ9SNnvv6v/z+p
unajNS1IDAzh1+UYY4yJvRMYaQJWNkbMSEMqHFurMnz0EKU1zhISlD1F+D5fUvtVUDg+dwUBs8dn
tQmvEMZ4isSVuk8RM2A71+HyBDk5MNAvgFpntcKTwSX3fzphqNvXlXjQ+mNNCQraoL2Z+N6cp5DO
tw4R7+eRYpl0A+TMgU/cf6ovGCXzaMU/tt1n8JRH2EMsmK83EVg5L/3A57WwcciQ80P4RfylSDjb
fiYr/YiW1xzTphcghMGmGMOYDOrmoklBo1+4v4PLZpWlTWD8tFAnnwLN6OvQXK1VVJoRJVddMoXe
qJcU3RiXBZvcY2WLPTY12BE1uwBW31jytynLVLSCnumV2uN+kVCGOPU6VmuSQ+FJycoi84jwIwG7
C6e4G+n1HR8Ut3cZz4VbDUqxaVSKrCu6tDXSxw0c5p8EFMg7Q6W0FlPzej89z4ftPCYRYOr8qC83
nEJigeCiTLkGshu5eHlBRlAd3nhjpdMqJ3/ImMhTADnSehEk8FhruVtGdEO4g8+2uopwuLJcql9s
CTuuvrMUvu6WBd9U99S/YaU7jEpWgecij9MdHe/8bDpWKrSaqI7CVkdWwMtIomDGVRCi6eWCH1IA
4dxzMmnVylsNNAjTum8RVcPnT5mWNAW2Mvj9oG76GXT4Jgg8RusMjOoCXGeR9ExEVDIlITRxXsA0
iZ+5i1Mj9VxiCP7sPoRas6N4eeHhZA+zB5rAPwFENBUpYQGctG6SYg45+8a4NDgvL4i+RsZgiwUa
tuKyUm4cZEQ6fB3wz503tvGxpWWQL6oEbfMh8Qi/ePnVn/t2KykUK1KfGzO3p7FNXXn6Oh3IUi5j
C8FPK4CZ62Ft/l0R0+HSoKbmaSM7IqR6UwNNGd5I066AVT1GsECFPUMLorVpRjnipxDRBa5EGs9C
KUmud5lSWRSJHC256Hdza/cCClXN6xQsfSu6ADWifropGkiUf4U3v3GujxH0gm9KORPw3BWvlF0w
T98FLLsnhn+hmYrBMsaneq+jVSSHyIwI6yvoC6r7+YBZ4FF0/azRhNjkqJL347nO9dK8auTOh2Fn
V6CpINprAnP87nV4xTYK2F0FQ8ghggZ2NJAKfeF+CJMuH4PxlbA6WP2Uv/mjg9uPagszkEDfcL0s
AHksRt+VdLD51uEh1GDODDoGa209MyLmyqIkuCph89tgJXiUetFi8FyASugIAkFN1CgCp4W7MtRl
yfzmFQfG7oz+3I4V3dui5I9afoA/jBdNdJ4hiidl28kBNtYl9zm6At+sJuEuBNPpvys8tBjWO2s5
ZunGxWcOe12ZJ7qeAKf+Ivb/y+Q+nDrgsZUb01sJ0JlrsDVHAcCVXLvd/jrZrYE/eU7Mk5yOyIJs
LBp6QibJn/jr8RcTA2e+r6pU+jLApoh+YSkdyKqr1SUo59i+egymPtdMsOvSunu9PcHHu4C3WM9l
o9yeTwYMEwHG/dyB5uqOqd5InObWOnmXt2Jn6U5UeiCL4iSqNE+ZYT3+rn4i67hu7UJjo+YA/hBY
E82GPDJAPRxR8p/xZ+Z7SpPR7ZB8RfHaUmEWUv2BG88ZfphspgfP31t7zCspuvBocyeWwv9+A3jq
OYGt79TU96CBQRTjGk3SqUxcAb4RiHkxSEspCuuLLcodkwy00wNFh7fF85EVvKWTBwe9rEJF7BsX
4hIL4ZkJaaaVmto0QJccaXFW40hSN/1n9KbbhZaI3wpIyzuF+uvH/R31RRfkYAPPw4YsGC7sBDoh
Y0HiNfy+4s4dYKIQRxTCFfVnooCaU1Q3PSXuAvt5bvV5v3Zdq9Nvr1XtWTlyxPa7EDAxJ2Toyag+
72ru24c+QoIgaCdxbNI6o/VsK/mWhL7AKJU14Brl2+P3UJyJ2RLIfI9MecDqRUW3P7FVvMZGJZOX
/1SH5wtUKHat/wfUQTZCQQ1hWjlNis+nxo4efbo+vtwyQFEG/yFKDp4VGOIquL7/GRGT26NO7Q2W
9mSTKSE/58bhc7zC4rEfv9ufF/D/QLsX6agWOEDGCz2NiZJgLBY/U9gz/mpklnQ3Vq/SijQqHqZX
xIXbDtKDKZNyXEqpZUoCEn6BwKGa18Nyd4t31DpmlgAV6dUMIuc8Yw2Sb/gcmMjXYzLAxoP6LfHh
2pQYexRmEElW0GFmVoHCek9J2GoS4s07o00nWGIZ2u24WU4WFoU06LMVf8y6R858/QFMFm1R46J5
MH5kmnyyRIYCP9/a0orZz0ueuMyNsP4t+d6el7+nzBfNlE7hJfz+XNjft73+pml/2R9TTr4I1FCE
x76BqyzjAxk2jdD6OZ3AbQJR2M55vzJ19vF7iFnQuiORhGn8f/q7h+daB892H7gQ5zJ1ZsNaMW4m
mYXJhAvKqtjbIBO1bpfMygJn71MnSMCWmQUXWIdLdavvjYeFbCi3dKhrTpQjZBvStiJ8Q4s2lDMO
5nxUhYUNKnmnVOfhAm8SaB3BiIOTschFnSn4204zrTrP06LuOjWLoCzGHPqOk7rzDs6EPfOtHaAF
9ehwQ9LHQ4qfjo7CHYF60JOUCf+Kmy8vVSv3ed5tRcTc2NSjCeuaNR55CqKEOtEhiAZwrN2b8u5b
tsoGzrjTedWtAjihwAKk6IsIZ20Br/bRlL1DsZ5icl1IMTM8QRvJQhmF3Hyz98oTz8T69EGoIGa1
M5DxY5Z+CgKtO0l2ze+qC00/oF7T0tR0frtMn2ko+xBCle4eGo6411zFW7efCkh8fldtWQ1+dIS8
jdHTJvTwB/tDVn49C1pXRx5Yyb9jnC2rHQJQTsewJObeOH26v8UMIQ0nufXqkwOBQi6ByS0mjDzj
QJ/Dhn2RPw5O7uHuzXlDWv7XRgN00yzboil2CE/iI0ihGRyqone6JCmdnwQsj052WGQE/jzuBbmd
WdjPmnQeJ8/PcAmtlbP4/85f93sDnYeTbewTpveRdZE3zldyQ0IgYCIMWHFPxDIpy2aesxpnRQL6
YWSC9qbg28tKr8zwstk35A2AjFCA39V5Gplm9On7eWyZGwhz2t2vuteVH2H5c4YB4Og0t9EzSPWN
2LFzG4cFguDBWgp5VXnNgrLS3vKPUNcgEA1kFB/2bS3PtpT6rDe14QIk5z5wuBLuUqsTFZVi5tnf
bePyt310D7cshzSQBtHJThFOjdAp1m/J0Qe1fjnZ6X32zHY5JBwp/aCitTDTkzD4ieiqtmSmNJtL
rkunlusjwlDgeGIs92XHlU9xisyEb00o/h2yq/uEdhKbcSRIFW06RO+qHkP9UGqQrR22bNgGQyVJ
WMV8h5AUaatPRzRKA1YyJ9CYYjIjhSIVwKePLnYUnvoV1vrNYm1NWlEmD2h2nMlVvYDG8oaaUqzX
DmKD/5NPS2xYyHNaYRhqWMlgR7JKunyNePylnrTX3Hh93vXYU4MQpiFRY/q2TfbupirYZ+sbBZbq
kpxz/K6O0cFpYihLDIAI1QCHkqwiTh8SemN3TMK05DKlQygu8bG152SSH8k3PLSVSiAyTJz2PFi6
+pN8yI8fzrzJkbamoiZ4zCsCnTjuYp80p0pHbwnZza9+KLiKOuRfERFQPBpfNcn1buEJz8BiEzh/
jo/jfuphpkcEGoobjEgOwjXHqeddh4nMNVXq6dSjOD2jPLBf/+igeP+/jpTsuA4ukaI1ersskY3l
87YwmEHCAjk8+sGlM+sQDxx7ZqAEvvxXChmKf6CcAY5STWRGJbZD28gwSJAlUPADKVMHyqpLrAc1
QS3UtI2rbnyfQk5GwSdL9OmsXYTLU2KfoCDddJ7nqziHQw==
`protect end_protected
