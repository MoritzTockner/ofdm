-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TjL8h6FWuYT6onKqZbKSgExJC+zaIQPLmPSuvIJQNEUX7ALlVDelBaQU6xH5y6wCp7/WPDwMQ/Ki
HIS6mdBVFVoPHug7vWHkjS5S3qUFpj2CocDIct3aSOQfd51wQCLrdtRl4FYEmxbsXoODRBszyegW
cvZHC9EhiDLz546uWVP72MTwZVlKQT/61KCrenD1n7o6rTb+pBwFd4xLF2/i7baJuTZeDMu2sCG5
MNkt5Hx0eoYUdR/fJq7LkWgsuPYXoMcVGbdIgi97Cucd2YWAaXPs9/Z2hAJ3G1d+8orntB2DzEn6
0x5P+uJAPi7Z7xouUyAP/T93vzGJSYl+biBpeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5744)
`protect data_block
szgOmJ3+/ZaFFKnTFH535ScWw7vD5cjp5Gv1s7jaCA8m4ERN93Y+wOL/fOUrEQWeQPsqwGA5xyMY
riFe7gt5awo7wLKGLBBGMBdbu45ScEVrqrzdpF+UratIJltO9soHgQlV7P08lTHqTrC83Jkt4s7M
yeqI7OaxAZSR+/Y8IzEZxtFrbt6sx98eCOMWYVCw3U8Kl8lyuY7jaUR/zvZRMTKMjUu7p5BwSmui
tHvzXnPQ5xXWfom8I3WJ3+4PcX0Y+gWWb3Mw+Y7xrCWv9QRl0KsQuyqEBQW+aeCJ2q/abmsvijaW
bjlbt91m2HBsOf7rmRIOg8uirwsEcWeHaUrfSN4B8GMb8BbgbY2mizqkrEklwXUW4sUwIh/Zs9XG
pxXOwcb1hC7c0q+65rZeAr69ORpSZuu+4+TTJSH6yet2pg+aNH/t8QVLyOHoH+TcwBqeiJbDY/Je
Uq/Um5SzKZWsZdSPyvuOB2SrCawdhUJccmYIaqBM16RGPmH8e4SpS6FMfoeVxCmk18wZXVG5fSpu
2mxWeuaGpnWB0bv22gtPj9EPZucK4PiYCKtSsmklSK2AP3lBERRxkj340ZT+Qg8Zi99gVvFnc14R
uv5JZG/zawp+VTj+9MgHq+/np2+ZFjSy1pj4lzMYNEG+nNy48D7GJJhRKyIfgcuV51oRkj6SjvCj
XNcI0US752H4MDhJ+sm+4SWXGo7HbwsJOzz/j77pP+e5ctNbU4VRT9h4Es2/R/Nsm+dA05msCKBq
z2OgBX3WNUAkg8f8IGRd2saoVfpanfRKMeMGazO/U7nduWw68jqzsBw0wqspxc73hhUDJtCzFSDK
5itF8IQnoMjmMuUX0n7UamO3Saqd4LMjj4fD5Z2WtyqsJlcxpcLvD+2jPnF1qf/O9sZyYgn9dXyq
r90LJkpR5wOi9hvNKPEqH/ztOpEVPymvp35hO/ttHqvFbC89NQDP+yCivlafrHUmtZ9GUtfWooOH
s+nrtYKaD5ayjI0mbb3U/6OhAB1KEaqHdqL0ROVbyfttPcPE8fTkyttg0hGgC3ggcTooFb9te9j0
kRCQkU25M8OaD7/+bK/3UWhqt8MUI7BG5S5UEHuJ9UpduyuhYo7zUNEI0/NjbmLqNvKbhNlFGMT7
oN1zXHfYWzzjOxJtY5jaz8vcEqDcR8HEWE6y6AmfInflVW3bV5kde/zhIIAF5v5J5lpgbjXhz5/0
ppRSkLpnZUpg9eWSTSBSSm+0hIy9QxMgYCYHPkkMl9IG5lF6qTg5RnawUHny6OCPrOQm9cTGuzyT
jl5+ma387VlHLYHVfehYv6afSDDvJXkpJC6yuABt43EGSmBAHqEIRAX10NTPLPTm7140PSFcTt10
uftEPELjS8SEC9bRBtesSMU+NV/NlTegJsn/FschfZfhpc2UObUN65UVaOqw+u7z/sXcMf1ivpvq
73ydw0KBMSoRS+V6kzXcLoF7FjCF7Jp2epzXdl0HpsrHz7G9Bjs37gvj6XWsA5dI43nAaWDnqgvB
d9yKrobfG4MOnMukDdDLfTVjGU+GWeXMDUDPPPrDUB2CZPkAbT0IIvN2dvgUT/qSe+gE2DLdM6Sv
7TZ0kM8rBqSiBQkS9CJybLjq/fxJfAiIoJw+b1qOrlOlYoMrtoiimaa0A2Tz9Zp5mnWfZsjyDyni
1XDpj7lu+nxmcNK0ClO7fYSR+APG+u12sWIegUvSWYEZDogMzCiu8N/mtFFqNgIf5wOhsnqQ2e8L
3+p+EDxGHfEFx3yQBoKaVMjPIdMh9Rf97Fm4xiUoBjemAr8C1SLHex5cknvcgW/VkpRkxrvoUqNs
q3Ol5XZSzTWUV8jnrjyMFkIZurrd9VPw+awL7GLA4fcCRIB1Uj8ruen+Eg+/VwKjxXFJN9FFpF2T
BW1AiygnHdlfQpYFFlww1/6NgJKMiSkJrDUU35dfPBEOdjDrQY4tOag1yiAFbO2Zq5Gd/vwp2AGL
rYniNld8CibrC9MVx33+C5SeesnbV58cU0vAtHEnh69M9D1JzuBVfEAhfESuALX/wArjG5tZ2LaJ
0mHYrHW24Yc1N9vDqWBdGDGzWdNJoNGMxEblMTGXghLpQ7W9TnA5qVJRbQkUJoqKzhjO6myhGCI5
jWsn+DgBhlT3sWCehPS8+w03QhHH+1Pfw9jnIQ+FmQB6+2bOVh2c/w/o3dHY5oz3/LQjvWWTklAT
272lN1PwYwmWH8XkTeaoMEZZtmra//LPWnh74e/bDjO3vw25hBwM3u/2tNWQNelaSYLxHq9PPAHP
+HiOw1GvEEVGz/BXVhU+I9G+DLpmSdAysHwjHF730gg2/GBXPtGmpuGQhnUWpjIcI1jQ24frZ3KX
Oro0HJxoe9iUwl3WB29vr/lcEkFaTFkWxazoABP8NYDXmqayUl+AEjyaRvwS1L17p54laxRge+6Z
fRyrOmRyNmNC9jphey+u8+kSZIehEYgQp4yQxkT9wgzlCMeMpCW2VeM5lQW8CFGGy9lYIqraxBLJ
Tsh1XkwvbdBw3xL/gcYtStsV+LX0OKc1yLW96Tu/alHXBl9fkKhDEgF7U06iMLEtLCyQJZHcHCUi
3uMaI6uW3ju5NyF88nuBTAmqYfWj83QnWD0YQo+Ll2CMqFZvitB79J3ZbKWRd+vxj3D5xJ1RbF2k
s2R8u2sMsUq03ht0t9+/NqQan0TCPVMiqSub4dV7+pzDLjiaFfZFpWKeBu1LSbpGqibUVALv04oo
eZPIs5vsTz+ZK/niTe5G7+0wuh1WMpriMFgKfdbpCJYsZE1rGsMwZHYD22vfZb1VIaDBYNVtERZk
lXlXduRygKO7iRJ1OgTJD2hv+oECZMS7JuyIXawelDHY5zDUplWmILB39nJQt2ENS75TEVpGSva2
CilITIobSgCXFaRVww1iyHKs09V1qZqLj4mbSvvOemuyQtmiNJtZKLbU4xqMPkWZsMpwuZZ6gH7Q
XZjykg7L+qfBBPi+vkt0vZL3TYrj++BP8n0CnJy3CFwABvQEypadUsUc9+LGym0bXRvXogYnhEB1
8MUQqhX6fevfE7SyJBoFzlP9FiEDSECXKr6zLvQ0I3gc09D3vzCnFero/n0CWomQE6zuEdclmOJo
qS9fx+2mniwtabkRxQcGYQCYnhOQNrOEzVcNwd7vqH+a93dtHLJSl/BcUhzpVhGI0wNBUgYv/GzI
c42phJxOa/qEB1aRyS+ECg0F0ChbOIjbJa45i/Cl/WF86pVV1pbVnLBXgfRhVg1XOia7EXwuXrIE
MHyvhtH/uP0SZdDDE9O1XptzlTqzHWeJQli0EuAM4nGWbtLV4AfklU3li67GwvZLtVJTEhowQ2Jr
m/VnDDZz3qU2EalS9r/wMscKscfDBc/lToue+ttRuKLyMXpAGVDXXrQBJJnk7ypmZOX8qpMm7uZg
ORzAyEs7IolEACnP7KDx9HJTKMwRuN72E7ipmQIwGKzbwN7uk3nYkcIS+idR2IYFpyFpvPyTjnB5
hp8yqISlLgXTDibFNnk8+Kbg8d7iwO5f98wGvdzKeKcSwhkoKeDuxhqoENT2zXNt5pLH1s4ptZ83
eSljj242X5vR6v1GTnK4XCInDoXocbKpEeUESQc8isqIfHdffIo/YnMJSLJKT1f+QI2qJPA1hi//
2l2Cx/PTRnXfAN337jXe8AbPIHAo6p0vkyhZdSlHIfbCJ7L+kqioDSbIus/hLxwzDSzaXbSCksnf
xytOYBJP5j27t9pK+05asseY6moOvBmU3UoLH+QERZD5fIHVP16lK4v20tjQlmelEc9S7HTSwMye
iKC5cas6sYAlv5NHCdC4Fu+jrhl4dX/i6SSM48xwE++FQoRVBGab6Pj3N1CRSrbx3eG0m8MTiFHB
Com2dE7dCC4V82UPxxneoaNzzehL+gPpaHa481FfPpt7rQnsXLgTtTG9oZiek74vqA/ESDql46jU
bMG+WTtxLZFukEWTjNepzfM/z6f+Goa/KjjC6gEoPKK2Gxg/Gnm2uYGPL+cTCe0Wq8hux8wbENHR
xT6pmiCBWysi94Y3ftGvUYNNTdMGcmnbqRnvPtIMLVXtlTekE3H6xg5gcmu41Y4lh8DCni0Zkfy8
TOfpk6m9fzMsYhY4MRg69QZf+N86HVT0w3IMmVL1KWHmzUmGnE+f8dVnM70R1u0xj/6FAAGms8Ss
sMptWYYCcTwTo+xa3P6V+YDdvQ3mTQAOrtUU2QAmqoHSxyy1Ni5a+5gDs4CKinmSwNQFC+V27GgF
w5NtCh9rl1tN0VXI+VYb1bK5hkZTqKfE6TWFPmiTLvlvzIpODSAtBf5H8F2oegWnmxKMPy1/IrIO
UOGjYIg4xNawVLxDIXHVajEuX6cNb5xPbj26tbkFtowQjHzmU8EQYn2vvdUIeKAB5NM9VTX6KaId
O3nU8DkRJ2o/w5UmwxP7Jp5aShkDLAVW9mwMCbrZL19kGG8k4CU0XuRqB9M3kZCpqPBP+afsezdg
3oX+1IaJwDWvw3jw6BKsdEw984eiUdg6ceO7wMKTEL3FwVpsGkQxivbnJhgEGCqgjpJHA157uykr
PPOAzyHynyrOL6pSTFMCpfMvnr5hemvyqlydPJMca4ApLcXwJIbtkgeBr4FWfTBXEC4DjBti3uS0
/Z1LhV/mZTA9AEm7sK2405MJlKglT4XP24QxxcAfuTzzmOvdERwNPyOCFCcnMJDWo39aIFLZRFDg
1Cbns/o3yH9/a+hzS+bkUUMG7jEqmkb928TnfylOZL8NEGJNoEUDFqjg/M0vzkRyAqw4EKzBN1Ue
qoH8/PCzokpjMrKVvhTF/Mjll50cyVJVbbBcveQZGF2TrCw6hlwu/fMzibfrY3P8wV5k66B/MGlG
MyIxnKDlQZnZ91ybDCm3DsSiRxZgysE9YXn4WyLzp1BJHYAzUWqZW2g25ZoN5L0CedMbxvAbT6WE
x9bqBeNMuYgEJ2Q+e5AHndudV1k+a5JG36XvrSitSis1aCnTKhVa+pk1wdoYPUlZfmGibn4BvyL/
fOv8YI3uIb68/8wHumT2tpzKvdxB6qRrPAcGHyvdtE4djlI/o6EraxvvsEfaDHM6DXT7PO2jOAy0
zG/Ecizx9KhkVxFOlVoP8rWfgxwFuYCEIYHPpLzKoU5qxHRvkEfJKnSBf8nRv1hE0boNukSLPK13
2x8P6Ys2IkT9qFslBN5/lfzJCi+jkfSg/Kr0GudYfsjnK9AQMqudL1+26EBFRecCdzdiFtV8So1W
yzXrd2Aw4Q9PMVXYwIUy8A2EwExcG0kGwTTmBytSvjC7+Q63xMGyOoG3u40L1Eg1FNMz3bhodN43
mdGiVxoNwk65vDz+d75yurpn/Ra1rPagHt6l1e5szkvGBnTc24SYcOnD9OoGYbLQFGOY2NalbCHy
ehfXjyUUbdYUleQlmoqAeqhqwlOLdNuFnFuelq2OjIB2BcQMWvVUcZ6X8gxnOQ93MbTYv2sU2QLy
Ze+2mVOOsM1MLGrVHICcQ+4nneZlwKlwgY1fo29PMktBaHjuabG8R4Vgjh+dVAg+csG/HWiwfP3O
BDl2JR6z5AEoyo0qDlVf53cuDAL+Y7f+BMCB0Nw8HEbnEnfT8H2L3d+UEL4m8jMXZYf3auYGGtM2
S0Nam2l0jw+21RULTOwqYLrqigQKaeniGg6l9CWX5xlspWaWJA4C8MZVndx5S0H2FXJO/GCqt3ka
i+ROsCVokrnIvS/bnxlIIrue0i/R2yF0nutsLnl+mi95UlBAzOy3HFtnZRyB388SmyK2CDi1HJCz
hL8OOMQpCN7Q0SyjlFyWHZs5+PDdkZeX9F84PZmu3tPy0nxpKkGBidxH1/d+6m49IW2QortHQBpd
kWEoAkeghiY6I1j1n0y+QhbsXUbFOi48d1pt/21Xk+ArtwwVMMN7zk739bydoyuCOlpnXQtKTmvd
pMNmn9zFdteit4vPR2XgMSqnW0tYfJTRdrq8xcEPxGV2q+ZBlRXDvag9eESfk20vlviwi/x/DYCY
niYHGQlzkrntp2uSEZuRdmW3nWQETQ1dZwYuSdzLROLmgV7XbVd1CjGBRtc5GY6X/07ll4MF3PHv
++1krhKZxbYi6UxmKSEsZoOukSwQyeDkQuFL8FpIWTRmIH2PglLkfR62c0G2GemcSah7aQ1U2zsE
Rpn+HQIhN8HCGBIEJDLIQysQNpSkPOI7720bogQ2Be6B+Hg29s8pUSoqjQJCoEgkdUV2qsf9BAe9
3ljMiyrHfEVbyM1waqKOkaAs71j2WjD1gmjgMvOQTqoBDjsRkZwhf2hB6Yyuwe8xdKdMjdugBlDr
day34sFGFz2cMyJHbkD/eYmpBztAc1taOIgOMVoHAbr0JtxU0gBAQklgt/lLwWYp19HFdrS9u5lo
BsUsPib4mfFr6TPeDmo06P4RnJn3HNU03+qTQt3/B6LGvWqFAeWLIXTnFMyS5It2Fc0lFL6vGgPH
IAySpqM6l60XG0ui9Zq5d4egAaOYYliiC7i99uiCZqErndbEIEZvybO62Gero7bcYxu1nNuWN2iG
k7Eaw0UHKmAXjfKh88dYYtzoSLCoZq3Q2xMZUuzO+mwRMieKoEh1gVZujbhkZpQRv2nzHCu7OmW9
5IXIb2DPUuMgAJpwxag9Uyp+7xy58DBtT1Q44NLku4t4sArwOZpKiEGyRmWNtlH5v/NflZ5B10GC
/NaqTubU7ndzTNKCx1vsLNqIiyf/OJb+BQ2oDbpRe3uB4M4LK/r4OOkG7RekBZ5dP4pcLsNPgyPw
OzhEE2w1f+qGiuUA1nsa4lf3vbiQWanUXpciUzGgu8O6APMh+kYTYSRp3guAESdQI6OIUdZNsDzd
mU6+hfKt7YszrdSRGClhG9ogHLwumMC1EIO0ZtD8raHqjA77JxFGgUn4E9AenmsCUMx9dnEMEqYO
pgdfTK7/cczncw0NpUuekLHXm5i4EZ3fSk6B5EfhsAc5P7WgDM31dHmDEj4I4NLaDVoy0pM0Whgw
JwRMr/PByZhEEum2gmBS2C8/vMfav2ixQin6uB/VoQwiCVmHoiYgf+Y6bfOjHktzO8Ddjz5Bb37C
7zWCRvR+/QDLXjqhWb4fCEs4coLQLzx0RRYN7A5YrPVdMZ1fjOa2731z3q7IA9l3fyeoNxv9tDFP
4qYEJTJCpfxtq29knjV/Ev2bWwAKutB5q9Txc8gbudnnDZEqRukJSuVMB1zXSNTIvtOMdrThqC51
V/RNzDVeE2gsUPgPBccUOwhxEm7JXqoukXf8a0IOllpYJWEsROgwDtgEiRGiIDWvvGLm/x+L5Fmu
VUYrRnZZJfucJVN6WAxshSfl2isURCNZJt+UvPpApiSXyiL+MzH0AST9WPiQNQ8ha5t0AOx8/SVE
0gz44j406Z4DXUbOoF+QO3uVUqJQ4HahP3VX8uwxOUL5YgW+TXuMGyhd6VN8DNPXU2YITsGNsHRu
lpSVtjicPs8Cy/ePkvAQMAvuBdxSA9m5AM8niZbs/TlGmQAf+k4/o6wGccPuTysIFUL4ki1HXCS/
bjOg1psJbwXNCabeZpm6M5h6IMCHPJZRz7gbgD6gMOz17G6/O5J6tynzdaegHcgqLJbEiCQN44Jh
4zGBrNl/vThwPoYUyU+HhpGibPKmH0E8W17SgtR/ZY7cL7dT8OpkbioA6jM=
`protect end_protected
