-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zYZ3Rw8C0AC4PoXcebIxmuLyCsoU2qcdrEJ6AD8XosrKJZGPgHcyNAOLX/Ue/hqp9pVz+IYtzi05
po4Ti+xd4mLEC1EfadXt1Lsgox2nmkvlb1BHp8sSkse157R+KxW+e/3I/i53/dfc8tgweabMUNSH
nkwopZti4N7b6V5Bvv6VFGlixIwLI8hMG+Lvx+tXOMUYBC1ewYSb4oAVyWzHSOJfAC8VpNGj9K1z
ElRQmKPSlP1VWE/e8GPrWqeqyWsRXAOrV54sFUopOli3VPcYJSwBK+q5UIaN8PFIVhgLukGxP8Yb
wNPLOcxTE9iZCSjDL2AKKfQ47B31Qo22WUAGAA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
bZ2HdlIKa+sr/XrQyDtAguq+LPqhuEBHa4fMPtBEEgINeE8bwDyjqsuABYBUIqsvrBnvUd3Fyp0k
mYUjYaftQOyvY9ra7PLgK93QYKeHAs8w3AzqAA3VRDVO338Ie4qP3IYS/4vbhTXmqzqaEWBDvL94
MMUMbY5RREX/JSxaSQFn8mkuvLCMbkrXFaWONGniMHY2sU+S6g2jKkqF3VxVQiO1kQVHGjtTj/hv
lxc3okKaaUglWuDkm9Up+R3q9n0jnnbtHMjtfAjVtTboqAmYiXUmIsc+KHjADbYMSJ18LR3tZvYx
vVRKRsX8hgptxqZjMrh0YUiKsxEOcmYDm57QhmUY8HwOPN4U/aQC7QT40tvC1b2oLdEBFQ5HYJw1
c3YeAHuZQQ0wGss7iaHOlul8EESh+Dpk2yilJe2o4zFlp8x4SYBpTNtYil+/Is+TSEUZXoWqsj9R
jeyQPoxFuvQN3Jx25UL7ELllRXKPq3RfzOPNjc1DWQEPU2EHQFH8/4Q9piTKpI+CIAu4gIEZxRyp
cHEs0+vgRTKmHJgIy5/xi7ZrwLRpy2OLdMzUWr+C+0OjLrds7E1QYlGvhq/J4p/nd5WqoiweihBR
nh6Al+6kCE7Cg6gW3oOCqoqhQr2gECY8kldZH5ZGWwA7lvY61DeaESTGPbVsrJkhBdARFN0VMIJF
RpAro4km1uU9ah+Qpi5o2FN1neU/FhM/Fo3f8/iIXDQWLbGsm49NxiJ7Erj8KI7MpqychVGqGiZ9
9ULGl+/O1eRl8S6EKYA/De14k0UB1aGK/0yo8tUUXIazwDiBTiVE3btPc6I3d54k869yaCnPcWoD
/i0UsCp2hes/cE2uUJPZ0t4/qxK0dg+NInqrTkSPoIAFbP1EE+BIay5LBFX5V3svjeRM2zSsSZlm
zJobgU1u3ET6mctdB7LvXkScuJ03cKSPLv0rfrPojJ3g4la7A0peYBtB57O61JNJvBfY7yU7TcP5
hoUPAX4FHUqEFDGlcmdsfgomRIid+oM717n5u64749oRmuQbSIkpfKyDaM7KZ4XOol3DyqfZebb2
0gF0lw5NPe51EXHI9N0YgCjNfc8OuNv/A0V2bBvr8EbkM7RQhZr/1taeZCzjAalOAUFDWrHze15J
zMrzVz0ZeKzxRlm/TtkcrbZAdGJQqYkQxbZEqi8lHXY6pAmZ++PIjhPOkyzzod++HRuxhvo4aGra
+nIK9hR7s/+58FZj91BAClcOLNx33wLklL+PryHA1SeP+dQlw8prsDvDdEwGdl2E80ZGPk4qX5xO
5lA/m3NpEyd4fgTBMziJC08lQJTrf1rDxeL4ahpTJeAQswAEvyQzNWZKjigu6j1HnBBzw3Nzby7T
aVpmJ0IT26vfa13bNeYRvOm64S5ArjWl01VQkkPgOpqqv58FKt2uqEdybVr6WvgUqL7hBDjtrxz4
b+b0D9vkLojF9OJDVSAj4NpWu+L5dOKAWbJGZWobfSgF9QZ++hNYdd9xk2diLrC1FmUwYiUmOQ3t
HmJgxEI/oyx0O99o2/CMyuv2RmUwyLu8/NQm1WXmnhp3KcKWKdlEtZ9VKaO8HwMSoRsDn+9lQWaH
Zzvob4Hz2OhRi3SEqAEUo7JZ9y7Qzuz2bq/yK2nEhYBObnrgR0d48J0xSn/1Mcqgs9F6kfY0K1Wo
cFJp62Vfvhm2UXxp0PjNJSMB144avnOwvsTBsnfuI0ercJXs5BXiSkg1/+jjok0pG3csyjBPGdez
t2EdYNEh+1gMPyvMhLbzhgwUJjWzxvlqpRsuRjicU5tOPg5rSsrKxhMzNcHJStADKVGJFi3Ugtxo
QClaCnsnUZlBrq9zulxoteVqoz4rwNF7u6asrTSRB8sqnt09AOAZ9E/cRhvmnwV9uJgl3H0y6fHs
kee3G+OxVU650lELFZj6zuI892bFwRzOhE1HMg7XY+bYUeufnecDi4IO3QZliIAJfMkOSobk15DM
CVL8juLRVKaudYkS8xCOHHqbFve7JsvJVOdVdoi6IBtwsWmRTrMAXfmhSHqHNuyqgTGvFc/8E/WM
kpOLuQYiUyXJos5XFgLGoEBGtHl5cl0KxuG+bYBsmdoBuXtz21uKngf4Ywn9qdYntCRlFA77J9HR
4ZRxWi9BCPA8IbSVNxrtVFnhMxRY5Qzd0yZWHpQMws56tcRb4KxCESbbsI2Ztp43oAOVF/EMeF4U
mBK8IzZ6Q42gA2uuW/N8UH2AkxEmueBNMdHRDC9IY9KTO5lsji0l2Q3j/h1pWvzpiY/GJuscmNCA
DzO8Q/exuY6ZR3WrXibVphVfmm7Swqs/2BNcPtkQY2NDJ+IfJoYGcvrTt6amSgjCiYuIfRq4H4Ra
GUcu0OkRv2FwhlMZMnlVvP8h7Pw14tD3ahCmC4/sYIQwztUipZbImJF1uAvKsBBIs4y+n3AMqX/L
v/qtu2m3MrLP7rluq+ZIua1oL8z1+eF1wE22Wqfv48ArbRmyHBwunPyAGsChnBS9/RImzpFoTute
l82Kjyc9mjpxMNACxwk6gGBu1qRvyDsX9/M950LYaG1PrU9EXozZcccA6IgYJP1C8BybqgYmE4wM
prwJ/FTk94x1enApqCrXsFfNQCDZPmr16ekOrqZx/iNDtGzupJb1O/+ZWaW2WHimRkmDrriptL2s
F7zUxhZAOHGfl1TiaQpPxG1m8CYEPS0sDaIpnhqVdeCNk9iTpzhLA8PYYtgN8OjyakE3wBRWJOgQ
VQdowlO3h8vhQwFguR9fiqsBirIoOnRif/WmLwMhMF5sMgByN4xZZgescxYfCiu2P5IsIXFHxdqP
9l2Ibe2DRY8wecOo+72ZS1FJit5OkTbnDmeX92IlDQV33c0XrFc2iNE4UM5QKHMKH6MUNjlKEU2I
A2w2rtEspexWxI9coG85jL9AWAZ4FPKFaBQd1UrXxS0vP5DhswMh26jcZs4ka1u+SEkQ26+0U1d8
O357/SzaQSNFAea6LRHieve2KBatKv/FcUofmHi8QISYo6gCWrrKLHM/qSy/H/HquNdgyBVkiGer
WtnPY/U0n6dWOn5T/MHd38Lc3rZ8Hxi1RYIwFb33ckg8S3RBAD2rbyS4HadKBk2JMxn188C2qzh8
jrPKdPemg5XHgZ9U2G0C5R9t716awZ+9fWhTROIOj3gReRL2r8jEpRwhvTsz9uy5RWoA4swe9SiS
e1Yb0eJGGP6nMYRFY2kpSWmQCJx++WhgwvDjWsAuHCDJh0rP2A/OPchnURVyTI6iAhvAKPiWQIo8
OWnMZYnpqm/tnq1T9dk1BedwEaZErN/xNlx3kVWIIUuuj2badkHuAAKtSnDWQxzludUHAxhU/Gfm
rTZZJPLXXEQxUyREQFG4g0XN0IXa+42xq7oAU0Hcu92rmhLynYdgK5wvB6YbUW7ycth7nBhZq9jj
d0Xp2hjZrqqlqc8EHHWigtJlwQdSNo9XNohluweLa8Lg9CfOM6+9PTYH4Mzb2cmZHnB/G1C81XPl
8FTWlLvmVuhK9/jx+NVNKvNmpY03pDlIuwm81ETnYjlaf4enPoHiDMWupLq3w/sBUEBKz4yEfavp
Hu92FRE2WX9mznio0gDbSLSP1cxE/e3shdkQZnlLCwTaTD64Fc2UdMVH/jz6uV8OkDtrjo851wWK
SZqR5ns/PjgD6o3PNZxVazxsyClfhG2bpKOtFUXs0LGV4PwmZIR2jF9tAmBCAbZL19BH+gezDqN8
kz8KNxydEWjjbyBvi3Giz9693WjDQWl5NWwXzcYe56ZX033Hh0xko4GI46sakv75VQ47/ja0ngtY
CKj0+d5BBVlZJlUP25EQsscoYc/7tc2wFbsgOSHFPNZTemPCzSriw1B7mA2PmN+H5RqcalgHqe91
xrh6SLUg+aiAKJPUETHD71abOGICl+bHlqSPndAvfKgZZvxvh48j56hRqD9SLbMLq+FtWQuyD0kF
5MDwHTCJjZsBuj9vI02gwveNIT24R0Nrzl/tjaJUZsmAD7UTcU15xqgQBiSClDGq0RdKFVchkMa0
G7bCVCTK4uFZ4Y36XoXUnIuS43ybFZbKWwjuQmTogMch40zmtTkQQnRzti2yJnowZrEmaHjqmDhr
93f0JX629U94lPUq/05LjRUvdNA4rPFsf+IBckGLy5+6B1XF4AjxG8RbUSrmaGWwVZVk7ouxToGn
aQtQTN/niRgEoRbN9N2TZlc7qBEc5ED9yj0pXY0Lz+m1heBU6dTamgN5gpfQ+UOZCoM92tnork/4
t9ALPGcjzBeBJqBgHLhW18eMTI/BnEhbrtEAfe5RPZvIyKAbmYDe0f3WRXFxGj/USNbdkeK3Jsp/
h6UM2V/VXp8qn/7dmtxzB2AdZ8apJy5gHUUrYdiHoKwlIiFHzz5/zSMeq8Uf7j+bqbVg4nWGC5fV
9bxv2SHHBO8UDiysqB8ixLi709oA9MC+whUsytx8TATLGlwEltVHFF3Vd/SOjNoZIxYfTdKHvZVz
5myKA+bzdDwEjWh51UuIWLqLQzHhu7e02r0q30bN7gcHBu8ScHlERcvzRcTV/B8kka/VgfYzHPwU
7Neqn7Cf/PUtysiF5NWtOrfKQAKFuL4NbCemZzknNJbOFKkrUYxT/0n0VQUVZ3H+KeWfz+xdZRVh
PTToUeFU9QCU189ixcYS79NmByEERyza4GrH7jYzsIbcmPsq4i5ULOKlNTNzmTvoYBrWRBST5UNk
1txuvuYLcjMxKwo0auvEd6ub0PER+aQ6Jli0PD7hckCx99DKy8omJD3N8MeHkwvNPwywX3LWeqkI
snVO1dKeQjjJTh73T+DVxPPfKunfI1FWR06mTLQuou9uHzuQwRkeJEDBzWlT05Kf2VgivN0zO8nY
bqwK9YQGHUBshkDpLKvbQXczecICP85hLOQnU5GEC3G7kyeaoP60H9DUzzt+/I9tF2CvTOMlYzRl
3XbiYSUo2Y+SDEG4nOWEmXBpjR8Srqoy0lATCGF6cyHoVW4uRFJzAZ6aL5qtBBKWs8HHfnrZ1AyJ
vct3m4uWEFVFkSw6Ezx8SdS0RNknQME2Bs1Z3hX/7v7RkfyBZaaxTM/23k9H7HdXQ+Sls4wXRiTs
yebVT/YJkX0JSaC60fDB/pyZPJArD9NBoJSXyM4CgF5KF6BPZBF3dpkGf0Pf3Y78UwtzZMod/FfP
vt2bf5/fg27i8drxkjN3qQz49bHPhTO06bHchGY6m9GeGD/2G7f2DcpCZXZgUEpWAtX7TjXMf3cj
odhX1Xe12OW/odpEDKmhKfsFTGQDFi3HY8IkYWSs5xnzFzZwIgOYPtIf0+Oi7XD5XchfOEnC8CP3
LEtEkorAJCyMQGVDWHHjMnj8YR2+gPyFq9DKfDcjOoohk5LANJV8o2dnn7SzQH+en66jkAwlrQL3
dF/02vPxOAFUuNR+Fgs4MF96RPmigerwlq0zWKY4t16yoDLIFatmPQzSY3YZ0C3QjsDUSBJnu73I
1CiwhmxK+iY4cigerk267FUYnYfi3ITfK6s4AbUtmiIysc8yJjoz62WQmS/KfkjpY6xKARHZgD9v
v+Io6M7QiT0GKNf9ArZSgM3iGZs53VhqtICUPU2xqSqmv6K3rBCKTBFq7Vr2HeU7lHvBSaCggebG
FHicTHHpDjw2XJ+fRiIogUz8BSA6eidy1y4mf4ufYGOOjoPb7oDmswuao78gql2ZUhIqjYstugll
CI+3iEreHL6VKqY5FkmE/EOgFQwLr+gm1udGoTqaxYirg8WwF2iUBwoHYH3sNLLhuvivFvSzvVP1
vl07bG0dY9upXk2PnE7MBlPwSuRAkIeaVqiKDNq5eZNar4uufeCs9O+gFHTj+rApkRWvndCf15Do
VGx2TAtUqNFx5YHfv3sRzR6NBsC088fvEGolDfri4nOinwucRLc9yRnyF8TrgIreyeWBNHLZeu3h
Bb67ztNnZu5XfX08MYqcSK4I8JlOyFMAGUne26ki7ygqZW7Ak7+y0cImDbZnvQYIs/Gq3zk3P1qg
8/cmoWXct5WkYfuI1azjqBgMj1BF77yg1aoObevCAgjjhVJpAHG3JfJWUOPofdwincb2OQMp61OY
XTQLvC8L31hPYKJKsEmUTHeI2MEynDMLsZasAdQccqp9CBT9v3eKkeIo/bwtYooV4+ycrx4SW1Jn
mPDJzAJuCjQVpfgEGFqBApub2vc9tOqbdjnAL3ezeYqAjyb2bGGA/lamzj15Fpqu0idx/I06eSx8
DqRkx1+nYLIlvFlTWsftD7c7PDMKoMbvSP3a5TY8nd7gvNlP8lbS1DVewiUGrlj9ipVa+snPBzT1
Hp8vyC/N7gjavjidyCqYwyhPC91LAUhpcUU0xr9v6pwVYSvevx3skkyjrfA7UOX94qVunkNdcn5g
Pb6T6SBdoWGPUiSNK/ZWe5sIjRTSNWhWILFxFbdz6+QckE29euYumi3UyhFUWA0t+WxuYuOlvTyw
uEvHEe0iheNrRbNw7fXnQ3kdrcYl+JI/ZfZRNOzyofCKrJ9QU4bWqJGrtFEAmZ94MC0LzZJDz/IM
JjivbSRHmM2RuQwbdkWMlruKXkX+t7uuV2RMo7JHN5FO8/3OwxodY7pf1j5I2Nk4eETIVZkg5hUR
6Tl0yUXZQRMMVOpyKR+VE20pfnp3j44828HZZFenYrygdiiwUMjFxv6QGbMmYTNCVqK8WoYrRpzw
lek8/4z/hcBCPQtjLoROhdYIREagcR9NRkQD8dN+3zjw5to5hDBek1MWbYrKA0C2YOdXsyqaFB1O
p2Mw8Em9/XHHxghJeihP1aM3Tm92FKP1DmfTuoqgU2xa4F+7IVLP5vh415m7+yF8A+FnqzyBY15V
TwhLttimXG6STUwtNUudRVabFvhNLEg5dQxELbZPS3fLUGuI1lJKt7AKan5IWSLRB5R30vty7TXa
Bzt5yFEIXAEovfRCTRsBPHDmBMcPQwiLryHKY3K+MYi8+KTHWB2SQuVsAROtew1V8cuO5mco5W7n
HcigmtAaebp00skKe8gSCxYE7T8XyhGt5ERxRZHp0u/Hy1dYw4rQZpqY/EDZJZEl2yDYmeiUF8Q8
dAqXVqCPV7+OFZaxpdD5ew8quIqy21Xug5fuPIH1WOx/QedEbz8Y8GDAbUGgPPWU2YUXaNVAXOKF
6hez+rrTfS9sRFQmsXRZ//CKCyrgiQkXCYJAA0XEgj7XEAsVvpmNniEF4y3H94WZTqYdBcvVwThT
hs5sUPTb4dh3IbLlq/m4279dm6+5MH5yCYmFtP0gS3WSuWIM4Zn0pcUHWHaxzJovZXGEEgGFk1UV
T7eYOgjPBGBvgeYv80gKTrhoo7hOBOtaXFbfre/Jq12A9dmV0bS47sMmcCki9BeXGynBNYta4Osh
D5gWnzSbozjuBSLSq1NS1mhDbzZIv68wn1x1eB8yollJCB4bcqfKjtaH0mHEnpDxXRn2hJT44G7H
QdDVV2aKnOHtwXlhYAhM/vJJXV1p7Mh9NU4hc2PkZKMs8mDXSItb3gvRonjwZ2PewH59jr/bNSGf
t4O4VwNVVMS3dv4OE8F77KhrfFwFvplIBpkOviCPjXTM/NxjwI1poDfHIU+tx4GK306exuSGcNtA
2DEymX3Er5re1wlFehj3UAQRzeU+NVdS+5enkL3tfLdIpvtH69hltR85MAbZjNXrh6xXLQMFRxqt
WWeUxGPIsRvEMpdJYqNxHJM02Fr4b7y6DaUP6W89aGnB0N89pEoX3PMvi07BYlZ+DlzJ/pgPN5FH
iyuDb6IfgOpAvc9/rHlcMpbyHKxKzwhsmE+IBJ9BgNbV2edK31ff5xR/PNNL7mEhEYxG1Xy6ACYR
7gtgBCDiSFW0cjnrGFnb8sZ8dcTMcA+2/g6AWsitTlczIFDDgZ+CwoWZb62RLBkYPIxtWjVLa2W+
BPNHHrprQvEKIE8DTyq5x2KZJ5JTjrWrhWlUkkMFjbgQyopeN5GDHN4oEoIy3iHzTK+QsUebN0bC
rdknS/J3HNyGEJBjGA6wDNsOeExX/oMJhfkrDdm7nGCCUKR1resH5aIZleyx23WirfwUNkGNsSk7
HaTOZf2JL+WFPH2FYLKAK6znEeObm3F6I07zJfXPDtqDe45qV2mko3+8S1i/eIIW2/1TySzcUWys
3mxOxcDV2zW0mIYk8R3ch3gxHkvqOVbvUy5u1BKOOAIryAmZRe/Z3IEJf2/snnCoHwv97D4+hFs/
HqC/hooGgGiakWI6b2e+fGWdndAmrPrQcnAtRRNOKe9Z6+EaIyfJ8iptQhBY8rHsvwipHmsGwxCQ
RRaHmeXeBPc/3wl1L191rZNf/8EfgRmfnrkeKeZlHnQOkht3otFgoZBVkTQTdDeJN2n2wR158fsR
HOzxN3cgat5Kl/OLvIN6duf1Og8fA3XNyiybAsBtvsRrnQGBfPROA4jLCIYPjiCPn6KtnLbeOk4O
F66ge5c2Pkfpo1vQvk3twhzVs9nzm4P2e8RTXX5tHIprkSOoUh6zNAzq7FCD0PsZvTpQy/znfIUH
2dRwWSlB2JzaIAnLr+zfyTY2lmgvNs/RFMqJMBStnOZdokjH0op61Q+ejf0gJGeTnErtLF8LcHiC
pbzK9rlF9s/UYmBmmFsXpQkCc9H6cAJTCjtMVDwM0DqaMsqUW6ORZd3eLpw5tkSgvKMTzLmmS2d1
7q6iSZUeuY0gGxAwca6zKmHguU1eGH77cG1jlDcl3jNwXQmAJjruyilreUxoSm1GhASdTCa9SAxA
jzcOnahGLNAUSadqoVciynd48/hZEhH5u8cUdKxvTMrlUCSzJJUi/Ab6V/+HsxqE3QWomxrdwF/+
t/RhcgOpKsNeTi1vplWEtLz3quY/YsJO7aSCcFXP2DKf4aCN3zEJj40+Bl8XGBlRjN3JBdqwlGmO
05Mag/INgJq/MEMx7i2Y9qVmYXr7B4a3fT1QxUpcBjk/VYyHhHQpj8Wc0jhRtOWs5/ytwBYRZzYR
CGXI6gsGmOCWePPHwH+MhXQfujDPWYfSb5lmKK77NlK8ts6z+Ks5fHMDv7ft5u1ypWhpnkYeYmy6
rYqIVTTog4b/OJYADGA8fA/sqS5XRUBAlrOI+c7wLsY5qoODXvqVsCu/ySX84ovuIUrnsXjhrmt9
/Q8qi8qhHQo0qTrLnq0XwVOVfqqkuM9XpAtGR2K4Uq0DkVpJgjhAUfSaSyeIxtw4s17O+0acxAdg
LvCPJwcL/4Ca7fywPX2fd/itigSBZpOVIEO3Vg1O+gz4DkLDgW2W6AwJNra13Y45OZfKUa2/n6nd
c7+Ocwy0p9ui0TCNH7rCBcX884zzgufPqZkvPm5JGP4avnbsRAp5iksL1Z7ffX6xiBPksD46hlxr
8RUW4I28YdMVSYg7D6X4Z84XPdc2rM1YyvkpUNFPc1CXN9hAAFgyO3an3Ezk/2weJRy6dDAnCWVx
DNLpg63Ymh0yg6GYLj0iT0TyakqZdNBZN/gB/tK+PX8odeDVCRFUI+1HwQIfQgmggGRZ0Me5WN/q
5qja4wz5jcx6m5NxBo9uXBB4/IwCFiwd1clrQci+QtQgctCp60zmjG7W3FNb4IWYRgd/EuuW9keq
kRye0IXe0mD4HcXt9sJkUdWK1y4NDpYMFlUwG6r8CrE5tgaBXZ/VC3JKQPr8Gffk2jHQQ8ZXcisK
SJ/mABGRhpEdnhZy7sagr48bo9ELciCXlrmynhuoOgG0HlSZ8E9Osv3u4WmWA+67rwS1VZOsifIi
Xmh8R3UIcWCLohaZAcNQ7e3APAJN7tfrC3KzH7zxXUwbwBQSEBNTzOmZTAuxACrbFnSTm6o0NltG
Gwg+kmw1yw1hlAnHdqm2i+BgDY9I1HtpxiVdvHHw49kqxaTEkuxfrq0Pntpkzs4cLQIJhbRqOzrR
wqpyjs8hx26G+S8w743S5jFFiHUEexnJ9vduA5gY9h65uEFkotPtXjNSdeS7ik+c5cLMDTp6wmP7
YU30fc6PeerTb1iC9r9VHm6CkvPU7K/pPmyjyRUVeTTOqabTEdI/hYkqQxBj8edbZrjtY6yj26bt
H4M+cBfi3ssR8RbxNSJRto0zbDw914uC5iErrmLX3rgNmypmv9ZkyShbp2Lr1KujyvIgNrXp6GHX
e4Mjx45LnDks6CznyPTUHXSqCDrY7wm10C0j+gHvxJtT5ZC4akdJc4ASU35tsvkywlAObqQFnNc1
tho9sPPsAmq/6prswYHN7+liiiJYCtQ6Oq16Xb9O/0Im0k+LBk4z0XHaz+sdeDyozZtPhOSoCAN5
/X8uHIqHsyKvQLfxV8fhOvGclENdzlzXCCAhr034gkpYktp6KGI5HIQk1aiqDxn/J4nFz5fnGjHI
qCd2MNn5zZatN0Zfq3qSZK5jpW5Qd6sEzAZ+kgpUIQSKfHYh/tsPpxJf3RvYj3N0MpC+bd2/v/WA
QsGlxrA4iLYaOmWHoh2yRVCEBtBwLwy7OPUIOeO8uk3vI9VaH16KzO5xOQyQTOc6gxaedyphL1P8
KnO4nZBHKOmBzAY6Kc2/PK5gLyxsS8jfMYkG7XN94I3R2J4SpDCmleyQquKWqS/PIqiBmak9CvK7
d3gksCRAMzWebwPd5wO36z8FsQAuSMcW0JPHEm5wpWr090fGhA9pb3ql4/aDL4iQCWx/05PbfemO
Dv1LMKrYXYcR3RoICUkM+jFROqxTOw4A/Z/yhUMv6U4cvCRUKTWfQqSKVRKGh07hJjAosJuimUZ8
/Y4C+xCQbwWyhtP4D4DZswHAH1cXrpbeDsTTziJyure8NVdi8A1aGTCUi1KNhOI2E9toXtC1wjpi
op+WJpX1SUNvMZ3NIklKJtAnWhJcxGBOvSqH74ICh+BEwOjQjFwpUluNYZmYz9C9UTm0vqVglmkB
SUuAI5Mb/FYWPKqXCZgX3/aip8RREkSiCW70/4QTSHed6tjWyR+tuat/AbvoEk95C5Bv04ldKXdc
jcqhnA3VoDbS5Meniht+OgG4T+a6ezjk3aOewnkZVW/hR7Wv3zIRzIGD1/R1RVS/McjuikGxOQwA
BwjtXpN2wV/NAQm79e++EEb2639S0Tu/eKsyqKce/KY27ftoJMHYVvP5+ntvuwNgvuqD5z0HRH6X
DNksrH5oyaVKsV+eqqJaZBGeZwm6EyVvBxEjUx54hR8bCl/B0BhkPWSnPR4hDpM2bJHUPeNFe+B3
Y4GSoi4sZFOB9xVeppi4SX5G5JFlB8okb2+kZpJsiIBpJbu9s/Lg9ictuUC3Qjl9glbyowtLf/QD
/5s6YkRsMIzrdLwxrdZa4wfFJ+/WiWOlPuB/mlVzH9nTfzVzdPiMYjW5jKq3k05ToPz7fgiT2hOP
K4wa9ilLOzoB6KcB2OOxT9twxEjILmT/o8/6RTWGt8/abJsMP3glSB1k85MPe2M2aRyn00VXD6LY
6eITYETex230FFN+mLdK8Ou8oL4qQ2+IA6Dj10T2mGKdCO88NTYQ+F0C8Z2j0NpTr3V3kQr1nXUK
pFdYDDjNSlOMzpE9e8Ke3obMxSrbCUMc3wYZJSkYn2lZ1fH6OvsaEWiskLNYUWlWVZR4yFAI820Z
Y1x15tL5n4+/8P3jzsF0Y9a7Ic3ir6zgsNDIZTaBx7DwfiJ/ozZ/frm+l4xHUmp3C5+3UNkc+KfT
nojz0z8kB2pYOcETi0UgFWp/23VNZAXNLNHAAbjPr5m61gH/y81y6fbI7rrp3cJSTOY6V0UHjR8H
fTOfPqzl0BJnEOjcKw1RAp1V0p8s177X1Xuxaxmpa/nMKxUvg0fWRfScsFP2A78+GXK5zX0rKfe4
tV9TMFeCQyHeWsrmAj3WHm2DT+BRQsZnlh9A/FZdqsmaVXBvVvz+iwsKR/lNbvRUCFMs81SVVuAI
nCo1G/La9PuyIdqFXcSBHnNzomGPTgDiQJU2vGhdnBF2yILKrwmmTVdWsZ7TAlN6CM7sK1P0+ut0
9i6nSbVPT23Bc8yfyI32lcC/G5MZ1P6eNjcPctIBXx8EpEqNq7Kir+/fDKv//YWPkGszNYDDoyZL
f7NwCSwOFpswWsR78L5kw40hXpn8umAqfJZex0EWs5ZPdOrLwDmiKoq2/oJA8qEqTbX/GmWH1fHx
lMBvXyJeiC7/CbX7yirryl1q0s9rEcPXm1Qh0tPWZQaSh6IQOH/uhE3FYlES1Jf9DxY+X64Gr0zb
zQd736CNrJw+pgsogdwoDf9M+rlFTNO9qxckA4DsrTq/igKTmbLOLuinsqB//a5/91q6b0L7f9BT
mafNXoTxYxuTH6WWCeVkJK6ZRVs2TBXuqElWsL8pjJlH5qjLfukUqLHebTnhonMgjkYRj0JMgwdi
6q2iethBz8VydPzYHZCnO9I1tjG/+iKl/D+MRz545BmJWV+04QeUF3vBrl48c4PdFneNPzqIFITf
gOwRLle2YPC0ExoC4N1sSaiokvB7OMFKmoJiGqNVYrgxXhuNOS7MfZu5DgY+Y9LppxztV3x2zLyP
reSfxYNUa1wlVD0+Ro9X3GEAz0m6eWDk3hzkB8CM0VdBYv1MBZ8ZKkiovmVi0tW/KApT9Iafk39V
dXYQFHEo8PTJXV+ABnjOg+lQZneIUY9Nff7Uj5KAOQ0kAlET8zpmmkT2Kn4HQ3DpuJunBn1BYTZQ
JGg/uYAK2jW8DeHptbfM1S0sBJjTwMHEvLp7dCKkHq6YyKbBSbHTZXrRXl7WP0IoC5osNmlsBPcz
rBBLwVnNCcr2EYG+YyQB8Pq1/O5qwFL+UbCnVN+WpB42gyh3FAkcEbnlKLx/9ScShCnhfCWsnODq
5T6uA/C/+KxpzsSsOtQ45sbUnQY+WR1tvibU4N2XO8K9uWwSXdN3fCHw/FpjkevkVoci0cwXg1mN
i2Fi0dy19gX3v9wavPhEpRDe/EjFE6xO4/bOtIqVI+geUHMqZ2aKkW1vBnPK0LYtPm1/yr4VyWgi
YXfKEFvnZ/qSWP0pzoqeFsq79f7XExBR0yAlAbQEpqY5/mIQ7IkoNAwUhboRhBba+GcWUaQNgSRc
/tQ8W2dLOurZ/ij2xST/BJ0VSTVwLSB9rFrI2zZro6HOA18g+3d/U/XmJt8ybXMPLPLfXxPiH7Xa
v/fD3+tTZQCDuAwMS1GghQGsp4Lsj1pwjQDbxJ5CL3Hplo+ZR3XlAOerA1aJYKct/hM1dS+w+rK9
s/LaFnwPS1HKI2tsG0dba6RSgeAoLKC7CIE2WbqQK97AXeN6rjh/SVdxQBZ5sOCqbx+/k8724r4+
auU/ntBM5iYwzhImQaxQ1X7LVC3aFQUe8JVCmGHYYWItiLZK9BITclLfu87WH0EWxQKEbhmhqbq9
CNbmYq1IGAlYCwpTAgPPvBXL6NMv1J+QLb13Yjwx+aXAe2dvmTASiDMvhqd4jIWG6iZk+n3+Kj0A
zX5ovRIapJeREqSc47VkqlGtXvOCThdm7plIvw7FJijzx1CBIGY8AA9G9K3QkBhbRYgtQCeCAyR0
/XUOrzmXxWNbbAC7S9CMqJ7mAI8+fjz1QwloLZ0T9zqTiUAl+hbBo6XDq5Ky6rUXbDeQczO6uBI6
hpjqZe/PdjSD8uZxNra8P8rgoNgLt6jV4ebY9bXrXZeJzNv7cnk3sbfItZoor6HjQu12KI3lahaP
kB2HU5TrElKAn5DrSPS7vSvM1oVDLQgB0Vq9MsN6uu27KSXDnRYLtRpzsb2uXzhEQatiLOYJkawt
qPxIkk+TelLH2P2YTIXowpQP8/p5GFoxG5E7gqAK86+Mr3qy3WsX6Dc86Pe1PxxnBbgEF9eSz3iM
IuZfWnyz/3QxtlVg4BnjjCIQ0eyPrrekRjs1Dvi0tAfhgJjzH4eRiQMDNceDAaUNzC4uALITk89h
eMF7bmwhOa2qSauAbhIN8fAOqBf7tzOPxX4PT08xmPdhk0/l+y9KMmN0gAiVxgm+GCJj6gTOpvk6
K813B7AeWsIpCGTghFMwvIclr36ljTYEVRPRvYcK6kvAU/uNwI/ghhfBthLQ0+H7zsrZERjNMqO9
wODnxj/Z62hNNVpR5Op89glyyfw25CP/cqX9YTROPo9j5HPujw1eoqpLtJ52WoeO5yrA+6YhPMgH
R9q/iF07rPb/SPEKr6JJX5aDQOXghQhuLWKIjnAgp5QTchnz/m2F4QmBrBQzg++oAwey4y1rCyQB
XLxy/+VgtY4zJGB0oUHFxmwVS7uRZG1ty/s/NwBzTtBv+qyl2vJNhEPNKSMb43tgesOlLL9u+tlv
XCBlj8aYC6n2ifq+HaGux+GttRhtVMdIlMX/BxVx1vfJPfdT3EoarNs2n8jbDfe8y/Bng+smNxtr
WrmYnXpKMB/prdVze1omY7P3PJYo9tPYHVLC3Rzpa/8sIuHrkpPI1d0859vuGAAPwfJhI/s2upQ3
H2IZWd5atq7c/0mqm4xIUnSiFUMVZ9WNE3bL1LA8hD7v6UQX/nd9lPBToLZmumDgBUJ3H4GGNUNP
kdsdDa31QekDeaMRVzFs+T5YKp6DCbrIoi1dQ5L4aDiDPTRjPsNTzZch/XBi/JQU3rZSYFa/QtrY
NTF4/T4BR0ABb+Qtucb64X4SH36cTkfigXzX26Ty1KrezRccv8hVKiAQCOm9dqnQwa7t6bpZ6fQl
TxNHdaODJO/62XAnu/S1ljzvxOJGHGOFRhfwduXa10Fqp0hU1BlYWIzkFpZxkacn37ygtjbNUKNi
JyaKN8uWSP4ELpVzwq5LP8iqmfOuXTBYiFctpbkJZNy8+lVddpfE6JUBsfwKL58APFBwYz972LRQ
ngqs5Bzc97DUMgwuSzqP7J5k4n1NNuZsVoWuNTREYcAlU+L1hRzPZ0f9NBXN47GfrZBomP5ntv75
qTYWiEJtcu85y7bPR9FPFPxATUspCHAcAOhWfXiaru50gLECGdo7AKhhpziZCVVnNw5wcPmtUnlX
LCFH7n2kUnwCt48PGDeNSvKt2k0hHzrRAbZJNfglp4jxM/Gsed6TC4MO1lBpd7ybcSg+/sv4sR47
McLm8RdL1wv2WruVjwxHNXTRLYFryorrZdZ17uNyI9Y1yxXKGwDO6enPW28ydS14lEZU7MlPJeHW
g89p3kc+FUkmFQC4OWtg0gudQaFGPtho8Q7TlgbgKPJDi7MoAvcOSCA1iYM9zINNZn4qGhYpBroV
zyecccU4wS+g8U2jA4sLzSWPPdFcwhJWTUhhfHIXVyyU5YtIrlnRE3VIwJT2DhB1+WZkntL0fuiy
h3OKXAdQxBvJv6Ymeke3zT7qTOAtHW5h26BgwigYip0k5QstN8FxRWTqf+ovzXyB3xGvKY1iMsUb
igRSHP6ga6H1q74FGObYJfuEsg8ArYz0/NdzXD1vFWFqQFR3XpuluuK4XZCTLCNoNYskMZ04TX/+
4g2S7Yx35lhwGJnnR6tswEDgsWERjMVNlolQWFrAQhm1RMG+P83aQBGF8TAMDsf7+BWLwSSaMjCk
mB0j76FhVg2DNVEX8SmJUZ5X1xeXYHmUJTetJN4rKVj8b8rpuFfJWmUTbnnzgiT5tv95pvouSLkD
R2ygmGfC/mpAkusFXlku2cX3WCMiMJ0l/oDzyTZAu6pDBDI0cgo9QCL4KVHeS0A7HhJYtinmpJuA
Gj98IPcevrNfs2/N/pXBs0oXrLfhh43316U37ytZDFg0BXeIP3ScwZdyCRVc44tLLv0KURgYQfvC
e2oHZV9qNc8MrZYxWiaolaUqXcABqyU5Gcxq7657QML+AvsVLe+mhXuCxDTtwRKonq/yGyApM+t+
N/qQjKpulVoD2ch6iT8KumrrsQveIW9MXbQAeRjg6c5zhJ7m6rUhtR33h5gPNxZDtwtmmlq8sGlz
lgRqF0VkqpvqjVAoaiQGpdLFSkx/agRt6o9xgbQBq3SE8A/dRKrO9Jkd+yISbysJcbbUVCOqrDjz
IrOqOVS0PsNmvQMPoFebDaJ1Oyp2m/ew2n4vJUfAiIS9AUTRhhRJBUr1VU5yECSIKpa2OcVUvuCn
5rx4B5Bmjbx4bRUZ1FZIvNqGu0aoueiKOXHf6w/crB8cxjxoA88IxjnWqMiUpDNAKMNjRbzriRHg
wH9d18G1wu+II7dM2PTXQC2XMSLG3kYbZqVu7oz3U7SFGp//o28cMhVLaptNw6MLgRYkfSM7bOot
b5I8us1Operdc+CxyASLqyZvUsDnQ2Gh8jTmn2RaYRCoiOsRsjf1d2UWpx1PHFAd08uAQkF++ZkY
yI6TSZX8Cm72/Hqqc1QuVKbtcH1e687yP8gaXQkwhnsvmcPdN9CBPrvyLIv2xF30ZFsbDlNvAfYN
xPtJYetA10xNrQPKwujSDAOL2lDpxLOBdKwxzkHKEMVTF+o1FutlOv9INDUVam1Vh+uXSTPy9ix2
xxyTWs4emavdwl3iak7pPe/cGUBhKGn0iH7dmyK8HknsFKTULj9Xk5qUGdtvjY85fngjQXuuYGBk
6AP8U+lYmPIrS1FacFYwPDdU5IoWw4sCB3tJSXaJyRn2bmDclFmQOZYEcuiEQiAuEtD83tDOhKCj
HothyDwx/e9yUnrlQ6JANq/avM2uuoS2xdpaE6pdpKoliyz2CTyJbER+cEHMDqDPFcXF6kIX3e4K
kJEka7JTvPCqAbPoh2+mj32fAln6jIG8/LUtHZj3zJ0EUu256C67LDZLGwav7cavG084Xv6yUMX3
ewBeegoyKph67SXcX1UQizdqzdNS086PTyfAB011q7Kw9rH774SBZXbnQFX+REzVfxJZSt2JLU0L
ApkmxptJ2GyRV6ys8621GmTO2W+MzoFTmeVKwVQT24YxOJATjDXcAbk2cEKCojMtNhMZPXqaxLhI
KcQ/CSLqmNTd3GKSPL6xbepFN+OlIDE3UJS8OzKggsJNRqMRApfcl8G8XC1kZ4gK8+kkJv9Gf4zQ
l5AcwplThz2DbYuig/uNa+j6fJ9s5d46ftCOwHYB4b1Lo60eY9YLti07DSTNA0xn/Jr/KELSnaio
rPPZ1xWVNYOhACnjLEqHewiO1SD+daXcqKyNhnvEbqg5hzi83kIhO260F+Zpgl9P7ln0qb4W52By
X/82cBdGwF+xBxh35DMPoaUjVX1J3JsGcZ1n25hidlNn/bOewcfOktLppnAk4meJDXoWiFRS644s
jkPoLIa83R4M4Z6sAIKsLbbPEnivqnX0uXwLhhIMOSpNQp9aU/bowyiKyhrtx67ARBgUFqm0RcRG
nEPbkHViJ8XCJYt0yreB9P01q4pxHvokXNQ43C4Og4YtQ2CkfZP+w5LdXpdVnoJNEN86EYXI+JhM
6FQmSJuxTx8kC8C1DkOCGu7GgxLMHaFDhED0ZnP642oZIvmMAcxRExB48VMksFbSYRxPabvHCKki
f6S8MQWzmljNEryh/XtJwHvwXVhLfzgOGtFAmictLckZMQjFL6aREcIZbnajkmuXjyHMi5T7dGtW
HuPaEt3x6OKI3zBrMQwggm5JVNZ+GJfe7wlbb5VVG13It4vTylAlht4sovVpBX5aa9C2utX5AOym
97VLyFcKHM4CEF11v9T4ptNvmduH26ycL0Z/r+/D9m4043O4kmsD3FofXpeu1ezvjfU2Q3NWy9lu
vJwYnECJ519ovfTcsrevr//9Cg2YVEWfy7r3CGD2ix0Oxq3nPwCTD1RN+nSpZo4iBea37pcgCzV/
BfeKC8u2kDjtbjK72pOJljASflBascT9eO5CZkHNURD8TcyuGqVyNxqZIwCl6I/0J9X9DQxTgMOy
kAk7eNGMgvJBoDSsTnr+Tv8oORXOzazvKDKPw8U+1d7vFqG0xOlG4Ntrm8p3Huw7MuXLvKizAjYi
gOHIuz1gep4UjaVkkLyO/mmtBNiYeXACx/QjJe/JOp9YDPTX2cv4XDxkgPScpbHDWh15+gSNUD16
zjm89K3zhYNQ8oCyh2CVaYdgZjScOxpUk4KOtlwofEUDXcxEvNNqSqtYbX1gLeJIAVKoz1fufCcd
+3GRPwmFiuKllAWuPf6cUkTBW/4W0219jrb18mzfi+c2Ouip4Zc6T9Egphx2UceIn6H0MtCwOLc4
Ij7ffux2QOv5X/tebFOC5kOo0TcrtZEQHsNVQ0RnMhNLuemtisXCI1rGnt/IzGKUmXE04PphMqwd
qfEgZUCsND4q3FY4EBPD3iNnEEZGntF7EyTRrIjPPgDYHjlcl0igfsQkEkrxE8W7SkRS89G5PXBX
bTE1c/Mwj15LKZpW6cHW16UcwFHFbWv/PhVYyavIhz/TRLgsqQXZUhQsNLcb0ZLxPELgc32qWQcE
xPCAlgeovjRtgsvK/oJNouRRZELpUERms6OyStXbPyt//54IaPkQeix+zeA3ZeeoflcgSUZCcbbt
vyl1jf9jgf1Wb4omT77tu4EJ32lM9deqThZfo9xTggk3GYR5KerS+9N5mE0LpcJLU8b5vp5T5iw9
KJMRPiVxoG7SzlhPXRGakWCslkhR0PXIj6Ko+RfMq3/guRXkVosWwYSVvKuqbxWxA61aluJT0nWb
G5JPsBBcMb0bAZ3lscE01IxI19TOB6B31qyAcANLP/K3Kz2V09cp66oP724Ct7ekWSHfDgHtZXVa
jXogTB7tSrbYf2lBHq/9pWELteloLvhnGL/DqfkPTxCNqi9P9Woq8vj27pAGiWlyiLNYiIvF2ByZ
tNTsrmnvuGHU7OeI0kJ0TKx0svcr9f0A2gnA4V1POphdc4+guTFN6NvW/reFSh8G5SEMONsYRNkQ
yQJZrP8R/Et+lY36D2soiGXmBBrFJfySeeuVRI73q8j4lbib90LGWf5Ma9KX8oD6mexlU+mqe1h6
rb3V/UVXxOWoMyvY4GpeHEBEOy5Anpz0NL/Y9TJNWQlrtZ0lWzhBdpxMB0UhotbI3T4dJFbF4UrE
vAZunHwKdkKUc8i2RgaBaSF4t9saDRbQxbMLpU1TrwKtkCFs5WfAcefphPjNLsQIotYJ6/4x5Wg1
PxsIL9YH0bJsr96L0kGFGAKEvAYYW6n0pwVJ0W9xWvf4f2pivBCNgOrbarVZBAhblWvSZ+cWYULk
9rBJugAxx4OW1AZyMF3uFjPVOGh+txtdwsUqeqQNX2Si8p3VzyqUMVqVm7NBQPwyIzlJ9nLnA56I
B8oOWrf9SCtM8JYI/K58mOhO0OCkr9L4jVto/3wYFHFgu3Xnh1TKx4xpdrq6e4hprF2oYa3a9CH9
T8N00A8q0YQcVCsuS+vH7cvRk3TyHdwqw1GkpS72uInoJQI5YkjfAcupS8040+vu0Sw6PqUJeYfa
NLwEIvQmirmuQX5LBVIGPgn4IiM7xnGUeFB+lNiQGHv2nmWoRphPNcdZuJjOKkbu85wnBSrYoYiY
3I6zfI4rbKp4ws4+OOM10BrMHZMxFyY9UkQjyQYC2WWWE0KQIxlywsc38ig1uLlOv7vS+UZSCzCk
6mH/9omPbOnst4xYXhg8P5r2/g2AY8Nru5a0GLkP68o2rhhidwnwDUG1e5YxdOTrSZE0yhNPcL3y
T1MM1p/RFzc0lAUKiK+6oRLra8ZvPScRAtDDwqUxrzwtdW+Evn7Y8A49Hp4NXsDVujwVqxPFYR5E
Q4qmpN959nJI6yHNiLPbL9LNaL9GkCSVXK71WMzI52X2bi3V/3p2ms9rCEbQlc1+cTjjVQHvnqL3
Fc/UNs7/4e3AgxhcVdu6WoQ5a1swyNhKVT35hTBJig2/eWAZP/LVXlpNj4EWsjba2/Td/A+Lm17i
1JkM5UPJLRWvrJ0BzitfDRr7HgzipuGpyz6yHtoMlFud+D6KsA/Rnz5cy6r5W8AvXkDunx5uozun
G1/n90wIUzV5gD+3oNieL+G113niC+nnMdoHQepJLsiz+UatQPd81KZD016iAghw6gER+F9nNKvW
mx2cGWxNDDOfqw8geNXTVPxNIUD9Dv+9lTYYR3qBV0c9Je58exUUmdtuJ9qfigNAX8BQ0u+FU9Wt
YoH1R2bkjfdZ9aSJstt0GO3QjzN0WInTSv9hoKB6AfxQuWWkJ23kA5pFBrJCglm4x9FWOXSrYAzr
KW3C2uNRno51r79pqdZBmwm0Gp4unBPGWntBpmivq61EAbsKTv64JjjduAv10NsPmaNMgLOuD0Py
gls9+SJjczAn26BWMLsPahAgV6006f1XOihctygqqvh6UEhXAJSKmx1YAyPpWmEKZPlykORqpJ3t
vAWR2aKJzVRobnklsMiyp3oLL+BOPXlKVi7WdietKHFFUCP1rPSfJx5hSuxivgpiYaa44VLn+ylA
dRM2k6VEV5myBLf6FRSSnFdEBGt+eVtzv9VYFCUSztsWROwMEyHE5QB6cigu1wEgfIBaWdjfcN11
12rqvotRubZxdU3B0Y0SXyX82+V+spc4JcS6+3e6wr9ZNOu59Y9CJS2uc9Bs6mMSBm1prOzR7nKE
eGB+TD5TiOHtOlW6nmHbtAhMMGHbUa8CtZFk3mVG2+MmeK1oOGlKn+ueslQLuVg5FMczqa4/d9Qh
UdSFzaiKXPvK9FkM83FSADmW2Gftxwu5p7vcm6dy+SyL6+GrwlbZ+8Cuv61RfcjzfWIr54DF0VW0
xb4OqnTija7LlPjApm6I2JBF7kT+Sf/xRWVWlFpeYokVtJefgGretfu9kLjdTO4xFF7icb/oydac
8xjx2AmqDbMQ++B79LydWXwmcuBTtft5OAm7MFPXBH0qbn3vAS33F1zSmSl/UZtRma6+VvRfKljQ
e5Qo4mJ6MNqGHARG7n5SoBYo13t1tXAgTZBO8OgHTbp5gf3MTpI5I0EJ9Q8wnAr2pTwlrDvZkOIR
2pN0CfPOOrAp4bV9Sy/maF0o6wXWxc/GrgXLo/JeYvkY3pdEe3Pd1m+KFIk0mBeXwSlHIDW00Czz
4KVpTd5Pxo9zU7ko8VxOSB9gK4sVHnWkbL/8U9ZDTbZfDJ3XfI4jfyZ/VcuResSGqW6eYtz+5iMn
u8DLHziUwTIZP4uD0TDiim7Scvih5rX6puDSsS8VYcfp9e2k9bb/68G2keOMpBgMfcTk0rOAbpHN
sG3SZuspua7TlMisaFOdj3wp7Alf4VzXDkFNXrjjs9ELNR8oIkHfZIwsMv+slgmt4dbr8txSegC7
FLRWyzUuyCkzLa/lYErhmvon4XAnsPCFNSmCkMdTZ7RzCoafMJREoUFBrQDZ58R6Ms4uh8OTqrE1
f6SizBVwUo7ka+5/gY1OeyJlMjH5nguFwshsd4niowtpKxE29bHCz9ywQ0bOal0wsRReXFOs1dJD
H2ARP5mvNeWIo3Ez/rMLCprixAI+/H6U8bh02KGSVtdKLZYAk+tzu6JoZv+vA7H6ItpC8ldg28Zd
az8w5PIu60sX1c/dYBDuJ5yHvYo2Kygisjune10SJ8PfdB6o33PdvSBpvos/yGKNtj3MkczDXQnp
F9JWn/vzEWswOvlp9aGgh9Wer+RRAPzkQrhxgFRwEM5aWxZpvPmR0YxK2mdYkvJeXTZvMRoH2/Go
EyW4UiueYt0bzk3WW0bB6lgVI+Yh7MP+Wc458iKBofzWYPRVXjxsZybPbqr2ogunpOm1SZLOjNmz
l/2wD7qeNMPtafSEL6NCmd1zHoUDVtPt2o+fsr338ZzoCpc8YX4ojQ4jJfgZ/N97c/lFpSdD8YJj
MiZuUvNhPogctMteV5q/IRS9X2ZQ/AldzAu5+SaQa6/K8QUfptqmFRyuA0vpzuneJwB6nLvDG8zr
V76d/CqLV5rtFornEZCjxo9W514ffuGSKxbUWm7ph1UmlTfQjy8J/n0tlGMHMoo0OxOAmJ8P3+Jh
/51/oMiLzR0/MHB9lxgntk+k3n2G0H1Z/IcBfZP5rewbV0AgJSYyAU5YPPf1g6rGij0Qt99Rk7Ve
4lM+Ihn2nTCd1SYEkTCyxoezy/Xbpsb+LozFjmZDYYGHcY5B368g4ZatVDbxpIyaCxPUzfqJWPkI
joYNTydMYY5TUPoNhqIY353DL6j9jh5CDZn30ekvN+ClUkjVryMJBSNMRO1XvgKyQAmLsfR8zG1/
uN6J1rl+ImT3SA7x72fnj2GF1YOnHpaXfnPLLX+OuwtJCKtdv30ZKgUiaYET/YjAwIBVwB8Ct/t/
S4r5S3tkZjrShrCneDfCP/x1bDIuPVQfWk9kyKbEpQbh7wtGUYOdatBo9QFZSga4PGU2jxUD9X1z
mlRKjFyJiXgPRz5z3GIBgdxAzb5wuwCtPB3UVF8RwP1eO9xxMLBwsc8o0FP7ut+xrImMHcOpXhlw
KFuqVsrlHqOXRTka9UJgbWWn2d4fXxcBdeG6dlsVIDT2JrVIZGHgu+gG8NXCjo42sBwn/BNDz6rI
fM0Wxv94yVOX2K5h+UqAL8aXOJEincNgEPXkdTUTyQlhBd8ldgaYRYnySWdW3RVCUoVRHUrfKPMc
i8h0/I7dsSyFoN1PiY1Bg52GeImOJWa+pFDMAr6Bu4pbsg8y1wKiEfHjIwpPNdBcubXNa1eGRz7w
oV2J7YTfR7nn1izRlMbj0nG3GKJ4U/kzrOzcCVKDgJ0jbVYGeIh7TZ3EfGsLCW4zyoEFXGUdHZgZ
OWgeF9tuZjuk+oh1ngLTx5D3X2Kdw/bD3DP9GAzMzB7eGe6wfTIO/WWO3tbRxM4r/FzbyYeW+OWo
cOH5yt2mGP26pgXGXegqrlRBKPXNjdAT043BzLSKggWdeIyoG3K8shBpwNmBN72OnaKzoNnSzaLX
y5Ttls1UsWUip/65Zlexcyv3cYkdGBmq3w6KxzbLpalG6VOOccGO24bsFAj6Ku9a0euPcSNeb4B/
HWBfV9ENyKv5JD1r1NMDhuvHVZ/NKl9ULk5HkPp8TSw9eiHbE5xpk8qSsKGRbhurAUGnfBtitTy0
4YhQLlaNqRp16ut9NM294r2cM6eJy5TFCXHq+1yYA+XR6Wv5IQ20YSrJP+xUYTKBkWFCK/URix3u
F/kNl2gZdTh0vNzJbxQLD3GNQLSz98ir1rUZThTHfQc8V6xzsnhoE3yRM4sHMxopXCluBOr4ACKG
Yb+7k462rwJ9JVDGZznDOtrzEwmZHaTH1942oKxlag1PGcbjOlRT0z7b08YvR92SY33qTcAlywWm
SGXGvTONkYre2dC2zzB9JUcEa7lz6rZJRhAxTU4Mf8mQXsDqYqAFjWEukJE8PjPhtMFni/abjPwm
XuYE0F9mUxFuw9Edmweo7iFkc2VylVXjphK+DRktrF8XuYP/lbvlcP9jvE6DOFRgZM0022hu0YFF
j1/4ViDOxugK/F58W88i22d78X4AvtxaCEmQ3SC4W1O8DWSFC2YiaMQAvby2oNiPFxzJvbQuHXr+
k1PTcGcskExnlFPvbNEWCTIxCgQECAo0hsXfOhf5yzjBfN4O0IrgWciCHgR6EwvqfDTwFBYO8gVI
tUPWYEqkzMmHtZQDHfonisxwLct7Jz2U6IsciBvS/Q/zjyUwdwAkSbsmI6Yi+1/hQmk9Li/UL8hD
8VCG+5TFMagJkpnXn3vkf9hPeL0Pvee4cX4KPTkV38hGJ+HLQdaVVdjMdv8xZ28/9/1b1w8pPGpc
aGyPf+8kMR/Yacp04W8fnR8LPgTDg5sSgfAlRqUrjOgy+0w+fyo9Z2mP70jXx9ZKbnjUeHrIoHhd
DH+7Lp+UfanLXNJYuAwI81rrFKfDgkcZN7Emn0XGa6poe5WVBAZFihguKvLGXLS7LX2ZGxuIObjK
vyO9FtEWVr5XLRyzHgAu/X9UiIKhMp43rJGKLSKMJ4wXQBM/HQkg4OwNAAhlcYJw7X3P4YibSFcb
a5A3iBz1QF98XsTpbnank9qLjY156WwC3CFt5FrW5jj4g8SlnEoU2rjsms/7AeuF6jm3lUoqr2Hh
18dMedQu539CmJp59ESDABcjdBDE8LczBsIikDZLEaKLn7vjKS3LoNzTASgZJLb1QVK23+VrGAoQ
NZ911sYQwF5nHZZcbOTQse6r3nC4eUdZ+11uDyfzoBybf2JGb6W8elbrFqW7uDjfvfFHkWP5RY41
4tXAR/YjFyEl0dLEsJ4rUGyPC+Va6A8pbLibTfIUJ9QZa1LspOVjGkzPUwi14I9AmhhADILWkfCN
e6DcAlX/xMf2Qh+Y0UZFrFa0qbRErJuWQ6CDLdY6+QAbufEH1gdB3VG2kAs2OwKhtX9xgDhSOAp2
uuLM5ponZORnsnkEJx49229ig3RZgI3kULFMB0YKLfJK32A7N6rvnM3WXJTsO34S+yhsGkbf1H8R
gbYnGP0O8yiAtUvpNxlEhqNjo8BAH8bDpo8GP+s2x5mdbu0Qa2v8C9Ohitk7Mvrqz5ezd9rgv2Bc
tG9BQS9jmaAo2pdeBcvoqJxaPkmLRrO5rreHoSyGXg436Fr55E64dfHZh5AKpMfYg5xr8b5palft
O8AmM8EtPiMkuUvW9v8L6WMnmUriXcKqaAf06QYCDadPkIAaVFrJsxvs35JWZU1OlMk/cPJoAssz
SKaQCPRzZMwanGv++B76tX9DYfOzH3YYGoTep44sN0jMnMYi9At8Q9XsSrs7yobzJfmi+5rBwnXh
bQWBcOUabxh8vXrwsh56SeUzpKtSm1Boo+lso4PHLJpQeZDKNs+3YqLxdV2DPUmY8nOmG1m5AHd4
6AqKf2yz5wBwFlyxhR4GWMUn/3z9OIQKHuJdChJqyL5oRORj4LXNUHNFB0pN3h/mn3oZ24H5YMb+
onjnXasIsg0mouKi0/Zy1UrZkEJZIa8v5FwLcR9DdY1vonR4LVZLzga4hbnWCXgjsjKUdIcVb8wb
9aNfhr04D1u5zXFddx3LXAxk9Fbi3NZ7Y+xCywaq7YH9VYUyle12QZDhLPSEGtRZhAAeyzrsypcN
wd6oFsYFGl3KWCqPlLMTE51Fa7D+JDrrzjfqeRpMdvfyBF60u1IKiaQw1mnB+4hwt+EN5dxncb4j
zZ8/sPMJgldOk0dCu0/5Etmy4O2o/jGsIRcieFg8WDrOhEcdsqceS1mNAjUWVF4mTLNqBi8Sz5PC
oAKYjbUaZXA1O5aeTN62jBg8nVeDoUR86d9DrbJ4W7g6sycD2YKR8tWt0yoWumCo+mhEm563yWr6
/yS7Ntw6jZuVzj3YbC+yWCe79Jn1Unq+VrmqdaCCQR2dV+VBPrZ6/zhazY8dfcgSHvsTTk+EwZQB
2kSE2NEEf00HJ92UxjAWXlMfPqrxvJnxHs0NJqzGIGYJ5g0yU1vWTYbCvwYwIClxC25iV1zJaU8i
SSc+DGxXhXR0OWu4EhWpfTqSQrs5wDevfk3K4u4EHTyUlcJ4hkazZAEx8US3xUaNcUyyXxp3sJXA
Mow3lSGZcPyJ1PRcVZ3qXoIKbq7e0ZN1PNuJymNN0fTKtGdKgxGz8SqX0LqD27fPVROwrMZDtG4K
+1ELdciuTHM664qDLQoVWIQnQKM+RFnpL/FvQz2H4kdSOGFqYIKpanhBVpIOFGWUKAvc2PFrgnkc
BY9ukChfic4X1N6g6FqYB/gF2HnjaKiY8BxfoQORbCfzqbx+15HPkDgggFl7UmZnzSx9VeF2d5qa
BwY6ZqYOap2oMCdaTF2W2TqHy1ej6bWywil3Qp32pk9L2YJDE8NOIoQb8mrZFVzGlZedPSmjd6If
ehFeW+Om+O4urwl9J8mBWi8pf57jzHdIFvpyOydATTGvz+NT+3uz9IaNl24UEPG0hWGZuFD9Uyfn
0j1J0e2mRHbZM9qAizJcG2NHh9fGmlDiDgwViTRUVtOXvRsPZQ+DLb2w4d4gFl7MKxOOOmWVhjsL
8yXFd3Oa5IU6Un8ywPESDGR/wi5MsyA0wyyU9w1K1qKRICNfEvOGMkMEzOmKF8YM0hpkBcs8TyYL
51K89QQ+zHF0CPEafYEoZteA2bbC54PRCKQgZdJ+O7Jh62rGZN8DQWB9zAf/r3oCoflFfWyZuLhf
4bwWOQDb8AuVsWfApp31RTWuWap9xpEFO3HrnjYESNYNG4BHLd5ZFI/smz7XtGkbXh/yfccJ6shu
EIMXvJaiyM8lv3keL4JIVNBZaHK6uAIDqj5bdLTyc5CsTOUhvaYZmlnovU6FGfDovrA5qn4P67Cj
+XkdhJZXRiSW7Hxh4rj/qz0OEGxl0IKoIMxiSD4J8LEy9bRS3erO7/vnHgO09NqoeExdgh6X8aNW
T7NQjQ57f6T4qI4IujwccFtXecv7HxGNjexpbO/q8vwxNgw+xSuWjLBO2qMYxJFElPcQIF5JycDD
deCgAV2CU9yHJvm+MD/tZV2iibJDe/k3b9LsYmGtyN3QqFWt9tLpwhqJ+DGC94wsORV1nSwh65Sh
d0G5+yNNYbQd70a/1MvsdtGH8SC9tZ2+vJrXoFwGQnKbAhRhZBYbV0ZBz3maOd7rhiCqJTndmbEF
tYWc58c3brjtSDH4dk6AYtLa1kaSkxMPVfLbsN1I0NEFYES0O1fHYR9p7NpiSGy6dsti4cEqMG47
JWBsiqAc1Gh7+H1DNlgmWP7gfu3s3TtkkSQQy1eaRrucuArg5vzWj3LQAaBtFF/4BVGT+WBQIS+B
njB/X7iovlc0/8QdSqFfOx0KDE4Q5y7dp0hprMAYx97MgnXGccNfFFEBzbPnZjDXocDwWc7W9a2K
BHNC436GXB+EG+D660j3DrXRa/oNBLX63OIz1F00PSZm3sgjNEAdE50Z6ZURu72zOyLFi10UO4Ni
GlQVADsoVjB+9eA993bNZIwj3EcHb+j7WNganRVQRsUYdLWE0lrVbjg5leS8saG+c2Ydd9DDEJea
98wSR5FgxcFH+W2TYGA3J8Yo4AgFpIR23YJDvkHflBfAlkE7P5juA9qfASu1jsaA3T8tSIcREiTj
TkaXTS0+VCjNkc2dZz7skBCtT88Na2ztoV0ZRUtlbk3MZ7msOreeuYS2LXSYFsZNlDy4WUIeH94I
szSmjlkg/cOTUiV91Hx31UQ5kHf4ycuX1EPNgF14d3220Hc2iIqOgImmwrYEHcam9apUoZpKJPxr
fFRcGRHVi4PXwVBh0gAbCSKhJD/jsvpe7t8rFKG+z0DXZVArzu8EsazLBEJefQix0HJ316Z0+T70
5R7aDZ6tqZOKF0dNYfpiB2S2NjkBu67C/98p3CrrvMfRpDACGJNjO60lcFuZs7T2797DBhV0ZsoQ
oQwuxsnGERn9aWkoW1Or2bY7X2akVeLWC0iDfLaA4k8vD00DaSqIcX/H9xdNqe3aP5UDIslZW6j0
c8tbHxSvQcu+jrPDERuUuSNUuswzGID8SWcMjNNC4Vv87K1DAS/L5n4vBf5pQ07FMpHes+jYqqdq
4td+3sjRXuWm0TnAoguUdpPBoDDAPmpUBiDXPamBc0vf4PNZpiRx/c7NjuONfLC90vtruhXUt4zT
NHUW7pT5G56bv2hbFYDeoOjKauK4ajKYcAKytDjHPuOzMJLlfhZkjBcLEcDBAy+P3aQcFMwER46c
hGzpnrA8wv5/ndYQQnoq+IEm+orL5bh3/bBlqzL8qpVoQsfnffGrhrzP5OJYT8ED2amKtzl0k9SF
8r7cBCqS7LpxqNOB1ChkNQU195+D/9jsFJWX6HpdGbJr1azFd/seW5cv1Y6JHkeSmLD5LlXX1V9Z
aVViY1P0bLr84WlpzxGsyQ7Gg4zcdr6HfCk4eGjgik3pgX+681VUpjP+hpyVDPFfpA+bvYrHh73H
CNmcum/gmh4X7zGA3bvk6k+Q6aGtspy2vdt+kOFh5mUqZsG9PoJ3Z9PHM7KiTNpDBO5q9lpPHN/X
40b4fAv+ln6/v/LyFx7OEHPwitcd7565vZgZJdrG+5B52G2OR+vJS2Fydj4aeFHZRJCYBz7wFA0Y
Y3HGkb3l7WdPAe0Fnrx5Agr9XosGoT2YXeLbk7F5x1Nd3a8nPC//pEZrkBOU8Vd+FB31TUf/J5Zg
OAaHURndPdYH3uhwILGWDoul932bJ2uPozKnbmJZM57CJiXmQKR38EbRxMazd01i8hBquie6+y54
iJ4V4h9F8RbQkLYpvdW/opskfrBFnXabv4kx7nsi/KJnjnL6C9ZNFCUbIsNC75uGDw0tt6V2Fcuk
9UmtSx3aUGoKJSSC0DgUwin2DDQflEcbodLqkGW6Oezor6y8Ps20r9Ja8w8lKakOfLex3OWmYIEe
TH4azoZ7Yjn1zZrZy4Vh4JZDn0NwsGVxImX5P1AYkQtEp8EIhWVNO3SqwJEJN5ZyTABzw7ob34kq
MKqIm7kKSbBiMB0bH/cZ58i1yq4ag4GaZyMw82Nqu/X/M0ORn6fgRr6gLvwecFZoZncOnNu5USLW
aeqhvQMsL+Pfa0k5IaxIbNyjEOm3xcy4Za4H+SifvqeO6yN4tiE0SzHp1J3yh6w/Uj97hSjK83CA
UBZkHjdMfNkybilRqhOBvUKSP8mlnrRX9IxDvQkOQRO9QjtACb6sYFKIsMy1byrMBZjh9BNQ6SHT
DHhAgQW6RP2Cupbr/PyNMnwDdHifqEpxANhyTjxThO7pmJdwAQy+pLMw4LORDFkPBw+0JR/gZT/6
MWr0HP+k5Y1LWfrzvUTt1aYr6i79zOpPpiFjD0GIKgMdRImzmG6WpG1pmcLAtf0jsiMqVKdGwIaR
jbvyDlCxOBF/Dho30Vo39/2jpFIuYjuI7WHGWFsppPDAschRv3r/gg6RGwCDQF5BGUbPYvpfBllN
j3lWoSerEG9ey3hmjh/e8h/fIgTDDAgY0qz58Q7lLd7fT7BmF5h7no9F7QtekZfD7z9WGC0qMM7F
RUkQSr0drQlQMLVUOPhf1fujXvdEs34GokK1cADQTiFLzx6IaMyvylS+i9a7FtnE1rx6mGoxegCz
5V1XvLRse+5mcN6mBRXKY9JinT8loyyWfs30h3al5BZj1aLkU8sQnEhind0j2SCvzDn2tS2FTJGM
jBu6BlYlwF4WD0xyjKo/otZSEA0oDiguwW4MpyThv+7iqgYuPRd+nOBKLCnhsI4roxshW+c5K4V1
FK5OBtJlw3WzeUduggJU/0X15Nkq89EXkqPWFcxrbXvkmpscdfmH+gMYTVPgU1V6kl2rhhhNaJnc
2leUDtl48kznUmx9/K/sAU6R1WAxIicbQ98hl7tOyGdVvtgsAzl2cLcLPU0Y+HXRM2dajbG0588p
V/4Jh6aItgHF79rwLyhEpEB7xnl1e01y6J9y05NRtwtCVJXm6iW8JxYOZiz/szqNMaOHnQbSMu4R
1tzCirryHgp+dZvo9CGdIpgbd4K4i5ETpPQClqLE2aNY8mAe2K/Z+UlC+ayqAqd9a0Vd2RyD3l75
H/4SaWk23w6XW4P9Fh8TH3Jtuatkkop1HXCgO0wiJvFPd/9PtjHPoVYCptid14C09T/lqjoN/D9g
9mfGJTVbp34CLS98hhQOO6LtWkJTW/aTVTcI2n8wACLWtHHgle+LSzHHrqw1wFR1w5+DwGP6WnBJ
QmvNG9i7bAw7s1Zbs4IRUrd4Ecj3Fe0il5bBqHQSRQBGmSc8ZFIsToeFTWrapegz4Tp2ECT93XFl
ut6RQurPF5F/2WfpAVxz9Ky17dmfz11OJRB/CYnAK8jFQ3CPNaA52JWhNxlkcASMeHYt0FBhOTUI
EE2LJYZXOClJLWSJrrrMQaNBEaYhfaJeFSZwffnXGsgqN0ONmNvhTys/lTwzUAv10tfRIlYjZDel
7LuRhXhDf0n9LYrsWD0/dS9smKVeSSqW3HShfvaoalNKyi5dSvA0uiZ/azaulIN6DR/nGsa+2r9y
DQ0i1ia1uAbaKI5lOpUWAdMkASnQVDp+RtdE6cK29l+zMmqImYO0XAHoTOrpKXljU45xa41ed3DE
sfJJvedQMErZ8I0K5xQqWcnVkgaj2mjo8WGn51JA1FcTPQHDdVHF1eByRNXNLqgMRXsdtHnaYS3B
ZrkB0Y1CAGrlvINBZ596rbOr2NIQNQYMJKmkPS/0Cr9NY2KzeqEpEkb18ixKHO4IHVDsQTO6FO3u
OCdQYVZ70gO5JKwkHfLQKoAvOgPqeFS0hj8IFn895ACyhO74guEajYH+8sLtiBldohgUxw9bRhSy
ieyyu8npWrd68vLNFUWX2zvpUohpiEdGyv3Xp5kHaM1U5eCJ77szCW7YJ76AntCRpADbtwPjtpKR
5tNWnk0LrJY6/nEnrE/70OpCqHRSnWQRyWr2Gi56qNUSVEJnlvG5gWwJCnsaV4OOPrf0A0aBz5Om
cWxSup02rBKiFOM7h3Ga/JIxhbjqDeDbbefit//6nD6WRp/GuTaVYn8LKbJkF4t3qaMLApoPnqw7
TbjRkFJwZAgUOi/cVWkx730L5HxDCj4C6E/ZnWN4HEMMPFII5dorWyc+QRxChUFeuyei8GJZnDwq
PHoTLCioja+4kwOgooAKz6W0YddRnFLi/YQpYkFXUvdFslsZLLECNVTXeSjWb+8t28BacijyaKEw
aQUfYz7BNgKr3PuzC4ATHHAU35ziHjsLa0fgNi2v/Iv7Y5iKlAPlwRtIvsBp5nurJp4jy0/qQGyp
GiqBT4YuPrB2vcyRwHzAWZGrCPc0VKOn6Cl+VoixP0my126Z2Rb/pq+15dBQdlkAqNABD7Z5NbQb
vJ7dbXfMU1LwwcZMKtfVSiJy8ny3yrO+N+HeeKzebht1hQHkmQgtMOcPlQasrXq2gPbc8xA0uwm2
HWzTbUVd9Uq5iDaKS9osaMSMYTv8++7dO8QWT9rjWzMq9zMGlg2ctUxsCGYxreVQPfn/y316ueUF
L1yJmkjGuZuEJnCgiPm11zLFtLa0lEzezA0Gr24JxLyG7AcNB4a26Ma1nQvwQQnTIT3vaTfgqEOO
M9FaheUVpm0PHIK2TVfdpTFuK+Ejnv1JAGxGH2dl9NiZagmkwPx40i2X0412Nz428BitYlhtrQy/
+61qcwAjap3pom3NsEPoVho2pO4XPEc8PugZxrf5GFr3uROxfqMycTqmhICKTZDf5cggyu7qmBIm
wbkGBwvAWVQFfAmjDvkV2xfT3XVdDuqilf1xZyO/z02ArBX/NenZYjJ49oo2qz4UV8U4HdBdKroV
lesgnnmkgYu+hBr+MgQAy/RR+ZUH9DNVKozhWHYqk+DLJ6JOicxI/Icy7zo9msLDK7/SHsPF+ake
nIRLnFOyz1cgwuy2zso2qM/CmVz+9uH6oz1hYVBi1RXq1ryUyoL9qZLG7iaNL0GxEcncF56RWldh
ACI0SHW+kO3JRzno26d4gBet5leTQfipD/GiWAquNOKs2uw0QTEGojnhVOdXCBZroWtCsvRQcp68
8iaqJFaHD5iV14V5DVsNqc35FQRrsyxnlANT3ulpyfm6D7iH1g12CJ6Mn9KQ+w+wCREUoVxT37gs
WEs5EH0fPF1d0VBWD19/ppKlDm0x2N+OIifaWACM+rU+aMCNejXmT2muBj6dULTN1Ez5yDW1SyU5
3HwaZua5IbGh6+wksj5AvIhwFpRrsdvJCZM8oZ1q18LfyHw+Qq+Z0E02O8At3weF0zscg4jWLBgS
/bgQelB4i47yDk8uXQh7sssvTHVYmDRDm8+23cq1FBeKOK6mZd38Zk8+AYKwr19YPUZn8Mf6SVuX
EPYUhQ2pbjR2eRfz408UTYIrQ4LjXHNI4qK9yHVcC6k2stp7Y6UUuwABUNF3sttBfu7Db+BMGifX
ILgiAPs52+l6CMQGFacG3Suq0gEHfTQXLu3ocM5varWdeJiATNCMb5bqlB5W5497xUD1Uvdf5NFM
XfgM4oWDOXsELRqaS0j3L6uFJ7ImtgrjMYP6fes8dHK7PIiMepPmZ0TXy5aPHf7n02jWkSwLa7LD
FyZSTjqA2lOEInIc2IkXygA899u3WAdAq4kbTJHIbsg7vwR02wU5vDbg3M3zT3jQwTqnG6ua+dZN
YC1pQr98TZnVN1d+a0e98kQYhSEfQhDhC8P5Y4TEEpfVl6jDbiU76q5iTQclfFxqwJpen13bMvsa
yNyAjyQSHIonv0rTDbJDlgSKRavtEl6euSjt7hC8y/VfnlZ02leLnk0p5qnBVevJaMbQ5g8vuGuz
B+D7ZSHvgN8KpeWDMeXbWk8Ib8lkNDj+Xhz0fYqMSZJq52CWlOYbgubx5P0PVL5HbAk5vNE/uxBv
iQFi0fUECfaYCVrASP9K4RUivpdnchb1EoYGSKHWTfQq2O4ZAb6sBdnRgqfGiBbPXuQG2YtLTGaP
yA6LQFPYF82o6Kx7bifRkuTl1iTuwuR4Vhnc/BX9qomc0aMG/V9gRLD096JNx7tHlW6a9DRhCFRL
Ra42BB31coC497frLnmbdr5ES0X/vPgefwB2UyHeX7XnW6fKarsT0CK6uqRopyav4EiM3WbuKCvt
iHy/cfuptReM+Btjti4MITpiV1eI5Zj6hxf6dpEVK1y4HxXgiqfUSt/dyi1CdGBxk7Bwfpa0oHXR
t+3tPWPXfxiV9MxyXw06e8WkPFh9dMhLzmZ545m34aY5jw7T0W0aOaAiauq/6p1CcaLkXN4peH1E
gt13FWZtUJTrbiQObWuL5uVI2Tw0eIiVvglZtAqsjIPjE4Y7XJq4M+EDYshiv+UbyrjOu/EfPPon
thIjPkSnEs+eEuAVPgZrCQupx9fWDiAUuhoByfGgeVi4UT/+B7nmN/y2fweOu4H9LpZXnjkDcsN1
HtqDLmEhv4F+aHoAON5wELWCTAJRfcJFr4ur0oSopMHHhf2z5CXJYEpKJChbMIu6pAY2ISTt2h08
EFwe03AwnOibPbhCqkJu8xvsNzgKcskqipAiPJRmzUOn/YTrjdA8oZzBViaqi6QnVkXO6V2p8UEN
VOqKddDeCdJx2HIQ+61sl5bUjh0W2x46kOTKmgbUY4tRs/RFozp1hl0VtSt3H8xxL2wR1ZpVE3OS
oEojl6KkVig76gd6NW3fTmKyUmDn6W/1UOBnXkXML8xnBnC+d4qc6EZtWEIkNEi5Qb9LBxvs5Ab0
8OihEQxEfDCfTVKrGcBFKT9iTpVXI8rs4NIjOFgtjKIaKREgeOb0aOEolI5W3tg3I54bmIFvT1IG
P3YgtEqpJnX0EJqlKyyO3TVrM/wCPVRrkAOu57JMk3C+SKSYeGahhWoeDwSZjwtm0CsZpCHBfHJW
ePCAx8V2KGhlqWxcTCngpVVrL0htn21acaOfY590fIKf15J6n7EOpHSTy5s8UEjpyih5omF2mlDT
/rhwPmbSU5gASvdTuAWQMh8wYrnbbNTuGrJSwA2WwVzFJSUeeP3d9Eg59JITrDrdXhTI8nt/RATX
Sfi5Oy8Gf+lPHExsXxbeTUhwZf0T3Cfgy9/AuPkVckdCi5bahswVUuOId8OnS1l4d5OokEyK9iTN
VCVO50v3vO5nrESzy4JpXRFCoiRe0cyExPGuf/NJ9pURI8gu/SKV6cM/UczyMVpUV0nWMqHFhkIT
UELk5oTAR3NhISZxyHKmT37MJvr4Q0RDGB2SoiwjqGjT8arsVdAY15Zs8kRgX2k/BZqwA/MucM8L
sSTyvPCsghJVvHanp3k4omc6y/FoFYeRC0hj1rJ7HMa6uSkI8nD+lOnd7IsZrIbEb2lb5MZpEw/G
n5mLVvIwQ7Vd7HMxElbbQ4M+AbYwXClAERUrYW1rK4Jwlk2EXVeZR6HYgusZsl6NUvLAbtJiS8Xn
ve3gO/Urunze/LO9L81yIjGQ6u6kgsx8b6Bs1p/gd3rILSZMqjfHedJfZTZzQseVFqPuNT39KoEb
+nDqORbGDElvlE1Z0wKk7Ewnvwr6HgRofSpE47Xoct4VuFuWhcdCBKwVCfGK4aFhBkmfCG1hpFrJ
CKvn/PEXBempqB67sUca9y5kafDcdcSz1s7OVfwfcGsQfH7k/iAGERiTtyrtRTXvP03jX12TjilF
QvI/wZFfPrVy+QCWJpvmMxzbRPvE4bR+x88DTGrp9A7jjTc2QpNJSG4QynPD4lZj1i3X72QIWKeU
yBx5Jf694ZoVqUC9UiC0KnMmiIAtOnFo+e8tl/RvXNIBN0/n/a6z2bkg0aMJOP+6mmVMVs+D/b89
Cz7LEv9/e/y5qiqv2pQBg10Z9jpxJ0z1bYOEY05HssqTB2hYZe2ByAmB81VgNqO3k6mlfC4FHIFi
Ym9tXgKPzp6c/buxFR1FlCDc/ns6GrjPEMDTrdUY69SPBYKNCoWwI6aWPycDmYk+2n1Ap6b2Iaor
9pGQharLBSch7BUxyN77lejS36tGu07rq6xLN4a1H/JPt+qyXcU0HQvsUy5uvlmHUCtQqKXdXnBQ
I1P6y1xYcMZ5/wjZSOWJ46QZvNE6x6UzKYXV0zHeBEAl4631j1Xj9IDx5ZhdJ/kFghke11mOZ5Ao
yg5cd5SyVzW2hcL7vqEI/Xa5kXG2eFuAAkhwqab9NW/hEgcVdAILpeXZju3h8usgqKGKB/uoAlVZ
eWWwIfmOrSwadkqgZ9ZQ32/1IzDjCiQLUrgBpayDDnvlRPo71WneZ+ydN+ehINFJBnvNXZPFMbIb
YsCPCDiGZEf3B5ODOqG7aU9t9cDVGKFugLwfPwzhi91SZejdd9K5VpLIkTi/quIoMTHFITSF6mB/
6uaLsErla8HJZ5D/pN0US3+6JvvPbPRd3U2OyPMSNtgk55RiRvrLiBiTUAcUV0Z1bd+C0Vinbh7C
fUkfFeiPoXhqxm54++e2hcykCNWMdByDq6MOQjyWRRHgycnY16nIkluUK4gl5wHdWLwLd6d+xisa
L2v+crPkI8F1lTgwNxVVab81XqJLabon5IHsJQuvd7z2wSzLLmphWIoML06J/EZgaIVkdGyAgZ2o
ThfY5ekZgXX8/iIKF/iD1p9Hvn8hheqw3FzXlbehpd2Lf3CSKLo8C5rbjT1iEEGVjqZneRLHAbgC
AxhWs3Dq5fu4uZ321oznGM4MsYJ37gr0PKUYc5oVhqtKi11RQ5Z9tQdhm8jY/wxQpnqUnW2PnBJU
R+q/Mc4fbaJKGIbtsCA7mAXnrDVfPVX3lHVazn8OogBuC3a/aOfLVi/M8cdHdFsmddCtU/iGRc/C
SYXJ2m5YL6Fx96N1hhGBPe8gX5JWeRLq3/2MpcYwgt9NLAOD+mb808eBTJqZj+Qi0egCKmNdcVzK
BnX5TR53zWz4kVlDonOrF11mzYEQNq9gQ6eE067xjn9tiT+JV2vJZJZHf5gQIVwLz5W3RvUnMtCm
xLs5mHxcFe2Cfnrj8cmqmrs9wb4JnKGawRoW14XniYCg4dP3buabQmUw3dCXpWJqJnyHUW/2OM5h
9zQGKzCccMYzLmL0KsDGsFcrlCAmOaOO1PI3ZbE7NKQ2SXP5XwVE3X8+T120/LCG9das/UTidAfD
ln/onzzyNQmm/VS6OutsIcmy/nLvr1t5JGddfP6ruuLmMaboCSdEk3eM/h7BKAEZK7GSUYXohpB8
2tvm7aTHBv7y8XosDXUaFfAP/IxZEaIeSk1iislDf3clXEe3dIs+u3ukCJndJrR/HBQt8jQAHGf7
vqw6NpKIn9bfOkU2IPfiQ+3k/8FADEUuGXsVzxmHLD9aGTCmrCkZsYqj4Y4jr43R1nkDJJy1dqlC
IpHn+0lT4ITlwnBfVIpSsunjwpOYeet5ul0WBMSRDIr3CDP+iJxq0wB87HMs2X92rtcDerhf3kY4
q+vKIKbkw386JK7Iu+qNrMj/C4f3ESf5+zMGG5I3PvSCaQAp3gOu5K1HMLZfgUXql6hK+LlM3/ux
9dp5i7RFj0zV8zlud1rtoODV9YZolSs65eMP0bLE3FwTNrWEu189Rz8pOsX89QE04sSl2b6OQ8gk
LiSf4G8uEQ55BhWddEoMHUrunDJwbUaKLprh6ByxT/GyS8katbnin1rJKQlJR/jims6RCaTczO9A
MlvOF1EjuINAStTysHmAm5nU/ZzxkjZH6CANt8qcDAAMVlVXHc89heSoDaOaKPF9wkhriCmjKzEv
wflR2Zpt1pB1m+XzjRhXZBANWl0sM2/e/rk44Bncn0PMvyymTMgT0yfNxV0GwKIb4dlHisW/hpxj
7jq6RgaPkPNvo/DS9nQocbO8uztzzBQPH+MTuPjaoiUsNMOqWLRSnTbpe5dGnP/O9akoDgEgH2ZI
A2+AJlMp4Xw/Ht11uL+PiMCvJ+Ugp/yIty2v7QpqG22W4GPNmiBGP6GlUK26HR+T3o3tenV+7c3k
FoaNHZ0dupsNjCOgXv7gxg8oc1XCHr1Ppbvj4jZFgqBUsYvQfwxhAb409/8wlfMLzqFuy2I6nwdC
IGktWYeO2YcNvZoVTZo24WAeoSTVRGLB+TbBCvDhyjgL2gHOCK2Wz97tC/740vKdm+nMlVO6e/Q7
xAyOBlGoAxxCetZoUaf9ATpbjVsgbVYZPOgKMWHZeFiFgSCLdsbU3QGpKHOHGZR9tSNdwQx8fgPR
6qoWjlgrWcEq+HFX7HsauiTerf3L07vh8udsjOVJAwXt9o80Sw+uBcjXNd6iVfcQlU+ZKPwS1s2L
Qnccry1lw4QDyD29LLx1xsPBxUCfK8HBrXQ8Zwbcuf6BLr3itJoQQWE3vZxm4Y2Hr46mjknIktI6
J3/MuLmAcKMZvGDMrfBtjLO/iZaX/ZDvdhQ3r+TWC3NxucuxqrZ0rhz6J5AlvUxOY7myJDpbYJS7
WkXu3CyWzhZsZcay/gcLMWv9LJQA2SgC+SaF1MqxwpKxgwY50k9fG3ThAhcDiG3xj6yY3jiXLfx4
c1dDEt7X6f4muClB7rOl1eu+/2+qEAbixbqmUl6UU8Qj5uu0j9AqEO9Ci/J56WZqu1Ikqik1fwnL
9dicyPaVfWwoos6soen1s2qPDehztfibhSjx/JuURff/6jONbkkUdYU421lbzOnXIQuC2yMHHewW
H/n4znMG8eNzUfkVo1kxV/FzOf6jnq56eCUqfKv9opmW/lgvgU2aWPp9Lz5mWQGxF4/sUlNiM7oG
JeA5357/iz8I3TmwXkKP3K9361gECMt1tGRegq54eqi7cXtcVNEO9Pmv0uAID83lSWj8mJWVjTyx
0Ku0IN43r3m12XwRtIrEO18BiVtsf6LS04H3xP2d5HHssIYmSNzGzLbowR7I57Q3UVaGoFtdMLg5
4FtaIIuUEop9XIYkbCtE3pm2BqYgGBy9Umy7KlKsFxBLeea1IC5jUprL1c0FwE+HvprZSIViZy8l
eqZpKTc9xhopv77tub1VG+hLEPc9Ct7h0mPADG/IyTkfVqMIsCTfbkAHZxHcL2MEBWOF37iWBCA4
+/tHRvHnMg1Rocz2G2Jj2OfQ+UNMH4c8XmhHKRbukjsIcDyU46BF5WKtQiVGPmEveqHU5DVsrhNK
2EwwsPFe53xK22r5DJDyc/tHUFSHpA1WyLa/vvpx0rFneDtiR7TL7p5kD2mixUaiHm7MGyt8tQyF
B3vn9lQFRqd8lABhwMN9q+9F/GqE3W4otT2c5Z1wh3CrZOWRkRlaT8xqCBCq6USe3zGkgYZAeuva
W9g+2Rr+bTdGueq2H7xmVkGvPhQfwayiUGP7bqdc6VUyLwX26lEX2CTex/tNbRHWQdbcQg/+D2UH
T7CPDPBx8YeVfspAuxxweT33ywxxu44bZFgii++i55Tpk9rXfdhdrlQdm6/RN4ZZQZ1BGT7yYJcE
2ogd40uvn0rjGDVEoKsvBKluQCbOvlACz2x39Id5dyh2k8vytRB1ZLFxVPwzVR00suupYlZjByo/
/mXrZJwBqqL43PAfvDxDoclOD1tPd9dm/LTkJmvcQUsKR38Cjip0EvuCkWorf9fFAB04fOKjQcAz
uSlAZNCmL1ER7+SZ+lm4a9wZy9ub8qBka+VYM8XcPXUtZVd9n4pnT17G9Pi/rIhZjjR6ghmyYh1k
4wVd+4pkuPWy1joZ35s4jpazzPoPDUbIvJk01kPv+scyJhHigDjpzjCV67euTcAlYa5OmR9kz4ba
i8hHe44dn0O6LqHXvGfo0ZmphAgf1lQ8eR+vvlNinmkJBAQyAdd/J6q3MG5SjtIL03Dq87qQcChX
sYNVo31/agB/5fVVMcQJYQymiy4evyGTSh3M4qJwXebKuhkJtJowIHsGzFctmdMgE8ehtdsOprlb
a3fwykf4XSK55FiW4I7fHDFTGZfD1cBxVnrEumrg68/SDtHczM3kbHA2Uf/I/Powf+JRXh2C83Jm
nHHfFqtI5NoIKiqqLN1NJudtD4T3VwxwieveHmLyNnmn2KUJg8tcoHgOVcZZ8gZn/shig08bwjkE
5SAql5aWyAP7IKvWLEvXh8w34o9Itm9qMjU92MQFCiUJdPcle8un02qWDbD0GF3OG2yFlQ4usp5H
3zeizS4lcXySQOOdbKbmMQ9zo81PrvPPXPOdkFMct0aAhSiM/IFVNdNqzNbSMAvryyth2TPhMrMw
DDSRZhVjpV2/31Pj8AAgFQBslYmKMj53J0cEdlii1erwsWsSB7892BK0opIYdxcDwInmoPingU4x
Qvfz0PXwC/BgBXWiNldEg4y0vV5idNjvo0gpIFYL1dBG3nncfJqcW4RbkFr31Wd5avz7KcQCGgvk
fi1+WXz6T8Co1YzAOyCvKP1O8rQCQEpJq/v3HOY4T5pGJdhQr0MOFMpCL1pqYMIPJtFzQwiJ2s35
81P2p9EUPLtEJGuLUFNhwFryeGD34Fu4IdB0RZRdWj6pT2uVJJw3Nq490wNo6AMQ5YCXnDmL0nX+
afFIKTkqmbDKkLZYO6BeOM+emhuBSv8mpLRGFUMnxwL1FQJAly6wAvGFnJ6gsp3hR7vaIBoJmyc6
v47/xaDaP/OSQd4pvlkJjAPAQ7I1byvKKoGIXgDXq+IyHk6S1s5iQhM2ccvMIMj+6AMxl78tRicG
k2mUeWrCCgSDqqHkay8eSQJK3NMgNqkdyeF2Sefl7jsIGi5YXvRpnEivwZ+f3obgdQKo1woVWQDC
3yFOR7N09XC1Gc8gU5VB5HF5MmgT99o6hE4mvT4b+tiCob7VTJnBOzTc6E89+uNExl6xozH72SmI
jIFU/Nzm0qy/rFiR9+PPjrOPlDHYWOw+GCG004mclNSpAKn/aCAPl35emmS/BmFKkV/1cGcD4P6C
l4tzXvJyu8ipaO9L6onhsFbrJvSB6wUuu9LwM+Ei28xnJQBjefvM8jbrEkg/JG42fikntXMzlQex
8hH2Ls6IgkFxcjQlbNfmFGlP6JMU/uq7LuH8Xl7hDQhLzpCmqB0sevSKPh7+pXZP8mMehz7XyRVD
y713Jf5YUmKhlJUuuq93NzDaYZgbQNnymDljyrRnthS6PBOtWrKhZ6penZevMQ8Ujg14I6K4+JK3
oQx2v+VNVIYIDIzuYCK79m8IGOGDir+rJHnDpTH3fgygcqor90opePPrnEPRdXMRvO/2AY3gJuLV
k4NCjW9aPxm24AU6UmRO+ls6le57yPlug8gWwW2J6gNWuPS0oM3xT7aYDYFWJMnOQtxyNUWMJm22
VeQTVs49MmJF5YCHS3MxndKSZkOm91elYhAQW+2CD1IA0v/DJbO2fqMywMnoir79vt20ZzToK4pb
jxlyos/CAetex6Qaa+KDD+h0X30NQ4WBjKxmIJSjmFvlIFJ77mNTEizPrp9/i2yPWAAfLOVsxBJk
SztVGzk0hwQQsxIw1NonXv/jh0KlZKVpfGgfnHTpE/NPPCI557R3qN12ybGgyRKTr6lYceHhGJ6p
l3P2sZqmkMosFYOEfS2XWpJwFgIDSw+ZPMXcqX8yv0wXW9jMLAmHY4b7nQCKzAEC6AmIBCub1tx7
ng4romlJ2UuI0b8kMKqpG6f445LxP2J9H41q0InPglgMjWka/9rp4EMFqzkSTIJCOPsZ4Uh1cT08
pKHQI68HkX85q6AuwiFRqLvOV7qqMzpjoJ9K1sRJYzQH5C+iv2xtyrXv8n8WUdWvU6QLeC6jPLvN
DK9KMSjontDnzXfY9I31MS/lL4wd4DXKfuaVdKbZZpJlX5soZgU736huWeH90TAyCEuG1a5O7p7V
goM5RNbhyVffaOSvLc3COskWa8oaNKu1YqYInz90JhMt0g8zKIgNPNa197ID1xGDUvX2vsAGX4en
g8cuwun3RUsDN8UDa6POdE/E4gd2mXTuEdAyrSRdbwJ27ELGc7RUM45PTMn/KhaxyWWMqHY7DZjt
kKUz6Wk7sXKLx/J+DDY9Ocg9rMPpR4grfuECY8ACLNc2maOxX6IpHEAzRIF56i/aWk1Jorvfo9pi
XkSTDjmsILaZohR6kcdhLJaDsxLgKGXNwjBfDnVzC4rrdHEamcw9jrAKF1EfYOZSK8B+PRQBxDEH
OM8fKWQbKrg9p/G1Ej8hA8hnyVcF8GfXFYIYED1JTVxGp5JCUHNzq6pFsWrSV4Ygaf/Vj7caQ9nV
o8XfE593srCN5C5nSXAGCvpJ1gattHlazqWeBNgPPYP5uuknNNFrjFHwwwQec7XueD4ZAdltrCNq
TEgnYdljBmPuU7UrmHz5S/RhKgC5mOm14b1YWD7P4gYceFR9N3cSFbXGjZGkhoiNzRMJ/NSqawLz
d8DGuyqEYFo9CRxEBw4EdmOQ1VoooFfISUfp5U5PHvOcMErEkZzdo9Sba2Eyy6EgyND8JIXc2rLC
S8jzvzlaTaI6PfftY6gqA6zJSgRKvEXZzrEpzrbz5VW8nRBNlQtg34P3KzPYuP+oZTOIv/3P5/Ut
rbo8VUKStJ3gCaWWdKihWqI6sTZfNEsvB2HkRxtSq7ikOR8wNYvojPwU349STZuvHd0Ks3iQTVrj
Jmpw/znH1gtYu6Lto9ltGmEQACld2qYpCPxvIxd45PxJSDEdLi46l+6nq3uFNt3ujtOWr0/oCsuj
pCwhulyCGscKDpIF3s3ZswgVlKFMXrg71ZISZf5/AuLGm698WU3KkKaGsFjS3gJqvBYnzgA7DF4J
3Lhlv6DiilBhKJ7rGQYOiOqeIBXoNm2eqlCsCK171kWBVCdOa7oDZw6pZPThvZjWUOf0bDwoxcn/
ch3bglJwX/ZLQsglHTANm/SoQodfQZK6VDJ/JFygS5IgFad3/OD7ICu2IpXLZ2RzA/5uGhNE+yPl
WxUBAWxBq4AnaHBjyyOI1Pu64PQqaU5ljfmcXu0iQG9Ym3MQifruvVndle4qWSNouytHmgW2AsVb
gTthVFlgNJnYtjS75PV6isvDNxBVTTo7MrBQsUuOXiiTlqk2JSaSfrM/6IEV5K1TCi8fHdHRHnmq
18H4oOQ/Z2pfa48eMcyIhDuAwwoVTCeR12GEnRvy9AFMuTo4uomy52+t1IyihBryL7lGwyo6k76R
I6WIqHgteIy4tVqkgf3euQz6ZW5jR8c6m2EFvPvf8oG8UY19oh94khw25ECMWPq3Zf8pXJbNrb//
xkNuM7EDO2vRHCRIzTRTAJBPWEc+GLwZ/B1LpKpRR7Wi83mxDHR08z6GaKPyQvLLKz3wb1PbMLoj
jBgpWcxiv0vZvza16j0Rj797R+iSDkWWpi7lRgEJ0z2Qojrnd1nGc7FyjFAtoxcumojGhZfetSfZ
NVnEpox759yDXRIIIIot1CPEiWsvyXBu0oNlD2Tlv1zwbt5SLjyIPQRR1j5ExDLC1S7ESYBKuv29
0Om3JyfKv9YBPsrvIFLsgkMvJdW6u7jZBhQ/Aj6HxHJ0o1Dh6VePv56HwCVuzvJSwbnxKRhsNOgF
KeuS1q8q6ik/ah4sQ4RnZWOdYnIJb8VEuhYqS9uh/2cik7H/cWHCwnqdnoTnai2PxcVhhsWFkyUv
MIwaXEB4SHI+dLYf7FPgDRUH+0jD/Xt9+djNACm9SeNWeVOANEq2F02KPSinaGu0777qsD/L4tT9
YANJlD5V3ZZwas09FGByfWjg1NiwQQBP9a5W37XwJMoQ2ytwYSVlVBBWB5+hikVS5tmDyvX48B+3
b9rEN4Ep0m7aU3BESD/jnldFDGA7py4sEGjM39Mpyn4ylWjLzMV+9SjebWAiTAxxK8Xxqo1qUaan
ZzsA4TJ+wQk33xCaFA6GcZyVrQMq7Xe2/vFDSQtCJ3iggHerpk0HhaqB8w9ntTtbukLdOaWEFFSo
Ij5qal6HoQNOL4BKvQvgFwtdZqmAuZwWz1/i2Yh6unq8OqhKy9m0cQnBBrRuZwFqk6pUFWNoPv7r
onos1wjYry7onqmy0YOY779jNyPmFDWPDIFVVbajoxFflGXyWYYdXdz8kIRMM16UQO9K5Doi8miS
JvzIUq+frB2xrgnS+mN5h+gza4pysDdO7m1tB0OBuuO94MXYIkYI2blsHUKIYqkgfSc7jAo0i5r+
G6y9aID3WypdN1CN8O6/7tvdz34QZ5XdCqabDVoaY5EN/YTZdwatEbPU8+++fj3dycwlRV/rDba5
4JVZo1bOunrA2PxwDtcLyA8OtgX4oJ9oOqMZ4J6UgcvpM0GR255LYX8rnHV/VKoJ2nX3x08Ma9Lt
oUzO5XH46+cpLoYGvHBRrv6vIAhqIfGaO2YShSo8oeLtONPmo0DeRCbebknBzz/RgccOnZwh38bx
zwqLDSCkqwzdIJJfbcb3xz9BcvjUK5xD1PpRl9uG2pvPcYS+Qnt7m43bLQ4nWk/uc/MubbgNLRXG
nS9hopputK4UGQwDwLuwPh8gHSQXInzmgMb+IyQzlzneYh1bAtkOGBKYLuF7+b8AGMZinhU4i8Hu
GnsNzjmn/BY0uPv1ZS8hNYeIX0KHXqAQb1gcXMwsYbi2llp7HUBQIlq8PapX223ZFj8TFP41FqEJ
gaWrMaIM+EsQQ5UFOd8Scz/dhANOwgaiBzdWDmeR5SaHaCWrFSqn1YxUq/i8O+arzF51wYBwgWfW
aOjaHjfrKsvNVqGNIMk2liGeQxZe8sx307K8ghGYsoFphh6YrV7W6bLq4auXrfz8a3x6z16PJ7TC
jfpp1gsCAhxkTxTJebGt/kdhH1QttUQVYpnHiwzETp6ZPB/c+93XmlLqdAXYtv2vJMoku/qQb0Lp
OO6hSG8j2sZliLxlda3SxgQpYyjqHWgkPGq5bQHti5Ww7RgFYVgWYbfeECBANTR9Xa4MomHTGqQv
NrPmdttfE3mHgD1X3hLsujmv00/YeOlb5veh0i7ProH7OqasspcwkzjLeXi5cYIor5APa/nX7bL8
VK9k4hizCTA6UPIu6va9p6bxFHt/Vb2vN477T4WGHk1+TqhVvT3NO/V5ZJiFxLt89N2033V2hQMU
QjoLm1g1KmpOUMiLQenBSjUJOdhKM3d53yqEifhVVxN3YbW9wUy/vK8pg5sPLJMCGqmSoXmVpEP2
r0n5EJFcu4uOs9epxoRPpnvidIRVHm4T644Bw3Mav72AS2aTMbcERNDY9PQu/SRv1Sn9+VKgQQQc
jguPuWwo02DXJUKTsA5kqPY9rDlaD2Bg7+i0+4fwKHWMFKG7ywHAq1utAGahmrKEOnnG/OPLMMdI
tnQYrbr8+qEPnKxICjtP/xAGcKXDwVqsPtHtshlf51ReiF+tFwVB3KWetCRN/0GfElvN/xr78YtW
nWLzBrabgXnyQPDBdtgDkVna6O1vtvSgGKXBnxsnB0hLWy11yvN8qJfR3DClzOGOmC61lIp855CC
9fTk1QZAgdUZccqET+gj2b5xuk8PIMgHnjwo+zTCZ2iqE0UdS4R/ek7tfGvPFecwEnYdpAgZorLi
cj+ugj5cMHMyZhaU5jCfuPsI6j3bGInzFYP8jxuGfkHrnVfqzXibhRMmbCSOCLFfkJC+bVcwNSXJ
h/3NX4G99294HqTIW9HPaO5AB+Gd4bdMawWTUhYVbMRLQLxZVni1UiWpcSF/gkxFMue465WfWTwM
FU/qL9EKq+x4Nbv2EDzUEyCDOWq5jYb2GImQliYA0pl+VjG0raqJgcDVTIHEfpxZr0/9O3lpwTch
4SJQza2r58uvuk6OaqhuiYdkaK3VKSEJqerokZsR/EX4Knm5FsltFJbK7CZNZdUh40eSKxA9C0Fu
n2XCk4iebf64GI9YU1zRghisn5SrP2RYkDzrJ5agujnbad4oYENUzePNocRdxYF03rWiNXVizEoR
OnTNE6t6geOy8bgePak3D1Cn73NGXUN+8/09+4+H0GlHtZapebPoHhorNcjv83P2kaaUrL0/378P
1EdZBsYYjcBZN06ZFpxEBdmFKi2y0YOgmd9RluJF/WbFTe+/W1tcBhIb3SXwp5NuhuMrNtHSlzj/
U2SiWchDhZX7AxKjm2K1YSWdJ4be/seL0IB6dBpsgi5A3uYy9jMuqaI4HQ+IR9AzwiPMf2KXhIkK
131dYpVMKUSiA84Qr01yBqakYuyV17FyY8u6IsurC3czpPp2A6dOYTqaEukQnhdrkNsVOQsw4XGT
VnsVui89GUdtNyLgqk/JLOp/Visa4rggaa14smszMo5FkH8m2UQbZ0mJ4GsMF6z6pcJ85AqBkQkt
aMxXr0EW+ZXOskrG6p1R2DhmHimLYaPvsTJS1Co9/xAV17zLnlSxivWIfK2QZHCw4DjVbms59KjC
CcW/UjLN34fRf1gT4o0ZGNjYag3+eXEiw7whS1pg2/feaB19Ac4WF6y+UWacyFjbLonZeFAqikez
awIVwjdsEC9Qd6hoOdJxqmg9MzKWY/CDC5nABQD6M4qotbajb8p9H00fausACwQjkETYpPaU7Lo8
fwXHLnKmO7qY0lVZK7Kb0LMnGMxlMaCs3J5cLWSRj9LnFzsSLE5SoVnyDwYf/CznEBRki31GAMHo
Y1sjxxxj/Ly0C7Mq+/rCgDw9ZWNdmr9DbamqHzS6CBZe7dNtV23NiX6xl9tiw2eb1oz4c2+MhJYN
Gn/dVDHm3uHL+EmHfucTwEtFtlCre6iZ+mA/u91hYQn0VmuINafoQRqcktQe2/G67Jj/yY82YY1z
91uIc4khqDL3qiV9kjKUdhXEjjlO2dddpYNW+AkaQqOHG98FtSazQQtYKBa1mwEssJTUvcod5RXr
gxkw3bzWs9LLDk78nT7QvCajA1+gnE10eD8Tga2xQBxeK7nNNo0T/t1VnWQ6NrjKN6H82mC3WJ0f
xb6y4KLBQwnb7ZaidSUPnuAqu6UCFSEpfMuB9xzV1UrSZmEeVzJcHXyvZosUSMZTSSXgamP22yTY
qBx17BmDD8TFiemaLizkBUNl62NcCV6kqwkGhzY5oZ/5edQ31vicFE0ZYGuvdzn/vB+K8I1958vo
prh+Us3WUbDxz4e+e9aQ867n+UATQPbr43AeL7MqQV1XnonX6vWugHu9B8VPTViNuv9xhWUqCFR2
PKw0LtKfEbgNAJGKXqt0BB6xFC6XQ2SB0zqbrQ5jUga/OmJpEZIVDtPty+EunplUHc2I7ychMRP0
xTuG3BfhG+kIItMzF5QtPccpJkGIFPnOCYFClkZMDkd6+H1MibO1GHNXYg7mCmB+uyVe9rc8Qsii
Gc3FJluUTjGKY5qckjqCKuOS9wEAbpuMhmCXWW1+RmjUHdm1kHPu4pB6o2JH0QPhaO7RWTRQdSrC
dQxG0k00BWiCqQeL0hIyxf+86NGKuljJOmYajOljI4Lsbb/u7SVH1w9wY+k/KH2CdYjFg9713q6t
Qb75DfA4k6Z5zpY0xAHAnVVNAQblmiHBa/k6dfG7Y/pDXkWnQSXWRx84PCtZsbOiqN+9yB40Hqs3
MlM8EODKPPTssorE5eVba/MTjb5Hm52uO5ybmXg9l1V2tNYCx2K37pajk3Mp6sdMm7VHkeqZvi1g
1693roEA79f3O63baC0ohKRbt+k5jTsCEIJ2f1g15SAO402R+wFokBxoeK0yVRqMlRMZWp+ddDOe
NUTkr3U7pP7k2gEU+tJIxUcwptWTNWeem29VAaPd6bjnb0EsK67VOMtQnYo6MmmYfI/hdIPZ9Eeb
BTOZ3Xnz6jX5HAcGDXeKuh+e9eI2pFf/qKbLrnx/m+3Odl+BIlzaKpjeOs8bjPYRQofm63U716M0
G/9jGN73gdNJdoubLNzEpCchORigRi2DPTxVehjAZ94xkoC2wz1gbdhn+hTIylCM0Fg5Fyxzebzz
zClz+BEhPs2s8Q4lqwJfKD6GTvnJiUmu9UDtEYWYsz+HV+8Lsf42182cOKCOguNVYeXlApbiOMvq
EDTMlBFjCg+N6P8JkP1WPmNKVrB7KCPmwMANPlvnHcadvEn37fNempJglI+9gErWUHqx9JkW/XNg
fFnGmsKIaJehp9IfynopxHmbCSaKHDItypU9IBUxS3imNy+RkWEh3N2WdJ8ojCYU3+DWQpgNgPO7
mtjVeaZVRsL+9lMEHR4M40c3MmT4JG8ymkT9Lb/G/gXooiJu9qWByudpNj2dEg9Ij71WszwmAIzm
o7DVkP0r0dnH+faSPSXTfx+MWUNph3eepauR/oVoDTnV1r4zmcYwsW3brfBiD9qNRIcfNrP66dgP
nF79b1qHvH3EnCh7JGscy3NzId4v24ahxYaKc1pZEELxzdjPpnHKQKp7ksSwfbD9XAaK0NHmBhiJ
m0nl0pW3bT8GGoyqIBw2KKPVzy0333qVdwm0/HmFjm5A/oMgVfPbursQypXd0XjtyQWGSLqzNQIZ
81FweZGyZq09/ChxnyB1JUkLz6oZbBseTnj+hhMKzBjzbmh28Go700dLYiXBnSKlMCMvBy9lQB2w
q0JgniWqWxRkekLJaIKOf33RSwcWwz4GRJuB7Mqh324ASH424jmh91vVFH/tGAzgYL8KDwSBKBFV
5DLINGwqwO7CgERnUpARN6SMAkDeepVVhgSAsLn/qBs1b4L1FLRh0RU231EEvTAoihyY+TFzSdmq
Qa3J7hsGVBe8Bn3ZyirWF9tj+Ojlugng59a/34fRlZTP3ZGvb19zN+NpT7dqZG97WhKQX7pn+4cM
9nqc7IlSNOmcPAvB38SN4cZTu7Iz43RJX1QYQWgbCTy+CEd/YVwBiVngrlqRmFUIsvyG3KC3+lqE
rmbYRgfffkG2/kry4QdvpgEmg0ReCFlSX83J421odTBsXq7m4lHztAc1I85A/bIl4ok+oa3OtgGD
R42D6H1aMijdsf+fT7ppMOw48Tzs5CUR70a34sB5MkzGbMYaq2ktp8LJB2TTiuvAjFhkFm5fQc9I
dkVcWi97ZO9enydnZyE19dY8HlTpvRVGB5f+gj3SnQOen+gZq3o/18mj/k2XvYH3pGIvKM5EjH1q
vZYZ578A7hPU/UwJbBrVZ7OLzxE2a1uWj0ErqmZqAbuo4eM2gI4aqYkMHM6mkSSsKxi+jjl/4ZvD
0YqnE/v68iABuxaQZXsSc5RQr/pd/Pn3kZM1k8TCE2k7Al4/ZPDsjFsVrZxFAL+m8wRVihIoieH+
R7GnM3m5HgEqUoIjSVEC5oKkdzxJDt/jsNHlPLiBvdiNM5sbbaXkfn0HXoZeIW91Ct1pRg3Lqh98
Zx3zYX0MdhdSJjNzmdnQyt3pTEaqMH3PuXnznS9ptQsGB2astpvaxyeLgWVI9eQCijZj+Avb2Eu2
uCk9iA3Xjom+x8prpqur5RhG1VXiO1RVqX7gnVZ8N85lJJCgI5t1zghkcwCmkJEwsswIeOIqwdcU
jtdXUBs9Arg6QsrUwb8OC1SAPp5Gpl5zZ4FnEji2EGPaOj/50cWWRomYU93S6bO4JsB4lIIqPIpM
hWYlgj2xlN9aa4DVYQ0FU5RZIe74FWV9GiTDnXueZOjuOVLjIkQ27VcbdQhe6ogwnZQHG3+xT8E1
7lZxQjXVnxSw/kz6HW3vb6t7MV0NScP0bX8VSIpqwxu3Esd2F3dYGVHqI6ySP/hURAR/766yB88t
Gkx4F19+tNLAgw8VnhLg6jRe5sYHXorjIiCWOstvG/Vqz75IT1CwSXDGAeMHKMjcmtSxJLUM8DXn
60swxqwNgjUBqGDRbCFUZ7Qgue52lZ3ykban7yEAIHWpgLv/4/TWQhqhNmHPzli+Z1GQWE255WGN
W9Jzf8yA2iG2xaMlL9Rv5/3GXJcRcB/alTk8Tfr8VMnpd/JiCczsDm/ZeFsG9yGy43uTNfZQomHc
2YuJu54WbJFrESjWqEybFH1atDAmpb2YaoniZTaalmTqoELG5exo4riZ2rYw3SXYnmrxYCud7LqJ
0WzcSxL9ROrTfT+UHKc5mRPmEGYVjymCon5uZ8EauCOo8sEyG7b/7SM1rEKqUWCXHPiDlUQEUC1t
aBOUZ/ponMb6lBbbdKKq+dXW6Ij9qa3HWFD/4aI4k4HWdhoLkNSruqfzpvGqFQI1hmXFrsfF6sCX
g0qW8jiAO1RWymECClGNVmemDG+sOT+usszSjd+sLbWsbGBe5w0oBFl5Z9gEKB1qJmApeyABhAwC
Ww5TZ1RYsfwyE3P/4dvF63Au+o/9mVJsoWXUhgFiD9ALHyVTDVVws1m7yy2IroTfmPl0NNfUjymb
iWmtVhsSh71EWlnhdR6zdOJjN6hxv377Vta9wh3Ti0TVKsEuNAnQQHHL7SFTOSx7hImtQ0/W/F0J
fX2uqrz3n39GB78An+dXoQ7HMibblWtzfW/OtGSlsO3HBrFD5W8qQmsyUCo7oIM+hbODRrVaqVJj
vz2pgrboZclZavd01kK2XKyG9P5Fz6SYOca7NRBMsyumtctUDurFk26vazXXkoL/5cQQjKJuI+3H
bp1oJo60xhJDRUOxkJ5xQtuL3Q2F199ZtbEM9ChhfDc64+lDShtQ8XJhR6YoxWBI7K9GBkybXGTN
bQa/5xLxX3mA7+hxEiFAXZznHeCVzojX4zgfpnxyh+BUIOM9QRqXCVp7MQdcubz9xDGMDI0ltjAT
xaU557ZSm2TdcPIIAaEmix7R0bx/jnQFv4gSswR/tjVfNEW9pFTcl74ZmhpIuxQVsDr2zxScXihi
+cl+LfAT3WME0q4CuezOoidIw2F5JDPPSA/jWXelIsVaNmNo7v2+RgzQIHJjyZWgxazBAgS5bKA8
hNrYF1lHw+oCqwwp30Q41tnY1IxqVEkHxr9DIqKnix0RE4wBuf8wIvQfBuq+itOpBoJjSZ8dLn4a
dMB6L9rLftsA+jP1COQgCy1lPG8ovn0eAYuMRY0fUozF1cTmcpkdJtwgmTBSZRtNoWpSS4GsQrMe
JJWK4gwYfe+JGG2pBd6JIShaA5AEORPmpf5T/0UqQDwmmaM2msVAWG1xTssGkbWUlfRXzsP0BWxV
VySMZO+boX27G+8tw0wiRZH8hb5SqzdL30b1BIac/ZcqHx022GoNHvqA5PonXO0LXE9/GGOsr5vD
VbhV4ZKnuthxRRzZ1FpdPVsPkSW+B/KQOh0wDQJXi/srJSZy1hT5TjFtIK1lerNzKQ22TrNNmXld
IRDSXuGDEEdeCzKh6Ek57g8v/jrHL6+0swl5X1YaWoAIoO2BxDT798oHOSoCeEolxqgLC+tqAJ+K
DkH5RlmVgYZbizwIh2TE5GCqoFOYsrxegmi3HP0TgHX5L+DPXWQDE/g9tgS9/3WcK8mJdvpW/pNR
z6KkIprRwscSC+nhojQh8dqyRNOICTZPkLlf7KSaWwdGu2IucbQNIN+LkfRsmhwpXbFUIKdXs8Hq
kwFZ7J2kDgdC+GYN11QRd5Mxy39UUrKO+8KvdJDF/rXySfKyJegv/wOfFgeXLAiYEFjJzUoaeyK2
P1/NnkbIfWWo4R4jGG1bpaiY39d+jsryWNPxz7qozI4yEpn3TUrq8TSwdu4kcXXWBHy59xOcEMWJ
OmU+FjTbitBbukpo51lsg8BD1E6adjsrOfzfzCqN0WrAozq9wNkASEyAATHQlBQ+nHZtuFUxSQV/
drJa1Jw98dNWUS58ne/446TRmSLxbczT+IBqBBUpOCXy/UoD+gZHl7Vd1V+/zExTuIOPDA3lp7Yq
mfcmQxdJk3T4+cg8ppMMz8RabdNXmFLPes/qu4IpsgzWfJQWWJ1T+Rw/3PJCOGuEftd8ME7o6sbc
nDEMVR6RGMeg7rLYFSL/3wLh0q+q89F4m5sX9Ak07akNsenaWjsv7HacJwfTvJymzI6eJ8/F6OZn
uCEI7tcNs28DxbobP7VddzsMc92Wk/HImXQYUueYtOJ7HSsqjxLE32CuxrxElDtHFCpmeEkMfbyI
w8Z/R7TDMPlfxKUfuevpjPyKCSYloj26r2BOw8Ex47NYtAVgtNAXErModeshZLDofScVH9vXk4OB
Fpvr1pqPaT09I0vdaU/W+srWMCr3KZK4sqIYy5lOXfmSDiy4nCVlrQeXTRNAheQNpJVaoJw/9Hkq
DfNMMEqTwaOh5qVXXrHDsWSglJxtvHwWM44lk3F7yojxbffoGnMYQPgpgYaVCEWvkcUb5+Q56uHQ
9grBum6QaAfYPpQ4wbiTMWJ7+rtjEJ/sflQ3dd7CS9hsdGKgN8p2ta6E3bHFq6sRI6vzHKNLa+5/
6ssahshbGRnNcuU50PbQyhufYiNRdhrOWvFdkEb5JloGmjjkzpH2GFkrk7P1kd8Vyfzt/hPMl/7c
NkHtsIy/4N15xZZoS049VsmUTxIzhHoQaPF/Qs0lKwpqAcyuVtwXKlTqdhsejnfqlOIAdG3ZEocq
QY3c6Joce0Wp6gK5ceL+aZq8IqgB4c/jUhnTkdU3/MvsjSGXehzzQul5859bAb0TRB6jKOTYSoSf
xgdG4rAoZa3yHp0U2GfAwaZSIT07sJm1WL6skxtXIc/0OzP5mk44LpfV2YUxWU0nSmd9Ob5HMWfL
wVVrYYEnxFRXDQpiqzntKKd9aYBHuugrwCUdv+tQRF9uowDxCg2xT/iHPM5Jgbh5YdHQMRi3c6jL
LwytIPlcIFA+eY0MtZoIk9gVI9m+/+mdxfjTD5bnAZuRwnf7eQH4wcdB864Nr+XCNEHOxhmzbRQn
mKCEXgWW0AREu/WwTc2c+J5xMm10rgdQV6V2d15MAf/oad4AjObwGyxAfYDbJdv38lSk90iazfNN
mnrewNmzz5DncwzbCrz+iAzvoVgFLX8ZyrrKCF3eS320ZDU9jExXCdIC0JyPNaiXxPhp7/68+nlc
hc3V+7p4JcKqPxBWUdQGbMBaz8BATljD58r2fWg4lmx0mCsOr1S7NC+Gld1zBxOqWHqV0YGjyaHG
IrdNqcROC7azw0CGB9pB/se3EcHZI12CFEwydYPoXpXACr/8dLN07M9b5umsEDPz9eTDCOy1E/1A
Z10B73MAEZ/u1ExgVIfct4DGI9h3uBI4sZYnyrnKMDpjbJAF0x6i0ZnUT11Xo+ln7HObDbTL9tNt
AGEtel/bPLX/OrmIP2+aWWddyFDMqAXc1SNA8X0g4h5YquDyD+lFnApxro4vc+iSWUfozLBGbEO6
4WoIP0imrGEvBAuLaa3OS0P1TlZfad36vF5NNPUYyT0Onzf3Z0aC32poRd7kTrssU6vvSdwKh2w1
Y2+o72zpxuPOL/hXsnGZBSP2Ht6AEW3b0dtihzY+7doYBataJAqjaHwPBOM4CZZIGb1fhuDa7mbj
mgRQOoCd2vH56Qz9m7igPjLBJG6flr5hjqOCcn2VvuiJipGTfHew4jNdUW3NwAU9pnYy3jel7y3l
WzS/EZBhSyYyKPLUczWQ9sHUDWZhpzMlPouF/s8M7MXt5fs8TaqPoYTfR5ol2zoUH143968GhW2H
QXA8H3KOodvD136lpD+S1uGgOHKcF/cT7EzZkZaKpQgR5JdovZFgZUC9hiuisYsV/CZS5BMTaC4f
rAYH1BNDb4KQ0RPsq7QKBNwxzKrytJ9E4HMba0Gb1v8ApeVZEMsCKhfz1Cbtq7spspiQVwBo7EgS
7tdchr1Y4Z4/WgWp/oGeWF7SvpLoH7Gz7McGr14N+IAAXcu/CXzH8YgpjMb3vw1A3TUlpnnOrMWf
Hbo7K8iR9tItS760977blRJTEOUgioUeO/v1dn/P/D+UNd76mLUcB+arZDSdmjfqWpUyFmQ+NZh8
zbefWxP9WlBdmNndRCozZpB/gZqj9qaQsuDRFeoRLr91V2Rb9ZAAw8cOQ/+S7mIRA7Br0v2+wBPo
d+Rslv6zrRJn8vLkIkTc8NRkRDQaLWOxIz/obn1hqARKoi6jzDbWJYwLNzxuBXDvU0r9tFJpEw5u
OD+vDSiyCyq7I3hbKUFuwCCjKlShplGZV+19ta1yhD63EMpMDUl+Q0Oi6kGyw/PJQdiF+egr6FSa
Gf91G1aRrWRzrKcaQmMd6sZUaibvvLNDfCmpqJUkhYxkRNy7ykX8cz76xSI5AI38abIsZIezYAiC
XYztiPmAurAffDlvDzlh1KmtoKc+mSZvb1ij8ogbbMljxGufh4cqmTJLZWww/byeYsJpNAiKhMNR
9Z6do3jbcauG3/EK73uwTTYKXWRJU/OxvD+LiOBk54iQ2OkNpOdqxBD3+5HqAsGYrflobCORv+z/
l4mrPDRVFBk3LEm7XbRdMxb01apSzReXBUZJB8olmvOTwktvDc8R7YD/cLvMtxlI9KpuPdGKAWRj
TITsIJgMXiJVrwWPHysf0DmULME5b2w3HbsNZwsC/yPVa9dqyMKNZiL9RZjCdnTFt8wpsj9/R2nD
jIy98mOBCWS7KF1FM588W+WF54emxQ4gSmZB6DSGn5T+IWQnrhCU+wHBRVxZC9gAEHsTb5n0TsSE
fxvfX1jTAl228+PJeYA0Dw46Ab9aKRVOo/bH/oXzgHUbtal8nDZjvpTVgkr6hismrIq0bzmImRSo
6yKoQXXGo0rKPpkQYfl+VbOFCKQN+mkae4cANVy5FqHPCGlGCdBolHxIwOBZvSPkVsrMg9WkWftS
WErmMmdAGo8hM4wBnbN0A2cdleX9Vok7Qosixj6fEGQNaEndQu9JbwmyKP4VqqwANp2N+qPYXQRd
U0m7xvoBaaXuid8K4MdrijnRiFgJK2LRotGYdqun81SjZl6QMj51NTSK2SWEyKXDrTrphD6HZ0RR
G7CcR/XzWPomY39h2xOuLD3GMHsM0ioM9zJbK2zGjvSKsFFpbosyY6WdOAb8vXpRlElDP2lJbfUO
f0WW5c9R7q14NGDWNTTVDMK+1GDB3ej+hhTG3q3XdBZ0TTdCh0iuPTQbNe6mo6TIEoP+NLmVkCs/
P1YR4marPDY2m1+rLwsLyQxjtGetd5+YTu5g0Iub6opxQ10GEmjsrfOJS1blhavOMfGjwJ99tvRN
fDi47QxmtBkTMDdjNwtbnAeNz2cVyAdpByN2MrYJTBVqxMI8dx4GcLv4U3gjxntRODGPmlUJ4cb9
3Vu2qsVoYZ9jwUUPxIjpSptO6gfDkpjVYjShonxL1HevsnTqTjCESnNzlaGQl/QQwyEXVjfYdgLf
Lw8OcvInDp5b9GoXaO8FLAtG9Qi/d3VnGTTrPc9kTlI7WZEi9XimNdLWfFBOh5fwL2eqSugYFTQg
0pCohbV8W3lIHv7kKjTI1cpW3LlaegFFcX4phax7a6GHEGKtHlsLTIVM6xR0jzETa8CLK6ZEiGpH
5LSY3UycMPhyxZOTdwlvtQ0Th6+WdkUOSwTi24NSkZS/1txo34C2VbS1qAbTTbAAMOiOrpLLpntI
MxFp9w4ZfFOW/XuFOoA1bWP0AFjh4VGFrhHJy6WVPYkW0MUa4xVCSv0cFbq2JS4gXj6ADGoGlHzC
VSCosofRlAMK2aJ3ber07CdozPqzLG0tXAfx9kl1BmypqkD/dnKyvNM2xGMKYV3WT3m7sUHW82L2
vZJaBVw8iRm0kV2iIDKxzIVMN/2kfom2+1pY8LHB1+gXEJQLsa8y8JcCltn4geKmA8TJXjuLV2wO
sKih28/F1j3JMZ6hhXUqZd6/lKAWFdmVV+rQG9PNnawp6PC7qY8zxuPwU6ilOrV9e2rxp0wzbZzu
nyPOrbQ9Mu6IbARLqrXbh5y2FQ9znHgfMLpDIK24bi36SjM7uz0MFEVyQKjhaWXy+efXPtyliWcv
JoT0tWxEe+tcYGc+fExnsHmB0WIp1xrjnuHMRYsINYXjmH4Aidcj2IjrUQJAw7hRrjQHllb4YdlZ
dCIZVHKxTa9hPAsp58hQhn5tgK0mCrjdksErpxAAOYCnlHMTNQ39jYBVNJRsbmI8iI6YUjlU9r9i
nqE/0iouqEEAMSDkef2GbyAm69CVUQmSfF9kDk5CCuUbrCazaUf15JfJGFFmten43ZoT1fY7y0FT
g8gLa8laznKECkCHVUFsV/yApZQRT9XTP/eKENfPCIvfiYFes75sIyxbUy0LiV6h5Kki/+vnca3M
HstvxsZcJTms05Vv2RR2r/6qCeC7RKOZvGR2bkM0yd8ipiZHnHzrUcTqoqtdD/e+MWGNBppYR5TJ
9TyqeIRZO7QGSQCPMrfnJYh/Hy1wiB89DVAYi59BIdubgNLjeinN3C7FdRlrF0t80oyckkDy3ISe
ZbBgW7cyThqeLUfKn9YYkpdRGIoRzpCP57s2cDTCMCrMqFeuNnUDzfQPh9LvYAAgCFicKZaQrD/q
yZCLnjF+8RZf4sTeGxgpUtPvnnoqXpgmrX3TFw2rNk1rlJoIpGpM9NlTYHbFSTEVnZYgWI0r8cy4
dBgeFvCHtMUCcshxSGa12Wvpg/N2T1eW9qZCeTtfSkElnfZXCukyYEbegPSj4jRGWIWpC17j2VIx
M7EVvKEb7drpGPPN7pxb7AmS7/KJUK/hOunlaxDs5uo8WJq6Km26TJ0uDuuohD1aLnBbobHQZ2Hq
FXz8iKlU8FlZpQIJpUil4E8ex3dY8Gk+aNDQJ2tpFhUBdFGRrEvELZvpsuFYWc1aXcCIjouCxegY
loykcQ5tlKEkW5vmDeW5zucsNXDrxyj4pyinZ6RsW2n3a7jUQANEnsw1Qe4zhnRZR5Tl0syXirkI
ljMJk5QS40tj7hjPgkQvZVHBjWAco0xs7k4UbNpz42G5mPUk5mJy4uYcBIjl2zls8x1lM4UlJI+0
dLKSjMbJcPSwmmebolIcWReGUxG/kmtj6X10vDFyYGOYX3NVBke3ISR5XOvbV2OKn+YBB85tXgE5
JZ3kYinpG6PjBW1s/i1HpxGD4tbEZOVKKLKXbs0MeizvmrEqXJdGg7E483nYMTyMYwBuqnF8i2yO
nUabYzrehWCtXwe8Mc3T47dKMi/BVn34c3eAlH0idJlSYfFgjBsQHyZ4MrGyVV9CP6FjC8Zpri69
FqPLo1sHb7+3/7aGuhOYAbCV8YTvwSCOrqExkEWZDPantI6LK0Fu5toUuyfXFvbNYDhmB0rSRW5e
xtSn+0A26KfQ8fFdkHuxdWjMCTn/AMHeiInq7UN5Gcrbx7zRpDkKWaW8rihRGoQksoBPWb0mTYaV
jI0E1ZH36q84nhmSHP/fGjabtcQqzqzYRnQv82BKd0c/Yfan79v1zhgBFpfggsFrzM+md1PRqauM
Mb3HKxstvZy4ixpkB+SqDWw2CWuMVFrcVcDLF6QGqveHhZxJp9OburW7gXVqrgnmfGzDnKXANHou
I8PbFzHfdMuC506AAjJVLx7WphNkoxYKHojzoKeqP3mxWAn2D6AFAj654VFf0h4XPHZ98Yt21ngp
4xIRj07fsZ50Xv7A3gn5HNqIauuyp2EjpI3X8hGz1cKLzbYoVtA0/8AgmiAAcOfAft9N9HSTxr7X
0K6aS8AsOfLnIQzesgRtFPhWAgZ+ohGD2voHeUUdNLMMIbJh115AKJG/pQB2+kSjaaJkw26OLZXS
+9bgbqnwemMrEOqmxuJOJ+t4JJRj6JewyaX/2HMkEHm/McsbSHeuBLaBNtDGiVd/N087L8m4Cv3F
PAEaBlddh1fG/WqnuiV3+yOp7b+DnyR29bHdPUc2umaUjQJAnCZO/LLaZV2oexAXewtF3KW2FpNY
KC6jAtmYn/TpcW9MZkMxjWSwpujP7N3QXckaYE19FFEHKTTvV1sip/KOBMO1vnQiKep+m0M643eW
S8/eS4c2n9hwxfGKC4AHfE2NjjaAMJJA5COva2yjGtIdRAqVfROlhsBx1+xXTofGaochNb/slALC
2acFoddV5mZyFpmd3JJFF01MEgXhqn40Qo/tcYRybb7nubfeHukKD9NAgQT1gDfY9MvhKp2Ala0e
njiTXRBAitEojnonXBG9q4WkG+96mC678K5biRlCYHodAC1KePR9JWt4ADvip/qSllaCoM8IvaGH
gORsMnRgjxfhRYW5ndGbl2cKgyiKnKEFngxBvOTqWbPtGun1r1Yg67IzgVgJgzRgdiNc1dN3+1Yx
bSBuQyrczmEi9ljJVGHyC/wmWaRRFjNKnMnUUYy5Nx+GiaQONzSviwahztQQiSrfGxN3E/uYrJqM
C9vJ+7eaD1GlBjNg0qPmwXnb3ij83Nkn2MgIReVsOneUg4Jq8Q2zqa9o7OyhHgOYEGkwrZ3B0zBM
NqqFC/pCq6qCaZmMwT1TmB53bnR0bB1/125CCCElZyxoQ1XGiP05tSMLPSQ3LLXoHfQzmi2yzYKD
Fpixjd3B+9HJbZkqqim71OyCJvfokQyFa7HfL/xML0bgw6jUSnevXGeWo6pagd9NU0XNqy0VZEyv
cF9HH5dcmX0K92qjmk/4Z3KFCD/gKPwxv36If64ZSUYx+8P7twMB/MApSYBWa15iUtdcUs4WsGJC
NljQvzfkpkGFqryOKDhLbR19ArsND6j3Ec42+ELQmXolAYYxJHdK89pNaBbw7CB2erZZp6csG/f8
VPS2MR+7m5+URJ3cib11E8WCp6iOdxyaGQdb4W7Aomjc8deYu1LNuAucVzANKIX6d2fbE7xq8HxH
E0a1xyMKpIwqaBjJOt3M/2Se6oSUPMvA+ZPwnz484OmcRvs7UyrwDy9sFpFBn2L98hUWtJD/K/2H
+ntTsyxRPmg+C8JEmukm31byyWNhv4OQRSN0K9eWEkQHSDE0X3e2NUFhGgv6TdA7u3Yji/A8WCW5
gIlO59gRKkhYjvJIQ3JXnc7yBRkLXJLHP8/Oq5WqRtealEQkvfEPZIPfMcRJlF2CqhpRYKN+C5L/
DswmWvW2z4Rmndeciz+fb3IpqOWf0sOidwcugqKMHq9dxTt+uD20BwQS4BKs6PsYfiY31sMMCcTd
lZpgXbHFYUj14Og+S54/bxv0i23QsL0hFsQD7DTKPvLCbOu53nfJJg4yJQyKp3XOTUB9Ezb036Li
mnaz6uEmwku7ctpoUxgk3TRMQiCYhTCPNKZTk1Q7UXn437LPq6uRgLBDX/vSzlvR2c9bZTPJKZe6
qHuRX+J4/f4mSIyDxZU3RW4xY93dI70DjOsveZBa1WkKA8fUUS3CLMPkXnnSAH7oRgWWGNLJ8SXZ
YBsX2mydhZvPj15GnWB08dbFvSYbr9JMZQDIPFIRwD7MZ3V51shrAFmF1+DqMlVZLQSmZJfvIyDn
K5JLTBc6a7e9thdfdN+sPv0eBX7Nv7w5QZKUvzvGiZUkOBGNcX/crQ3lXgy+Oqv9Q+A5Ru+z/wwE
cA6vEkvJii0TqJRQ09iK70Og0Mv1Mt5MvAgRDTsC9WDjUG0MJN5d0C27VzuS2NLMSjkVodHW3Nf6
Ir8G+I27dL02AxHo9jqn5yZIIkyBGDZZ8dYJJ+krnuv2nxV02HKqN0kFd/aRQsdXu7d8eWy1UGfR
7Nqlakg+CUCXPmb7AnFGEF32ywlKx5hY0obOPfvVr1qKgca6HCwZFvuOOVZS0pZ+nr8grZdvL0kg
DXzYmaiwdU9c6ZmzTjzkYWDl3+bdWYO28PXZ+kNpeoNsDZiuR0Vbb8S+P7njzXGSPXsHLGu0BWCD
qNBC/BMj/Le6uFtznkVZPwTDJQJdr5gKzlAuZ548nrqzgk0pTIwWa3NeaEwKz96OxC/yLHlnNon/
xvN2NeEaECkpV2tWS7nCf3fW8wP585jntTjYPRmLIN37EczANASuViqiMBbuZmFWneYwZioLxoeJ
DIIgFe3J7FO7eV2AWIuNX1Q5RqSVEVAW0A1onqy8ZdaKyy9JgqEH5WoP1lXtJUSp12Cum1IQBAtb
HB9aZ3oEK+rDXd3hMbKw3bHVhrSekr3xE8pkxxHCYUdMKDSz8KnwMYm7j9tmDj//dKDmMcEDCkfC
0/tarsH9b3VzEmL/g8mnzCpqcUuIRG9v2FWpQtEbSintGBJqlAwPjZ+M1SQSsRWVScD4xHV32dWo
+NHoALNO4Op3sKe9nrxb9Ib61HGQYnX4IXpoB7Kd7O/bdM1FS29RsFOSOZllRe132XowH7p/iPm4
KN4wog/tP6gl15TJqUdPkabfm/S+abgJ6RzGALYRf5I5PJ5/3jYV42CmeyomIz4WqCXN+J6F4f4x
A9LH0k77+4/ysgkzG86DliYVrfdN1sWxygWsBtBA0xsqXlaM4LpTpQHAW9mATSauTBTkcFvpeCUV
JF/4DE0DDu+R1CbRyOESc1wb4ow50tHmPTr46bTV5DeQa/M+SCyskVc0mjbkt0u9kMQMjxQTb8fe
AX0QRLHa9DYIEr2KbyyNaIfuLPl08m8IP2QWdVEk5ysp3ktVZQZulqpzs+ZEfU9sVVSa3609+bpr
HPbYQDyXdCcLqVX94mV5NOCFNYkegLdLirS8S1gpwuSDN8QYsCZcQMWAURoYmrSyy883KdwqIFs8
2uRF7ojtHbmqs0ouh9OFGRMRJv2+khey0m8K6yrS5WbuCaq0KBXVEcSkw+pw/w4jA0be2IzGP04c
Fo/IBUng32mlieoCKAJiiymLWD6mKpr2MSw3MZk6yO0imySQqJLrDaiGj1CpNkZ+fsZ1XPNLxRfg
7WY7OZLPGvUZ3vEnsbOVIAmSglDMq9goJ408lu0xO+bLVKU37Zp8wiEFk45Xx2YFrwduDuFBC/6t
M+Og8rEjDAMNczrzGT82zQUhqt1Dj5RHf5I3W81caKnfmS54tsDXBCe1n1k4l2fgIBAayjeNQn8F
fK01nkSnSYq0wDrd8xaNuF7wOQ/dim8mLIsCC7MLLsuM28DJ9IFb00Et4yDsIqQBD9QLkvDgNrqD
P52BPUwfsW8DXr0AJpXB9vnarYU2JAnPharLefFt3HtHM81vY5my6AImAo5NPXkIP5kMhHfBRAqc
uZyGCc9q/GRzHfxb2IZ6g717oNoUlQU+Wy0/LK1vft2VcrN4bJfKOLMbJckOjEjaauPYuHVniwRg
fGARpeIiVIcoc4Uzp7/vJOadz4xQoKO9nNhOYwS34TtNr7+RkyVA9E6ew6ZT93cB58iTEGb3/6NV
97zAAkSBvQjgXprhsNSku6FDGpulk2d4yTeT9YVaF08Y7FHuoRYizI7UAmP5r+afrtU06Gnh3s5G
VWGnxMbNnSBPdqPDwv8zqo62RyvrdOopqqf5NfmH7V61fkHX22Cuyy2hqUs1nlUQNJcInSeet5Wi
Mx0KE9HnriDlDntVPDDdFofi+Db5ncKsaLwskspQocNCnWxV4ga9P+gTrVYhGSQXAGKkF4xj3uS3
VBlrV0sFqGbsydJ6c3d4fsm4QrQnl2pV/tWDxNrsy2d+aIQNwTqheKnNDzs2OQYPkQfWGvII+K/X
pBd1oePpn+t7FqD1WYduEUl+8IadwqVIYkg4cAwxZTjr0W29njXhGyag/8LnBeWUdDhCwdTwmkpD
4z/zKgvMIndATpWfIr1I+xVrXDNQc0TNnOPQwDhdsl+ecApyt6/rxf7MN5RuIScvkuoRJwTgW89q
wpOcRsCEDR7kRkF6JK6+FJ6UKrDouWU05y3846zntyaKZkKBuiCH4GgMKJJLGDItg8QmifesJvAJ
/HMRChhV6LFfuVqhX2hpLbQbgbYpmziySMgOPj7M72f0RvxrT4rEr5J1zlMv1FanpbaRVbeF7r88
3Vfi1ck3Q4cfGuQJq68nXJWjiSVB8AaPG5gie/Z9u+jT59YACRaU3kOzwLKjJzTCfSvMhxZSWtr4
BWgsE0s4MTKsRYFbtqhxrX4QXchrSg+kTZoEFcY4VIIFfd9mT0bV1Et60kkKLudrD5a5/91p3Apj
kI+NYhRRxaxaXEfDE1b5S//dw+OPNGH+sdB03PNmCJ9lUE9BPAUxQhHo+9g6sWlt7zgRUnEc1Sub
oLXULUUnJNLLhMBbdoTBAk16maTjLwzfKADaqphspG8FoTLE+zZIcJZCdv3a8LJjaUDvCty+kL7l
AAEJY+vd1vhsmkvw9FxOCqBRG86KQx/pTSNZ76vNjA0K09oJm/Nr2YpmbyXFQg6jltVT0f4i6h8O
eI2C2BBL71icXkgLcW9qT0YDLpH2GXH+YET9Ardkw2H39f2UysjO8cWI5bQ8bHSHWlWyiyAym9Wl
LFQjqQMSrQLa3lF59IG/hwy88hYJbxdegUakEh/yYZE7qB7mMR3doeXBZ4+MHXpuDiypBPnABdYK
zvCb84WmY7MhEuQqmFYmmVJtKJzLoqWTi1eUhZwRbN60QzhMk+dZ43rISTLnwuT/JRp2k/tTmfyT
X7OxjEUkilW8D+9Whff+GN5X2L3Gp+Ruir84Rhdq7jvEoCgOQZbtZlQt9ksBOR1KcYZgEc2fvalI
cueoDwwMgdqujLjY6EagQnPq/AaLy/vadU2vKuP3Aa7KDkXXPYOPPg9HY5j1Y8QQexACdP9Ky2GI
pxKjixxCyg0iIa00/3VaaHpLa/jyEBEKfL8KlOub4M+RHzY/KKgI7cqIc7GLJu+QJnEqgh+1c36C
ux0uKRq+WAT58APBwrtx1EVPY1nuYBDDIdsuKhprBDYJgSQPAiZdmqLKp2BTtRp2uFFluHw9ypuj
dBac9kJXCqt7EmDCADx48Qwex4N+A3NWLmQD/E+bbvCNHIDk5mBjEn/PxNvh5R0Ts8o6af/AR2Jv
6C/zhaNg/pxQZjxOEGSXoZWEWF+rqvrSBk7HprVm22nH0k4J+ki6WKP+K+NUO7cW3dNPxcwGwLWE
3pRUItDbT2+tSEza83cX3OGLyINwyDQAUEfmnEod1eHHIMZMW5QLofiTLG7nID5SlUNLK+GYxaqk
cyDoNbnVK1W+7QM2eIZIai1GdQakhB1U7hFlLXrdQjpBVPne73H2U2dhnZSUni2PDRVpzKWNLmGS
r4C2Ke3Yt5WknfXpbay8lCS1GDy/CmstWzk37xqmydE5jsSWLant5mV23SbH20pAlvVMltTf4Rwp
AxjwMQKvGQ0vv1CFzhzGo4GQDjG1yXZ/sSzwon9gt3EWZz3lXuqQxUx/WGnZuF8IJFBniWbqMBMt
hihTMzRO4hsZcTKk0gBFMxKqi7tonAWc6HhLML4oA2iN8Q7Y0IX7SBJ4PP+2FrIo7nL3BlHMAO62
tXk9g7VxhLWd9h9Y0L1l62n9VmlOzk53UFrFV1B0VmyH5UDNKNXzs8he5lSe/lVzn/3FNR7ulAUS
Q9SVGGUPLwG1HLoPwhSAdhslScgIBnm++gkHInfuIPUxCkT3ns5sSlP4nFOhxWOBEyG31JnM/qHq
nQCy6N3rtjMZ2zSt6o7camc5qhK6btfRSwUOUD4o2kpebUVX0R6cOOPja47GGZbA1FLl/d+rXmDi
qU80DI9G+vFzitmQUmLCY+1Ki/M8a8eh8q090QrinFaGvcJZrKEGpXF3G4MuyxqdZLhSfITg7GK1
ijZS+MzLRhhNYU5aS7bKZyOmTF3ImzjG4sl+Kfsi2ji8vgjgo9tlE6hHQoPUp95acrS6slzO8L1q
nX7G8CAynsdLO44LlX1niWdxSuVBRbM79nICVyVTDCGxFDQg+Saq7hPEkGXIhboej6hKOsChPvuy
8FxdLsq4MgFbwnnFRmqb/NjHlqvnuQNwlcq2ADmQxJqhNfustFZI2UKWyLp0sn7BWg9gT+AoO8Um
CVu8rrg/gj2LAp+uFSwKqTH4ZTZRbUqYX3RqjjnvIuqbRQuxR3HQIdLIwRy+WO+y25eMUCXFTNnq
wXI0p6sIY+cOqKi7HU4Rr9ugsVJAh/tCssiWfIw1p6hkKxfGt23uhyVfCYCycqArymcmunzDv5YO
lTEZJLlsdKRKJEFMJr3Qn0dBUxQJPhDER0FZY0LFsbHaZQCp/JE0eoDgebRINtFgWj4AYm5QkNSR
4UKEeNCLHWCyi1l33/ul6elCEst8rFW6nlCA5B3tOkfwgA3CCYElcHZQ445Zn51lOnfB3bOuutam
Ezf9aZ4T1qsdXkGqJaL0d63/YXpHEWCQvqjwK1i4UJxEAPb7rLfJLJkJ70hQmZ2t/+SPAO3GQobM
QYjOjzbOi59iZjwJjuj+dUGWK14b7/R9akEkh9Ajm4KCaRFUZuFuxyP6uEWzWXF4MNOaNYVm/9Hk
7k5vsT9bHn87SUr0eipqvabwY88Ttz7WX5GCiM0yt0Q1tocm4fJZ36JD/jgatzYWmELeyVD90lD3
CEpqNNdB20RFGSNIgtro/0/kXgeTw8uPmvqj5JqwguwJkuZydQPNBDUr/DRT0ICa+d8Mo31PbDNS
yNxK1ED72a1emM8FoL7qYyakxiHFEazTicKnMZ9mvw6z48T0ux+oZouTyUBe1bTewpqDI9vuoqry
qAjfVQ0LJZ7xoDnNx2SWs/nqcIFF4VNrokoAqxY/jjNbFfsWEH3rtFEDebyI3fMI3PKYaBAvOA3H
BAGo1rXxZVEdCrjCX8zHhurOiw7um4GNscFnYuyCJrDFM2dw4h02xMP9P38bXQ7hnNTzrkRN3oPb
FEjFJVDb8CUAIxsxgNdhKy51ShVEPdhfGgChZ2Qya69XQhXoiJVLX5SfwMP0XLyG/e1qjf2Wac/L
QkNoGoz7NlIyMwU4XIDW/EQEB5R2/jgnYSgK5Ig9cgVynZrCWz32Ng8J9hBxaIVtIp1SgvnN4ayo
07Xm26tl+PFhGrXYV8/mVy/6TF7mjGmpYg/3y/YTnEAt2BjEqMxwwz6Lb4ElgGT58Xc2Ni13/Rom
/9bbVpt7QZmi6v+Qbz213e4nvrRCxuHjtm0VHWuYWE59icp8aEFMW1qRur+NX/3otxb1OSf+L/VQ
Uxh+KaoczK4/7TuUwQl8uTU9tLmax6Q5KZsIBV+z3zD7acd6yD0QU9aM/Td4FUp3QPFmm8/IvHal
iK/5Emx4Qn8KvvoezBTVSZ37vYyAG+3II8jLi0eJ1j7aH3cBUVD1MXT2C+3ACUvz4pIYr2lvDhvB
REhteeGDH5smCVBoW3M9JlAX6fWF6BZpbS7UsCRZAxWZwfEnUwq1qU61iTlf0BvnI0pvpGS2lRp4
+BydGVQMmvqWD36hYXikTOlsPovqTMKR8hsXi88/dDipB1MICV2IV9XUdABMGrFP3sRObvzu/BSL
NdwUOcEzGIZSfmjSzhNY5dQUlEHI1T6stO440QzYxIdG/BTm5h1SF0N3KpjoAvcv4GL/GG5bIOXV
4y4I/BsF8lvHltHqco8qw53BAxHNmYtYNBud3ILhdjJi5Zpr7ymsMFrVcwkT3b6x3om6Yb9QxqzU
uyV7OeboecA93QJUMmmDE/AE2xSLQNBfSRXHHwcyEeHajhjj0lDm4aQerdEY7dkdYqNu4tHACQ8m
5muP2bSgRiQLxtcQW5i2TGnDShsVgFS5INBgZ2rMLrDLYFk3/IF0+2gi7ug0HrNWT8CFFd8WXqWd
TCgzqliD/CS3dcYelLtGOcpIXSlO7KAVs+TiC0H5qCGpxnytrrP4K/c281Q4KcWKQ6BDPTcfgUr+
AMBOEFfpvRbaUNHtIapiGneuNEYYQQ4tCdbLziZfIHP+2tSMQSIZIX0Lh6L1QuEGSVbgTpjMt+KT
txH/6rCAh3hkfNYhxEAHmatsvJ17Hz6/zdzEMr9dRydTQFWMZiJmWjsBKrlawe6KcbeicW9AI3DJ
LJI/6kmubsv5RCjpTY7g+zczUpfd7ggGcuGk+gCLPG37lR23n4ICIVJtmL2rroYWG+NuSisCSp6m
t3Q8VhCheLxThlNj3xDsOcNqwd8dCcL6Hjj6zA4KEnE+9k6NwOAdCtGAgd5Zoa/mJy9loV/eSyQq
bqc01IRDQh2xJstou8o3gmBE0LEEvcCN5DAmFk15ATstRZmkSowaBe+v/8joJqzWnqOY9JHBU7Ub
rmspThw2NAWONLSnpWzhnxvXnmmgmC1Eokm57G7a7txY7zwL6aiMSAOxHgdQl6fYwd8lbgUIzP6/
X/Wf350DVHH3C5v4pJx1aOFv+k/TM9YFOjneEHoHdlcWnh0pbby1/nELvfrznygtcGzQVfpLJhXn
Nfn030SD/jD2bN1DZfkq50HUtgSkvmm+bg8rR7A2p4QCe6EdNzVMfSs5F+UkzAQHRnAgLB9NhivO
XRKnSLHtHI+2lQS95BMDjmgJRP2Mi7qkv/tOp0IC11euCrQRm0Tstm5Kg2MDoqcVArV/oQMPoNDC
Y3tDXy6b5iSvsIOhi/Dhey8X0GoiwrZ1lZ0SVTy2lbMY6CznEa+ECcGV3EDzNFQzmKQBkU+Ty4pk
uhuAfxPr5VH7lbbXSc90/Nksd06dr9Z9RPl6f996DlZNGVofyM4C8mlupjUklYTricurNnNehL10
V0TVWngt+PZYpmYNa+AB+T9Igtg6xednx9k6lUZNWrJAqL9/AqBnKTR70eZTD2FXG2LxqtcFlcR3
p4RLHY4bwZA71MszFlZs2XMAe+fClcMoSHpSTHc9BF9SPXbHteVMqPrOcKcpr0L+a3ZoapYKdoJu
pMI7O0lTz0WVp4JH4nkwQOcBEmQnldsMIJ3mHxJit8U53C6T6LlLocpOJLb3sNSepjIMbn6IqCW+
4gVs+u25xFv9wRgeCi/WOOGMvsg9SZvmzVhnRaDBHpDZWbz2mXXv2P1yrKRmTc11ASSeTv2GyjqD
+PuvUiCWiD8fOT4vFxejz7sB6K641baQJgyhk4uJh62AZT7XVuIcji5LdwP80PnnXxOEWzochdiY
HsBXMm+AJDQbRM0M90pebmLWZHGo68AJ/V4dwPkaLlk9Q4pCCECTdNvxbuM45Rm50hmT/TqiNeI1
g8FrxwppakovHCpEn5OsT137XUaRy3PdOdGEUCPQASlD3E4owmo8Dr9ycnR6bCt/8m5vS/VbYNpL
tzqNxhOFGpe/R5yO5xI1gdrAbtq6MEwUzB7svcdJ9SEQ+0dPmo0tuAYiOvKHCsMCoQOPOycNoY3h
cW5hTtPNt/DOkxl5DOF5T4nvtd4uwOqQ6xz5TmQhpzzvYO1gCI+KMEc1cJOPLfvIiflBKwCnQZTI
ezHPZ9eduj6qhpl2mLdQzp+UHVXWwAS2EmS9FYgdbOnHzvkDYQ5n7SQMZCoO+7xzEXt/axdA/6dF
hAz0bOZzFq1rUp4vRv/aHpCiFjf49bI0mahZMq5pDcAnTr7IHuo12e4kvIL6cwNoSJyRaveV3w8L
PI8WhGhi4T02QB4fv1BOxhH9BnHzZo3C7a4thMR0oLwO44p59ekoXj7yLZUqfaSk12NS4Saq9YEu
P3kE3UXtZCHirt16tA0r7cZTumV8rMGe9+lh7M9eh325glx7LzNn/SiO1TUdEJk2k9e7f11R5vyR
u8i3f8cIZ1PPjodCCM+9kznc2ui4rTyM/MhY/jBZN9khgnLKXgkXucxsAJsquyrRmyF6TD5HlhRu
CDfqFU6hWUjXoHflTAHhLvyuHCfUYwFYPIyVYUt06bEgBBjB6XCrqzmeM8pPsjLrqDzsJMhFeEvD
4NKJL92fSXbc7bVgh+IyfTZIG5MqbW0I4+Y4W5dC9Kzu+cEXRWjAYAF7Pw+UCKt/zXJdoA4wiGy7
g1dogBArrxui3KxKMAIKfB8YHpwxNd5D39vWFmzGF7Z6PSeJhHkb0UEPKeGmj8JcSJHq2ypjfiqF
+7sypMEpmHH6a0Tzyc4N5XQdxkAW5dKEZOPt1HUU1GoPoxwgQOXSgsddB0lbndhQjOpdpcf7+bFL
FsOxIKgDQjng79XjgERPhxadx9wr2YAMp1kz8nb90+L64BgY5d3yYx3Qrmg7faGFAEDZ8Y7xO6oo
TDw8W27HyguwOJS8g2YoJyf2SKeMlEG4Mp+uF+WzjQjc0LidzU0EmYh9p4DPZCtabmcbkgRjHQWe
mZaKmkZwI5vdm+fm7axEHFvS90zgopXeIpffPlaTOvp7ytwjMwfhJfuvaFTV7TJQxwdcjgrbZ/mm
ZLP09GTyIzBuOhVx1l2iHbvlqgab0iBVLCAb+KWYC3EQtuhOTuGayYO+ACXfbPqJDhmbnkpsMmzt
JdTbFdfk1/CZeDJz5ckBzb7Ld9TAkK7ZU4KsDOPAtg7e6R3sUGziGpXHo3O6AvfPaS5vNMbUDOy8
qAizdfJsKNlFbScfjm2k7ld1DsgbLgHuvgLj97PzZvTCAIf6SaJL/zwdMTtM/6QI4qnkbheZUiVB
ZFSX7oWdQD6/JQwcb/qkypJshaXNWaX/zQzFjAtZ8kja/gkwBJ1x6l8JNGT/znVatblbMZRs3bqw
No7PyeT+ODnYNTKMwsvm8yVrrECR7ePvbOY5p6Z0hB+jfmIpBxlFHiKWkz/cg7yIKL3JPwfC0yFq
zb8h0vfmRZKyRNAjPdUpaC1dw+kkEJbsmOUjhY2hG03I8O72u33ZCZ/E62F6Ryc2v9pFU1pkbp+R
zGUfkGdxnHzGpxPXd88t+JhESWoQ4kWPyB4azDKmz1oVD9BeeXWP3wwZcEHvgh5bmKpPlepAhitb
tYW18yW0nOd5QlJsTLs0X2+2MD1egEeKavUYPm0Frrt/pKmTzyo0E2XUwRP4Ucr2hJCxFh0kqEBT
W+39NQ3g6GK7ZASrTLcJV+3aBE0j7L3GhenD0r1+HbawnMF5Lk+WxkRLC7b9m2199DXRkJVM8N6a
lSWYZuaPOwUA+cNJfgw6dxjLFWReWokDOSwV8jnAg0XgUR0tqN8TrcM6nuUURg/b8r3DdjDN9Pss
Q7kHMRzwkXfvQMCIJ0kr8byDkgAa6oq03cVw4onhSpFH8FLNjazpVzipfisVFhZkq4fa/UVGL5UC
So3ufZ75GOfgpN0wiMcFpZevAqRWGa1YpD3AZu3BTJp9PkT5iGzC82lNBNNCeUaWZtn5gVUW57Mz
bE2I/DtY6D3pK7hc+H7OSTCWaOoUEcQ8NRFcl1IlTAVAwJtnYDduTwu7bloy/3hnI2HX0ticcMEB
fC9KbzV8F3IG+K3Z7g4yabF+i8a47Z/NGz+h+zKRCajBbKyqBLDhoP0cUVzPZM9Qe5gtlEvNoDjz
+sDAiHCMqtKZ6v97J+OGHC2runPuXAtfrG3o4JOsreiJAVF+Fv0o47Cg82X8yj1G6anokUbRURkw
QZ+N+l/kWV3X3xZGROu+K97JL+i91wAsed6Hgaxv6Kw+YqEZNKiaEm1GFmXXbijMoQmxKGYgtU9r
euHpkfmWD3HV3+4QTfwjp1v76bWaT++YtsO2w3bZulIoP5Fa7HyqPLhvP4kQBPEX9Nq0EV8fZn98
MW9IQ8QHCeQ0G7aDfkHIgyYh8zDdtzn4q3ZH+Zvsat6PVX//9MJl39HSncvbeV6cTkFJBvKRFcOJ
RpHtfFhJHFyDc7H3i4PNcNVrXU75KjLsmvYesMX5MOtcNv2p3X8c6L3zgxavg7HkNEvGWd7CW1CW
HPpboK6KK/6blu7xjsitKF1TJ0RZ+CdwBx3YL/KsjH31mx3eBgIecgHGlnayjU/FxPdl1KIyqEbs
IfP3KeVxfwL45+dlX5uG2cvS7rpEcJYFvqQRFjcdybybe56ASrCmjYPBGCwu9qEdHDFvx++AbjT3
Y93QrTImQH56kNnSRf9YkGuGqWqPZeZhFjP196HkYAtdFmObbQrS8rA2Vo8kBxf8VWyhOVfYvF4a
d4cAj9ruQf0qxvnJ55apby1BYURXHsZ4/mz5q1shm7w84sP38mRKbC7Ke1TM8Gk8IIXtWJR4u6So
JNplJLfWiRP9SKXznQ6JZXRJBrtzzfUFWGceJ22IVuVLRA6JM4vErFcvWvQqkk6NYOJaSkfRmWoa
ZKGC77d/nzp+rlPOBc431deRZybwrni80u9GyP8n4vN7K3gdQnco2UFpCDXeCEpSB/k/msoSJPjx
2yYCFKH4ObFM5+O29rBtASzmaoO2Kd7R4wcVflrh44Wp+5zWrfrpGgd9+yDbSjuD72wgLfJ7J30D
j5QjIc9zjuacKQl3iFCvAm0vEYbbtuyR/RTS8kMf0r6pF2FMoh859qRkJjio6xkoYbgsbXlJ5iUA
ueD1iMN1Cw5GuIUx64yPqeLnCH7GQVU1Aj38th89cAYWBUv1Py16+0oX3htPczws9CT26btt5LZE
PSQ0YMqDaMVh4SqOtktx0cVuWjwGHz+arB2TuEViBS/24FSn4anuHv0oeRbQaV0qxnNEYEiWli90
kSMaYB7wblhFsMvUibY6+j/f69pznkb7zmg2UPIVoJmfpw87GD5Fi/n34U59orzZA3syi3rcj/Gj
aCw0y8WXtQaE+DNvmiwsWm7muMuZXwaQg2Sm6lhQ9w31J8+rN/PYZb5mu2JuLWg0I1SGmTnm6Lxi
h+XwU1rCXu6uNbVb1qKnCzn/2DasLrCLFOy6nfvLoimhvaD6YduhFbPmuuv5UdzA+uW/Ya9NC/0/
Gl3uwEq3XLj2N/N3a77v3FTdUFLS72scnQ1egliKdFo6SXUaF59hmYgLmKFYyRdma16A5A/JU6Bz
+XW3e88LQHhPEHguFrZl0IG/pPDeYFtL0i9p2H5Pnm7TIHfzQOOcjAflTlQRfsOS333cnoMCgWBC
B3dJg3a6kSpwvIpJOd3tDzA/48O07GG4q/ODavQI+Z73XzSI1sgigZlUZxHzau2AISK4kwLdswNx
4CwnfP50apvKiLH20HJrvcCSyJR0uJG2VMgq7Kk/GQTORo/3rIo9nWbrZK1SJShM2G4BdFDdmGM9
QPGiwahwikWSdDMhnTnp4Z/IpBk5J4v1IAYq928vmET84BT66DdIVdHoRXrmgI92R1TzFZt8kOwR
wQe+G24kMAGzYnu9Oq7PRpW6IDrEUS1BBEdqKrJCpL97vZf1n+ZVoLC9KdvSrF+27cr+jqyMOuq3
uNS7+V5nizZMLuzQrJNkXXRvQVqXBUz6XbfX9tvv2DS/rXx7r/Nt7pzSAU9P2ruxVmFlFqZwbeJ/
JNqqXAsj8U4eATOGIB71y54ut9EnNBqtlBO+laMKamEGXVXv8ASkWQ33dp21nTV/oQTJJhZ+eKlN
inLJ+EQEogAX9xC+e004ja1ZHn2JM3mpKCLvyP1sz4MCBqgZYLb4ThuesIpj7tx3bHj3F2D4IUyT
BraPJhQpE6p9VrWL2I5fcYF3JboTCST3lb1B1XaQEqCS1CnL3D9iefsKBTtN/VcvMBG8GRNkRx2U
AEegzeNb2koq8dXa37YTg+J94myt7bF21QvurzaXlGR5LfDpvCzg8/yr1QgBjzECLITPqxFTW5em
TgNNIwkcTJm0UL+AIauByRGUlM3GA09l88cQHlCfvT+tl0m1q5clREGXFCjP5CRbHAfjDf54g59c
npxNgQeXXGmQ8OSEL8UC3fX6fRDr2O96XdjXYRsFAnAEbp9skjEaEo517ccw+oN8e7f3/ecR5dSA
91cDGByN6xchTbp+cTyJ+JA7zDetzgoylj0eapMJoM2WxoY0a8lT0Y1bykEqBLk5MzLePXutLvjC
5coQxk5O6BO/dXxrz1W1vJCPR6iu8Wki05LlhnZwQH6lBb3+VTU0dU2xf+gi3grLDuNK6fd3KPAy
xYHj2aggMjsIj+mmBo0uHJrjJ1Be+ZqmAW0zTNbp/bxcVdINay16ijn9wmqlZNc4lXwlRr23NmpU
tfns2tJGXuoA22N2w7AzO0O5xtT5LJVlXDmmctv6/foqEX9GwBGf5811I7N7QubQCZGYz9EHuy+j
AKGb8J0/p/x3sfYO57veXW5uCRPaVY8PAnmnOunPGwv1OIxBuxnJ7GNyhIm4uZL8GFX4FoYNxHnn
0I9h4BW+kdDq8qIPE1yTnxURgt+EEXrHl7O9r13gPDQjYevqk/QNqoEn4W3KP+mQ8OAEruABGBer
hnKq7XvAgzVIfYRO7tje6Xh3tYYofQOZjfCwfMROnobjZxMHiFI7xuhVyWuVFQkKQQ1YczFVHZh7
H/uyEnY/fsbS75DjhX+r6EUjPu8mmrWrbAOiGFnYsdQb7N19iLZ8lLEOvdIHBTgu619rEkig7MMA
HXz+gXl0K+AmlCNjf8ocrrJ9BdnRHQGfaFpg2wltsUoHADpyESY4ytU1NUbousO2gD4lg17WC46/
iWEKeex2wpU97GZkRm/vU0VJnFsesaQH0RK4e3ZORyaPWANBsA7++ygclICkx/IrkmJRbbcTfFGM
IFFSjU83VYb3bFjIYwTRXWwVHBdl3WST/g3YU96x5IV32qwmxE5hrKSgB4YL2MFmVu1OH1kCfm59
CiSf3szZKL7cQmYIrrf5ja5QiEnzMihJiUAUOKopbSulQZmY6nVmWZbMZo8lGZqZp7e07ydUwkIx
+vRHw5gIXtcLeki7fmC4zn4WM7Uu7VTNH/ka85xI7a4X0Dv9oVHqdoO7BpNgziP1P+Sjfk3vbWYG
r542q9Z54qfEZyq3MCA4llbFn8M8xGrWf2HwBfiKrTqLBXUj56dK/ZAxkI3jtkchZ88KDuCOi3Ty
fuSbsKmrmrZiKYo0ni0mHRjpCI3yajfms1Duu70RQASsGk4heC8D5EFex122uvlfO6A3Wu5+FYRi
GTsCTVsH1i8dK9rD6LUDr9D8OvGN3yxsV56QjhPYzXkCtJtS6v6LthECC/FYVNySUdvXABqSqxuf
hrbDqp649VK1hkSrH1n5RLpaYHj8Bqs9LLO3C89QFpk60S6Qeg29hv9xuZTvs0Yd/cfTF3JnQ686
GPel0IYy1O5hi8oYPmOLe5+1HOdt+XbYAPv+uBwH1+U9HTf2snfCv54juAt/6mDvHwHyxdkzrqa0
SM5gJv3hhDA0G2R58NsWrgPPmeyBaO67rqRA00BU/yOFhmPna+vLa+XTiIU1d292UrFoB6LqLRJG
yvvSeMU3QvRn4BK9FR/sc7WQ8fZtD9F+qKyQcReyIDwiFBvIkNeW7+k2UYGHr/IQhYEeqxo8Q/C4
GSZ45MoUU4M3KExNxezBvRY8zNB4Wc06rl/c8MphzO+so9Y6L27lD2TpNqQGgpeKG8M4CrVCYPOy
/QQmoz9j5WXeOShaNoKIqQUPllNHOBiMxzar+wQOEu88YQBJuC7dykneEPEOZBHFswfbOWC40+Av
aeLV0ZRjrmhHej6t0UXdEJuEgYYFEWSrRW6JrT469NSRIx/rmpY1z4s5Gelb5g2hCn4G12e5MBKS
B9ma73paT9o+V2CnL6C0uG9KmP+ZScl1guolaqgoeJeQPwTHL/7WGcIBqJnFCqFpIa5UlroLWn8Z
rTJJIqPOlbDD9qOt211dWvIQVs6YasOmjKPNxqVaH8ChoZ56Zdp+UGor6T1JkjHZu4cANSWy6/fo
7lJNNvtsEAVT+bxapST5sK3l+pRVkNeLHJ/RqQPSdcaqc0LC99vJnlND1ffMqGuGBS3WQZPIFWjr
7W7D2x8/YOqfY8VOBVyjo57GU6EDNk2naZdyvkn9c7xZ1ozryOIe6d9wKQtwAEDvGaE20X7im5QK
tt7dSmeevoLTdMyVkUdqzFHlCtpHehsNAh6u4wmhpbyLOPMbRxYPrODqsnGMK5gy7qypWT4U70bk
rr/QcAqHi6biNslIa6jzWwTuvOfv2ZwZ9ss6jEPAKEzwIHlFVuoTVFgyetHKWqiIAdI+V36cBRCU
ouPVOQl10sB3MKhfxOklk074iFekKU69ZdSMhRdfsSxdy7Sb88uxK+TruJaGwzVFWFqz7+DN008R
+luADC6QAQuOzg/McuaVDoVupRNWDtgpG7SJr0IvnqNzCusKsWr+umBLtxqAI7UvQ+u01/RLvCA1
zslg+EF8bkC+DTx3waF3otkwkBxcfzTIvUCUOIZbKHfFOPgClE7VYVEmPnX4PhfcnrXG1hJz5nZz
xmyirVqD+HwAOnt2tdfKwGxIW4Pzm1lnHDMRVKeKLbqzmM58gsShTKNguWH/edvwv/CrdHtnfskY
v2ynR/G89uTqXsm2FIMNSCUEAWzVKlyktraE5dndK4wDUtB/YZfgMmyV/M18JnkhPl6wBPy95wG0
6r5qK8IREUUQqMI1QDBsroc03JOCn5ZnfZxj/wyPAyvFtBOegrx1ZZZ1JU0I7+mBIkSdYwq1ddoc
xeP7ZS3XyVPlTgZyrAb8zQQVbnPMt0OukQjmHeHoUYTjtS9Iyi33u7fgh64THb0CkX9SA129qn0U
x9D2N59KdK55uzxBozPIsiD+T24/xH7kO3Z/tVnr6EcLyDUAjN3qnVjZb0EOQ6+jn/wTG5bNfRKw
/hqk5rRCxHbVczaWRDOh+MoCryaxoHGCg+DxUdcZWL+Xytn6FQ4IQDn1vDQoKvYfiBcCg5VBoi2m
jjFfoZq4hMItFma8nkYS6fcckWrlPb7PQ0GrmWHmBY4Fk1KKXqB3DbzoCWCJVtVUk3OLdzDnoew0
t6P+iO76NsOHokGMiOA45WbuC9S7J28PnJ2q+RSYsnc3XaZGp7S7KjTuyiKRevJXx3kOuJsHBfzI
sdJYjSd/CIfN6dqMZenjwC4NIFK+twSiMT7u+PJ4oi+b4ufXHspLMBUVrqqykYHU/YvdjmxbLGU0
lZdZXka1BOWS1JN8vfmtCTDea5A0OTDuaf0zQaZ+tmxlPBw2Uv8c2m8SN/GtkJ1O30OGXE220xdI
hMbZVIcs+CYqNQ7BinArcZPMnfnFqRBwBbdqvJ7cS00C+EbSn10scJynQlLQkiBKpyWErPjsQuXN
LRoeTDdz79O3LvdCCc5SC0wd184pQCBlEt3eUjIyT4jjishyyrUkMxMMjkkjjwTcI8zl6om7nMz7
weVIg5EfQosyWQdqKy9e2X3c+vtztarMdcocvmAQe6O9Xlyz2ZfDzOWk83iRRDGak+mZotN+Nt+y
z+2iHOrObGdrcnz8nPgv1C5rD7KBFMX7uifuO59SZcI5LrhzhbJ7VdEA7FXnzVmyNJGUHxx25p7a
a2B1QMXUw/6uFhYgLmVJ8gcBy5t2Z8xLEkHYYC5McTvHb9NTV3UVcRb6EZIzknGwXDxb45jVGuUF
JCMMYvX3CXGI+oxIgriyJy2msiaUocR7WHnua40zwCqi6yHBWu11qXsQ1gNrMzNXgthQkRIzvhGp
f4yX8URyPO+Awwd/3n0lfAcDcs4atG4MDpslYkybod1bOi9SPRd46ixvKjlD+J++cv+eQ+eHB267
s3tRhpY/uigaHwsHRnVcb/1XRhgYcHDscSkpnrIr8PyFSDSQS4qkdfEAEGeE+jkZ+9WXqKUkFbQW
9+5ncn1GBY/QJRYwy92sl4W3M5UOimN34+UOFVSp8psoIAdnyJQUxPKQSRMKqQFD6hrdnftgb0sP
TMjAy7dm0GfyWZ40yqOPFTltWuMED7K/j8ZcuXKaBL7tsW02Ofwr1rqTGQFXNQRMgQb2JG9ZOBfJ
9wGN8U+6+I20Uhkw5diz4czlrShRKQcsCe+kA4gvMJSgJkIcn1ab2ssy5gpfDk+SYE8yQ0k8S1NS
SmQO25i7GQZvqR5N9uEINEblhcuY0wk92/cSJf3Te5hXlKC6sH21FUWR/0eEO0HRrfde1xvqoP+c
IScxvd1umuxFw2YcNCRcIFHL2BPSrR745lvA7mw6YuRH40LTvIU3cIzHL97APbqXVO0n6IbIH+FV
VF/IeHm/Au7r5RBVnxcBDKzL1mPlbw1L2PvOmE45QT27RnxzGHa/u6/3gFxhuiqNYYjxEH+Oqoa7
z6Ib+uGCQaFyq0hhI0eqcIVKU8cmuowWOXbDT5ZNbHvD8aZn8zq3cLbiE+z/FDaQabvMUST1EfFm
vKsUp05YVjFCpd0kjBfNrl5M9tHYjgJhypgZDg797FZAMASCad5GCPB1WdJFoGTJzaca4D2XPYIU
Tou2kV06ycTvPzJPwos4TSACNqCVMGhM1MXVniqj2a+MfezmdlAbZLRIBceBSyhwB76CipiD7qJ1
LDPmUdp5S7qRFFOqkP+EMjQF9NKI/m8/z11GxQtHx/IPN8N5uoju1wDsutFAZu+sV/64zpiiLiH/
De6nkJuoqnxL4V6p/cmb4p4SzC/9ff9hXAHt8tpYnNeS6n6odChlUiWO0D9/BM7Lu9jkKaRS9aHs
7tkjPj/XEdYb0jmGqMn9Zj8Dq37VMTuhPQEuottCYeKizC9oz5bQxxF4yG9yXzZbxgBCX7ETMcqS
wI3xageJxUYdPAK1ayP9DOmy5Jvj9A0LFvb+tRo4eDU0s2D4SF372T4J4RpXLtKutjU3mV28m12M
0dBMF96VPC8nX3q4I0cqTfFkWzAhuZLQNreMxl/ojP9uhzDDzqd52BgBKj7y+nArNh0m03cJbiX1
QZKZBHc4BJUp6zR7RGooxXy8mFF+P2HMBygebJjMopxww10pZjXdhdqSdSdTj6VM9HjZsTa9TYwi
jyapmprLckJEwUIfRZe31vMj/BkKBA/V4lWCyF4azs4p5P1hl4kU+FxqkP7dGIZR5lVc60i9zc8F
xcPbCe6Vcmq8fZsT4QSpCaQSv8CtpKVvcViWb/koIQljHTFpRmfdyxREZe6FYH9boRQgMcFULHCe
3xeNX/oC7oNy0Y5Ro+JfdZ1WgAizi65WzF9r3oWsz+QF1Tm5Bd9+qf0XYp+i4iP3qmqzJH3IXkdg
KLeORfmgx7/PMOtw0NxlHxc0pTCuBOW+x9400Yl8xz/g1exTKjyRme/WFCjg3lEEyvlUfzyfOB5N
6dO0tOvMbzq20hD22kTgb+glqHWRc/g1mmfj5K2+IjQv41cxP//0gNzyj1x3Re9nuJBwze++7Y2W
irSwzjneXejOxAWt71B3+JZRLVZog8I+8bZDggo9eN9M0uamZ4zDyKiQndZC/7i+CldLBfnGTsMx
Jr7J07djZ3+x3c9HQ4XFqJ1SAU6kXkuqz4Xm9GoAPgnwo9xgoHnAkuqhCJV0KduESD6PjIMhMrC6
ePUTdTZ+5Jupl4OQEDN82NFKPetIssoMz2XeJAOZh+8sN1j+ZlHCzR15Acz8UrVOv12Yaf2LPl+P
0rx+52lMyXc4QqJaBzcYPNyS9rj7zNfgPCulVWFf0RLd8YSQtL+2JA2oPxL/C63aqJ4vPI7PFnxI
HJlkI6MPm/E6wfXQLjsxdwYY9b71EMzDudkxQjawSschi4+x3F1B5cFjbYPxuOpi2K6FdhCzMKIK
Shj/j2zmExRyd8TEjYBCqOWO7QcTyMrT6tdXujPxFLjrOZuVSOobHMSy8mr6Q1emIJRYozEfn7Mw
+15Ns3f4jLJU06HdcA9V4stw4DtjZxWPc26CpZlwIWCedXXBRY75z1Uuw18HBETiMNxU+EYpyeQd
VHRkANrW5w/1zXRc+Q==
`protect end_protected
