-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nIWrM1RVkt51BRSdyLTaMPd5SPk+ebhDAl47ToWak6xqPEtEUxpHABPGr8wZwnN/navajuc7zj+y
slsYeiO5wfHTkVaRCvqtOeo1xnmbosBEHBKFwNyyZORqso0a5SNlemGWfgsqwOErmH6VwXhZPqCN
jAupAITswnRtBf8TE63IwM9DzCgtOCGJsTce8dRho14qT+sue2KI49bNjwUYX96uLf1NiJZaKZ5m
ZsV1q0fbmlZ4KNYSOKqzgXxSYOL1FfWWxfGMfQJFa9ZYk3Pn8Ld1xF7dEeXGmSMEC74NlYXWjrxR
HIMAB59CNIBpTmZXAhj8ZnlecIZT7ona+L3DpA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14528)
`protect data_block
vcvnZyhAbL/Rio/Zu6UIOdcj10K1XISlLY+jxO7qMsy92pUKjKmB/02DAJj3HOVkQHNPCYCT88go
zxZZDS+pWBj6KM/OUWMenEV3jMuHNFxdnorTRd0GnaAe2xaN/knA0uygQoa4H4ObwBNhtpuCxTW6
HyY4EVQ1DXXHNUbi2w9HZZrrlbQ+AnkiGGYgAt3S4NlMtgSQV4bzntErT5FZS98IFhZQECrgcBOa
6ZCjVQ7EP05VPLLnffeRFfsaWdkunTBpM+9SznaUQvi1KlIlbSV/E2C2qyY8vYLlvSC/6EiRAq+F
0ffjUdoJaBHQBlX1zWaN+gb+n8Vm76wpSE8I1LN14nt0D06kec6+PrV/nDcBrv9MzWZQBZCpuh4L
lDKtK4Fb+FMTuDPwM92ScGiXaDCLlYbOyXbS+GlLYLLm9wbnA04QwPCz2Q7g5iAWTGB69eawsarn
OLqWs8Ba8Y4n4fN0YKMNG9teV/Zlt4igAm+Jv9RazFtEiE/hpFzdt22vJU4CxkImkGFR6KW929Ay
mcG/RLgD/YBoFruFz9hSCwvY5cFv4zCFRxaAJpd7kXbhy4K+RNNCLCHXnvE+XwUjBWf6Cafrz8C7
py6e18LxGd0x9tWzTSR2gmoCC8MLEWx6Y6aVkHzQydRnagMk9CnrykE9thgYQwb1feVwj/G4nCFW
TFOpZ4iKUxT74GEYUXwX7OEdikqIh19EE5KVXZTsczBbQbgvYSfSFF3RG4Q5ju1GodNhZEIJBnBT
8gk8vUToT6z/YixV8UbVRxggBnO3Gv9sI6oyiSbjgabGCR9luH7kIrLRu6jAI5V9k1AAJM6xDOxo
NAupp0vKqg9J+UaalPc6vzckj0mPKEC7JAOcvXdvsYPPGcTzSW9nePOCjcvuDvnAeKf+XJb/5wyj
K9iOBoaG5XjoMEnHbdzlHqwo+4cY/aBuiJFDZOG4pFQ00HjrE9vEr29bmCcQ8YR8nEdoxi0KpkqU
KdaPwgVhO9WJTaaKOI6RV4xl7deJQQWRi2u3OpLfNOpxtarK0WjqNdnYmQ/oQekzokBFPNOXvEtg
9iH8HoLa5PRaGmZIzqtPfo9dC7zf08lyCpgFNASR8G63AtO/z6XtPH81fPZzB3SbbgnFObfodMX0
0nhyOhMmCkZaNnQFxBT3jzGTcOgeW9QozWpaIKYWOkw190MyPLS70HFXETkLoUZhWZv7nBGLcX30
LH5aVgdwHHzej1BWz4xIyanuQ1fUj8lImR/tERoKd9fdrkrsL9H3Aht9vovrt3guFXDom317I97v
lwI/HZsSbIxKyEP29dx/HFsGt5r1ZFFg11FhvX7iDrHV7p8CptcnrUriWUHCVS2EopIJxe5ahoSH
xqS8NJyvwAEqf67lKfB4d4q/gyv4nWE9Y/Tf4auskVT00wJWEP9nTymmtqE+aF8xh8ia/OTSCZiM
siZdbpaye5uUs22OJGDnjlzKt6F+paGcdg4vXwZBIUfj48Jb3nsqxt6BiAfh/L1ITGfr0WyMjdL8
uDXs8y2xTb+eq/RRu7hnshb3QjzIdgcFi9s3wT0wwGSR8twuuEndq53OMQYX/IQ7PXiltv7R/JTb
GxAPDwcmtmwOtHJI7HFxnyR/2ElPFNY/DZDHvruRZEw06uc8d17AW8cE6yLY2MudDtXjrSRo/7b+
WxScSAesUk4a+8XjixqAHgMd46FUjeFhDSTEebYpRCnYsS+/AfQkTgsI2QNCVrbNSpWu6xGv3PRa
syw4VQrx8QPPhSUud4xbR6lAX984+fGvqKQ95wal1ImrYP6Rd/cVHk+uphvhgW6G98BJKL3vM2HH
bbnLrimbyXL2whioclFMil60P+cBVRHMSLD8RoDz5t52AiFNJD/JJt5biItSScxoOIiREy6b4VGc
2/FK3gN9u8M2LUlzd58QYeXTbNmEEvW4P0M3YkDytf64saDm+UGNKfC0BVLTJi9uXPaGDymMpXvY
l4HbAkZJZ7TfJ9nHUBJha7rdJDUC9yogN9QY57kYglrgbflEv2g/vi/+xlD865xHuTSS6SPoKPUt
68PZfnH5ZZ3j9kaU6xziWlLidBRFwLQWdmJ3PrPrdDGDA6epAAsUnkp9Y7wdqMN+of9FuGxuLS2j
e2rwpd9/FzeHv33kf7qJozCxoP275Z+Pxmg32OtN//cyQ1pUyFx2Q2KTuVu9Pd7IElnGEaX4+a4p
jd9ch1G/22Tgcd03CYrfYEK7+6G77LAaODeSRzJDT0DtvOLW7YFr51bPg8lFw3chd00FdUpCXSVU
6K5tQQ4tWPXXdM9Sq5Y8SLL7tkK58FAG4r6Zf+XGJHdcVaViN5liuAkzppKNpTqs8CUiD8WHsPoM
9N/cRZvbb41ca2Q9c17QWSBbVhvMKpbNB/mvi/jU6bSsrycBpmf1gBeMJrTKeJFyeBmFFopKl2rW
KXWsHDfGjZTB8XhEDuL2CAQTJbo402xdPeEyoqTibY3JMGClb9hRsZc2EV6k1EJR1tqYBFGWoUVB
1q18y4ILFYLAqvN3akfRNHhUIzdVmSy3fdRc0wk56JvD2NJ2+xRM/UcRdbJk0AlCwko1JjdvwEaD
ae0wohn0aTE8SFDQG5OZ1OVfinS5gA2QGl6kl5mRyCRdTGyeVyHlwBs9JPJDBEJAMpLCe+3D7X9Q
BN1IwtOVFW00AgtXDmid9QiusHZwUL47BcCf8MyXl8UWYAlS6PMFmGcU514J9opC0U2nPPwn0QST
r01B5gayzYkOJFIXf3M6ZxkDk1UrklqeI6S6P06LBfS9Xtyvg4QyAsiTdpEWR1GQ3bJqXuQ7LQdR
B7IrVlwOnxXmJdb/C/2ggm5kZkFJkitPmQbGDE4W6T38Ie9r3eP9nMdqtbrea3gi8z4fLtKyJi3H
Afz7QuiFVKXPHQ/osn3RCyEz6UnBpwYU0DtTlNpBWKMnhYPQkiXXMRvvK4yeM3CJzjloZwQn6E8y
JHumw41/YML45/xg7hg81NnHIpOlNAvJT1KK3U2UxUs7EWa/CvcsIkTTjMez2xHIHi75i/2m6CPp
ThyqfFSGuuTXCbVkKOkTZxj5mSRWdUHLdLjogndKivsGlhyt1PIjwcwO0dtBbTYKWyRILDSBiHzl
Qlf0iKXNX+95PPIW/xFxfIhs5ONH8GlWHL11+2fI/8+C6md4vvNJ757BY/237Q51B0mRBnpOjhpt
rzDV6rUpFLAC8CUO6tDFvSvzfo/zERP/yeDo4H7a0vzCqVsl2bA9GppVTL9dXdOZrBQVrD0GttgL
UOyG6qxOU3R3ixufigYTn6sbbkay1tHyheZxSC8j1ySCiiNXKbGCdlBAQOZUboWy//s8kVXCA3Wk
pBVYhwPl/xWhcTQyy6y/2xmYRO76LYGF9WYgvv1u2BVsqLRd8OpEekQLA5SEIgkEuixa8T1HXYAT
N12A+2uMrFNH9GON5zhPal7aHBKEnYgEemQ8U6PamOYNFLjNrR1A7SItCDgD3BETx9HDlhEQFMyR
RCvRyzS011OFGJza9irZgMOPzwNgoyaKDl+7HEl8hU0csEF2ZX2sgrQUb7OQWVHaWjInwxdwsf/F
vQjWYjfsX4HUx1NCR0l4xgUpKfT7quH01AkcQiFHqcbrRngnJORjzir3yyH6k9by+zGUDlOoIC7/
0tWpjnYAKG0XQTleIS1HGK7lRwLxIlF8V3VPFlXz1XGXFdsredMPSsyUNdDEOxqs4VT+R+LOvXcX
ta+jbLa9QBbvpuDARVEmt9+qJ2n546iYhQUkEkETHnSCscztiG/lLRUgJCxyQ3F3I7ytAs/GRNpN
LInKfVeclh4CAfUWxsO9BT3+JV7kCgLSeDLuOdowBgFDvbCW7BJUSQpMUKhvR9l00weJiSLuhTFc
rfyl69bsWYQ0m3pGm3ltKPEAZqAtzp22RR7xst94C3hh90tN3y5MlXlZs5f5iVcK/36a+fFmDaUL
c1BgZy4KMdH4SIRKF/aFHnktKJPBwgcXgOcaBPKHmK49N7Xfc+Xr4cAQrl6byirPetXlyj2krn8p
J0lSNMV9I5xkxrq88sDuoIn8xxmK9qcifPDqazjQuwZuvuYjCMG9F3/bwAJSDT94BZl1DzSz74Pm
CxTG5VytBfJx5qKRyavEl3FPpyzw0hoqOm+fNkhMHX3YUKW65asz+6g9jaOea1V8M2bosikGJZ8G
AAWoYMHol3Buni3RU+7h9zCAmPSiVWvvm+geKC/1ZSLjVuay83sDjwQURRSf/hAzuuY+9A8DJV3t
I7iS3wHVEpm/JT9lRtZ7TjACjf2PkI7Ha+4foTB6m4LQulCKYaAOymLldXtyYNtQgd5kL2tnvOxK
QHgdvCUbzKYfpZjhMSj3idqel9SG0DTXZcTDF6DkyKoNxRcU5kLe0Jj3F2Oaxl6Sd9DDxsGAuFMi
v4X4/1zYm2RRF4K02Niq+a/RVQQ8Gp3rydoyLSWsV1Vgb7BwJnaGwjYYUSg55olGBDo4XnvK1D7G
7wKzDVurUX8Sb4eijILxahkWwGa8ftQ5bOTA7XrmY5t4XaDy1muWs4L7wiX5lTRSJGla792Euyat
To1voYgZShXyTHc7YrN8WAlyYHW9hYoC0omMwrAxB86Qz0mq/C/Vb1WOXvR58yt8C8AOAkWBE6aL
Is92OSW/2R+zPCJ5czfA7D8xXHa3N6hb+rN+CIPteAxYKBWV18uMV+/EREwK8wPuNIKsnBKWnyID
CHHh+hBcJ6Oww1PCMW/2PQaxzfxOL97q456akaGlEK7HudFKYsO2pXjMLh4fhHcn6Zwi9uE2IjVF
sGx07ITeHNoKRVjPhaHgXyx+6bronM6LmKnc8Yzl0MwjydpqOLN2QSCaGLh3eLXt4b3CbgYs21TD
dmUNnnZ1sHMnfHHzUWKPDy0nuhRQpRQo5fq+a5LVAhMA9J0CqfRa50+g7eSP0/VDsVH+o4UyzVX7
Kh+vXbliBsF6h+wRweUV0MDYdIaSiUCwvnpVYFFioZNL7j1ELiBNOcnOou5mLViWXXYQO9sD3eyt
+LhaX8AaJY9kAncrGQ2cdmCwASJocK/qDcmbjPRxC194cNxlv1iF5cxNyikWUYLZeEi3xBwrt5YQ
GXKl32vYK6BzBpoOaPcxhMzIwZmt315ovw/PLTFFizDeTfTIOW2dFksiPn0+qZkFcCv1xSb6W9KZ
TvAqpJiw+FEY4GRPZ1EnqJK21cukVjAjcOdYIMTBMHYFtxS5BabwBuy9WRkYP2OTRDjKuQ593WNH
orsmkYvJBFJMr0Sz7c24FBAVZ7J0D674JXqlXFi9JGS+44ukZIP3zc3+BHkhkAKJB7/81ng1U1U7
0080own3VD9YHJ2RaCh6TpBpBXe6KGeSdX/OB6dy2XcsugKFusuMp6GCD/mNetxFDaR9EmYPZmFp
0laMMCWyb/Lj/LJGNoD8xGa+2w+ATVg/R0EK858Jp2dnSvrmOxS37612I8ljeiniQqH2JLtuGEKp
qo3/P9pDtl3Kx3Bxx7E7Mm2HngHfuxMaEEYnB/yEiUzSSOVRb2KLmytQuba3KSo37lv5HBt9W+7T
TsaVJa2uUfj90JiyJn0G/CvhwaobUOKrsdbh3WTneWke+SEWSnL9JQP7zUiQ9CFUpYW5tyO6nO/i
9+nF+zCGR868LMoHGQxdpGCNB3KsfnFFRd0CbteDTFjSajfghtIf4Lx1KDN0YCB3RZknUUzQDPcE
KA/ufycpR9UYmRINjTBb/KJo6jgyoj6oAfqMPQsoe1kyLeEc/DxVzIGP6uc9c04E+lwR/sppGTcN
L44+jTpJ3cBSiLEBpZ7uVbahgOlBOl4KmtBH9UtIAXFBI5nZxtte/qOAGnf4jtdvzw4nX1XTMddc
5lAyz9MCtqFlyGf3LTL6Bqu1pB41DyDejQhGSwTPTwpC7Ok/q5rDdNDmGC7N3B7zm5ycsugWzXFv
jNB1HJE/TVxank3dMVKCLqNS0rbNN3tO+HvuHSfranvMN9LEt4vdXLMpI9ea4LQ2YSx6NJnEWD2p
U3flIInUBGWggDL2pF+CST3v/CTERZo3gsCM+pASiR+6OPE3ffHWw5tcQncW16ottFVczs+TYyre
Rke5aD+jbP8yo9LxIDziYqN1PUBF5SBRlOeCtFWpioJ+suc9evlM0LAJVnf2kX7/nEh5KTU8v2zB
79EWDVU0HPXhcNmXMbzHiV4iYYVzi6CKpu0SUgPAjiRPBs9zn7XIqgWXLxFHceNLLz8XW5VS/WFG
F3nhhwgvxCNqGQSCVCd489EGfVivEt2Bg2ZYkVbIC8AWOy6rLwbMD+2a/lNGytj241jpYnBZRKwW
TqkOGMWp6ibHxAux1GQloF1Vnl/B6IIzemODhNYMKTSz6hIuh1zSLyVz3+GsLc3KJyyk/qeYtSYV
5QfbJHaplQfpTvx3nTkCWYJslrGGSYp5TlLmEyLCnIlakQCBvyJdkSXcS0Y3/tu/4G/sWDXjy6YJ
WRav+V5CSjePa/muWT/AOCflQ89g3L5QynMUyui9xXIHvfULZWRQddHWUKoSc8e8BgwnlbuhHydy
L8J1QQcbn+HMB8dHWmwzeZ8jg0P6L4q8dRgEhr4hpRIiBSQS7O8JPVDb/vI94WuxAVc7OBz9+2M5
UhlGqLCxR5h3zLEUmED77HPXvIAtM4osaonwXVoBPE1QsYzUHy8X+A/Mt2GypAlQ1vAueHN5gXYD
cf+tjltxBfzD27QPqhznNidvscQSvtDd5+iQg2kkWSHifoL4N7YVJuRVYcjLtL6vQYwsn7oiDYtz
0SlWlQ6ZHRpcK7vgoAtEZ4tTG23ieQ+8FiboX2VfM3FNMH98qWukf1NAvFUWQp5rSRcPiG/Qrcf1
Z8UEUVo0v7qEJMu3fT/QIywMlUFesVIIxD1DZLN7ib0jvC78yzOG69UgNrc8xfOr4Ip6XQoBMVsN
3pGOWSzWoaA6ow7eJvaD26EIk8dXi8Lz9jTZUJA3JUMW1byJ9CbCY8Q10bnJpvBAXdJnEx1mye9W
+qkg5qUFrDUme6zLtcc4S1vdnyfRe65xvhyNKYVjszgJH6fQb6jxkmH/lDSAl/RciT0PJs4nsgwk
VrsPdoQ4tUKCIo+HFYcb222wf53i/JxkpDhPVgR1XBz+Umk1dzftgSzqxFsGvsVlCT0pD0O/wS+7
Qa2i3qjbodDlmEt9pV4/bEoe+sdvh1e1tjcbNXsUQK1ClxQX5dxZ3GFRwuqQNzJDxDPWBS7q5x+M
dH4CN5l+wlhsCsAQjs/sduFhJfQ6+V3dw/mRTa/6ZXEgtElQyBe8+c/yGdJXgFz/2p/v/wp8P3AQ
1Drg2SCPswmgY9AMFhW8ZvsBxPRaG+LXmt+Nx4oBtsDe2X9Ccm5759Us0uscKkxtxqCUXsbRr/T8
lhMYohicFtTBexOpMVMBULQu1Vc5shTIXICteOpujEAt1NjWfsXG80Jyhlyx9/b774ON5My7U0Qr
OiDB2pnyew0NgRCw95CpmVsAqBhCghTkcsx+rH4r4WCkbgepGXMbHm7mJ5luCrnAno1MKduCkVVs
PeE3R0lQ7MFS59y55lKokqogfNF4S3C7R2+5LokmPZ7DlLP0vcXBfU+V7cY4ri80xp66GvRAnAzm
g/CJYW2PFmpIX3LTombwKJv8uIQeMQfaiWd7wcB78875sMhUrYEl4X/XeuD5kF4YHDUc03I3KOEN
4I+6M7JaboJGv2vSSiEzk6E2+1wbya6X+sXVKXwvg5bQ0PvotJwJQg8/fYlevIw8teta46o2ELkb
28crwjQ0Uy5F9m1waYYpirx52yTYzJorfIbKcU9Rf/F7ZZCoJ4+gqt5XzmSwf94QaHUVJM5PJSUI
jI1WVfOTy+9S/KtSxsWRp01TIXPLg9ObnM1gmFqOpV1sikP4UgKhz2rTQT9RyQ/TQxKhybugTplm
91zQTGZcsPTo+NIhdO83zegb5W7fK3Ha0pSVBUMFTMKnvgTj1vdtoGXNkOckoEhMIXYceDBB3bnk
ftoXVHvPtM/vOj718s7r0OM0hs3lQcGTnUa6B171xRqw3WV8GLu7qDQgTXijXMiQjcnHvu7JoLu9
RrOsXPM40Ilh/DmgSOSaCpi169pjpm4r7V6vXluS+XEMx+rxa6qshQDZgAokud2aj3zb0gBsKrqQ
HiYm+HmgZO05v9fOLfQoT35I/QHtqXJ58UYf7PcZ2nl5x6z0sSSBHuVVPQLFFg3Gz0mfdAsQY02S
/sjTrs98+k1g/cZt6tbxHp0sAieiEIaUczxkX31IPecdC+hqFouVRot/2F08FtAhw/k6c/CG06rg
RIMS+HO3S6so8N8QvCiLo1efnihSLnWM4pn82GUJqko94HKMPsjY/qbHmrSXtmcb4GY6qEm5wzTN
cBfEDbj0Cgc5/mdCYCO58H5A2JzU0j9vzy4e63MDG+TuE4Cs+RRbx7sXbE0H8N3IZFl1XY+BUY96
PNy085w5WTVo9rZv/HjjVc8fQtdhZM/ZMC38AxCqoMK4EpOuExLopdPAkXFkJ06U0W+o9uCJaeSb
XF+FqQyFuYtyuoOtu7ltmkVUeoMahe5r7xxd57GPXMCjKlBBWzHewczbJSadsFq2mWE5Im0IGE+v
xOuwOpKwRcQQsXm+KezL8qJ0RmIQgZDojc3nNaBoStZdW4FZPHFIhaloAPcnPbg9QvcrggYGv88k
IkQhWO1L3RJIYjsri+rGY4weQ5fn1lEaajAiN50kGw3aErjCH6imdbR/g+CH8Li65+Nu4mHZ9zqg
5hCAGmojRvk/atKj6N6uO042AkdwOiTKwjbmj85yJSCwXeAM2/abupYhbdhfa4TbUifv1WLEUd4D
z1bdXN1E+Q8jRmETYTDteCq7qxcu7r3jOCMFPoQQ++DoL6GOyJFFMQFkB328yxtQUqBHYNctketo
HJZyQh0Bk2UlDiwSQ9q7K88z7prYzU8wXrqb4bea3og7GjSdWDh7BGui4xvcyr1lki9x11+kaGWH
5J77YlNIIdsDx5j4Shb2m4Bs9Ey/mOickxQOZR1haCTh4o8f7XOjntxsR439SlWJAcC4e/U/Xp6w
U1XvdezV1of7DEJAALGVgRA6beLOwTvAqKRofXkZl9x++vU1AFUEER6tTqs7FBcAvQ+TkRIUzdUF
XNRpuanVBLaVs3yLlOVqBBuQ/w6kiHSwHQdEd7ZfQkLhm6FVKt54QF77/h7jKicGxctf2ZZxVpgR
JkMQSIIIIy296nhYNOLbzJT2aqE3KTub0U0wyPgT5REJPEHGx2q856YWMMicA5PgEOjNMcfAmh0o
WtwgGBYTpytjIPz2L7DcOL4Y/uq/nanF6xyyJ4tsbF6iGL4J61aeDFi7vC20TbIsp9PkZ4ff/JrF
WQzcRS0EwEd/gGjLWBbRdAf+xMQgmquU9gIyorb68OF3Swb6ZvrVTzP2iQJaD1R0D2FAso+FfYae
SLyRhfG2c9xxB+tgbqvyX6Rt8Gc/HbV+Ww3jmlenDe2dwhyoOIccoyvUQBl0Ercz2TepIUyKB3+T
NazhKa/1pKQbeveaOw635RkhdAON9BlOQhzNVws9rhO8nZ2b7814lzpJDxjB//OTI1ud/FrJAURA
by7t1XeZRgpLaFW+Z8LiH8QQBZXxejguX16X6PZ0zv8haKX4UUJgNpdA5nUelRV8XyvcnX+ZUQA4
nsgaIvfPquGwuqyBMOjAxpzQgGaDvTbDg/RgSdoAt5quqZFqhFzBGXdKZoqM1+5+nPgk+MRd8OcY
U1Zx9MU0LIH8qt3kSjmZWWNEsYEa2TEgwtB9kZYc8fjrk/Meb97bfI+Nc0WG0VTBASVwJDMRECKn
DQGFQcW6iNkT66Sbx02lJhqXOpym5zMcpvoXEtwFPB7FrRQrki5u1L73VWUR85Q4YRr1qwdfj+7B
eOUBVVNfdeV58BzYXHyuFvLBrJyVrth/RsA4P0dVVrvv26nP8+EeEVWKY2bxDjpltaKLF0sxw82B
At/uVr5fi/INQHXdf/vnPXTIdlNaTtIEYk77k1i1awD0/Qw+/68M8kF39YmZ+DXRNBihi2O0BZvt
FXn7aRewDyIVcmTJcaAyyAQa1/UMCHWE0/o3a+oEiQdnGBEEEY++NL9eGxZv9GxCgGDV7YYo9onI
I6pyaImqQaMJb3SjwHLkOHpHUYUvy+ejLlUgAwqo3JuG7JLrVY2q9uN9xmk5RBHsBNP4kHR8jISF
I9vD54Bd54YyqK+SgSqFjcvEeawDUv6POluvfVTCcKv2GCATLuwxyVrdWMO79qxuc6ydb1O7W4J/
sp8j4bn2Kria3s20Od96g9V9KNDQ4YrT9181vZEzERvV3ji+CqX6WCt0c/t0ndFmQ6DmH7blZOBM
haPQWh1i3IIcHAGS9KKCN1v+fcArFx5YZcHjKa3odz1Ai+L7arLHgajxoXFoo2/hEiA6pLOB1JLC
m2OCzIaWHEDYpK8ocNcSQkNG8JnzyNtcMy3XjI+wDgQcRIFfjn+YGK8MdwDAHIfH63Y+/j5e2oV1
FrDIK7Ia8C+KEPQdpp015hOYpl3tz4HD3WtJSENKTdCjLW+CoJc5ZoyQbbSNJWx3JFjV0/hVFf5l
ywCpps3T1YeMbVWX6O0atQC/UsQg2HwzAhnW36bNG3dNTh1sIwajMExJ2bDaluP+FzB2eKVsQvaK
4Wz6XxMfPy2dpP4x0yqSrks43qD4w5BBgaUA6ptVNrLT9ka5FabKxobtkOZwEt/NAgwEtlBalyJP
apIyjlZgziEVYqXVAMPnqVwqmOMgOiC6olzxBQT2lsRyaGeSGQSoajKpSbf1eMw2I6QL577JITRU
naXjXPhzffWMmwXLC3EK0E+SJwmCjjaJoKXb9tAGY+qR6MlzG+o+gyA5TLMuFe0CyG46ypnHA36c
SKcUdhazcMJwrtRad90rXg0pS5pONtMpEsgA9+JZADnC3MV68NWjm+4IALNJXWbkjYvQX+qpdKkc
o2D8hafcKh+e6BWl84wRwxhqyx8TmpTPmLwea1UL8ijbFQVfhm6S2hcsz+rSmpWNrs8PT/hBKlIZ
8gccgPQaQFu/tyN+5j6271GnOMrxzSwYBAJW9tOk78rlJMYt9u8SjW0CIOPcC7ItE2h1w94wKm+f
qihjWDqm0OxPO9wddYa7Cn/F93s/rqdv0q062qWIKNp0rFYPu816oNLjp/u+P6ZUKwKEV5ZFHAjY
Sr7psY96tUrrqmaIPFVQiY7ohVpt9dygt/iRHBaUxwkZ7ya+U5MTeuPGnxmPwG1cofV8w5Hw0JMk
rt1io4MTBC/Dlfp5e7DSrlr4d6PN8alz1S/Imzu/JwwTJA/qXAk7tbsCsgk1vXmRLU4cvlwvpaNq
4oYl3OM8FYxuL+61sIFkOYPdbVXHhHg7o06/QaaVeJbOHXPoydpielG7YKijJ8VmqY/AIFfeHvPF
zbOLw8XyjfhKMLFj4MN+t9FFoHJFMXLg3mfFR2PoARPK03r5uRvEQoW9AvMxFraBoVwoINqfkNz4
w+46CF40EoqY4BHEEBcDr8WrLr+TxJD24spjR6AglaxTsSWRNxIs1CYVGSI9xuyaTggtPoykpwlv
J1U9fBJt+M9+UIuY8CI1X6l2xY1frMxGRT4iqrkF5Yf3hD+8uhk5gcY0PJ2oKfeXcIK2e//It6N9
6ICJFRG5yk2qwTLTLz5BmOeW8Bxf/+bhZC31R3d0me2blJoYwH7dcRCXEEA4lgHS6jDjccj4Fh41
T1k16yJ1rqpPcQSYPNK4HSTFbS4zO9y46p708ilMFOnM3S8tLnaPNmx3UDdIALRUtsalmWXPpsRJ
nVgDqUB5VDT3wrdQc+6tOQ7Ouc5+cjd2zX3WFkr9Vwp+Gvtm+2eU4ud8bPT21Yi0Y8veety8XHwI
5VZk2d3L6bq3lfgftX8YPmfSqCoXs/JafQJNasEuq4eXZFzV7DlybSVHx9LG5M+9zwE58TaG+pfg
OlgBZNRdTDzfmANLMM2Gu9sEUZlV6FshV/1OfslQXiGEVpKTxkutnkuiC3z5zsCKij0OaftL1QEg
+KmyRK73y9+cvceF8YxmLuLukhHUfmqhdFu1fztC26YHxnsnd4ZdRtvHMvFa+Q+ChbZY0vv6WsrY
hrzNq6zHXtQdV0MVugq3RF/tTaMI5YgAeL7czfiqr9h47wG9STkXpedhP6ZKMY+Hhx9vE/8bSOJZ
kuS4qK+/ifaQSnrXY9lj5qgMWtLjhK/22Ai3HzWLclR2cC+H96CDbOHonRxNTuIN4hIYBTQTHe6E
zuPDrFMqsKCGj+jXOSB7UJu8rQOc8UXKyewbRhpG/72x6Eq0JhSVBl6PK0VLiTfEyGH2s0IhJjls
2fzAjhXWKyLB6KNqILi8Sacgh/d2yt+yWiEm5+L8s1JeAf1bDb8hGvVGo4ld0cLaMc1q+vvBkbYJ
vnvnRhZ/x/0ukTrrth0TQ0cGZpvdohLY/dBQXE6tgV544+A74A/pfCsTlm9UJ8PENYFe5esav7/M
/bTvYP0LaujyKOCa4WExydy2h8olcmXFNujvMlJDxFKkQmNSXdf1TraLhWpdmKGk0SugPDcTjmpg
rhaePYhn4x+zkPB1FykvdWQ1w/f6l9Yv1oXESGwJPQRWj5wF7Hd9l7CUSlGZbkT9imVdSf9dZKS2
TzA2nQ9snKDpbmz5KgdmeKqP0LVVs4+1rpNofl/Udna6tJRz6svXklhWLlAceKz9m9gb3S3Fqj+s
KEXlGFseKyHEy6I5ojODCrACv51fxkDYiUoN3Gs2uGTuiiTzClqKgbwp1cC3aGU+0LFSLqFaLnaP
2UhZJhDAnbi0dusyqiTFUMCrTyAZCPEah7J26QUQJ5zb+05MHyahFccO28DlWIb0L2wXPCoruB7X
+Sg/jpH6oboBPHMA3x+6z5qiZQolJGkQk/Fca9j9E9FpJZEdFdC9n2hBxGPYyLZ+PG2JpeVm1U8w
mG9XgE8Ofr2R57z6v9h8uGlFt+ueZ7Z619j7pDM3ZsXhkab3K8IUEZylru9fX/oJ9k5xZyU6b8Av
w1U0DDqc0wiczUQvNveKLnrIoDvyhCbHEoY6Ia9BuLL3d9B+mESqUq5YLeS0YLSin3A5BAzukxRG
i+1oZPgl605A163PXLlaXPLs+tZREcvP86huHMdY7dMAf/RKyXixiEinXnYV8+gCvgG74L44Xw0/
xlnPdZtvGzleWF3BuGiIJqSK4iubgNYKzWQFzsmxv3TvwZhI7gVJC0rmmSs4EOKyFhiGJAWmXTWD
1SDWW8hhEzqi19qqHJh6DAQ++utzb/5f0/SoURMV/mKn6sakwmqaDD8yJ5ZQKqaDmsejIOC2ch8n
94owheDh5PmTLn099w+ITXZPcP6gzzEy7bSy/Ab6pozsHKjrKco343Fk/evqP1lggrb6Ba4VvuXj
jOgR/Ld+rUx+Ivxqib8Iu+6zHaPxudt6cyC9uwfKURRsHDIHD9mtoecLvivFRvgWX2rUaVkIZDg9
bXAoAuRzk8NcvXWHFS/aBGgjcc0exKc9nnqjtJ+Zjc2Ywkjon4WlnIUX8xtSYsfnExRJutdXr33S
blaSoXlwr5SbocU/xRiGPlqbilOX4XYb8plE16JWnWNyCMBaXIz2njGHk44elU1HnHQ9bNMp2/TY
pzU9A7xxIOIWuaHWNpwCmEopFRjTco8Hq+7KmeAsaFfMmzrnF4vsMg7NaIT+5oLrVTrImaF/MH/o
L2fQbj4GqzDeelHmtrrE1bnfbLq6Jiv67Vrcp2CzRTt3RNt5mMfnDWOnlUZwHHECfx4/RCANIP6/
e3s4AodKB+HqDI5ipLvpiimYoMhFiqBSBkZ4T7dtgn5ux5kQZMTf/s19gemfhwsABuHAInynqh3O
Y8zGmH/8PBdApqPimJjQHnZBWk2Cqd9DaomMEkQFN1dnPoOiZK9VdtRX1JHCjzNN9ZLeNlxOs6zd
v9Q32NDNezRzwk9SH7oiXp8K2CkTxuHEpXJLQ6gllzWCTRZEdlkv/GeQQEBRw84GWUezw3HxsQB9
6SwfqYg+BWIuEQinFVTXM1J27qpjoAnMJ9xqJGArnH/EVSEqAAwc3E4U/xFBcI+vlHo65dwts3vA
dLePDf7EA4Te+Am7uxBpchiJNRdIxZerO5FKKXhj+qs0+OKQlnMy1hX2vuWP3A/3z4+LKH9ItIsl
wZUb9qc7bQqHS1slxf656FnzHfHzDRxFaOqFAPSP5WNQcwU5Kitu85b+Q7Q5frnJkBEBj1URt3cX
3fX60E38J3p27qu/ajz+606pNpm+xTuTTnnVACXK9oBNtQ9O51Hv3GMGeLQw47UsimjHys/kE5q5
Eg926V5isVTr+nLSbwc22s+Iydp3vx1S7JIrOoFgquHHhcnyi5r24wHaYMEkkA2A32L4cj599YHN
1g+DLcHgEKXeuIm/tVKKiNJ9UWPZosJkyN7HbvABnYo9R4amgcnqoMUpvlSL0iyWKwEJ6B28Slq+
dDxpWMXg2ZtSsSEGaRf4fAjC45rsiU/o+KXq0oDGAtGf0W4fvo9MyuT3S1zGErtDLugwCG/+yvZ4
OUIKJs8jeH6n9q6FzSI1WsFTKHdYL5cs/1Sywz3pe+ELQkAcQbwT8OLmvXuHm/z+qChpoulKi0Aw
yyk/E3Ymi4yf9jxjZeSQUAGYja9NkgDObIwAmK1WGWzY2evRuSRmAbhWd9XOwp1Sekk/uxUTlWFk
RxzDu066zCP/O17zgOX9Nl6IHda+FywEItsTB0sIERUDbEdon7kmcPtntwILh2YpQ/Y9SyZLvNj0
z9rs34NdyCFlR5ct/9a3kpoFegi5HbKnjy0TMj9MH6Y4zYpuNgAViBohPb/CpsdvZdAGq71frxeZ
uVn0eChV/idoiMaA2dJ+x3/2HaetQXsGUzDBhhnNepzTcK4U8bZb6GnrvGTWQ5O/lazT1/eWIUa+
jc9kmFaI+UB+tj8MldylKycJhT7jGuAOpnMh2raPuU7LCLJzA8w1G9W/fak623THlq229ecqgd68
WCbMrt0YBqh5puVWY3P98DO7bHbFLuagJlbQr7gDHQB1wj6Om1z5fSwFK+3L09/4aAuVyoMI58Np
p8sWMPanSk/FsT/1JM9r2AU6zbYw2yoGBKrc+2m9HnmdF8o5ILPbedHjfBmtw6FrRUL+HF75n3fU
4AUbokC01BmITQ7/SyZXOBar9CHsaJ7lWH04PRU0s9uszbqJ+M/T2pUWWZLUHSpoLZ6zw8Ldbq+V
Ch+U9vEzH1zVkIBM7ATRx+Unx8VwsIoBKjTLB1iTT3bvNHkCELFGfFIBu9OA2s9/yG0RJYXqfgpZ
6I8fox2nO6qRIbBzGy+CHl9vXxDxCo+aS6mALDb7wg7HsKUfkUXbDECU0vk0vTgvAx2fDdzWuh+d
Xvx54dLIRTJ0SOIhC09ia/GVg5It4BS+m9z+qxyWJbEVbNKxMARM3cstJ4JkFe0fjp8XrWiMrEzz
veXk/7FTZv318p/++BrSHJEEDuTLmaEcTT3FVEqyFR7Iym7YpubF8sBLdPAcu7MvmSd1wBZPeFAH
IxhnA8l4Gc8RBAhTZkOcf/inZJMAQorYCjYun9cWBjD+LO4I0iawUrz9qytaQmTXAu1WzlOR2sKZ
AuMBvSnpUpabu6g4zGTq6PEGMnXuyzoHo/lMZTgpdLXTBFMCLJ8Zl0i1KUgNf1RunZMOtSOiJ2Iv
TNyZCX8m1JqfTLJGiR0okSd6US4ssWDjrPCECGGgOTLzQ6YrS+hRlZSnZFy6A4nLLDppptrE/HSt
iKz4wuUdEr5h/lxKypz7vLtrm2RQzuUWDJ0EYlR/okFqFUaaYUvPSVeBsmuNpsoePfPgIPTrOcvA
qbhMMGwYnlGofuEh1pBBACPkY1yL2+VE0/jvfKrh0QaScDSuThjeOy0g1oJPqplUhoDc4Lmz0C6/
2eMuE2i92dW+o8LVBC0s/lZtF0rZoscef8XLv6Fu+F9AMrI0YF4AlGfLiQKlZ6JsnpFTZoqLopsO
zIAWOl0awA3UQ/z7U1S4F9HhP6EPmFT0RNnw8SB8jJkbtZgm1SRMheZA008oFBv3uSIl7Yi1zi0o
VUyoesLR6djb5iZNWCW35BAELMBMWWmOAoIPQW+nNFhrn2MEn4XkbHnhKeqxp8TLmHDXsR3yokoa
qg4hmafSNGgJuH2bCjqhrZWYvMP1jJa4DrxZwCPJsTSqh/FM+h+uz7gjIrmYJV5qFT14JHciwc1t
Ii8/Ec7yFz2rk7Ct76Hl7veF7voicziEwlvh3yX+l17KprwNN1e0/pD1bggImF2n/fzyKmZXbnXH
BTpSS3uBlGoz3rpPAeKakdrN4GmgJGtLz4G7gftW4ddCBA2yfbwim/6CHhux9aoYGnj/vBglN+me
j8G18sbtsQniajY7B+ZOqyBQJ8zz/VC5cbOWIOt2N5vO1HssfIXULrcVqS02S/7ff8Kuc4n8NpRi
PVblxtrS23L6GKud8R/DqDd1sFPswRQu4Mgc39jAsFwytoyFpa/sFUGB1HNGixJdAmuTf+5YdM7L
lZ8jkGlcTTBOZ/hnKw1dedu+crU3XgepmTeVBKCOsnkY7t070ppAsjCCeSyXLTwBmuitWpuTy7pZ
O2yeHUYi5vzI1YUar40IuPrt0xY2GbhEV4lDUU+3Y75RSVI4PVBG6w8UbQzdI6j1vxJtmY968h4K
U0d26cZOGIwbcGtzawmF5HV92JP7l5jvYsgWwyAoVAVIii9ksrP4MdhJyU/r1B09FAC8N02lpUsm
vXT1dqsoErqPflG63lnRKQVVidhiSvTsRW2jW9mrUs5Ml7wW69nrQGYA9aOwdFG1dZcuLyHZ9iIm
OAJjxmziVLJ5pcPlFtXNxx4hTfkMf/e1RvVF15fqEtw0vxfHaWaoeIp09p9Q/tFgX2vthxxrusGO
3LxykLk131vhywLl9gQ5pW187eNjFMgVTudU0w7BUAGJwmf8x2+QkSlqiL1cuME1m4qZ5oxP5AWo
mcw1Q8KDWaUP6fJPlr6jzNeDqWx7FB8xfHCicsQYJ6mCJ6rOmhryj5mKbCZpjj4L4Yz55/hgKh6u
pKquqlB64f6Rb0ZRuyLJNOZS2XpPpEo1KI+iXnFra7SpOEV2uoPWRiJoxs45ajQG+TFq9aUdX/s0
P+6Fb26U49YUOXGbKOd0eQA5ZQFLEp9dESdDg8iZ9eK4OcKqKIOLvYLyzFvJxZBbFoE1nq+TZpgK
W3CHYwvuJDR4oD6bD17J/9K1JA6P5/pqGfMNatwM3Epks0Pz7XxSCYE4clLFbw5lCOzLYcTeNKdD
ocM5Ee2XDcblkjJGN25h/dQ3HiNdgelNVKMS/xiaKX3A5EY4xdlQ8S8Yz6SfVonKDJIVPvRyIyy9
GRNt8DSgkezVYDXDG13CIAVC/iWznLnLB6sVZqfdOLSEijbqlccDzjlsHA86rX9K+ICcp9mCUXps
u606bLGdjIH0aSQHbn/K2rm62WoTgGauMH5jOdRZuFAuQCJBz2EyUrEPUPbkF9ofgvghmXZSJ3s8
b6OpPRIvQ92A+ewQd0vDbrK4aiWjeMgVfv1WWsYCJg0YBmISyBsmi+wla6AX3vVLYN9D0z/XjSBs
kMiFNxe9D8eqp9IqMmL9xe2rR9Sc+BoJNb2xOFOHZYxswwBFt9/fIrmeL0JSpYdtuEoc604ZoFkc
CMxD88Sup2BsG+iZJIQBaeQLuTPuhSY40EzwnWPBnaKs4yF08r+TLAxqc4Rhqdz31CdjS/CcO86J
FdDs+P4pO8iTPAV/Qe+4ZE2dIGJR2LnfoOjyzOsmg5+xtoec5QHkCrCR69BRNx60vqVq+ZQaitvW
JRM9dyzdUcyUjBUt/gmj3gW172Bl0gUQVE1UhWUNG6b6DRmML9k3NbnfD+Xiacnvr78f6oZnTtc/
O89acHNGCQkvRNQw5zj3i+FuJm249deWcbhgekO7r1VYThI1DX/g9oKEFBFbTdW3niPZ3sq6fAPF
zQ7iU/TVB9RTdQseDvICASsADveYhbzWv6ZLS7He2rx32b2h9TOXNwE93kiGvzElcM9xm0vaM6Zy
1a2U4BiWOtSpOEnRx+F8/7TO50DkyKdwhetrN3nMN0HbhzpanUyH2vusJPY1EzzuNJNSWQ3bbzk5
o3AJgH4aXoMzpvwafdgnuORufTdUxK2Pr3e/UDZfl1+T0Mg5smUVkqpKZ7xlN88exP/SkDWQRdtA
8KKfSlkbWeekEJLZV2Je1rtTj0j9eD3A5XXeOtmVkfZIP2MrFT6smIYm2TiWiXllOKSVMuDOTnFC
VyDuYskanXUlpFo1dMSscOwT9wWO5e0Vj+rIibgpAByB5qXF6VaOMDYkI5U8J1M778fNYT/qfNA+
tGrNrbZ7xADcPgMuJZsW1AIpcYtgsy25DTeH+DL3jB+xhXKnA1snZqAkDpsba+AD8hOcTL1DOGdS
8Rb1Oh3ncXmY5rWRntVOk90vbnLW6w9mL0zDPaSv1KXwfB0TGa9PcieicVX6ONTr0Lr9VdaaAXGG
Mhy23PwcZYemWzeFog/dEL2DsJpx02M2kmXZsQfJ9iwhHcjvz9fPyF2vvIyt9vrfCSvGOPTZOaue
NkXcu0alrlhuoPS3BYsS1uFYiO5Ds5WsIzvwkTkO1XSRx/5PDqA2jnVfcI8AYdUktzH/GnWXLFCX
6ycpVFpnW2fsjJiWPjKomXDkVfbZlnnsK0ltgn7KiJCDYJomiaxNS3F7CHWdhbNp+09m6ZtVIxju
vFEqEVbcfwOus1VsDDrDx0z9zzEYAD4qJ9W/V/fh59J6v+aFt0/LWyGnjW8bUD5vLN8Eb6ll7Ih7
bPWyKnYRX3laHSzvJ3+nv3pQqcqGC+ICfGyzNMwQPhdQuqXQl9RebLI9UeKvioneCJMG0TicafCe
18f6xRk0O6QoLZsx6QLHGFo9KKzBzt5/P9Ptozu660qHBSz3695OTT/kbDaNnWObA/Y6yDzbKC6A
s2WR5let1fkR/A3ko++e/nO9NSptg4VGfr2kCsFCJ3rXjaKDaHm9VGeTAriHxRhSASrRTfCuJV/V
0nehvcEIDoPAioTrRDfEbsTDVRpiCF3GanQgI61qTCx38sIdjJkEPbCOtjilho80qwUVwrPPrLK9
M38MgHJm8oBJIQ4iJBhEsMDGpNPZYWpIGVQlUZNbpyTxH6EzmS1/mRkL9Ju5D6zwUkzlPPWcBNpu
EQCBMZPn7FtzQdhtZBHSwQ9lIeWb+iHYklx52RnprlotVgh0lMiZPmk1GnaobpS/93uWB0jiCPh4
RjUQ4Ne/tL9rSGH1bynh77ZamTyXJV1QSNu4rOneF7s3UY05q0mXXdaJNq42eWNn9s9cM7g9zWQ/
PAo4Z/sF4H+UxzWj6ltpxPcb2hwklPuuCA7f1nkyGM5gX6NA+vmk/NpeDd/cyCz4kDY=
`protect end_protected
