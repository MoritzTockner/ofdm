-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bkfBftMAUZbWkVlmMXxl9nCClR9LT2d/LjF5amz0mq1Usv4q8PHBJR6T1Up0LsRR+0Rs/wdRgWmf
q6Kd9eJPkrcHurG11Zwa0C8yzWV6YWaw4WlhVWEVeURYTS9hzzAIyJDIlXNdxFS1+TQRE8DkEK82
fZDhi0yJFoIUqFiyccEed3+1tk6WIFPm9tfumMJxJE9CZadmi/1k6YgPjMs5SGXOZjAS5uQ1HJvS
42nUEpzkP4fhWmf+Wfpg3Ipm77jlTqxSG2EhJ64ZbLAxDkLxCOHcude9WiG6OXpFrD9U/bQbM0pN
x2zCe7a5BmYmqkrkt5k4mvlTHclSZ985bbZBKg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
cJwgSR3xbF5Bd+2PTDMCOJxyZI1JBF1q7lS8vip59q71qb8UNjA5P0flZ7jkBZd48JdvdFmc/qok
NYjMricFm+MbhNqSO4qa9FP6zsCjqBj1rKW7Hqx0cEIVX1eujTiR7NX76qLZXVrN4BtiBfDYKylR
69j3Vhgd2JaRZF4JvUUyROXv5VrkrKIRw4VZN3ouqmcEQEiFXcomgnyEsJiAdoq3JqnSSVMEzkQe
omZBWF6QPhxHu8J99fqFjj1B3xakzQKz3VvqjYibfCh8+aq8M0R/dNBaBi4UaZtuXqYh0937W14Z
SI7zRYC5fCsGBCjt1ubh0DyGgdX6wYifne1OIO0BAfBtzzCL8wGCy//J0tHHn36vbwyBsgTuj8oU
NQYHaaWA950rD6yPckwqs2k5Mnao4hnEd+vYcmd+5fjVkg4BoGMJ002JloSBcYVCeeCCzXJ68IFK
EMB9UpDqbqNPvDgePDbETC6UawQnmf4BSYkVi+Fls3eL2Mv8V8L1f/Il9mVS5jVlq1O/hcPuDzcq
AVb4652h0TMAl16RIh86pVTrgCztPfFVpOAEvSvgjWgmrrcgQ/TI/XJTH0R0llFYk/U/ceh6suNH
86stVu6O/n87s4Qh5Bzi+RAIq1TEwsh+TZ/5PUtd9oLNhIJ4Lb2UXWJYgx3Tm2lB5cJ9YZxYHU9u
j/n9su5PgvDh7OWCoHzAgCJ4VFz6DFU5B4VQYRVHNjVPHIUAuAoC4gyUgCmCHqVU9CD1gK3sRx+o
s+fCO0tfx+/wTAjqOq5BBq5oaxa+C/JiVhcM/Mpk6Nlukb39+Fdk47jwIwq/4evNGX2xf1v880Qt
DcOSAn3TQ/zcSVcEV51firbCt5u8VwP7abln+mxwlJexVrq3vlkY5rp0qMVww8gyHfFNJ9l19kOP
L40fMwlAiCOuZZJ543122Z7oKpwoKFrYGUuqoCNJNtgoNNBt3ZuFdpv4SyVS7dAhONGcfvRQbiAv
LYrVDFEXKtHVKbkILm/b+p4zd6dzuk8rafEPHGOyLSMjYMaf0/r/ImAuV1xBk3DHOwVyRXiHlV4d
dD4nj8b2n3v9ZnafrqWVRstZRmJJ7yVFmyZlOriyiJ0qrBd9n83IwaBxTb1PvzyAB/wabHRbe9px
pdYiJwhr4XNo6URluxgrz+0o1IbZ3b9ATgQ4QFH0EK1GThYUE9I7FvpJDodI6yL5lNX8CqS/HEjq
CMObDkfSxY3EcZX4M21uyabuLa7HthE0V4wQaPOZTiwUCInNWdbDAClq3yIk9nE9kd0HnY3JKz/y
6mOrT+EkYZW4RDKU21zCNklihPhExgoNo3arFswm8OeigTkfeXS4SGTa8V8hByXDFIOhQnO+dFjf
b1zoMndFxexb7zS8SMiAudd3lSzJaTDVz8Q0Vqt5rDnrbHWlUvpnsqvYdgpIt5Cq/c88HMtXmmDH
ytfCTApgkfDvTr2GmwWWsnggjSxrVl27zUxPB7/+FJjJs7J0yhUJT1+8W2t1c9/zjfX7jd+ehWyI
wXx92m9I+V6uqp0N/5mAnSmLVYylok6cIcVulNDLnILanVKyQO/QK+6QVCKVeNBfNqedGcNIVwIV
bnf6Cef62zo0TfVoYJj/MZJ+g9Bw7KH3B1xyCpfv3NNbJipP0youXxEINr5F8+s3G/NMCwVO0toF
KnYTeCw+rdjT+ggJ2R8N1CHVoS9gqjBTAESCbC74S3FgXzMibYdfX23XvZakWvaF0OqvETYutJ1F
QtGrf+IFfgBzyvbUfMgqwgnkfRf6EJNH3CAsNCtvI6Gxr44pFO3SJm4xKhjfwgK9e9R8JUI9DrtG
hG7p6iED2GuhFWWZOEeWBVVTeAktFrLScRVdDU3afFzq9BEuYIwe4I8b/h6Wmc2WdeyC5ZbYoeY3
LLAqaPJCxDvlii1rwif6cpVUMHiao5pC3If1mGBR0PIcJMBa0rWt/dI8K+o8wTPaZhK2xe9M2P5l
Rp69wxtWDGD+vjIQULUIDK78VYePHqLAD5DPR7mQXYneP+2gnN0oClzRAppVQ9S9IomhfiXnHGVi
Wdd2i3vny7qBTxm6VnuCjMJ2DKrZLP7zSWvNbPovQu+spXoBC6OH95+/fYHUOFezYuSTeK45wIhn
Vdqw3WomfzCK2fGSdh/ldRjNQl2CiVQneTjInJGE+nJiLCEODQ/FG0s17FbhAgb4IsqwQ+zDODVU
Xk1pFjCJopCrVfamFtAAEXxYDr3/wPcPxH9joa0vkWckrIh8Mh9lfXkOR6Jrlk3jtFoNJcTvSlxd
u98l7WJRyTZzcigkoScgwwaGv+qiEea1HM3esWaTIjMjkc9lJQ6jlxx0Wds2HDfzq6NTZQvLe6Ad
pPVxMOGru143C3VemrU/OJ47TIBPIbbgopxM3Im1esEvLOPiHkcinBPActev5B3ldDglMkgoyTHR
kjCPPn1Caw+CRSAySZIgXxZzJ/oS43ZuXM1PiuGP52DZRxehdjan6Fz/HLFtj/KhMAvgZCv3QNkU
0JjgCOh43R665p9B5VvztXzIPn0JTh5rx4NoRe2oWDuFZz06wCIM99SEqtxhw1JwMjF+KV196Gtj
wxNTFBCeQ1BBC7M7sWdj9viQA+EnMzq6ELG9uGa3Ufe+qvjiEulZuqEBiknOWJ1DByX8c6TnwqV4
kbWobWyxUZItmLijSWpE3mEFiMWnWfF+MvgJ/RdpeG19OESnqa3iNcITPd3CzQxc1L+9+qNkPWHj
dAbS1KJxpnwSTGuANUlBMa3DW5TI2U4PHULAuaj1Qecm+zKlZN8kLZ81AmSL16nipstISxHD51fh
hi3AwPH71ZThZIMmXEbNaDqNc9hZ3bQpw1lb44VUpcC/prn46M1NjyzKLq1H649NdfxdszOPMzqY
GC3AIDTjkURTu4C69JvF9mtP/0FJkoc5An9mMplvuHaB+W3lkXaarHxAMe4mR5gxV5deh4A4348r
0vxB+nb4dQ2szeAMGT2+1i6EszTJdOnfkRp7vydTipuzTP1ZgDHdAVhBhNjb9YtDVFT6uxrnZ2Dk
WA4BGUbbK5ubAuwcGHvqUIN/U5PBJ2XPfR+MdNeA7buE8cSOmCvD+qGM7DmBJMEOjXUzvhEcQs38
k2hdWUSuFQkF84suWTWaCNaZKTVE0/hIboCOJzQGqd5b7JpZwfX3D4+4F7fpxlOlMMG4HQh8w/sc
G6suFWwivS1k1mUN/HHTYcWpztelQb2VzoveweLURz9+OKWMtgLsZ3xhDV+R6X2QKWEKXGQGStLC
ExRSlSwKS3gOQc9r706KS2NiCitqoi5InenUmDnsollR0uPm/h3khIOxzixpQeJSXjRXRmi9WZEo
ZSOuXn094kzhOcnilsN0cBsP7RmwJuWuhtuKElTNhLofYs8ASYM+98p2xM3iuiNmtT3UcCW5OMyY
4NJ4YyT7odXgrHNyQ1iR3Cw2Fw/C7t3PclGUQef4knhIJC9tpV3s8lcbKoSQ6861orqi+C+QHOvh
j/Z/sWwNVNHKT8nWgmyBxZG6/scK0CzXEz3C+R2eY/iO9DMCPMBkDR+0qjjUNeSdP/DuaY2avc61
kPPc3Lto38WdzHumQLCRDb0C8dIrrKFV5O1VRlHbgks0Bhi4Nq+3nQto2PwQr0YQzrOZEz8HkBEq
k6B1GSC1wDij2gM146XJND3GJjyKd1J/1FiXI//lvdM5TzLBclO74Z3mis8/rhTiAhc+y5yH1dkk
NUn7tRqPKQ+cdEZwoySdx/P+5f88SwZrzieXgP913GNpLZ2aL+aexgJD9FqX1G0Qk6FEmMagaE3q
AUMJqigCh9Il6+kpM/wLUYYe+fFkbdRZB1pHKpChQuTlgB6OF4627OIYkyiX3fgJsmIA+eC4G0fY
HxU+RKWbbwjPxtNm4EFVu1JY7holLf8LA4P+xQiCDJ8Y3mAoRsN6PjFut4Crt6giexW8cnBVVzAa
ASJwk3tMRNt+glhU779nRENmwraApKU6f6T+H/cMurgvMktcFKEfFThjXFrkXpP/TmHk7PCy+do3
09VJIQhvyNAwJblfRmIom4Pl4OqULnpLBNTeeddSI7VlCMg06KeTgmRxl6TmWFW8JRqxQgU7LLCU
UcktMlkCo1+iJCilciGp6ktZSbBBVArwL+mo98lVkSiPWqGqFfDfX6nWwmJXw9qsBQVWjFBAV+M1
GDuTRBRvdEzKsU4WWuC8L1PWAjaA52v5AQk20LDJPkJSBIo6yt9Bx/lS6X5HWYP77IVOG8nWATPx
+1tN3FbPbYlYIr31YccnlECmgCeOApaMCTgp/teiEjHpI2u7ohzuowHs6qLDWU7e4iikF0/fAOBV
jEG7UJ7eyUysJv04FmRO8sR20p0ZSoq46HgnNztwe+DsrzJ01+Y4L1MGJmxLW2gwIKyToBXi9hQN
1TKgWMgYgSmXkFQs3Mbj/+zGY11614khk1d89pPW2N0VULm4tippWqBDdPkr1N4x61Ecum3AP2eH
1LmXkXmzE9qIFEhNoey7piLEzuLRIZTP44a5bT28zJNGQhacqQ2+QYEUgIaHcuThiogHjngfN6lM
GgconSMjzGR3mWUafNaPsyYwD6eO34Q9d7fpLRVG8rkOiIZDUFmAhKfHLr4xq4waCxGGeiM7Ertu
J9ncUWkMw8NDI8bEUtNis4J3VRu6onVS4Gghs/hBKMGfPKMm8dvaehoehxKAjdqOFwbbFNLTiZx1
OAi+x96iq8ftlIFxTJeqhpFZ/BMkCs5zj9A+6WbRHezidWe1ZFKzROzGxlTVFkl2oHpQA+1foJTF
liIWtn20fr6jpMREZMf8XXC4NKGNezevB3aA7+72Ex4rD+vkVMUbKVgsvlD1LNrnYSOkr62sN6GC
1nI+vi+SNTcxhQxPYd8929lP2FXeBRvr6X5zWKNmsluNSDWvjnB5TsI9DtjJik81jjoVHEHcwqS+
4O0GtCM0NiLFy0vHKMO/tZ/v60lRUtAz8bE0V5PEbonv+LrTv8hHaMwAI/i5mkWYXKgkuj5JK3FT
Ln3oB9XFind8NjJadBzx8FikDGIFGgIC/S6rIg9l3xu7imdpoyH+h+C8+/3Pj9Daf7eJc7qA91d8
Sr7e9hZUbEhc403KP80p0078+UYQk6Z0ZPvz3NmHK6aDWZPw8CGjphUNzBBBxuNBtJoNZSO7Zapc
F9lRhlpSMn+d/1hNoKZCKlhAJMfQkkfWJVJlEMUdFBT9JHVfdkewAvgXZPTd8mw2rT9NZVwLbFnz
3NRS9SkH+/hU+xwtn6OlyTsETPf1skK841OXut+M7TtnR6pnxMFDSuyhpFXb4nYVRa5RG15Orxq4
hCXGX+h8EbfovVH536nteOmgI4uWvOcZnqqo82TzZnT0eSVKtnvb9S0LTJ06i01h0wx3zqmONQGU
0ryr5RC0qjHJEkJvTx+WKGlJ5GvtkTGKYtF8khEeatX4Ojr3LvVz2Q07LIQCL/DvCXAiAXVgihbe
uZpXeukYntL0PqMKixu7qFH1c1QjeCF+iKdL2naJFOgiP8UMGFQV16SQtVQpQP6UyZljKIl1RiVm
xZ77cJ09B5SEgRUbl11DFHUoGVrEDCGPP5xFn3Ltd8UGTuxh6GL4xS7/dAQAEbPEwanEw2Ovowpf
vNTmWOy5cXoWqW0IR3SeGLRCciEEq5Y6U1iJPErts4LjaYiJOnw+F9wr9X9y9Y6chZpi3dvs4i0V
AUZ0KOPjQKaMy8exQ1IpU7s+ueylI7VTLX+P1HD2B1GhFk0K3L911wc4wZ6qbdP0VJiq33wn/ILg
uTkunlbqE8me+5r/UtQ7kLUOl++X6QQgml82VbOuBv7X9HT1EmbARz1VC0KF/N5COUIY1vfzA+kE
+FXV499+oaf6pylXQ3Sr0CBRMJDyBSThEHu7IKtUXbLKH+Ei0TySeIaF+RqdK39XpsF4ynApNifC
p9cfNkt9QeAp8patlPkoEPS7IjhdA25ORo6yG5LAyLGB0bRWMLhwAV3QoY8p3c3RinzRSs2avlyI
quEf7fl/IVl65Oqit279aSnl9XaO0zTekZZl/b9lwiMaOWzJtYBQhKbWQhuwFSDYvSy7wBDeZIXc
Wqzhefg9JIY2l+34tcD4+gXN/vOStBZl5MEd60GQSD3BE4RAMFalMssxsUTCsZkmZiIk4QQk78O3
lxeiw/h68JaQkwiDGeSfH5l8gCT+aKlH58v/zjuX5Y7HzXPppXza6aQOm4ZUi7cNE1Y6IufBHt0n
NQ2gX2CyJQuWMlIOZ7XHfWVbLsW+ZwJyZDSqvAPkFRbv6E9CRX0zTwJDR13ZEjyiWKSaJUHvJ7Tj
kF12GisNT9how7YWd6EogUd8PLEclaCCCACVCnFOF5uNsp49oXH/eeyzGcvAUZ9GP+thmSA/PM96
0lG3xorQWrupRBPdPbXd8WMLuAqAYI3caGwSSqd6yaIEyG5Z+1ZGAWuv754aix7Kp7shJsNJHyrR
UEBug4yCK3rE2sx62YSAIJEMCW1P4Qn7n6aMdWAy6TRURqseplJ0hyWRgIuV3qvEeOZ1U0hLHPYd
MyVYMyuigVW4B6xvijxu7FPmdvVtTsuuPJM7RipVpht8ahuXJf0WIqUP05rBHhOfKHRKQm0zSDTj
UtvJ1cKdbBYkjtgZLd9VeGQLBj0faEP45JXa+Y8bM1u2XR44ONB6jDQHg7W1o31i+qS258VdzR9f
OToRKzI9NjrRD3NJ6kKrdvXDa8EEsQxy5PMuunBcbNRKsztMZWVSyQDBU4EOq5MLXkEGQW+QTv8A
RvoFHOfZ9jW6ShZqATpIh3qwLzq56D2Ao60kZXpWBTXJyC3NYmi4upK6E4PSDL4h63R51g5yegXo
C1WsA2DyLPi2PSVhkeFcgNZfzJaM6gZGOng5K4hbiKQ6GZ0Uy0dntmRJmmCJYx79qF5pL9ZiFkZh
3R+zAmqycj9h77PErZAio0bjzJf6nWWeV05q4X8oZDcGsVKhAs63oGrTny+Jx8K3oNIOYMGIrtaz
f0roXviPQRUZYoiyzhvWck5q8MbjhGX07qeLsfpKHCnVcscNG65lmuZKIa+zir/brFOW6UpyhCfr
RwBRaP8qAOoME2QalV23nkzxMaPfjHNyjFOZlRXWVli8FwcdEjP2Jdrxu0VUmwGnn0yAm64cp/6a
c7mnIASZSjKFfrQrNUeaBpTS4tSBbXXOZtNDdGfOiYD1zCkuZ+C9KRXnWaLx4cMpUMBcgDmMQijx
uWgwVYNA8f3yM0F96mroyiaEXIOTs1fL+lYYS1z9auCEzi1aJq1Ty5pVHwLq7RU3H6U9L77y0xAQ
wdusch7VjGlr0ohiSdvoQW1wYFlrW1c3s41Nb7kxvYvhW2/oBWmyXSE6ActHzYVKKTUGrUA5B+2I
VqdSPwGh+XV4RTx0UkcO3Uk7KAg8uvHo08+vsRYSRHAprCfIZi32YiX4YqSwUnI1YkZ3QRatgrmO
vOBQ/XxZNAlx9A+yaAJcpXPGGFM+tj8D+1HEvlAoZ5cs9IsLUQilLhnphVeIs8kWcJlIxicCIzgk
N3jKtklPBsdoYY3FXuLyqP6lsjBlabwxOy2eCIJT2ZJAN38fPx0MAa6OSF36/tMz0P9QehMQeV3w
QYHHvy4ia226XAZ2JWMQ/WALa/LEB4xnbmaJenRzjCFnQVeWkFtESfuLw3UmbVWcwQrXUMPXOC9f
2C5b5f/9rDUcMXcjuKyENEOdAwYTFvTBqHj5WMZzl0cAqkliddJbweBmDRlsXhX2UneqPJm0/r/Q
PIDNe6S7cDuq1YqNC2QnrDV9Twsl2q5T8gcyCyTJ5q6JBlM/u3UnjQZgABPB70qIM1AeZ17RAOo2
PGeihYUk0wSo0yGFN04LSrPYPPe4LtbNd5Ths+DS5J1HfSBAmkoU6zp0jexcjxfUf7qADqQ4c/r8
ZRrnGuTvMypcgv6b4YvtPXXTbfdrAv9HZxpGwf8A7Yy2kl+/xWO8903jR1RaG3YwxYQmIm43GElO
wKOvY/Mjn6e0BqACKsJmMcwQ37+DGfsSf+ZSgGZiFy6px8J7sF4bzi1j79Mg2bGJ/FfmV1ai5CPz
5ehYENLiewGkztKFl9mYPWwcIqMwJbUKgf5OVhPly3WCc/ZJCzrWEAVKPEAlxr/z+qnf97sIPil+
Cfg2XFT28BVnhSdq8EQFj/OcMv94OL+k6YeEJfxowYMqaE+uH6XNniXYVQhKJAizn5srU8VrL3yD
3zFWrWXpxyNSbuUdHEf5IN5UrmJsH1fIJc/SfANFitplWvi+6bUGgaOl3oYRkaSkrQPunlHG2AA8
duokbHhIVLdW/O3ynkbbT655MFccUgZSAJmEZwAghnFZieSuBn1j1zhvhQYhqxamY4ADSeuldKIa
8FMDb2VBG89b/oBYd/qknWrcxmUNroslYD34LsOP6sjuyu9+9ftmZL15MA3bElZzF54I1RYqKP8a
vMhw1m4VI9kjrqL3GJiw0jYri5sPAK5ZcXqYz7Fo4i4iqsVo0J96RNse5IyQfvxhxv7eBUaE768I
tDw+UGpWjPQT3JfziC2ZbBlFX6W5rVT/ms6s5WkVs4dIlU/bn2vtewK7Z3EOq2qcnsJ82MzRn2Q2
jJt1hg4ICkSlGSRlR0EHunYX5rT1DN/PDgxkMK3tWd3HRxApw27b+ip1AvbuRoQ8nw8Jw39MuP0S
eX03hoTIfzgLZXEaJYbOgjJ+kAgenzO90i4+roydiJQRXoe7wmJBmjXykH1LRb0c6AFCzKCFh02F
9r18FTFdMZcDfSt9aX7rxhoYyGzdkopF/vHZPe2pv6KR1JwL8UNAUHX9PnqHhfuz+kwIMLMIjrEl
E/+ClV/JoHSBwRT0TB/pnBukHCg+W7uHwb07dz/EsTAyniVDu/dvEYikdvqVZGG9Btn2hO/GEKjx
1w9Sy/WkcV3Fx6YdX0KUAhyMVbEpbzDBC12YHYNjXfNSpiIXPqoToh+5o4/N3eoRwyhp6SbzykpV
aGWgx7R5KVyi818rvJTftR6qXfjzk/DWDHRLhuBXQUp4m1F8meKI3kwIjhfywZo6wxsljULw+Z2a
QaMqo0Qd6i/oE1iQseGWMABZJUmyEIB5sHK12ArhjY/UwNRUAkVmsh3oGngjQJN7duwVumXlrm7T
w+b6WRgSCr996I6Xs7PJi+5YoLhzMvfFC/pRQ9/DFVHVEh+N7fVvktawbXbIcQghr5XtVnGjWuXj
1UcnSqINsTcXJ4KJIXoM6y/bREC+eUDPsorFanvywVkC3YCfZ9cfXfFS5ry4gyIcrgqYsB5EyV1e
vvhCw2A/vqeRq8SnPy7IaiQdwxCCuP3Lc80U0hxYxacUPWks9I+wF8HST+X4h8XcZ2peVDnH23in
YSX94WAnTZCdwjfsrY/DgP2XJK1DK6EshkEzAKkUPvMzt0WE9z6jtot1yTxuX3glqU44aVaWSRK8
Ih6iK0+wT6+TSIaEG7kAH9Q54etAnxj4z4WFEgoWxLdgfx77myE3HHamC9VN0Im1RGwl5WI6yLjk
PgtfFlfq9/Un2pAjxl8BEKq2wyIoSnbaZVruGRgrNoR5nW9JPCLwtw4wKkSKnWRooHt+jjX+Q0xm
Lfep06vCTbkWrOkzgG80tZe3LZU8bqDdmLnfe8ac5thinhqcG3UDAgdZF0zD9IWiDYebtrzrdMfE
QUh0DYTfpWn+9UexmwYah0+4cShC3Wdrx2jNOAZqVrbodxCnf19ObZTD8KjwI1WD46T0KJGUjjxC
JJfdut1TqHDZjXmsJCGeuA/oepSkG+kaEGI/4+qCCk3hBbPPM18VAV/5RZSHO9DeowS+iqDZ5c7g
TT2BLvkfm/Y1WaB0hoTAOc9VPwueJtf3mzj9v5M42VRGs4pVNditq0Faov9WAMb7OOxT3HElwhEU
I/Y13VfJU34Qb0Vir9/lLK3fmSRIBPLcgLd5VcRap0L/LvofZarGx6Dto7QRvZDsMwzeD1i4uFAs
hWVjjntT+2+YorjYDT+kpBewrOZMCl2TiLfVS+Y7yS/kg8vi1nEyNFwj2MWSj33WhSVrhH8orj4I
KadPNZtvcsu6xjBtT/qNTTpMUUk7VKMNQFEmEEk1ZemTxbkBUywemYR3FXcW+J5oUuZDCe5azlit
tMCkncAhOaDQvbygnapfL1DP9kICzLO5NkmLVOXpCrVsNJ0PjAy/2oMRefXLZX7Tm9kiwh373TxM
9GMWqYLSaEoRQSsRfVj8QJwxylS1eqXdO97Y7UgK2Ixmd7cWr5H2VZs2ALGz+90UD7tJWA47ba5r
r2yg1G4P8Re6YhNY7VO9e+I=
`protect end_protected
