-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i9GIV3inTLnNaiqkuoaynneGdGc8siD6iF+DufoblAWX/G0mu4nDQOka01pC//6SjGA9R7DONsBW
RyhwjJdUfJoUe4P0sd6IQrUP1ibnOje4qvd0C9KhTfs3+Q83fTGAsEtfLgLWx3PeTloi0lAdHz/J
HU4kxvr1QfiOgdHKsgf1F9jsqD3AE6qDgOlgfVEUad073Ujr1YYj5FOw525KN8999GVOeiLQXUJv
f3Zy0msmIDp/7M92iBKDjHdCCKvavDhdqnZpgbJ6brrRi7lNronBzYu/8MzUBwbreZ3zUxzg7aCg
nBsDiLVk25iDqRTybtKIMhjZEyUrXzrmPiK0cw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
au+xR1k12QJZnoUuAE55H1dgwtSp3grBjYay6u0pKFc2YbrdpYzOiNryDO2OwOT5ZAmxZ5jwyTdu
pExDhlnpHdA6HQVk5Mvf+YhXq5fZcGJ6Rve35bODc6HkDXsbcOAgeJr0uFOyRdFpIcFgEAmUO8Qy
N3CE4DsYCxUVOLbm35qyyZTKowg6vAr6tyvLMltu0shibHD3knAeOxm7uALh/xY8ccolTesO1NaJ
9DS8QtwEtOU/DCZarfJQzzahxjyGTGMxElS5P7fhJotT1GqB+eI0p6WBkt8n3OIwrljiJPgXN2S+
dJp+dDV3NHC8yy5re88pAgeSGEOXLx1R5SpZMsuf2m7++zlxpbtzqukMarZRQYZK7406qIm8BX8e
lwpCJjpphPLYNlinnVjvhXPSYer1K5dKlH0trJkrHGNupIPbFCgm5vS7XTxt9g5xAmIuyyzcTP9d
9mDnpQ64akamlSk4iGqkcX9h/CGr3mcwlxVnbCce6XPh3UmTYbKBkNbifY9Il7jEd2/iVE8/O6Mq
U/LiMoh+qPMsk1uf//qhGiEfhmKIuhXc+IW0Nj6WeEr0SLIqcG6EW/SCWyx5oBCunD39zR7Rqect
6yB6TiPjqO2AfA6FaqpeV8CHKhuSqFm7UvvtKHAJcmpsCGxh0cUyV+LNgCeeuJ1jAq3yDEZv4dTJ
Kc1JDm9VXC+EgpO0uaEzDPRwt3gMNwT7SDLuziQrWMOykJXX2BHHq2qaznrK+OLry1IY64zwwpbw
A1QoR3SvPUmlZrsIMM9FFFbVS6bgNmOSSvRm0XOg/qCTkn35w6g1sUVhhdbaAcGD2FtozL9PPSh/
03yoU3cs32K1rtGs2kKzDDnaufRBWnVBqZEU10A/HNvRPZFcMzTTaROeATTrVcQYocCSZmt44OKD
q/L+3HfjKm8M2pjLqLSpHqvEmHvxL7Yv/E6Ut5dLWbwehkm+8ecL7fWGUkqRUqdu5Vgo7jwlo7/C
GdpSRArg64Fxnxfqr/ZMzySNLsdHJ8O5FWMfH77IupuVKZ+4V0WKub2ibtYl3ypcJ+JAa4iYsD2m
WktbSEj1n/ptA3nL3hNFeknMifl9nM4ZIWBUVjHnYkSVSViz3KyCN58UQIYu1rL3yWUJbCjoRgGc
NwSyWq9CeeFmjXRQkR9gqkbON2x7hn0H8A0OuDoc0ycYuWlnGWJeRBqc36yH+BOToq3T6sBQ4w3O
SzCOo0/knwJDIC3+tUxAMooyBTdvQaRVVQFcDMV9GctgQR/8zKsqF+tugDO6eU+uJ3MjqS9yZ5z0
0F7xD+D154E/IcM3P5ZhZ9iT1v83WFpKaVVXM3YFGzBSCpN53GWxkRh8ePoqxLGs1T5HIoBvFfEB
AfKNXxPuxeklKdstpgq2B4QdP0TqeQGeys6I0UNFjJ1r2EQYF+gvqMt7XGCGGK8BOgt2Wr07Ux+C
91KHxlWWr/Nh6hmuqHvnNmo7V9kl5tR5Z8wqvOrzWNArBJYZsY8bNGUTbO49LcyGJ7s/RL7KzILB
VaV1wLSPxkr2dn3R6ZO3ZFezEuvM9X8YN1dzRgfJbsB/4AXozuYF/hD4dqLtPjsxn2Lo7D+LQX5W
UCgni+BOxFDojDQq2nY1uQKTM5x5ntTRt8804RaNA12jawzqzQjjUZkuXL0pnH6gtnoDVdlxNenP
D2oBB0EoPHShcuJMGPavXHTisAFMIdFWdMuOLYHQ5JcsQroB0nG020YzUfbPBACXxILfM3ATK+qp
VenTjJw5RyQARBxEs195S6WLFnIi3+gnHUfSGgp13avTHRt1f45Vqmart3zuZFRh4Q/Xg3kh7GZD
dfaI2kqtdFKo2fCHEaHYgrImtPMyS2WEcc1PcyGhxKjVhDrsylyM6UrmquXWig8ZpbHdJck5caPL
Km0J+fZxYn+1Sd9SezOkfd9ePI1Mb29meZsa3LLop0hTLCDxEas0sgzfIQfnDMjnfzgQVew4Bcg5
CLZAyAGmFUZpR2Sy9qlvOgFhy6+t148iPgXvh0l/JEHs/FOkgZCeuwm+COCi08fbiM/ASmS7tMHu
gX6kRo5h5sJkmlW5GJnYEVBkV/279NRNd36curDSTL/Fof0PILRm2xqs6D8a0sOhYiHCo2RWqk8t
AJ30dmTDYVB6+2+6f7c2FUOX/UcqE7bCJCErBR+4ucugnaS1SH+/6Ax8kW0NAjHfQQa72KYjhcna
ZxTw7SSI5V8TP6w/rKdIBKuwHUhQdF1qTGw9cM/nQV5kSiXQ6osmhwcF29e88bjGgaJf507rn49N
DT5/wml4DPf1tWoqYDWrTRDCU75DFzRxwoyAtOzHBznLJd2PoZaTpWH5AcjSEUGTPYrr/8jHjtQ4
0YTPhKR8xgOTC/UBPJpgo6rt6IWn3xfgD8ujikQ7ye4giuiZQ+IsrRTSuOoU+0EwhTKtmOCG2fL3
+YSoDkEcuD5t7wysSNH5RjM2zZMrsSnfXvaGPU3pAns9UQi7q8ceqoN4TNiGOcTfrVfyiF0jAnq6
eGnot8rseyLfxXUEMnlozmUZII9KK+KGw+SEKOAWv4CMFHfk8lHLGgTFAlm3ZtbGUsAQ7zJHgXsv
0T/L7wkygMpDBMI/Abm4MQ8ZyULg/+tkN+mpYEss/AG2hQS3IupWznt8J68LFYioFqOE0v9mgYFO
1LLNHHnf751uO/EmtjbZ8hVbGPoZ5K+5/pQOVQn2mCh2mMwueeoKbZGOE3FN/ra19UYM7J+j0SGw
IrO+vg0SNohcGU5R4+F1vj4Cxcvy0QtC3uwo2++Gbrmg7bX00CD8LQyrBA76gW5dHS7Q4UzuMe71
vWA8jsLCu6+Pvq0rl4stm/CxxCk6QnQwHBanHaloyxCNdchYMF3SFxvebFowzv60nauqZOU8vqRP
0Msatgcb6vXnNWr4BmQ2sYkClkjOOi6QSeVZiKBSr1WU7HCyCPbNJK990ig40fSYoVk3qpOdR+lt
Arqpwr/bZuvOYYtZN8Rur9pDZtvqKhk3ws+r7qwqaB0nPaH8+rKEpW9DAQBnirAAPUoFDYO/Ej/C
h0Xc4806MSeOTelreG5RaaAVvnurjj2eahLJnb2DudwhUj3fMC4+eM5lhb8fYIWkxMqYRhNe/aZi
siIc3WdcnADOYQcBcpbZes5p747ls2+OsPN52NmTZ6jfvzVxpfAFe2ZvMERu5dAd++A9pSpGZML2
dkzfC2rbg7FH0lLn7zsEhtuZh1aA7SwjSwKZ259nt1mkm71c3fF3eLAodfZ5MNLstp99GzA1nbBi
5xQgVvcbigvAbWMkchCsoFAyXFCbBVdMD056L1xCiorBNBC9rnc5WrUEffCVX2NGVGVXPZO/rzhp
mHcPbBxdd51Mter6YulLVYl0fwXwnYGGlWFHELcYoN1RvqTAeWw/+2+OPdSjgDxmi6Oe7celIJ0f
7dfdR2ihPRJZ0h/F9PWzNhzzmbTfDHQ4A8Wkj9r9JuAA7xwGuQdehq9jTKJwsWVjSDRNTFhzrlXl
eTArNK8doC2FXoZI/tWvEQiWezQmECcu+sUcBUsWzgRQ22T+lyjX7WoD6+wCkn8z0h2eRGkKez3N
4Ii12Im6AYfwkyla6IZ0PSAaGxnQ8bj/FE2Vqvd2E4ApV+0jc0PBt1alTemlf+xU+8xg4hY2ox8G
e+dMmZHcRNtmeg8vuurK1AkJFA3Ln3njmG66mIMcJO7+QmHR2SNoZpj4sZKIf0mWLP6ZclXhjiPk
XGsVY/BBhnYyslSzf22R1ng22RrPLV9IwYt7kEInH8jzMSj5xbHXWv73SUDLml/jbKqV0FCnLt3k
3F5VzQ/qRVDG/8vyspfTZLXB668K/l9bC4JF2bGv0anMyJO3g2kJpD1oac8UsB78aNt0xWctKVG6
BbzFQlvOQZ+NEXgoD2Yqi8BbthfLfFgoSzTNNDpehlMtajXXCdvRxf8Ov2pDKPkA1jf+jF0OyRRL
X2tMyu9Jnsh3O3fTNHSDI+zVckj1u5iBpvLJa8ZKHqFc39HLBvrGUoWGjizDYygm7hyTirbGUYS4
akmZ7SSFxSWKNtnbQmVAQYbZu2FcZQkkZU+r3GjsmcIu4RiJ4QNRPKn8wDgXXwNwYM2OheFg4pln
GGTjVngz4mQTUOkDcsvTG+ObBSqDZcLEOWxWlyJ23lH3+wV7FFWdiPdRHLnjJYqbCIVADFlSvaEN
KmyMLxmdScru7ujynFJ0GVIcj4HId4EPUfC1vVgdi8pYhP6MmaE5cKV4eTh/auswZHrh1tlIi8x2
GNzRyEmTyKmzLhGPyCFqCWg98I57jsjXkJq/o/7HzFuFW+gqA2i92u+i37ILE4KQejb9jzYVRUSL
WGjXvQsK23e503FfnlktnJVX5T88CG2+3qc2M0L3ntZtJiRhG9ThTFgRYx3BxFdgMeyb4D0EQx3u
VXxQz+49QYW8Azrr2Z5nYa3R7e74UKzHD+obxVGtFT610NSQ2kLpa0IdQAJp5aiq9MUDjdJuaM4g
HxDi+5UBp69tJZBvWabTwAAl8i5BYKvyv/Qcge4WrVgfN8YuxwVIFmG8+GJEDy2+1zW5dMbLORQA
O8d/+toPeQCwpGNJLR9EHITtDO5SXZzo/jM7TiIdnfWU6oDGpiKFpq2gwW+oHNw8lOPWaxHYqA9H
ctcIqsXbhl0QuSJAsnYdw5apznQ0IbUcr8cXz8XugaCMX5n+cxRQ4RO8vMD0/q54nEQH514KoVNr
7s3tsJ/rQPa7XPK8IhdM0m7pzNZh2Ln/2Ecwx44EJNO+GBlah2gPWCq96McjD1BAOk1d5lzGh+ra
s1J7omSiILnhcqCgs88F/JfiQ9MziJlRLLtaW/noeKOTYiUlHGilF2GY50vWG7wE11py9PbP9i6X
s569QeoNYphpMv75rypwwB+CeLXd2BgYxwZ6u0IrTuR2SWwViS3lS/bAHS+hxA32GBvQsApFaRuA
oDIbfEu3EBXtWwAOyHolLml+mgKz5ZHhyplbiNZmgZuII18EwBkUOhk/e5mO1tzpt2uZEZKWGjb1
pxCSIzkvQQ9d0+RdMnkV2OjxB7cWPsOxvP6AnOv+5kInywQivptOy1X488eCdt6bHdkStqpQ9H/0
k0fYDlvQf3/nlhg8zt1C99t+2O3c6TqiAg14zMSKcEASlewGUYwsFIYALUev72AdijFDv482fnfm
gMJhkZS7Z5o7im1O4bUapnWi3uvL8pC1GRLG6HZdvbxz7znlW++fawd3q5/hFaAu971GS0hz4VVL
iZvTZmVlrvzxinLrdL8vQ8CfuI/l6wh5qBbkr9q3UgHKSwS7+Lti68wGVHdrCRc8/edsraZ5INc0
2iNd8iEHBlvgkclo6jMx3XlLECU4xGYZWf0qT2pc4TrctLE4tgHk7yr7FFX8+hPnjDdqRKi8imGp
6Tec8fGaOH/BrFAlcq6XVr2/cMpuMc6RWIGs1OozwTORg5cQziH1neM6rOmGcEiyASI4cT1BU/hG
yN4ISOV7Csk9yQP8gVwEBaC1K/ayOyE26rsljCcJZk8E1frFYaL9DNd81KfsvknuWBSznG5UGxmg
7ew2mkqZae0HW1sqTStelOhYohl9lJYOzrJvIk+XA71j41XMuld6lp20+sIbbdgaZDucwKYzVSIE
3b3GgE4wp4ekg9/U6/k2MSUh6f67rwdXKYXc9P16SMMOkHfzsr99X2UeVCYh8H3okzRgijG2roXS
tjg3vp9wIRMpv06C/nsa6farT3WH3Gd6bHJwbCXWmxE/HhJq5B8/D6xNxts2Sv2dTGoA77sl0e/j
aqsveA3fPKnzU24PHP7FxUKC8s38cfZ6bYmQI+vtGlp6vgD/OKc8lYKxDhgZccZ+7WeBuilFu32N
m/lmFxzTrv51Q/uY/ZxccPF6U7DtCigE/Pj082qQJI3Dyem9syM6CiPwvCws3yg2j0Z9eFpZbYGj
kASEamZfr3eTqK9CQtz1FRZiCw3oBDS4KYBnZwMPn7QPY9N+yMqzI8pCn566B9Xr+qsNg9fA89sE
U9rx4K7wSuEAk2+aVy9iQI6oHAMn134VjmAos7Lmea95JQY8LkEHjPTrqHiz94HyC3fZi4PPDIMK
4gOKmRRXLFZ55ztEzUsEgtgDWBXUPaC6jwgNP3YQ3/ODvbum/H0n7dJ9cjP1I4kygbJownJmXQJZ
mGUyjh1SPpWfiC0XEOR+b3u3a3YVh6SaCHPb3vCc7gBNjyb3CpyWxrwJuto6U3w/lBmMXXAaW/Z0
lr7wZjU22suEvGhq+I7/38f/2j3w4oAxLYs9DVxj6sd5bxad//VD2NXPcd8zwhWY91uKryRmNFGe
i/4xKkV5YNtS5nIjJ9Ij5dvb/AjOXK/qU37TPadw26F/IYjRp/XPzoNAXyiObibw3ADuMbzZovjQ
j4RfiArSQGSb+dwxNpu3dUvMhPa5qk1PzHwHfehgmTrzSmhHU9NmehwiITcTdBc5AfjO1XEtQFyh
8ZDkzkOFCSvFeImsIA78LzifRZ2i0uAa9L2ztldpkMpPfx+/ASAPDMi432Wf8nFrdaxJN1iOckl3
oDpNwg+AO5P8BPNVk+1LSw+I4iKJ3oGLh+yxzFlCzoGrLwywle10sbGwZgCDP6X+qF06n/KPQ/np
aT1tAucCxgf50o0ombVd45+pfKejyxWr1R6FHcC2r4AsDnZjCalqYFAJBdBWwPmTKEekNQCvt8W9
wVE1/NaoedVwSLNLRAiqvY6vrlLZUDBLlwwc1UfiEA90+BpdAkHgOa+2JCLOGWrMmArN+q0aIPr8
VMc/G0CjP5AKOpq1MyUCcuY7qc894rSPzv08CHw6FD+4zXhjDHz4UUXVHi76SK9aeVGfgP5AclvD
ZTYQpChD8fKS5AfZj7rDSbK+L5W+J0bLDGqqevnzIqwSu64/ARsvbGPtTlqYXvtK5mcgP8FFj6vO
d38HX0oYCEUbOhKNsI3atSxrb/lNrYBLpfPkYqVAGIlr/ZvY9wfMWG678qQimS3oSApigb01udVT
gXPJydymLUq42KHzwAXBR6uT3LnvBWmCsrDQTD0yULW7rzUu+5ySS9lkupvH3be4IY8220hoTLYQ
7Fw5yvBClbsxjo0ObJqN4q80COL2fTKNmY6U3QzZ39TDxmtOV2sZ07pWj/vFmncaCA86KW0p30tx
D8+dAZzwKM4gd3u0GGiz+l/8zsKLNnNu+dHiBD4BYXLpFRrJzW3OS5aVyY+AP4ysPXcnciniHKwC
BqP/JDV8QeO0n0Cs1O2M+D9pNWxZtqARz53haVk9pScJgwcqbLJX6hRRxEY7I9PphLh/wXvgxROp
caKpjRlrXogsC0kZFpbVQulfB16J02D1m/m2jUwcEtkR8WlpiGEwV8PAFlJuvCjQ6cqFYtQS0bmC
yEFC0OgX7KqHueSp/NCjg92Z2WAXjUXGKjkRaOkmvRiVy/OirKL9z7St37wlbwU9W+ERBiu8lUIS
3FDU8iel+kuLpoC+nqT294VmKxmwoz0R2UuYUDOdsy9I00hqcs2zQvoHlG9c0k/iae64/4WSt6YH
KHBG5jMEQ17BlAVthi7xIS50Omf1ksMNFUg8bH18kFkIl/9KSiB7M6K3rjQhMPvfChvFhSF7Tk+z
UwoQX14GLBYGQTW5+ZSqk4YxlzuG2ub59K+w3P3PGyAHYEl9+yjhjEsSLXxiGcfsbJg+EwZYzKoh
NaWag0R3w2GNe8C89NuMfyOeAjYzlwDabZolVL3bAcNT82Mi9xVqCbrXuZDsZ6W0DNrSiCELKZrD
TKUZuK+LWtY7SMTGxhqjqD0GKNLyx954eCeEk+DbVvFabN1xrs3y+YLJbWuzkP503d4XMTVP+1aV
m1zq4uY6pIIBYVziQTBL0BESA/TuRhW6da0peWAGS2TSdPaLpBY8M/1WnENi80MoBGE7xZuXeFrW
OBxqp8B1Ud91p/Jmp2YF2QpafLCBHZE7aY/uURyQs/oTgoxjigInxtUy7SA0TnPZC2oz3Kx0IezF
1HG2G7l2ncj6CMHTNkSdmbFQmUtRkRFoZXzn0Ot1g9ROfkTBnC8Yo4RAvGUO64UPcFSSAO/TDgOS
DNoDLtJ7k+2QlYD+GnbAa7ao0vAbKNtUD3uyP30ph7JJnD3/93gxBXTNBi4sOjNAJtp/aICfhqJ6
pd0luz6H/cEQ/7lSWEpGPKN1aC98wgtaKOyhgv0xhNtvwDilceQ/ECN+Q9RcwXT4iXit1MmR5pVO
icgniFmXSka+WeyWsKSDahT7UCT2UM/GPfJFBqHxLambDDLljZ3IFxaOni9n9ZljTV3YkxtjxjOT
dZ9FkGDCkV2OomJHWwhcOXXE7WnjwgskyR6bb7xcOn6JzRx3EbMIgE5BSQ==
`protect end_protected
