-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LziaRPmF6guUyPVx6mzf2O3xKb40dmF5jSmdklrRGYUnWLc3X64d2jXyNNe4+VNxNUSAetWwoMIH
Yipkzoe0XUi1/v2TH+zdw7JVgz0ummq4LMYqyo/jkqD4D7nAHIoAhS1OByXUj8LNh0uynX931H3L
hF4Gnk/HOWKswErE7YQxlc/3nwmCQVmyDssKqcscjousqt/C9KVDzB/c5UEkefbBoNQBUx1KrRrj
duaLPkVcY9SLghhVpu2PqJSdzRUq6OdwI6dhflrUKLo77cMshGLWPePLrcN5N1kd294piN3kJ9Lj
5V6hR4ZP5621MXkS2jpy5kfwPW8Mu1PDBl9+sw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
u34C9gjiwfyIqO1J0MCFpHmLQc24LKzN55XzTj5iZfKI7WWlHu3w8sAn6Zn0fjotclZRPTWiynMK
gbUMyrE2FDuImEMyOxvs63mzUv1CuY6tb6GNYDiXYUXM06Tk9QKgrwWX4IR+oxgc0C6rPLUxYn4f
TdrzRNP8YYXWY3OJu1RTIccBkCFVLpADFE+19uXGghN/8UB9J/XfXjYNJIz5eR4d0KvadsV1zpmD
VtwsmtNxNZ+lVzd1UsuXDKszdG0J4nW0K/U7X1ffussGDAKjV4o2zCWxjAi4waHB5CE/kESyYUDa
l9y15LMYx3d1XQlCQ+zTAE3KWcs2S9gs3ugELoB4C4VvfHACxNUBSPBPOr/4UG/+k3JramnCiYBA
z07QTBlcVKsaFWIgh7rtGEU4Hc8iSmDUCDKcMqHiF+QtjUprx7aovBTRkFKsK8TR2PpNMrvxxZMf
AQHKCJVyYfVk9atZz13mZLgLaxkqVMTiygEwIXRLpIim++IHEQMZ1/13iEro7eGNNEpbbdFn3v1Y
+42VfHaFRRRes09zpMb+GJW18ZK+oQZRj2LyDLcsA+CoXtbkm9RinjJnkvPfxn4PD1SXSONjEkm8
dQEUxDo7lNba1Ohb/iBLLlf0gM5lD22bgCdfsf8L/ldJWLXqQi/G2Rl5FLC9qO9l2DnRvIHFRoHz
e6FeMFYG2PdWabYGpjbjVZm3husIFM9pF8c/P+J1PJ93G7UM4dHTbIbc+SChzLhiyGuUA7gNI46G
5nbh6bO3q8SjU3+I+nOAFTAzLzpijPgnNwHabflyk2+QAmQ6TpvO1TxGWSDRORET4WkdpFRAcNJS
J2Tu169m0fGHe2CK2P/oAcDwcsAXM06QBRte9lO8IJuRIU+yYOevMBYjM3LttixUXPEy4PeU+XRM
ly7GmN/qJcYMqXNqycQPO22DFqSoQX33BFiN0VDqSYTxpDYQcN6rwMkdiUFIgSamDJ9o67zxnArE
axmy5d3krLO6BO92S6B5GfN5bVa7Tt0MemW7krq+AFYGJMyt1iFmEd2b5pSpGFcSqlOMHM1shIEF
neqveBje+lMfVQmmJH+wV30wHuUp6I0kObVwCtPIX4AdD2gTvHVghBc90nZDbmApV0t5qrizdTRE
v9dOa34Vy/xbuLziZD1DFhGc3lOVDIf8piN0r2WuYh6Xd0lD2mIo8spbJ6Z77iffDN2o1F0jMODj
tIeWI5XdjTFTrMuARFPAfh/clCz/YZHyByi/l5a6Xi88rDtTjqJyX88wDRYQof8H+rEEnyloK8OV
iWaqFiQYkzxBFd1vcEZRp+tyasKygWeXgyFr1Hw/cxSfOOsquCaRG8a/FLwPpqY+O4KQinAgmaNj
0H76V9TFRegbmRwiFvHEKGi6wTPMlV+inhh+fmTfwKRTAlIF9QIrBOviuO/aIUqXgMeJzhMWykFZ
XUeAT+qSpI47nfrrecaPqvGgLuI6IIU2Q+UHQ7djGNGHuyHj100KOLlGA04bVz8ZKlRxMGh33AD2
1JcKsD+knxjUIWPLym38Se48sD6PS1rF8PMzcv8XuxWVnhu9x9C4s69fJ9J7gJdCQJjNGPt6rKOs
RpI6Mxpfthh/bkjErckSdqjq06upZ+QGQPt9ItBWHpXJqm8J5w4jNsZVQKlT96P3NIGTKKXZz/25
++OU5sSsqF6wBySAADVRiuwmyywd2NLoBlLa9vzab9U26uVxYUOeok7E27dAAFNQAhpmMu56Z5C7
eh2jtu5dK6iPNFZlx0MDh5/Ok6DHrdgUWyhWz6pRGw+ofdaQltPoBWCDWBzZenXPYyf12uhQ11is
FGTaKDO8dlecIyiuPPz3VCIMkyZIsJhUjzaxPIzU/QKBgbY5saflL8sfjx9Sbi4vnt0Zj5N9cpmT
9aKXNF5NnyBkDatue5c+6KwftExdTW+UWPbFETJNwqtfQmxqXd08UXSNpjPfqgvI+8ROr0GFH2fM
2s6cM4IZKnWVBexghX5o7pGGGRYMNt9NBmKvOBxkUlGAK0Z59I3GUte4wMsODlJG+fkkhsnaTmJb
Ct2TisvVZP9rSiMkXSVXhqQWtLAINuhMK2rIJToUd5VuPjB6v8t/ZqxU7RWA/79peydzz3EVpCEM
Gf5Ekk+uIWJUPdU/cD9Ycxy8UlKtn9PH7t8HDRtVl4I3Kcf/jl78x6n8sSRr6vuu1sEieFhK0FfX
vdycxHwTL0IKJou5mqExhag1PnTzHqXWpt0cetVQ34RCP57KjGASteL7RMbisQog3z79oeuIVSam
qEvS6kkKxeJyamIexG971xp6KWKaBpjGdqL2XZtMQKDr3ScZW44nyWWgQaVzmv6BsdVATI5sGwrU
9L+0hlkZJhqKE+3D5eAZsLNq/+bVszunu+hFJO6zO0kloK81C00vy+CY3C528vFql5u7HwgOI5dI
0gSbnI5wW31xkJhSohSbtCTO+/0TXWQTQcMUCM+kep0YEeJTqgHff7331rjPeiBaf1s5goG7RVbB
k26WvC6o+l6xbsWqXPX8zsKvN76FVuUNfGuOIG4Qyq7VLRMgv3eEwCcfEBI0qQF/wzBxdzj5zui8
l6zK5UmnA43B/i0S1L5AYemr9XGLkmwhbSBXC2eQQ4SeYlHW3a2znwjp+9D7/SVAc/BjiWrFmsrO
KO3nUPJj63fZgYoKKAty7kJev7PgOiS+/XDnWEOkTz62lyKXxXhroeBWElNLddgIcOhh/5Mp0I7X
cvnrV0jKNyJNfuD0HT83Au1IzCFV/4a28b5erTJ2VxUIT4KqwqcEcR+GnJaCs7v4J9kDSb9qsLMw
VQhYQzXKo8UrNsXSJqAeU5omKgEAOET3pRUwSnJsRTzDzGs2uhh+dADlhOgZNEkdEnJzGjeDTj1f
q8jQii/j5xE7ZgdCJuwpe4K4G76enrWcrEDg2Su2Y6Szmoa0arLKwmxLx6dSpnYkavFmf1/rL6I4
Tnvbxej1N+lgrkQTkffS81bcKs3xH3/1EJQyYLpZ1eW3hW9sOMnRoAlCwi7NdtRHkvFqGgzXI5eD
8PM8y91Bp2dvA8fB8WP1iPbTkBqYqFaPUvIeS8zEYvrZyzWfTlCPVc4N+DfoRMPPDSUXHjo14Rw4
IFR3ukboKgJLI4zz2WdmSqUO9u0Fjy4icqVhlLzQQ+562gfrJvuiS+r5/XBw8tLg84xd1yUfKPZ4
5i2bcxhb3COHlSl6KV8e7fLtNVKUkQ5jZfhZimkQ13lnS1h2Cnbvzy8954wndjK9t4erViO+nrH4
werjltI43J5/2flU2PsBebFpqErgQyZqL5qqCQ5tO0BghV+UWPrH9gHBmnq2vCrD0qvQ1qdyQLZV
WGgNdEex7JDLS62SrDMU5r9wGHW+ZsHm5t4+CIr4hi0xEYv+n3cADceUDwuQPichR2Kp/oJ0l+OG
FKFmkRAD6oYQ2mn81OWXx7E2rbyGDV6eYTjD5SbQAKwTwhjOjhhRJT/9N8JPn0XEepAeHh/qpShk
3X8E8ttSWxy0neKL1NA31FmNiRKzgHz/6ZkSUbE+kyS2shLceuO6Rxo9v+eUWzU6O/tMud1wYBWi
05R4nuInay+EQI9IC98pbqEiE6wcl7c+Rskq2Jjvw/ZhGAcyVK6Q+J4lXQfp4vC2QfdHJQNQ7QX2
+3CJBeD99ZcpSuWEYj9JTd73+4aMI8tzdfyeRtx4NXSjNIIEiihZ6aKuMpzIZr8ilma5QPyy5obC
sJweqkG6dzh/oWQ2IFRfq1ewNVMpCJlabgTc5itobaijRoAQZmm9gXkrZd4s+AcShH/grJwhdASe
8qJzjVe5Oouhk1Qo9gjUJ8i9EFll1zwKg/Z4ha9IBRY+MrafKrZweicNvpVQgFOes/2qE4pmOXqV
BJgkGZ/UAgW6Ka+EcQdl4LGMOID3769njQVeg9PJD0AgfTyESBxKSbFtD+jt8/CsoIoEwpzfV2tP
lkgzdOL0S4xPxrk2oBM2LpHHPRsjedfD/9Cc/vLPMo9RaD/o/OmPj1MxUQm89HjfXXmWQzV8+BtK
mH7IOMbNGFaHbzOond+iYEEP0tRjlMG6q7fHvqqZjAgWqbKo97RWvCbFnLxYTVgroagMIWzbe/4J
CdmVcnDrJZx84Hn4mRO7WP9npYH1X2G02ZeZvR7ns8pbrkaw0mjmFCP+l4Kxa4XBgXWiPqNx0Acz
wMUS8g7AU85UKbo2tSJXDnkWQvltFQ+NwMUq5A+ldcWAg+cqgGhrvBio67j3Gm1t2R2OhZFIFnSq
Dag1y1bofkLrmVz39KBuu4Qb8+hXKnae2jssx80P4o+na9PcfCC6H2je6X2HU+wMEYHRZCQze0Je
3bwOIJh5qa1K7W45iW+iUbe82WYh2WshDcO06ggCXgc6RyULwyuJ39jEqBB8ZfVokiGpaXNbQltE
qS4uQCd2mK90/3DsWyCia2uMFLe6z61+Uvincmysq5bSd1oeWKC0ntN1GA7E+fVScG5Ybtr+qyMi
ZttmFJrZYqlpZnvoLEv+TRw+uzZlhACK+2CjmxIP+WBGCW94jNYPkzSFP/g2D54iKmm5LGTKSmjP
D2NzCYPsjbuZSLGtdK7Z7gLWZsl9tLT+6AfNX+tFFn2S66OHOg0AhpY6bZQo7gcnBaIsInO3hLGW
cLyv33MnZmCHuAyz6daQ291uuYPsZ1i9Tnt+zgIrq7QJDyio0MnB6m3ipxRKiyQJOdejbj5mMbv8
EtXvkZSSH9wZ+DYXKyIZGrWTrEwJ1xFq7ejsffT6bfq8tpanojVkBVYhgPI+9yF4S8ZiL8Eap7zx
fcxJjbQYMcJCoSHwlJaZjv7FmylL/PE2jPXD6tXgnuWTxrw3DFCd091/7YeGdc9cr8iWGuP7xv2e
9Er1cPpnx8TfVjwZ8SsQ3cdY+a/Ec15c6N3AW66e761RK4wWF7qGdHsB1WIpCwpyORohQIbVir9q
3bVaLrowbZ/eWzHh5gHZMrbX+IuDXPgjoP+iFdFhsir470z4Y6AQFI2tQtvx6S7CqO1O+uRJxG8S
/snApiD6FLnl5w4exEcZndAa0St7oYdHQ8K+eGwTFPwKTyD7fOlCnJvEhzlr5bMe1W48xMoB7MPf
vateh1oxvYNQKHv1/fus3upHI9aZ3qGCl1bjG8KXOCqUS/vy8DIiHzXKKYXjrtBugDSQ8XkkxtOJ
s+YBC0Vxtg56IUiNONhBVwTzmJ7YlY3zVQMHmk1iVt7GZmAwuGnvS4Xif4WAiPUtjBJEToF5OYKP
kGdfo/qCNf48d0+SrvYvdKl6QnRIFeSpISQn0cQ2wwz84243Tmm83K54uS8qq1gluWf5OFuBRaXH
0+/E/cYyMgf5o8qjUllX6ZUpRqk/Y+XfDzzAmDzlbnTbW5YQ6DssDNazm84D4xAlrO0X76s8lcKx
4oCUEU4peI6d1N9jKF62Fh0sop6DipZM6mbPrqbqYFXcGCaK0g+TecAlw/+B1kiO4BaqywovdXPr
eNRfBcsKRx12V1V3eiIpS78eVdimg7nw3vkOEqFymes7L4Ua581XqcCL8hvWPbCOEyISdMwhFd03
tr2r/xFo+UpPIh7xX6Okn7n8CSJxVC4d/Qf8P+5e66l+w6c8YAF4PVno11uY69p+DGKWy5QTxrtI
R137ePYITSiO/D8VEdOxveL1f7QuBKRuRxfhEA5LxLNO1737v3MgyLlLY5KRuRu7oB/ukOkXCMlA
t4s7zLGG4mob1eFHc0eC1+x4tcFHzo+kCNJBo3pzrIdiJ/Dw5x7/ORxsddEI8Ys4NvnXeyMNRLEw
s06gzzKpPoanry8LyR24g/nkw8DFCNh4c65HUDH1SKvbCUZOwfTH2JziHmBfW8lKZtWKW4XH2vPl
7OuVgxDV2GKI4CsBHgW0FXtRepQ3x0/B6Igk+RXU2PKnhfz+9url/rjTo26L4wjtN5BNrsVKLMFI
7SWjZbkvZN9tTqrUDqqcayJAqq448AlcSPvZI7W4OuGsDOrdY1uWbfIN7YgGBHpS4Fd3oAGw1Egz
gMhALaf9IQrqnc4LD19zjuWtrX8h5dvdR99LJp7AhaJGdVaYfxdVxFWWjHaq5HxZhexqE5P36g94
o2cLDFMydP2Wc7fB9rctZwn+lVErE/EHuLxbtOoj5TZYQgl9ylrA90mLu4oc3N4ilVGpTiX8CKFH
0eJVbVWhVgzkFEgDbHE3OdXq+rHaB+m6pAWjy9ZTIB1haI3hu1VwGtdGBuiaKwOcc54SK+4X1sy7
2ycr9a9c7ZWvbwY6aBhYqF5altz/GAWsboj5PkrtZ1Rb1KGAwqxtK5L2B8AoaqPCAbJqhxSLvZ3M
1xznXvK65iEVl5KeUHgPl+0AQ7yuLvMTudzjmzI5HALTnEi36CvhOHItfMJ/I0wLxO8HtI4kg4mL
Jta8ekKfV/W0t2k6pvaMj1266gPUv3b2/SDA7DNXsy0Lq/6QYZ/W3tu7798X41deXiVIs8PXMNyu
asvY5i6TkKtfDp77VWtxPSQcnhpOCI/m8ImmsdGGoK4tW6YIrz5GQrSktCOevLj+VeDqJ9/mGm9k
UAPxzcklHA+kHjs2mp21NiUdzRfdalfLvK2WB+xl4aGJqEMewLZV3CKh4TSYa+y8DbzW6YRvNzds
bw8JWRiaGy3Dbjzy2XaI0EfFQCDbKNyLjZUWP33WrBKCP+vgLF83kQ9kh9JMbPg7SmxfFd/5rSAI
kB32RuFnVWgJYlLoY4RXXIa75XwztqXuAqrjMRUlC+ZboSlazyI/1WeX6ksYwGxosxB5BoSeTxjO
24yhjT6ZiwDNJ7/mWFtmnf/JuCSehSl0zzfkiW+yubEGJ/4y6QVUiyI1lKeVKbnwuqbO/Vitk98h
jJIBBovdTpgByrZBRncH95+86tChpLikoe5QOgHbqpryGrV74/LfZATmdDRrS0ruzHvSg/1Fh+QT
PniNZZfNSa4awkRvvBiJdIcqPux9nU+GWQFvjo2GGuJYRghlim4LMlkgsqOBL56puWKr9Qst6wkl
cInlLp8jg1iNOUGuP56xVlHowMGnjUgpUbuw7tf8hNYw3NcsBSvueK9OTDqHvthLn4szADPIH5/+
Hp0XEcCT2cOLEGfXwDR6UJvVuwnIepFCOocGnEDe7a2AIXxU/eynW+mMkNbG3l8AjPMbX435g09P
wKCkla5skMpa9S3XIb6vxVEh7nffxKjl0XjU4KvNsawYiVzMxaQZw1HiSDWhidvtZRaSEVGPwnCR
Z3tBTT1Qr25t5PtJuV+6dkM/3EHhAvOZGgebQARgZI/4v2l0XS5r+g9JzqwlKUEwVuSfNaiP7cPX
YbUI5/Jp5dI/1BraLgp65wr3UK5YFBknILDY/b774ysk6HwbxPILU33ti3HIsxTY76VHw6gNes+9
C8fOJfUbb03PSdmAR4U8vxHb5jKqFXugUwA2ORjpBrkITGz5DyO/1pWDjqwgCXxWATuTn5vqaury
OV3p2eoV4WHv8Tqz1t817uIC/14G0TBLOWkC8KMGkmE8IG/I4wN+rYozwsr1O7kh3eQFREOAMaf9
B5NuCrNuG1RF8p8+j1kixd3nlJmD3AmEXpO8djCuehhQvJ5AAb3KelWOGzL+3SeGn0+a2F0py3/q
ZPvSjVrR8bwB7VUDe7icHEpn09HvzIbjZU36HKCPAfQ3XCZzdES7i/Uql1tLQOQ0kqcGEygAM/t8
Oe35/2d9m4nJeU7ZxGgmDSLiplxuvI/ZcZiEoYzgfPRtOiGN1j4tqqXeJb/+E1j8FHCIHbLzL5l/
LDpnhBmNFmmA8s4YgFR53JDTJUknIAX03jSqxIyulZc5judoM3GJk/heYnGm8dI9Vfloy+kf+Xq5
9V/VlmGlpK9zi+jV23lfJckGzHjCaWlbV+nf/O0DkT6tn8J8p6J5lsJnZNgDzf7WuRgsCSzehL2Q
JMjwmQW7r6Vgvz0hXQn+JhtMUqGYATJ8/PxxMN3MFVOGYpeRw4S9wigwxGEGFNyT2ovyN2AWpCOQ
aOrkcAD68YWjGLRXwrdA1WbDPSae4HGkfDAk1Iljm2ucfL5cMRAgcQtWNr6qvR6X+wCJt76c4X6t
jW/9mNLIbL+mXqQ75fyfvx9XMD9WimXYlasxLT1LDWy6+F1184dH4BonRfYEVIqyUZkNbnJ1JxPT
Xl0uGxwIAry9J8X76W7TqHocbVf9Nhi5BSKbJsMs8cNHTFmoaxMUFy1YH828MyQhIE1eUYbCywCB
Y5pkiWTCA6OoP2cEbFnRawn6L/Ul1kPv0gSRdJXEMhLzOuDffNij7pmS2o3+XIQyBBaxpWhuHbiN
h7xhZGi05VjOLoZfsJeEVQ6qWK6zRr0uBhydqyJdtJlvqDumcOsqKoPmJXiSRQasix1LA35KQuza
/YSV38x7b/HfVQULw3oytBnXsaDTMaOGnbhfxwfVPaKX1DMEiebE9cpSOBC4v0MhTNIImHT9lpp7
6Sxz0HWpfT0GRNsl3tu+amM2W5thDozLhZ2WVrSrPoj7IH6FAmsb4LW4g+iOh0IG+GUjV5L/HBTp
6U1+bLUgZ+3yXBaMst8skCllk943bW9H2ho5ddPZWHaT52uZza4EtudWZzmBBzh10sSkg/SnuDr7
xeogw+4cHN3wCtzdTO2zb4fFg5ezuwvstaYforfZLYDuiSsXF6Blq7ssVRI4ii7KBddrbr6AUc7v
AoWuYAwPOQ1eeOWDNuqR7Ziph7ZQf99GuNVpBpRF1uz95czofVNSSQt57T7CSly7HKDd9ncb11Yr
Q+nx9rH0oakJcTiYnSAeSHDpN2to4z5uPXFkBBelqXWNoxvAVTDifrkRpJpyn6cly3f7byrsA2so
xFmg5rIh7v3JenaTxUTOJBoDGuxRr1WvJBPyZD1mIc0YawlFLb7Oq1qVZ87o7kPL8OKep2TDbiJF
GqXwIVEegSHkw5GAPZaIjP7X9j/ccYuSnPwNlMWhtD2QEI22LZCCRRb4zM89YvnL+JUZ6KMBFwrm
VUhreVB8TBNhZNEZtz5K7bSYqMZ+FqlUbjhx2+TPN1JohpcT6A8SBi5En3bkakIJRUXlPW8bCVxE
vql5PAzNcS7IqNHRgVJeaVOMaHuV/TCCLB1I8oKdWaYE3se5S7e9oO96g3L6JLByeIFiyHNvn95d
jwhBjMiCIkSIG9p9cXEamGxqyFkHm1ziamVIFnX/CFFdSqHwdZltJ2d56+gcXJyYwesYtYo1iWmv
cJP1YmuYCoJTA4V9Suy3LTeLP8tJOIHmQ8X41lI1W7OxqGZSTZY3MFmQ/0WSaigFS4QXMntOKQsm
D10/sj+7BfhU0ur+LhLsooFN3EWTDPcJdXcaq4OQ3BJQ1fvFt+BDPibptpWSGvMI8bjW7VF+e5dh
7sNbhzUmZxeSvCI9QEiVYO9PBRvSPfTISKkaAp96/sTO8txOk0DiRVxnudoZqdnJ6rB2BWi1WMHm
QQizkduEZ4bNY0zOjyqJTlRKoEldKQkdXD71I+BCYgGI3PUENo67Tss5Xb9ZkzJrC515K7zF3zlV
YUOSgCnCkIE+63YnWGhD1FNxUDw5gPE9YdMJZWaWUhH368rIXVoWj2r6WyAHWR5aH8Zh03HSe/Ns
jKBA0tBjiKvE7KvQ2G9e4gUQxKWj1PT821S+iaWyiYd5CTZg1a4epjAvqcT5wa1osvEyvI0n656l
F+lUdvWtUpRaneCcNmzPiFa3iRvO6sb8Pi/BY4HQGfxVgCaaVI/cvgFeOGCYkf24uGdT/qHqzw8o
3JwBgBEibewsXlD5bf2W0dxftvadE9yBE0E/vLF2/ik7P1LjOGyvKHjBHxXRxHQzcwP09cQDk7c+
9AS+d12RW7cB1q0P8xpIt8Yk0nY13G+k8WAQvjHReFl9pPUsNmSHEX6oFVXX6ylxpfUFMKovtp1P
oWTvvLjwlAHnQARBx7rdxRqFY0FHNEg3BvuUea9bgHg1oS09Rtj++HECV/vHJHCQo59YQSJJ4AWR
DJVHvpykESF29Q3WDI/Cmzj37O7lfuekznMV0e31ez1Iv7yfIZW2+ZPsDkYuefC+hQ2bpCWOhJBt
w5ShkU+hVC0GidmYe49CHn2uMmXtZqPsRqSO+QWoHEjb82fiOAvxXlyvaDcTiLg6LOB5A5LZQpoT
BJsBDBr+s52aS36dRRah3reJn1+cduAH5c+rcqFEW7E1RA4B659XbxaOLkFaWRZniTVusqaWXKCQ
pi6+5VESHShSHdYrsD1qkaFx8RbA2nPUTCLrHXGCMQJx0ylcNeKzQVHN8CSUhMeojlKaZj/+haz8
Eb1d+JQy7+tizmkMRjGwHWqUjf19DDpD4sIPVbhTkqnF8vri1Ru9fKSkBJHa2MkktGe1EHAoqkR0
uccCK/Gr5/5iK6mikHE5UT5fZdWtfXJ/m0gchcBw6Xbzyaz3fN5fMY7bL6BC7Ksz1DSE5F+RjDRO
7V4KMT+c09yJRLL7SivAbzUTuuDuNtwgO/gxVj7ayaJYXYdnsgs5kOB58HBy9+L47EUQ1OIh8EXf
K8jS3Ix8WGNocC4FgiruyzCjVdkTE0fVAhRnTxLlg7PQjUH4KZFKns+l5LopzwwT0Ddu44YGlY2u
b8nW1ZG2MS+nmY2LyJpa+WN/BWy4YTPwDCug6drGLXiU8bZqT0RQTbUbs9BGgu1XAqArz0ayWStj
wJKeyYbRWXfGV4jg1sKgOp2lbx9YnnNAAEw3mZV/jq8fEKoJNpI2rC3/3vH76Z5tMLWyqreN5XdU
qMjZm2MkEa6mxrAuSamnzuZrHNiQ6fzsE9jEFdcsm5NDTrodFKUShI48Ab106d66Gn4/b6Ussgwj
RlJX7I3DJcfcjKKK5N8+03etjP8nZBztd9eY50QZPZMatFyOtqjBMdZoRZtvaHxk0W7ML+NYHsib
MuyY2zztf5TkU7jVoxFNGt+AfDdUK2rX+oaiPIq9WDmcnqgxSSqY1SuGVKe+VKRTewKUUlZR2b9g
jVuvO0MrZASSb/s3DRD4wkwPVzSDENyuemfROvRpXX5bvaYhsRCX/umlj84HLq0ogAtEg5JDewDM
4DaWK2cRWkM4qmr/81/3TwovOC20ekv9ifyL6l8LKHR7h16dKRFA0WKiUos6WTtF6Bw9m+j8r7Ej
F6kBX48X+qEjDmtH3QZnGWYnUtmKuP/DzNE9/4jV34ufFQj4gJFlrDDcHzVWIU6WKZop027tiEHL
wm8W+s7Khde123pyaSzHM03RE69dSDmtz1hM5LtW+qbLj4Myy4lR5peZsnqLhD+acl2BAoBqia6p
RAIzmcwNaiGiTIfXJDFezCQk//aLA79/VO13Iea6pti44D23Dhq7Jxr86Tw6EXBCL+v1Z6DYjfj3
bqElD/tGb4HVy1XUwtg9FJ3O0cq+N9Bqt3bBbx0SJUryeGfkmoxY+dTtPE4+MTkiSN63ZBDtNtMH
YB6TSpHeb86RoPx/ayBQzIY+scG7qQE7Vw8V9Y4VtXUOr65imz1IFyrZ9pslo+y+rRSqxsJFwIVv
v/TSlY1GKE2s1EEsp0i59pfdp1iTljt3t5FqorrvGI6KFUtOY4pimf0mGvr/E6OxMeaxfl5o5juF
tdFO2io5/ro6ARSVMmTSjsYZPnDKwYuhRu+iblpZQEeDewvSW/ESy2DhphYtL9NesqrYnFk/IUUQ
DEueM4DrlyAxUxhRCwIiBjkD2vTxbbBkuGs2r/138cXvO9Q+xxk9ImzWyatFUqumeUnZQ3hpKXkB
qObXv3kHTCzK40zCPf558t5uQJn2rOnxxm6dzMhrilO/eG86gHALhQFghRok5NWEoULnU2Kohex6
f/BdSNOSG0x1mPdXajz0xGvR7kRx6I6F+4/ZhKmKeeBdJrKH8YW5Dp8rzW1+Jqz4Ghhs3uDsljPC
C56KcsGaXUEm66XZoS323UsSJ4vsb8ZcCR85t6c4p27N7lUPtGTZ/MZV4IaGMxf3gx/LqD9FfhtA
Xd2reM52fJ0jdQaZsRmmuImdiYa3V5W3v09ZHLZeIHqznt7YyZLYb6tTUeNAiVrJ/p+1lG5EEgI+
d04HpTbDWCgqfD129T3RInxor/S8/NvHmqI4l36AalgDy1qvyCYs5QFE6F+rlZf7/e179ZxAiPlo
ZmSAHhWn90/njGf/3rk23qm7Rqml5ooxucyPax+EQlnAdViUSsHTxe+ubQTq3vYDfySQToLPvK3q
NIbladBfLi4ywgN9PBfuheA8LKGop4QSNBKSBojuh2CypJ4DtEnod8M440Vz8Si2PZ3QyS/vqRyf
hRDhRIJ0yUGHZx4wRsenoV+ORteXM4E/dwcmaJSHuofoqcBEmuiYxu4B0w9ncfHbmwKgybptqxkB
EEWvwh7YH3GWE2DFxbdhz6VyLyFSyF4qzZC0GqLQo5Q58ER2QfKqq7KmtLOcMJyST6hS0icwFqwd
RN0gRs1Csn9sUo00J3bJdxC1zeeMMWCfFDUkexvRY9c/20yFMEdZ5FPNrJIsBAO9llisTkOUkNX0
V0bbndh9EHrjeuFsh0pC/qHQU8lNmC1eXbMRiCIryU9oNgA51I8mwWhnahmw2+Vuoj0wYZfMpOZn
xmE/F5e449QlV05c/KeWw5oOwAYBIRwlBlx5ir57gTdfYESgakl551KS9m7mn6iEGgFlCXIOFKgn
8XAYQh8WD4aHJW7ENDhACZKd6+THXe4fb/T46i6a+sV7f8yy7BIFERw/qv3pX3WdbwcmbqVmYGs9
o6CWlHoTOEvSbGK3dG6Leisjyp/IGXOzCvy8/TG6D0H0VlYcsD+Iy+14MhjsjOskJbYFDLr2tgMa
FaLu9e01Q/Qdf54457oI8GSsLwQJqSxezpwXt7BM8xTKRW88Bct1XutKGbiMrMADR42+Oyu8Ayp5
Lv/P8+1ccAskNnKga9EMmeUYXxCYqKjGLSuyWuhH0gM+BQPDaD5FhFcpfXhkHWw6cMm35VNvcCLi
GmKchX0I9pGlV5Ejp0dlUS62gfL6KveYtffXGUmppr6kM9zsrLVJMsBsQM36TSLZiJ8MZo7c8mLR
yLHdzSZzYB3JraZbSTG/y/ZpSHW1q5yvSjYlGGbO+CF7Y2Pla/2AX+YaMDL72nS8Dykenp8DLd+W
DuMFVs7XGqp4vgdEUxRGAPEwjuAlwjwQVwYtCkV8jpFzZx1zqD1Et0utSc2ej5w8psdqMxdoC2cF
z8Y2wsTP7DwnoiwGD0NbcC0HUiHiLOWP84NBWyb2Fao+9U0cBL+pmWomiDqjVUrdflutOoX5OJWq
SxQ7XXei6PpZVEMmd4Yn2CrQ5RqYAq7VSfsNmYV01xfiR4y97Gcy0ASK39Mp1zesnAAEi72A5TmL
z2r+7ttOfCPJlOiwJZQT0oYi+PnzwgWlC/WT8uDnkTp9klJxJNGwJyyeTkvLnw1lYkhjVhw1L4Ai
/TPXRXu5YBvH3hYlZrLjmylDnW/AJR4JbOWl534X+ndSg5yyU0+LkOl3krQ69jesDTMbi3ddjWI3
f/F2c9e38LwmEodHiPNSA4RTwxLlb0nY97klkuNHLUrAKisYKf/vx7U43CdfeG8laMyv1h+dCidC
kngCCF6ooUTxORlUd1JVOVx6Yr4itXQSAKZ2bo+JUoSaM8MEoQ/G0DSwKbuWRN6/LGaxX52Rowsz
GkAtOVXn5AlUQnW/9SI1wRt79LLFVuDitVmops9MWhkntYCljFum5h0dQaqtvMXnpUtZD8Tilm9l
mhj2BuqDrLwribZGFQsGeEC71mCMRLZERsejY7rQSjIjGoyc4e0sMjN9g1mZk6FXEAq85TnLf/xK
QJ0h/Z08Zy4tZnpEouE8LKDmgbC0P8rgLGKq6qZq+f/5FzFTrL6Zl8qRzusEAqE6fA7VFILKc8WE
0EYs5NrZPq+XUYUbkXFgdyAWRQzr2jhEMVUwEC2iChXzR8u99WaOCl6It1bbOc1UJK00uXIx+hFw
nJ9xbs8KJnYZIJN9hOCgaiW2cNFgvAxjVmy7GkVbsE4P4+yrs8Pa1ZzEdh66C576nJtaQd3A348o
KjqtI1uh6AFMp0ESs319CmgOuFhcfsj9kaLK7mybaXm7NhKsHW5fDtPTeNHMmfnGgfHx95gJgAz3
MsOir+B6Y/Un8K/+QZ4zNXgsvNm105gKSDe7uxH8ZRdG/UcVbXpbe/GmhBo0WMtmgeyaZZCg0oVN
IG9iGe+dNM9LF8/Dyb/jWqYgqO2yRuCH39vKUjtL+URg2NmW+23OfzQLEgb9z8qV9y0yH+/al10F
RxIAL3KDB5AeZOXbgyAoiaRYg9yJkUR1XDITLAB0UXoFzkld6Lg018XdbD7cNl3nvz/BM5saNZr7
3yO9oDYWMrXqEemnN7/mLOOtczQSDaVPdKGMRP/arGcuuj59njsH7zt5k6TdQRc46RHgTf+Mebdp
Cg8u5IKkfR0cnTeCalGPLyF8KJgEMHXT2G/F9q44y4rLVc61YRigQt9kWNgVrcmdrL3XCaqH3ozU
kImXnLAI7ZzsFaCH0uxnEvUTirlqnzrl/pcIiBte4YTz1EzQN0nhXERpJk0qGmY1dYMwy5gz1/Ks
EYg+4x596ebFpdgrTGrlSaMxMn3fLs7BUZRNspyVWSs1oDrY2oxFJYwjOe62RGJYqbVw1/2TSZ35
PEHcNPlfcOKWit6O4jyWAsTgrJZuEyS/3/IiecFDoL5b1N+oTdcBRYsqPtq65R/yX6VJ6xfm6fT6
iZ2zg2kvCPaildF5aQFs2A/5MgHGVsdX7UVO/Kf6gT9K7RcuRo+bqEHTL1jbofm9Z5k8BqVBPtDO
Gnps/svC4zSy+5oJCY7sMzPyWyY33U/wYhVsWAka9u6OodNTAoMy6/T7s/ly1cRF+0EbP5+Mavpv
r3Ea3IMMLbykhohaUEQoOp8OHm4Up2l7TmAG2ZsYvhNhlED3orZmiuROVUbGbsesXhP3id/N3vd7
dr92Y7UB/s+tqLJyhmsir2aKxOqrWMIqGYcivxDWESO5F2nEsUCnvWwsS0NvTOOE0PbgXWy7DXL/
vZRz/IAzuO++/0xpARXhisPxCGXmgQnmy9J6VrnkXu6nQKj6CxaUqCkjYAqf6hr02CCVHRNTlQeh
hx65I137VYVJ3ovqhPslH6yaRQEGRzjlj6sNA8KkL18dxhh9TioGd6hK/ErQSOqCtCMtAdHyYdhg
gHgTAB8DEKOtfvwA6Y91Q7gCfx9C1E+O0ndj3KXUvNenLBwiyQZVv/1apzjaheAzfNgou96GDzvJ
DE57O3wwdMPl8wzX/eJmBsP1Y7e8Q27MXBwnyvgDnbcCjLvEqnT1b4ssCJeUbEVb0HBa7X2eo/7J
S/Ax9QjQt3GjKL2p0LadFDt6tPlymVtKoyN0EMCpiNiL1vFSQuTnPsWwnRcP8EwWwcUPmMIRW42q
NHDH1/lxPNWhBEBUnUTb7Mu5iIeufv9B+KZzuldw7BcrNwiah0fsGOEjnoC8Kltb57GWiEjmfbp8
sLdZ5SS8e5ZLRqSfyF3d7j5AEmramKG68OV8gAEFIA2eUQ6MWqppdyjjLf0uOkKkQttw+udjdozp
IwwQGeIOphTkwpZ8mZHIh96uL74l0EP1UDZKEBPEPAbQLbGiioDrI015OtaFtaOptp6mz+XpmdlP
s+jV4WUy5uMZ0ymmTGk3EverCxqUH84BdjmzQvuYJ3tA+RPP5qRoPCUENuEHa/q6JccDAhPSq/07
MYcp6r/rPqVDAVxblwyw3EcncHb92uofs3DsvAuyppWJStv9Nvw7HsfF9zyuAFBa6WgIygxmUR+L
tJoTc5UvEltPI0h0UioRnhSJccr8aCwdxAyH422gG9/VlFT3sDH1I10aEzVmXC3wrcuHBffqk0RF
JST7ifZLtPOYq4V1XhU8b8PXG0/FS7rCJzRB8wPiuxoQirGvXITZanpDhmvayFGyB4TiLRKtkvRr
ATTUMw5yTq8UlUoPUP+y4uFAE9VDvTuvc18MMtZIiBN8YP3U7BFb11Al6QzJBaEB98mk9m+egUdj
hblmy2TeXam+Ul2v+l8IJ3WxmGUKviAO9wwL7H/7MNmnBkZRqYQ27b0w7cHUDabk/isFCvarG9gm
YE3BOdr49FhcW0B6RqKlgyupTDVDotcrONQEus+AY9ZmV+t2STqivhXCt+rAzuFEbRIViDgMcXF2
r4UueBqfkHqWAPi7ME1+GVAd95SRsIdbV8r5EGqDIJcp4lOgItcZgVUWTNpC/HaenwY2M0pI7RuV
vEh7p5zhEPm9gU5sf9/6h2GnzeF5zwvru6ayQmLAcKwHCtdoAfmsUBNOPxXlNpsr/vE7/kMaTQb9
drhsj7MeFpMXEWK6h6MPkymJd2DnJpej8rO150eqWVrKugY1TeBx97+akgOEBK2eeoJ4VxdeC2B1
D0ArmuMLrc3QwOdSY7QGts+/jIbynRiNm3fFy8u7CT6MROIP+TtNrRvg7tVMQGJFQ8CFNP5B/R19
QW0K5pn6rJa3O9Mp4ShyZuJ/S1ledz5AxLRSPZxE+jj3Rqp81Slguzl/h/aj9HhzPEiz+3CyP4yN
BBRNi2Is1YJu4ZO2obZi
`protect end_protected
