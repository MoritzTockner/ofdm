-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
byfO28+x2tLIOnAjdBbxfUUySU1oFv1rr4vSlCyuqCaizUtr2JMwqqVsAodZGTg7XvG45A9Qyn/x
/KxLnc/NdzBIBvalyzjgIL7iBLcHaAe7clJO8fI02kN9EOZt71JY4EHlS3ecMdEAUO0Q2QD/b34O
hh69+lST83KgOjape/pldVCA+yEGoIE6AO4d1enVXNHSBNrlqDSfIjiEx0b7El+PlZoUSrDBVCMo
2VcAO04BFiNjB/E0UpT/7QzgPfIAXp+eRcrD1Bnu+TBHPOytpiWwZMycFMZFvY/fmEwAxoGr9JJb
mdXacDlz7K1N31JK4cOQ0Fg36Tsx+ErWiYlDCg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
cn3pJetYrg4knrkHte848LORgUpJphOUQ9wrckYUm8BeRFMCERa3tqpRTIbNJAkzZT0AlfsgSFWE
iVu7XbXU0+EwODbgO4hvXqnKMD1PVFsF6YnY4LpV+g+OzA/5YcSqTLDAsBz+XYX9apD9deyphxCG
OWqc7/7nK98qQqFN6wwTEutESYf+z7XiJb6DESQoOrmA14VNK7P/6CLudHRx4N78Xmxzf1TP8bju
BLcM1ZSyvSvnraEI/hQwkpRGW9xynkPC03osf/H5oEknXjfbsNLcj2gfvP95RW3F8vjkVU3txAF0
cipWLNdEY2gCX9qhbccMXwEuTTuD6Et2lcadel9T3pB7AUQ4W3JLxhwyTW1kiBEklo0Lm3fNpHkj
gPKhYSqw8C1u4XhAx3MyFaQTnNccoBN+LLsSJPrC1vHUaul0SZcTtlPVbQd66KGzvPS3zlhk+Jza
P83mruN9ZNg2hDZTz/fsSpH3fpVop4GMelrnxhj6mZeFCz+JwUlUAFooT/1czFOyb747vu2OCr/2
ZQMtTn+NlmSWTs9EYyUlqsnJ0ReNWOad9z9e564kV57DcqZYYtsMLLusDqzHTvFi0cw4V6FyRLTq
ym+I0sbkKYVDatOyLVDFIphwst+W+bxnXihhNb9cSjASHL48mq4oCDxKXW+81nIiN1IA0qVPRcB7
A8L0WE8CkestolcnHvJzJJDJAMmLvb/ZysoUcJF5olNh62QdNrjrwkceERQXh4YLozERI99SCtuf
jZuVwEU2UeRZm2cMiW8uTms1R6PWiyjmiFvP2PNU10fm92oxrgREM7BsU99s3dQAzm8TrW29ezUp
pVCvb1YRudZ60PKRtJUnPgrhxVLvE749ljgkckvCt5vfDd758nycpvfv75wxwPbHXs5izh5n5iEJ
9HxYGcp234UWK4jqiOhROUw/odm2la209TFPj3UKB6WO2py8e63dPLMvcDx7ao8Nwg/PnPGm7hdn
lnoA9kYrkAzmN5SN4F51wE4f4tDpql+KyLCZ8wgP24qpdlSCWlhzeISvZPvXZJ7XhosAdoTDZ+QJ
exYnFF1jIC6XtMDiuuXrSJPeVy4R5pd6h++ivJXVwQyxz/TMVIjb+OUtzxybM2fFuuIPh4cVH6Ge
opX3XTNhUek2AhGgzCHmC7aVCO9Bpn87q83JM6FuIqCkDk/av37N9NE550bqQvF2Ded6+tb96bS0
9M8TwWrbUB6riHOUZbPcywNAoGVU7X1yuO1nSQHKUZB75aO0k9EdFVOL8iGgI0Eq59TiGFoJu/Ef
7lldK3jCjPG8HoYOQfAi+oJvVShOza7hz8taCyjiBYpqC7qduDKlXzNLVPggnOERPeazUGVAUkf6
x+vzqThkBiUut7YBcpI5yuJCsyzi88lyyZSrBQfL7AJ1w1kRu9nHYCBEwcpcPaMlbjf3A15gmATh
Ak7/SlmGkWgYmR4d1KhBx963OoEpaFV/rZjuv1+5j3JzHB+38+AFeRW4PcmCGl8DCUcCxedJXxhO
uL/wL5l2vW1F5a5jsk7PyZB/fCB9sbTVL5W9p2jBSNBpbwmUgyYU+XutYEKf3VLWingj7zO5zyjM
27N3zEMf4CtYdqCdUkp9B4eLwildyToZZ+vGqXWnvmJa7a4dh04uyHMsKJkZtgKMCliqVziQDFf4
smskFCCKDq6lcgfza1qDFvHp6HVUDZGdtavyAJDoqLnb2tE4Kht0W6ueIpeuYbp5ezDBQwYVJeSP
McRm4aifD2yBCEplimkj3rl+Gp8N278yCCrfJDsm2XzHB9vzpuT6DCqk7E+JiNfKM/ipfAbkbjUR
SEhOXRcgcP2rRmfsLKtLNkvway1pj4zVJD6RnA0fzeWdfqmMhQPpqO7gMpMvKAAiwIM7YZNS6lxU
qWUvB0iTuee1svfjfcpOt60smSzNXfjnEhCPsS1j5tcMz8oKHxbJ9D5zi3pE+pUB65fF7U5elC3W
Uma/nCQa8o+/7Ea1Lk3VKgKSk1cdnBY16L9SBzsRQFs/0nWY6qDQc+vcO2FloB2RrIlK0PfXXPgf
eW8wj+7gthNtNMrRIbVjdr4qoYNRXLaXF4/RzLm2JMjiQeTDwREokpoYdOgJhrht60fFU/N4v2/y
j8i+j4kLRULKOXOjZYwbitcIG/+lUBakZZQspA7nF13vIA6w8MZ3rf5VR3x4bYyZSYRUMPFQatFT
kKqykCiWiAkYGGJ9EARABlYzFX1oW79IO0jfGewvOc39yr3EOrJsk8Mex+HIAjuYytOsOtKVu8qF
cNzIFAFCznQqZMq/3euRgOmZvpX/lTckFFbhR7nCuDhtIAneOw6BHVsAhvlbTh4lFpyCJoBifvvf
c8qlQ67brO0Azjio692yGhNOUodObeq75uAYO9S71nCOH1gHlgrf6bXsDKMh4B/C06C2uMSOz7pE
M91C6GzDiWO1CJfifZMZBsY1WgiBUl6t8x1sCzMMlEInIkoZxpaibQwbqpHzq9gI+pkuixNgolKh
7swq2yUOyYEL0TEaOrQUfIkb80KEgFe4HybFcmkMFGucaOuxH0NNRuu2tJeTd/mnoeroxz+ayPke
5/lH30q0vxxSa2z8NxUPe9XtQEsYKkqvuXPZQt0CW+xxs0/EyecdQ1TcA1eG/K4vQTWh8KAaabTK
XdDyBDEq05YiAW/rrpi3aVSDmLZIl0JxIrOyVgXG8/ptdnjXjm4Dzy1Y24fmagL/vbaMwqtz5Nyp
xmqvsY+YkKbwqessGdQ5XOioFtnQc7QAAgAfqpRWhd+xu9XgpGfi4QsnW/9s0da4vbkNctYiXfUH
fA6G+XA0+IyOYZwqH0OgQsd3gKytZibM++aqLqytfNkMTZ4OUaQdfN0uquRrHbFtSbq2Llkt6vod
9hSM6pXw7QouaKhc10fQkRh22NZWlc3MzDbPxxObQZZxdagxksUbJeCyQD5JztMKnZQEBBeNphME
gDnWX7emukS6yKSbG2x3ogd55OkmZAR5ccGoTNC6lnhYTeW33/KbncJMmT8Xg5SsO05KJ4lGjxqb
SVo1ltkWRU7f95YXZzZYeb2yKbTN3sZeqNrgQmnhyJyKJYQwn7sA2at3aQIwaGezWQ2vjlNRU1Ti
t1s9+zJjbiLbjIHrvifdPufKNrRJKWtH5z0NvVMT1eo9JsZm8CtjAbVQ13q0mVANAfvndR//faIM
06UdpAU4T6bSFIdwdUppo+kiNGBG5MwU4hzv4Md1hInVZmShdqynOYRprGKx6nOtZtaKko8A3VSn
ner4mZja69i1CJj7G0RJqnmjzbx7cHLu2wRyV3cLur8MUcoSJmA6+H0xs1N1/G6hhIyR0NxnbCZA
3ews73UX+AZ2Yi/fUHqnBDLyTMDx21uU+7sfyZiFFdEfwxtQzcFPbCalV2BRlRtf4tGQrr75ItDH
jL5DJVxYTWr5Xtd0uWWZiNhjPcqcvkDEWIlAKES56LTL3HycYUycO+NiVg5RzUIHeyN9sn1kbzab
IPjPZ0kqwUy+euPalew9aiIz64AaqPBIhupX/HdFtbss2b9z6bwdQ3J1fqq5yovXNBFB/fqRtmF3
pVP/NygXirdAO/UAU+5WLCBaxbFx5ngMXZj2lOOXmR/18C73X06n6L/oC++4G0xTbt9Z0oaOtfOo
8iH+N5q72sIMQWzACChPdfSVvuaHdht/4jZxkYiGj+IyOZe6HTKTOQqE4IO192OkkIY4XfhxxPiI
48xu8Rh+c0ymQMwT7MR8+4/7pUZSaMYFXOlvjL0pjTLNmh4Xsm7lVw449RErwY3NGhMF4mfyAl48
+mZaey/8Ygh28IYIcqf6ia2wxGmNrPCZD8xzUAS/J9QOvpHFViUQ1GyVu2/PhM9WFb/eGH0fjaP7
lLPTSU1ejd0Bk9WowvF1W5YPOHI/87Q2wG9V4f4bBB6LXr41tpx/rA7TRbnMi8Vyn+JVrj0IDbst
oSJfoxcBvrrhzSWDcJSgTPdNBIP2KTQ8Xx9SMnchHPrGRM09c5GTBz7heGyqIw/7iOVzDGsuKtfZ
TSdsXWJe4MZdFK0KnmPk0xvIYZweUij6qLVXQx86GzUrqHDUfmEYKKCfyvmvCWWpAbl3LOGHKUV0
Ej3/eNxGf1ah18ZpVopcoK5zIlhVsS1awTqOv6o56putL7dk1Cri2zgB16BP8Ry74pxOnA3H2jGY
6FSHsnrcGEy7TAbRZ6tSaPTALVDWtY8TkyaUCwm+B+D3KzHDTcJ3E1xDqFsA5ojJVUKynzCDGkAM
45psS/SQI2sNGW6t/fSJPuhaTNl2x4tZVZSJeYLjgn9+0Y3DvOn94I5w6+92DTYeCmdbTcDeHFXM
jpwPzdpl8GxI4usv1qWK9CqBtb7VZFUmtcnNyi+3aMZhxiWYa6MheM7rDyHnDshbuUwPUwyuQGOv
z1ts6d9p+mXotsDvnjHe80xgaWqLLa2AcCeh0ft0glCcmnksi1yxjsdlmogzPJsgTFYEjELQzw0a
XiowNAa2VODJTzEYJep/XiE6V9Sc6yGVHfFxDoK9ZAGcjfQZvwXTukeUAHa51Xhb96oKJfS6VMBO
ju4BSoOq+zA7RZfvB0jAkSZfbUnKHo8d/8xzqwHsbUqlnjnWWlBzYId/vxqXkh3KEtlKXMjtRuTP
zdjsz0cJpnJkEXfkOyhW4mMH99+4Ipcn4/MVVDXhqedPdSDo5dKuBCR99PXBX3gmCSAHXwBQ925o
y1pPZW16Gq39X3YIMzCnHuj9AwP+jBqQgYYqsy21Cj4TcU8exlyNO4Cht5tsPYT2OJHPykn1lilk
9+NtReCiPWBgZIfqZgiCCeCEmhOa93ZIlVqRzZ9N51rYN0rOmIhdndTz37kUJPED+qlG2/uXzvy8
hBvFXywNIH3QDgXZBAlc9OPt52iUjP7+fSL9rRZqKu/OVnXs0DU8b/ZTjURLAa4tURHUvg59/wt1
awdzqRGihde/mCvrxKLbEZLw20XhxDK4QT/cv2q1nNBxIm47WwosclUh7RJudSssSBv2VvdqxwGI
7pBAJEoTc4il7cxR0nAChwQwNzyY0W0qlX51iqmMCnycUzoJIcwrWWygcYsizmZ9cF7Uo8SQFZk0
b5BWS0Z5gnVJF6mbvQvwUyVBU/gR8pfUtTzQP2uK9IAJ2GXCgVC3C8a2FeklKouZH5f9i5c/wsnb
SSOa4za1PZP9cn5pul6qOP2obQuZcphSFldWVJ7U+nK9X2Y5Qi5T1BRWjIdWsY4J3xoKmOjqYXl2
RgoctuOdsG2by7H+qQwre6sy9K00w3nniRnGNY8nceOa1cYc6tn1rSm3jEYbm2W8crG3RNlaezIr
TZ/fKTcLu+kGtGLfJBX9yPdDNSslsOnzmVkx0e2CphP/O/Ra+XB5lD61UAtekKTTFrcX1I9cuDp5
9MYl7NmVzK/s7MjebTBRUKWukXYIMcsIuCezULdEAYwBot7+cGJCR3JH3IYHefKQHXGcFmVskpDO
7yxjxrvRt44U0m9F4TO1Zx02T5FPiBV30UTjXvFvt2PpnuH3FD+JZIyGJONwTb4wKSz/YHNar7Ou
edeRNwNSNIRUCfDDgQ+vWTeHcHW3cRD+oVi+H8Jtf3fD3HigXEFFn4KGtwvOczvfzt6Tb6vcvzWN
ahPzl/rmuBiCj1fxEV6FPB80AF9I94GgbPIcSLZSnW328vqqRA04FU1zHwKWDhupsxuFLep2QTXh
yuaknmwgWztABZmoACZlO7xRG/bkjjfvxH22U6RmyllbYFDD32LZE9mY2JDFKyD+OFVWKxkVX8E4
cC+/cwVtOmnxmZfsR+rsJzYg3R/4ifMUuvvX/CS1MYxEnLCm5ZL0wbEYu6662f/pJXfD+pZDI10S
/6TbQWjmbXNme61lBgQ8bIi7BUk4KPzjxZqktFzQ5jhQhpOn7DaGx6QX9ueweRSqA/IIdOMgP4AR
J1Iaslq2pVi+SdlNSGd0oIs/tsljF7T8xa40uxED7vkj2K6p2MxF7m9IttNW/8lVhyFbAUKbkUjB
qwkPWMfqkptUfTEEMsPPAwFV9AAkc4qEoIc/Se06DalCdc3GTb97ihESskNpYAcFfFgbqagJ1yK/
mIkvhLw6UjbXjlUZLEkqeMyZ6aahYhf4CuE7tfsMLFwuR7iBwRnI0+HLMDTZR5C+jzfd50eks0cb
lEdJIaWK/H1LAb2FgAvrNmjkbi/0YZ/xMm260zc2eAPYpMeGI8g5hfVcn9VTWu1DhnpCtIGRT9fc
0NCbjjJz4VnX+ndc7uHcuGwgRUavLLJHC/1/QUBo/MwZcNEigMopK1hxHSTLkC7cfr/jEaxr7oIZ
q3ERyopTjiMFDKfGQNJ99shlX7zCbNylYnS+1ubItLl+pJT4xNVh7/lTYNhS58ydMnP3Zlp3RFWq
N4J1XsdgJcUlluZcf6LD3oQfKDxmNYGU81yrHuncbzSnVFbQEEJ45TF05/qxohWPQlHYiRHwz4eJ
XTVf9ORn1o8Ita0C1qR9zbeAKKSI+SXiUy1ZRTOHTdfyRywqGrTd8C1IqbkmMNYPMJliPLQ0z9i5
yjdSwNFKKJ0/InZ9nJb8Kms1NdfELtiH9cc7hX3h5MXcMplAaNGcX9QV27Jd05sfAleMxFctmQgu
nWF0bmVtSSdgeT2bS1sofK4eAPJTKX5WAcU9O3HjXOlrsS4+Dur8o2Y5dcKd60GA1dqUDSrRV1bw
BU0hRhQ3EaHZhjvM66cBYp7Cbs7XI9eGbTlHdgNH2/cJL7ysnFeWvaBbnuHaIJ0bxR46iMH0hPP/
1Ojk8XsmYXHkDHLBlt4f4vBPFiARASrW3D/z+LOax3ogx+Vbs+MBsxATaHGlkFkuyxFp2vo6fDqJ
KGfr8LNASjMV/1pCwuWAQFgVWJD6PPx3xkRegsP/JSzE5aDW/5HnNYi4q8zgPmsjeh/wztNox0kV
mKjnVfF+fhzawf7ww44+vNR0Q0cMUb6/guT6aeglyxmzuGMm7V5qcmPuwMOMPgA+hRR6ugZPieWn
6isvTtyQoXgCvV5Rq+gmnQPmEXv18vwb1sY8RyH8kj74Ey7QUs/dZdQL4XWtqjwfatelQtVgNgii
X3k2zUl5+XblFKnUVBrVIh9XUN73IZECZI4TBnEg7hkqGte1+PRxxTIoyXtaa2tn5jzh7+qkvW5X
y8FkFrD6YGa4wrmnjcz147Ax3+xHUI8yhchmzumaDnhj7fxR6UPAL/4ZJvrNMDAfpMvG0ob/ESP/
Tb4gas2jOcyKYOrs+TWOL93Glye30wPG9YJuYruu7dYMCQYGpHM7eizc+Q0O13Ce+QvUXU2bylrh
zf29TX0TJiwyq57FnjFyd9XzNlje8go+2IDKkjmbfB++oiG1LPhTPo9sGwwZrFjABDjtQMNksvet
YBSu2jmoawnmTUO3axEu9teERBy2XqlOo+BI7wOT3N060Ekevt0SyrutPdmwxEkvrcLVJnTS6vF4
CzaIoFpa4wfXoxks9KFkW7fh/3KSNNWzSS9RCnlbbPrNkjPAb6TlCmqMI52bCMJFVK2Key+J8RG7
f0e3mEPAx0SllNGmlwn9TuurzNG5ffzVZADKrIkPVais+WlXziqPL7fbAzsqe0FGFhAov7ckmcrM
tU/ozuE00WBtjpBeFqC//XqSxIm69aM9Bxmnj0aZI+hbep0+UGK2imzwEKmrLkW2Vww1YfMw5hFH
1Ri9L3zSp8b6vm2pUyjdhYuNwBuiwfTV11MM5on4lLqHCe8ubGKC31rFxG3EsMxjQg0qijYYCF8+
m+ZyyGMSpc311WI7MJEhI5gx7z06RX6BvtICtQuaAxoGIfOQfcxHPHmAMJFaY01bSmR9xRhJn1Ea
Ire9kWMA2B3SJbZoyoZTLA/arNl4V5N/Pc+4Wsh3sMNX/Y0zxruEEWixyxQHGi9t/2Ut56PpcZa5
KT1/QfyXv4E8erce2Q/iXaC8wY1vdQhU3kkivlw4zbPYHGGMjChJx2gt4/+KckPT8OkNyUg5rAJF
mlimBoIn/7i4vgki59b8ZcRv7g2bdTK6tsRMxEMEydJG9zTkzaWh8F15TfH3P22tnmNhAN1Fvv33
lT9ItZTrzye0s4V5PTbpjXBUXBMKen7hYLU06uJINPfz+NkLw4wdHEJzzr7ePDNIlfNupmNgfh3O
Dj+5Ff+JKfOLyEY+1FEU0N3Pdk4eCGuek85ijbO4fpU18K9wZsvkyBAieAJjORA3yhwYrEcq2zO/
+tGGlCX765ygWJDvHp9fGHU4ymDofqs8sG3f2jEtppUipjILZuv0JNUc5xm9+dpWcVwNMOlBhOOy
tJkTpuHN1SCUsHRwIXrd9b5lCSb7sHUDKQMHkvl52k2pf0s6pBgMs1A2tXBoDSO1+7N7C2syS3zz
aYrvEIvxjFJM7J3Crw5z0/Izn8EQf4Xeo34I+qEkarAL3GM3nUT2RbIquQXkyBC4C9WNPDiRiLdF
jKU6jxUa9QduDkMc0++Yy+UCwINsraFtZw15bfvnoLqvk5+Zhy8zXj+x3NJtd+HqUYwkog5e1cjz
Ot2tI/Gv6UJMlEw1auNFgzlW9vYpAI88DtPv5ueX9pRhwjyVlJyPmpN2Sh0q5mHE8awCIlJBQx1E
IMHUxCrbDKBIemjuYZShf7l6n7vC8W8Ys4cXrWRU5HfSAzUnRyO4TYDUAAsry5Jblm787IrJuHm7
R/BPWHs6gVFzaNcIpTBA+NHi96ZBvK48vdmgZsAW7xcDF1JoO6OwHl7Ea8Obpi3JKUnoimzpUDeq
YPS82dUNXuUej0XeUO01UG/3uW5iLAHxdYNQ3qPwSs27b8kw2e0S42Odm066RyOWTlw4M3YJkUg2
kZG6kYAU2Jx15/t+7jIh7TPjUxCkQTlzKTK/h/TBef83tcZ6IkBHjIMMxHFH3gPqUNq5Ls3fDI8m
qWvqakI2o8sVwhY+72LkmWbHWXjRQbkTAHmS6KwkaqGqMty46n39wyuA3EDwyNRoheGQWzB2Jtqf
wveGDfKi7dj/d/z6754d4bzQEz0VHIUhKj4vyEI/P53AM0bglWDYR/PxPagIVDADnyZdKc8vBC+I
VaQkLc5DYe+pifadDESB1QrRGtcZrQicjnOCagdTSOuYVB9KlAjWLPik2+7OAbH9qNZave+NH4T5
QOmqzpRzhPr3xrb4Vd+1QPnG8Cm9Wt/ElUfgJj5WwPdcXSkFF+TBkH7FwkvyZBALMxQX0EuQcONt
JaaTfrrLLEAAazHNCIBJne9n5heyESEXjWtcWYRvpYvzivQkpM+VHvZngYj2WqCPwHfUnYtXvHPu
dSNL7P0JZ98/qyxt32rljHMDwDX9CO3guR26vLAUBA7IJk8VXeXRPb2JRX45laZ1vj9i3DYSqo6J
yVpDFjt6Bs4eFCzVn5817h70b97PrF7HGSB5gyF6tDafVAxcO2UvmIr9AlRlKYYQrwXbGlmkK6Df
UpcJv/OJRaOvZ8xpAJVw2YpIOQQCqqpByVtLLXuUj7C0aLStdvq2uR3k0tCS9HXkJUc85b9CVi+t
i3mufvISZfWOECw8pBp5mDHsjV4exD3nQmNZwcWxA8P3s2U/HbR0Pe9f7Jlz7SwTuIuOUULZ7gt0
9CJAujIPTojJljlinmU2GdSoLKZxLGhzcFdE97xnSSR0WetXi72hvaNv7YGWQd7k6/cUgIAyovAI
+9R0JsMSwxcYtXy+tRGsgru0jegGAuz7/Qufr3YJMjA3t/uq2yyxm4/OwOFYePqzkUiIK0gjYc16
FrF8FxdkGb7tpglbcWOa16B5At9vk8Qmd/V/RoODj7VMrI+3EH8owMfwxYKoZcBRjrCLq6LJpfSw
fDUdY8aYDkilSBqhNTqtowLTWiMgfTvnTNwn3bChWhW7diDO7Gjl5qrkWXXX6CUiMTekTkas0aos
+EU3J2miCO4uAMa29FN0XWpViybAs/8rz0qVYe0YZxkulQq5tWQcoukkrEAcXYH8RitGlMrZWhul
upP2M6jufnW7kK5ZYkmnY6uLFIUPGFh1tQ+h9f6MuZ0Rwv5WCbbIe6WfcC4afMLtWjWC6dAySi+b
zxcsTA1YQJjnn/Smg7IOIoqk5QO40k+OTSyDFNysk3muNCL0q/dM55nKSmZpypj3iY3QvkzAipFP
swqaZWHPIGMfcbCdMNaASglsNFv8wAyy047v4RBPyL4GOaigIMbZoqE7EEtxuOnlH3vyA0u5MoOV
f19gCBGfWWe9Vb+qvc3ZnbXe0X2jgfEYDRXOqbfgeSD3lVid0efhul4tNj9wq5MTc/A0lK5ZHeRr
p1Bmf+SZe6+LFbAlXuzLsJ53aL4G6V0gtOv6hdzYFdXpRZBi8berIarVbxCEhyfehEOJJo78lQ/y
GoRt+lMKtFhwKB4/HKp+LAzMSQ3+W67J2z13tJ6WTMFNSSOyAnqdb933dqO1nMXRB/2nED2dRJfR
qfUBoL3PlpfvDzsUmTF/l3v5pls/GRBvtOoPI7/iSatIDIesbTD22vDj1aKUIDrnN6aNXRokWMQQ
BfI5fMsZfL5q+uLyyDsAkaceJelq7EqsInt+y0yDXuRvozroTpQ03epdfc0xUtCCi4j0s0rNkQpy
rt5LSUMzVhQUNMxIu/j6XSadUBNIDt2as8UWsSnPdjvx3z+pq4eVsKh0qTXPLsh7Iq6bKZZLtDVj
QSVZ8ew5p8yj86comuISLG5m7ETyOXNd1uyo/enKi8BGprY5cXu5CT06BPVUu7Cm9R+YXDn5qgl4
i1YuC4zthNu968GeXkFnBoNT4GvAvLsFLc1FEH3hsiwOtlwAArfrDzLerZualr0BUINkjNRJC3Qv
uFZ9GmmV04CSDWojtvXdxKQC9rJybRfNjizL+lQqSiaTZKOnJviGWrM5bvmIPU5W2gz7c/FSLFPM
5ORKLJdKM1OAXJ0dZEzj4Ce/tgATq9b5/uKw7/6GjKEgFDF5Ne2LObP5OvTw5si3QBeWn7nn0kZi
37mpIvUzefbhKRQA+eZ8imp/LQH+NajtmLE0qS93smtrriRKy+lVRahElq3oOZCnr8L50ebrcChY
se5De4FhHs6FO+bRD3PbYqzIySLx6RR7Ewl808qQGtv5A92Kg6kOvzLoTH6pxa3d227UBLymalOL
EOrHgzDol62xdE7PbTOW5HBa27qa9cAJ6sk4avd8S8VcytlcQ5wV5Uv1yUWdO2UYRi9tV4gOpmLe
xkMz36Ksfd/UecqWT7qHA2lhXtENZLknhA3vwYBqKuNY4O/IcrUR5xX/aDR1MIZeZPJi6hubnx2V
p8mDqRm61CisaSIdXdPyOLHNYoMnhB8kam+DyyJq6QsKGb+ORzmoiPkX8e/HxPrK6h7UNsPyniax
xTHgabRlnVT56Oqo6B3iEVcAqUs2yuDvA5GKjqQ6pMmzaRMv+LOXVSemylDg/fv1i91ORkN9LuQS
15lX/0MNs9oWHxO4mSxuztRbTp0iZpGVUuKQfUefY+N76sdVowhaqjGjvhnLE5PXJSKp62s9x+Oo
n5OZ9W+yzR1dpYLKDHPllv/kplVAJW12bgv17YmFIj1l09jYdQFjO1KD1bDhTq1CmqBOxB3oVysx
/mqkjkq/MoWEa4MPqQHhzbo69t2zVRdEDKLFMF/eVQ4H/YjvT0t5csPsQLWLBBfDjcvuf5EtZw+a
W0R2VURvwafNa9Bgix/gVeOL4z2GaP0spIZpBOp6lSW6sMRHvxhvTOTX9/CjsEl37/wq9XvfbNhp
A+rdxb93h5TdVIDFgyiGb4ttDvlbA6Ddg49BzBkIEtkg+NhpK7rna9RPUkg1PsicXl7j4yYux5By
B1fZYEANZNAySM9D0IpXjNm2k/EBmbpSo7hajVenXLCGO7cNLVY3PXnU9sLMuAnjl62dyw/NpwH1
iywBPNQP+qGuFZuptLEgfFX25XyHv4P5O/0cCnX8rLV0UHthF6MHzflCTYznBte+HCyT2ZNfNA19
wihThKE3UxeQLm0wHUy+6wZA7UzW5fcVixLWHR6t4gwHFj8qInFSSdJ0hSIKV4C7A9w09un9+ibs
mta56Qw2XriMZTemeA6c/t6VF3yBUov7Qtr5cVW6FxczE4SHM+GeBQkh4i+t/YrnfwO8KJ8T03lY
WvcDDR9+SOYib01Vgj1LNHjAxnqCb+p5PCFR/dXzpZX8TvrSQLJAcp8NhP0lybRsm2gA8y326508
NT2Av0Oq3D0V8uRhkelYTHBxK57emrYN810HrVwGInjEMILnzQ08hwp8F7BUg1DMUYMzn1C3wgGW
4a46qRIA4EsLwwoxc09/a4wjBshATIODMlurMu68dlkYpT7gMYH+CWXZuAwNlNVK3ebQnDPZW5gd
lh6CBuVnSImFH4R5ll9OEIybu0MkMiVBaLvDcB6U0xl8j0oPmF9gwLgpT6B5ujrsstQFE3l7+zhs
60nMROEurJyzdCFjo67rmR/RXOE1o00MBJB2vu4NYlpwjh5rwq+ho/uzatkPvlp3Y8s+qAIpHJLf
Tkeds3p55/Ib03fnUZpr8HOwUUFvXYu2MCnqoObYcAyS9AEQ3twR+amVuckBnfdo7pnu8VaFJlNM
bnQgaVUAe8LdR43Lbtijuo1NuGSpU+yiqoKNmnNVz9T8wmmdPfxtqM0ArUTtr/p8CXDutX9q3duz
082CcQKMoWZYEAoL0la14tUVbQE6nGf/61HcQNh3R4V+1Z5L03pmKm3P9uSfArOnLFNDri9a33WE
iNaNsm7TXXDDeXwZ8ZYjx57U8DOVRZe0gCl6pwjuv8lD6KRklHBKAl6J0nqYxkTRijfTYRgq2d61
XDyY7c0+qHmYIUIN0ZRJ9C81dU/m6KdwL5KtA9/GtNcoYf9F59njltPGpPoghLgsMUuKdOMjXUAJ
brY47pOozz7INfCJBsevRgoKKMfbZxbILUhOsSE2jvzF70CxF8PwjpSDI06DlVn0xVdNpdGkknsA
+RmjU5mo5EaIvMEQU9AQwKcC1aHRnEPmaMTxS62F0l8/kCKMZyq9Zv6XmjWua9vvKU3aprRMwZJo
GT76qJw8V9V8AfSM8Q7ZT705bUMBO4a0yJwIJCehgt3E45Ur6QRU12wRO89RyEpoEToiG9RfXS8d
7FuFAT6uKZsPPuCH8z2P0N2fv+Wuhb1Q71BP2W0WAgvJ1OLaUrCM2XAcKzDNjcz2et4nJaqRml1z
jtp8ZL6DV4ZYpNluic146g2Eu0QUARdidPRtbvR3ZwG7yF1qZoBOcOt+OL1P9qHrjisX+O4Dq1Wa
d7zNpX3bjuwLj1oULWFJ5TVPpJ6ZFapR5/vIEyvPx4OLmxUnTylWdBbAmn5XFbIf0Fvc5HJkRMFR
5joLB1RfM84oKy59ttgESrbml1CXcFivoR8SSQtOfvDGb5nNNlLCRPHm8lza2hpvPADTDKlnB+00
Tmfg86ylxEkBmUUTTJ1LzN8KpwVvUhyEGX9uYfoDAjGBAbFo05UxTUJ3pTjG/0rpMXnSKb43vVPQ
VZgI4F5OYZdPBgMIUSuommhYrstmdSyVrPw3g8x1ZfW2gkk9JdY24KMP9DwdkxarT+p6BMX/IXdi
eptGRLWcrjK7QnmmSkNhLZtPGteL+tG5gpCdMU7b+owOZ6jaAmJFT0bli+kVocS6EldIvjqNATJe
JAXVEU19epCqLkfwRjbDuEQLzhUBuHBrjg6ZvCFILFs79XsfgrglDaYIvurzSzDVrE5YodOAWRYJ
UXzDcFOy99IIf7ascypAsHc+NIYF2DahUrN3HHYd5dap0YWTK48sc9OoRUf0wyhhAwv+YmamP6Za
+z7x/PKVBb+lteIQUtNVBbcvB13AzKFGoeYgSSq2W5lq3PBmx4R5IRB2IdmkwOKvVU+u1o8yJDHa
8Eos1WsHVzKhEH3iWQaWzqHBrUBPz3NftyTxBerSTiEhUrOkENdUxHzh0jxrVQB3zhnoZG85a0g5
GSjS+hkGFqq+JcfyN1LwLwrXH8RAtq8dg+U9RXQB78lAWWaSgQcjDK+aieh2V+Ne46T1KXsf+2oL
/tKDUcaXjqk3gzbddgQhrms45Pazthuryh4ybDRklhPEyn+IT/4RNieBHxNxs89lLLqNgGgIU9vu
tiDKoMFDNieizCF8mwJerHZ4kXmbhqTXcqCdrgBoWmxhTpY4lKvSa0oZNM9t/u9HzNun1p/BtGVx
mxA0wJj8N63Crc/85mMa312hvvAzKBujMWjcOdI6ejyYDY5x26IZpK+tvEzS15CWY4gmF138UINh
9Q82erXhYT2dLHT/Cis+1xTDrkll5LuRfpizPVfhjuAUCWSWXETZ6843q23O12SEPKKPGx0VyFGY
7snRKRWEreqgEosLX+jA8MqJnELEVxBsBCv0FuiP5QoXKEGUCEKRdvCGR/z5vcM5ZhXvnegWakcY
NhfqLm5fDh1vBuOgzoyquKW8yLJV4NzW6r2Unk1uMhaiQ1/aW+84wZpeM+7Jyb5yOwis/elxQ2Y6
9YLBNJf/2686q8+XkaOJqb4MJ3qjVGa2qEcdud0MiwH3INBKHzyST/dMylWmeVpj+Zz/5uHGGwJ/
Y6cAg2Mh1KLnKu3vzXT2i1XvwPFuzERB052hkHaocOhQ01jS0xyIdGoyR4Z9R8ZBgGbPWvmvJXX4
ETC5AOWzsJg3Mkgh74vR75P/ZgRQER8YeDSpd3Li57MGI0JVkI8Vqk/1RSf4ePXeeSilpAuJUDl0
jXVxCdKmdpjU9A2bqz+kY4ENOOUQewlatU8DJomkT2Xose1gjkn18Gn3n27Po+lW0eUdxD0PwQq1
w8H53i3+LN4yjLSPbscW7lVNmpUMu4wSP7+5gNKi60Co2dpTxzlqzxfQ9BMc5ivwdt3+1l53q9pz
GjqECN4L1OMvII7aicZOKPfn4YypAslEu0DYOdzFbC+hTvYWfBldVlQPMHZHfeftHVTKiwMi+icR
F8Qmwpub80qM8t6dGzb0SBtA/OGubRU1GIh3cE3cweS3bQpNQ5mUoqgLWdeeO1i1mUrDUWwytrW/
PeBD/78TDK5RtfIwmhCTrQg3YrxfGy15qELWLXldv+2/wrSpFQafA8Q0Yd5s86uZmKxW1dOf89cu
pgSFNB67bFmuI6SFjYciRgo+OCEZeYfrfrSWWkbMY8m4gB8LPRmIW909WVkBlwfaYZJ5L7ZGDTdV
8KV1Cupq0o/vBIwlv5cmgA6/5hmVJVPpach4aSdl63iXm1BAkNs32z4ZYwwed5tgskpQ5eGmzGsh
60mnTeLKluiSX258j6iJmXu6Xktud/pdNUWoe6eLMuADJ+R3MM/pFgOUNCg86caBOlUiUXRq+0lZ
2BHha8HEa41RTecY5WosmQtBxsHYuEk4teorhJWZ9SO5VveEqbRiEZ7o7OetfoAJgBmjFmzDqtKS
zqDnBv5vXr5WT9CxrmKpJj47sR+B/gZddBLyFH6pqpVx2VKWY9JEMOmPHhIRF2fqqO2xOk98l/6q
Di+TTe9DqGW6w6o0AXRbsZtsAh0vAtoTj8yGDn4DUWU8f3LtyJzivG0HEBGC28+IEtdeHThRX35x
W6HE8RW87qzOrPTif0krXOSCVVhkt+ChOW1rMbdjFnsET+HJzA+gCY53GupPr1kqMw1/8g4ICp+p
Uc/vKVjiAxWeavl/di3Ed27zoisDybIa0yOoY13z331TJ6RwNCoCvZpLsmGEAbvhluk2Lkw3L/o5
o+qgHvZT8nR84lG5kg+YylqZfqHNoko+z478wK32PwfpsTIQWOb0U/NxbnBPCs3F5I4MueIxMDry
mswWbrUXswZZpT/d9ReyG6R+zMXva98rEWVwkhT0EHWAfTA3VM9SWDRQwZ/4ro7diGuaKg/YVjgg
H0cvdR1fW7h2vwe2VQW3ucnbTdbVfxc6f+7duZd1KsEWiHg84LdiJtiFvrAGiYuSxeRD7cgl5Xl/
iry6LP92L96RtiMF4be+wbNUMU+9N7ul4RQZM8hdDliR2gIuZkteZW5vYqNW2ZHZBpzJfjFZYcft
meUD1L+0cwlH27wrfbxt0La0MJ22+h1RINoOLZBkYB4agH3MpKg52IYd6pFUn4JxH6yIubiDhAnk
3LJhDIZMjGUdr3D1IUNyaXvXF/hSn+Nb/7WcxW5ugRCocH6WVvK4kv7uckGJQAz0unGgQgTfhBqN
URPeRJ+zWQZtUX3dfl5Rqoqe6+81wHzWUjCMvjDBoXSYh8p04MDJADGUHPQzH9jpi5T+XmCFFTXs
wcuvYEK/GujybM9VqV/Yu0yt0vDmZetU5iOWIZ3owmmubhwwDapsUJUCwjQHyNG395E5ohuQV2cY
Y8bHMmGTNhCmikgHyTE6ZxbOp9Z8hc0GCS+najcDP0U7fvoB+XIdKCBV1nIJqrM8jcs5cy+b3w+U
4vaOrpG5jVqIh+ToUulRqUzuLh9SWdZICWxOCxYe8tfSfJiwL9HBIPHxvAbnGlWcD6KhPjDW5uRM
nslwbGRQYfEpeV/oc+sl/EP7CvjEMcPmRY4KjZMFhUqE5YRopRKp3wIGA2EB34lJmfE/1He+Nrxg
fdSeT7dateZedEhpm7222I4Hmm+TmR3RgOVMbQ6kuFLohfTI9dyf65CZHgWXQe16ilV5Kw9Nvn5j
bkQ3G0Szb8PZ4C6Eo2mm9EmMXpJcKwrYQgPGsFBkuw/u2khU6hCDi1X9cHWoDAgfekXgUQPUYE+q
aL3OAhAYD7V1oUO87nbWabtLIzPLYWAdqVAuA6YKIvJDG2GHDjFaai0eyA9L1y1NM7o6iXmxUda3
44cQS9vD3PJkrTIN4mjhOloTWTMM+av5Chbjuqzbs1opMRQWWc7A0HXNRNPSpLTu/H9nC6No7yba
lIFhY3JqO1N9D3JPQJxy23vLN+U7yktmEQAHNu/hOj9tlj7Uf3jOoU24Iqfi368BSuKvNoG36FaE
/dV9OTwWvLf5CZ/fWhkF0X1JOEqH1+KNx+PNPtS658eGIGw1MOScuxckLWMQrENDIlpiBbSt68pw
GlCQ0J461scfETrn9l6YAeAKNurW7lJHori/HLpe9k9RIqMVS7LY//GqeiVeCwFnlh4h0zo19cBa
Q2XbDMv5/o3BX+B37F6Dksv7wJw2JO/duKlayTnsQ8iDL/FId4wboTod7HeNxpGTfCqrznftuSdf
Yu9rdOpVzFyI7VGQcqnvS+8VDE1UdDk0HJFh9HkXdf6y7PxqYvHd2TFWklPzTPLdOdlwrw+AsxxP
YGhy3gF2LLNuei0VENCFkAYk8jmJV/GAjFwovjEI1F+1+l2s9ChEKM10992Dq1N8YFtwTrEBNd43
XQ16VCTBcVtBWWUhst/wj0HHAky8oyjMSg2VSsK9eVtnBgaXDxeNJDvxuAfM/EXmKmR8qgrNmpdE
udaSCzqWwn5rFkEBbp7Jme0LJIFOCnYvghVq1NHFPrt/zHnfujE308YWtU6gsOgrL1m49zZ4cg4n
0fwXGtah3KvD424HuNhbBjGoZyI8LVVzn2pDqLC1Nw04elXK3CzXgwLnl3+p1wZYYxn4ZzG/kbMx
KTQSCNZWpeD+L9IVUSgYGxAqCWfniDMo3+2Yb16BO5kjhDZ6zaQMdsxj6lQ978a68X3MjZJmErLc
gHdvCuZy0NuKQiiFMU781hTrHYCN5GZ9qaDbRyvq3XO7AzBdyfEUxZ9+nxnmraFEAZGxcSnZ6ccC
opIXrHDjNpNi5oMxtdL238kupDzgDdwhfQu7kqK8ZeQxDvXm17AK24rb8jg9XES9a1ztOX7RqU6L
Ex3wh5a36Z6owjR3PT2cHD9Qo7J4mdUtwLozwR4VS+ZJ5NkOqXs6ipEejAgCPSS2JVEEsUPduWXF
5Hji2QhdgJncQkxb9J0i5R5DS9//ruJ9jTV6W99xB822ohhzabgUbjRpqJ1Sr8Q7FoUomW2CH7DX
H4/GT91qjDpiwIzD4DGqdfesigg5Lc9WOKCNOi9xibuNcamC4OqtgMQ6R9fWhVMojqq5vrF7KlDI
JTtf5PM+tenXGtpFm18zJXb6djYPApcweOBBCIRKJMcTER+M2jwePQMXA/2dxs/LyAJyKBe7btfn
1ILFSrYJQTRCUvbjECysXiiLfYmapPwRdZpU8ry9LDMtYXuiK2w6hy/OhLoV/E3SGGy/IJPpqd7L
MF9ECRfQNobhYG/q+d76IOgXGGnj7Rn/u4YiMl2nJtyZH+6CBAI+uCUrB0OGSoeu+tQswg64Z2Xw
VVnv3n2q+vf8LT/704fTE7BSzoFNpWiUIF/EFqhylwBqVMqzYDKhUN/jHtefl/L0bQMA5VyLJ/sd
W84CoN3P5hr3XGEkmwCOZXXyv0qrZkcWegA2ptio3x+Z40whnFI5kpuz3tER/4XPe8j03smcn/y1
wO6NT+N12M10JeoBcRepXWki2TFhVJxrld+H7XGD6tA41Z6A2LhAa2oOk8eZ9Nrf1Z8TW8ph4/B6
2H6cHeoC7o+1NNft7KolMa+r2cQhAlWi4giWSuVfbRNF2P2hhnNM4tGa/ZLaWPjLQMxnsPVypNb3
Sr9nlR4uk74txojTSZ3MuPqekXtUDWOftj1072hF0lrImp+cQrgO+bfGV4+SSQfcaG9V5w/uFQJD
eXfEEwWHIP332m4mHvNjj49YpfgFJm+m/jSK3ZWDCuIh8L3rMw4rgVaFMwPU3ttKieR8AcEIZbjD
oYZV1BZ6GxdN0AmTFkPqpkne+oNWTIwi3lJTM6WusZFl3uB8P/DGLQg/MpW7Iko/dZXRJ4/wVG5y
yTvu+zYcQitLKK3j9g2zn0sKErFEtZqIhrdHSn+yXSBXR3WkFWNRp+nilUO+NFwySJ2F9HrxP+Qq
vD3M5Hff/5YjGJQDpz8jKYldhObPhgGnB3YLitFC2CHP75JM4J98NkWCc096UpMKk6GntSxBVYfs
PWBEI2vBJDzVZ4ef6udPVgdTcb//cUjTJ+MbMsMz7JdYBfaneXVzilyqj2QBx0pTY1ADTxksLaLd
NQYA8EaJFImVhWWoMaXofzdE/qS+pp50n+gpfcz8Y+WqooU0YwUuMF81RjupXXEvQss7rhvT3sJG
frFYlzrMvkmUB+2jsdWgNvIpxp08vq8nbWxBOTZfdVtvwFKMdgyuIgbm0I5/d6s6IIJZAzzfvSlT
eBbg8HU7C/mTDjK+hf7Qul75nHt+cahcuUGiOiaMZpJNExmF9QpfBNZZGnEgyn2RFskebjqJPntq
qWK4r6xNRD1qJXmZEpL/EfRGRvEKmd20GkrQSHCOXQNsYIP7efCIGIS0OMhnAO/SplWOiN1PTvMl
3p/xZpiy+oM8FWkoZH15wYa8sN27BZP006Bw6n6+0EKiTdOxBJo0kWEKDbkEuyQnaevLpa/q0z5c
9U4spBHOr6xddoNjMQ9f2xYrhxLPpCuHbDWndZBaHCjUKGudFNzjvzvwh2H8kmKV4QIQN9FkSgz5
eGCLSF/4bmS+AsbyIlV/x47LIzb8CLi/JJNf1fQ54LlF49tUOPKE8Ydr/KDcAtuCgFDj3QaNarVB
pi7KM5/pMMTOG6TNeY5EcETkg8b7iNBKeXM+esD7fsGCUJFVc0qD5nE4fXWdsH/BrFk8/3yqRjiy
/Mrh6zVSO0W7zG0k/sbfROQUD8wVLArIjGWBM2jd1qg1IMn6AqgCfvXicQ2XMwHJQv4BKxQr5vIi
32diE8cQS7xNS9hGWinJPe9YVAFWZB2rWPbE5Rb3usO4+wuJJAjkpqqpR6IlkNuLPnuIzPasGCvV
BtQ3/6NncwUtUvMoYhe60hhYtQWVyEo5Zvkqi4OpDtSN96tp72mvg48KwH9ZcDqngwyRA0irZSwL
1BBXOe013U2tLjaXPDx4S2bYVSv22Zt5MnPtrCSybMWegbTlDm87dWADPs7SGtRP8IqswiQt2IZe
LJxqR29UIGfEGXNUgGKMABMs2kzbqwl+ErK9pjTzN9NdbXafT9UOX3iVG2cDaj+ij7qPBGKKcMNO
faSDYZgoFFf0q+6ujVzUP+7ee40lieAULPSCkDxntmo7fFYM3xnYgp87blQEdYFwlXsFVKr4Yvtf
HlwU+bTRpfcb/3e1C0mvNT9l0F0C5HUT+3gG+paAID3Lka7akWRULKxR9kc51XoKOJ9uQMfW5man
NLXeM8tvSWatezmbdrtfZmBxnN6UW06Blgt/Byq6ChPG2YIs5cgqPhn5q5DrTCa6MBBJIyou0pmM
DlXK+W122QNoO7Ly+0P0Bgjvyp02RIcSy/C3nh1CXUD5WvQxMwQeAVTfr9qSSYBLNZjjwO/uua8B
P4/5KaAOg/2+ABMxzGD/HAtx28FqiKx1yI8Qh+pVirfZz0Xq/purrJlznZ1YDLV4IrbJePXn/lpx
O1cSaWdkUA5StkbITdrYwl+97QoVMtmw2MB16V+iwPpfjp3ws1OcsgdcOgkj4zyLUyZ2IkP7+uCv
aqf99W9sHwiHKIvalH68i28dV8en9k58BsIC8VlXGEVTuXjPa60Gci1bFcm7mpP2J4dt1cxqwmGa
+NMxwbDcGbxCAN6ezXP6OAuDKEk9OP7nZrZVjPR8DRY2H2G5fqZxca4x6/TIe0tEMJFLMxv7RDse
JgtfofgumbrI/FWeROWxL2TiCSQloszTB1MAqY+QjEsq/ES4/CiYHj4nngPPjDly91DyKTcaz6+i
31asPHd9fa3aAnT5e6Zpu4mKpRfCupVzs6OaGYYFcBEr1rHVgRlAM0YbIoMLNh/91VEcpFgqVwD7
vQSfkrIwU68bMX/RewUKvq6JrekWyafxNUdO/TSOGLx3sGgVDOM3aWZTT8P4skeGxp17fzFpC078
lnn/U87k33R1kPynRofS+diYhhjUGB2iBcHCgMfdzOLEKDmWY/K963L5YIUMhloMG/oIbifGegKm
EXQ65Alz8Hckwy6NADk+XR1WHZEtshjqkKtzmiwC9gAXWS8cOvpGkI98Vwuk1fr12SiHVR4b10L/
VjE1eQqw3hl2JBoSXwk7fp6ZE2d23t7vrWjYAq+pDy9L3NRMRYWS2yTl7GwCB9/lgxHBgKmoI2iI
LofzsTXCl2aCcVywfo5QVxYOD92cj4C/zzEM31ABCXOjOBleu6pICE3I8KVvJkrWIeopAZG20ZdP
9C7HKZu6eipuf/nK+tiEhLugu6cmlBbfTJ3qeEiNHGw+EGdqPqcLhUe9zpZSY1SGnrQ3h3/hj5Nx
6VTTYFAdJXH734sqMyFQTx+/cVrylGrqtRJzeV5oi1noYAI1mwe8KEb9OKUXFb4y7wHqPfdC3GjD
+CC4BTJp4d8gC1HCh7wBv5YvuFO2EVzCJg7dzmBSEGjoJOuxTPN0ZIlcPSXdspLIiouWaWGyIp1m
2aQWvMawuevTBq+d1xeS7CwkKYqa5a8pwUwO3di0YJjHsODxRgQEh3qN3Zja3daZJ/aXQcHZOKB3
LlHs339uaLMFsBO3Lh9zFP82HgSuE3CSilF+KK3kXHv8lRPXS5BvNbaYA0opIDpbdJTFvOmzs+VX
VBiUMDNHiGJzpItPxwAA0WDKmoayapMKcL1o/E0rNmY2UrwMMjL8uhwL7/w6A3JMr3W19xgKd9pA
sEexQo/+BA2gcCpsTLRR+JY8SDGsTLj6GSfRJNmsfzl1xp2jyXD//X2qXWfkX1DqmIHih4ovwA6A
IPY1vCJz1e1adFxia6gS5zrKSBHb4AAvlH9CYSyJAsJit76+5ZPvQa+/tnqrQORoByS5Va0ifIlu
0AAP8PCfgfMClKJ4JgD50NM9RZsCQ478zfyS+PClFaYE1SQ57/YKtXHtSuzMjw+52zBHtMk5verN
7NvOq4vBu/jJbIWytHon77oQPX6IIru3JyCxQVBTBuhZaw4aNPoV/wHSuqpzfFmW6Hu0PPP9JVP5
+wlxhVzVqavk1Vl9O+E2snjW2WfCLO60ImGQoVGIQroYeIeCA5n0tA7+XZyEABwikRX5MC/17/vy
LOWcVr9WVNfqVhCfhBwBUIhOX7feMKfldwrgDG9RgDkN78C4DzIWCwmwCFQXSDwqpNpuzKouXS/m
35TK71kAoKlTmrxw4q1OwbpZ5WKzJe/B2OdAO30h8DgTXZfwaCV374xEL3gVh8NF3a2nMwTs+UI4
cyLKi6pzUsvvoKyeb9Z/GqiSegE90GoTWH5m+VukgnUstq20+HVMHV2lMlxlAdxwQ1Od5P+2yQp3
RL5Jxeq3S6avs0KzGpRwzSsE00oGM2Flc5n3uYEqbINmW+YcjY1Rtfjl5YjQMWfSgtD9OesF6/eG
bXDoElrjaFVBuapbaNfGj9wzBYDqRLZ++qwh5x9CqOrJSh9wVs4XGqqdqme6/f7BSaO2JssLEnbJ
OtBrtJ21K8xvDdC4J+EKRHdYEiHQd/aIjlf8aMec0Pwx5l0mGZ3hWJWS573E1TGtpU92EVXqRYV5
+uJMBwrrMBxnBH3dMvAlHAzRTuG5FSE35vyq+fI1aMFehj11C6AdwprXmBS9FIjF0E4lCuPxXTT5
yErdGT8HEBrU4CQexYUZsmu5vb7PDYtkTk7ukYT/qem7Z3isYT4aFfYIBeOAFi75hs2wyjU1RnVm
a1pQvJGGkEGq6m7tT0tCj5j8JjZQxRce28GLVbVD3pJPBSI3sPSvjXx8Cv5bRgoGSHmGQPI/49Jy
gL1br67+wPKvezWMAnmhuMpqEpCXMqChXBt1BEoil2uCrn8YDDm8J7KWr+5+bM8M/OoLEo1GLHJy
u+nIup+Xi8z0aloeSqVAP++xVb9PJfFJzHDOJhryJ+4v6z5AjDFEdg+bAjfrZWUEGtYp6XmW9jyH
oqRdpqyI1cBzUkwXaKiekqkPMJljPy0HZb3DWsAgYuLC6gKOMY46fDdODhcBlnscWri171hf2VO5
4kc78HRlzjc9PQwABL+YYhTIRz8IfOc4VP0NUI4tE94BfTMIOw7R4esk86UjEo+KfekbgTKtzcX6
Ysp7CGaAERNXzEdSESg2A8C62JujgaGgYFI03TkhfKYFrkwlZSoEHHCjmr2IVt8mjsGYQ1rmSnZY
OxzZNd9yC2afVVrLhDNer9QoIbLwpUHqvmjCQHEPqn4ylq95/Xw98hCSNzsAjDUcesp7FrOx2Vy5
3nasyExISjipwtazrrzo22elq7ARA2A13Bs+deom9JjZSE07Z62jhc9ABONjMVBPqg2AMRqxo9iR
mfdunv7iHfv3iiFevlE8DyKBL7Br56kwy5Tpg5Ku48aFv7C2+PyWzFd2qyGvqlvYpmdJeuCA3b+F
g5qLlxWwvqyyG4xlrzxCsIImzkLYoAXGDHYLPmn/esxUtv4PyDGYlQZW3vwRXFGVzLpGE3kARCHR
l4NQWr2HYM2PXifrx75KxppoSnKvc50yzRUW4V5aZPJZEEA2qjJbuYssBHILef0Etzyn8lyI4H+T
f+HKcHpYpGV+/ri2Ri7rIQCLE8FMBBvR0jGi87EzJAlzyAPOfXOcphVsm3J6E++qHJR6SvjPX9bR
K3m76NZ0pE6jjcbgLHgpALgo4enNNjw0/8URgw+XLJO9Xlyf7ZUDZSgo2Jl9GKSIeDg2iNa6E5MX
DIVMTVmyVQ7oVogzDOrA4WplpaZWGJshvxurVjs5i/rIJNjjlADAdcp8lgys/vhBWO6oY2TRsI8X
s5kbB1vHR2Ln4ebp339B4R/XDjPn8DRjfL2hAx9V0QvBbR3JFeUcI2KwvMuV+9d1RBtXM7UiL/So
Zb6p1ApTvO+LiaDuJjqSXAI3gQb6bpzNC3XTV6KZQRb553bbLmiAM+S27zJ16um4Kdil5AEWsmMH
CBCcuA/72M81YGpIbIj9CfHqWnQF70gitUcw986mPFeJ2SXMDq24169ttI0OqXjjQQkIdrg1lCS8
oLZDHU9Fz1ja3Citrnpp2OrcB8z4onGoXCXwQZlezs7FeLfyvZ12dYpKweHy+zEql0ewWbb4SXV7
eOv8TmhacjdrZhisq4jCSP22hvVgXIbdfB2epKluNDOTn2A9XcXmHMsjSw16sfVEFLNKBK3isSa/
JhtVVsPTr/TqxVRESEHsBI+05zVsLHi2as22RBVRLTyqYvQzkDLh66zkJp6HYp84SFGDKG5HYB7k
GfpZoLEaYdCK3dIrXKxobJ/pBOjPhd2Kh3RnKcSLb8qdO2F/OnoUdgDB1YBbcMY7ZLR0G6UX1MwY
IIbySCrKqvLgGlOKfHCn/8HBo1xlQcaUdzHR48uTYXecwEVkPtDyV+8YDJazhm7l0cy9jTs3GjEG
iaVTp04TeMB69db/ZEZxahztNntoUBeTUinVlw3a4Pru7ARBOYUnTQ17z+xU4zevPBzQ+pRbS45+
KHhq+3CrD6QS78DLbAxyT2QGYeg69Og+PHqMKKlubV90rhaiYWREDNtsPbOKmLFb/Iy09qN516iQ
P/7nSyyxtEdmo38oGSPhOWye4CQJBSsxe4B24Sx0PzxGifLOd7WIXD5ha2K0Zl4UCONhVw8YSv5h
1zXRl4VEOxUCup06xpv2HGLIuFaX+yI4CEnwFEjcKeeT+51prLS+ibVyLz7Yf5GJKgQOIyHNng6/
zsPXGeA16XbgLX6OG5kApFeyiPADZcz7UpHTYl2ksoEMabZMW5xg8/GrKP+Xh5sLtAkTWspiQM3x
+eapKC5TAV3z5ZTiyMNG6621anKL0f45Fs5cApfZiLSKibZt2IWIlp6k24lwfQoO5lHdZ5p5qvU5
6EfTdpskgBB1AxMa37YizQyXeTJuK82CoT4ytmu68ipc/v3Y54QPWR5/uRsI5gQ+rB16TWOFi/MU
eo8mBItvrU+28yiE/1z8P2bbh1Iq1xv4R9uKon7myoOI7iHcFd/5ulJ5vC9H84uSMInE3uXEsyhW
cPMaHuY8pUIkMVg8ww9QWw1a+bF6+V+JWcUAzT7E9HWM7mWiW6lzESp4VTNCH3J3IWx1rwWaFcW7
1DJax4dJHtIHVh12LnVZPF2TluD6MjJZp6El2gNXDCB8bK1hRbAKbfSvlI2NmFuX11s6LcFfm8Z1
MYe8cv9Rtm7c/0B1IzJOiVUQETkZva5zrYooIORHmm2OGNXBQFZAKjhzxTgZ0LRAMgmYuCR1v1qT
WTsNvQOj1DtG8CZQHOkhIMK10D64CWnZZc+dKGn/HTAbkwCPBtFT/kMLvl2smnjBfkAKfIfZaplF
UkWpm09HkW0eB4yAtt6noG01i286DoMGYXMpKOQs2KPHgYcQqn4v5GY3/N9gJuRFLtlgcbYG81Ez
/STnmojzNCCsTDT4GzQodjqhplePJxrsLBC/uWKR7OldLSjbjedpvWcWdqdI0LJ8DA0BDgx0RLMF
dT88a4QTfDJOlxhjGPn1x9ntbqrrGLSA0+M8lEdomarkycZIrICD7Hwfs/G6K9ibZ/mnCbuTk07g
eXWAqJLj3+f6IiAzPZlWTu7JZvhNr2yZcpkRWKfYS8nsw3vyqGNOdXugucLGMU2GvGjBccwQ5Z6F
vgH+rA9XnWahxAcvLf3YWfX6sXOULlXfjrMAQL3uffKEt3vo6HmgjYeofKxubQ3rwKoKEwdTAxHL
+X2njxF76yf2BDCfoqJEDxUYTxTPQcRcdCUIj6FoHk2o53zaIA5xvB7Mv4shQHIkuWjpM1VTLDHL
dECQwpWjOugth+B6eBJzm+33PKdKGpoIw4TeqsIOnj3A7egaKeRwZRsLxF0b0YJFBXBsWX7dtwml
DB64NcGOjqXIU+prXTO1rRBz8NvuJRgL+WD+kCEqIqs9TNbFBUJycWwwNXxeu08aGhubv0vVE2Xt
WzcgNPCpaMNz1spQCphp26jaEI1tG4axWBxTK0gUoClwvVWvTjEVY4a0SazfOW5Vs8yx951bxg24
sjM/UtFOQoZdqMCUhmKqBN9mIg/UBmm1dlcttgIYvOxNa3SPWWZl1fizdhcTnp4rnhnRx7Tkt+6S
UtwRtPKTIS6cYSRCytSNHaKUE/gqRyXJWBTtNnKkFGXhN0RAIfJt6hqdt7B4SggWsfqbNK0B/7OV
U6YtmKzK8FAMnntxLCGlYN4QhYS7Ejz4v64BvtwxCgbLgn8D1xBrWzpkyPdKMrcPxJT8N4W6rzL0
OyEBz8QqDXJ8ArhvDY0nvm3m+XoDyaZRwMuM58LN6HQGzunAbgBX9TpcmwVCQLde2elQ1WQlntjQ
OeEq3ntF9Uneok83xqOiHI5+/sv48KIJsz2jYhubpBQbEXwH6JvgYdLnHim4zUR1YliIVf/es+An
yJ916Z0wx2U+unf2LU2yS1/joWMXOK8MRhC1kXgIEt/8zOooULoE1y+v/2RIA2F7djnztLgY2W+v
Hm6UrOEaHA6ftHjMMoXh3Jvxm8B97oeLJPRkbPgnfxmoqgOWhn0c4FBwsQ2TtlD1eeDnBWPmeK1g
R//VpIWl6nmmGoXvYmvQebErnSkLiBkUT6kWhJuDWAjdiYmUDXQgVMWR5P6Y3wmJCkmZ8cfEwt2h
Ci+HAc3Z9HNf/7zUvQx832CyxSRdHyPyTYwTTkASRSp9SmRNih39BqsgoXngGNRalZftyM41beuI
PpsVOn3mgxelQOqpTNxKYP/MQjy7CLmliyxfM5BuEAWsglBUL61Yulp2En2oB6CWZfmRVN/Khstz
wwSXGgWrSNJTtk135fe0qi5TD9vcLWXcuXsxW2TsopRm4pTOi60MpOdqQkD3aPhn2z0k2PfuLc4J
x+LFancoQH6uyoEVEpsf89uL4Yl6A8rW02e347WD1lwSiSBX46CNGtvS8fTuxNfx3O5ys8sVQsjQ
aVAG0mgx8NMru32Ac2P4tMIP3RmoBMs4PXgZkf7q0GGN9BOrm8I7PCMpVOPNJrYTPRnZs9tWfnqC
FgpvSzWRSZixraIHVAfu7AIdJBS3tQZcU9eGUzXO/EjxgZXWj8udz/98MODb9XVglt9VywABR3WY
3Rr4mgenq4f2x/SR+C8BUD872l1D6KrdybX9GWLtcdRcRpKBhuoikazLzrsMeGaJ65NWcjz/7vsH
fqBKjuCsHkdGl5wPwbr0ivnjXX1gLJDz/qla8J6xMcoakdZTuyBacXJzvKrVn0DeZEDkDUfusQxt
AM8ImBipfY0Uctr+Bmbpad48LoiDYOGYC524rHm8rRnMQZdm0vfrira3Rm1brs0yCUqVgIBtNMD1
ytcXyWkHswOP36uT7+AAO+b8W5J2RZWWd85I9UvQXudecW6RuMd3k8u0tZ7dzvq9UtAtV/aBvR0l
qFvcuxegMffsKg8yUg387AkGrFgBVOYxyCIfa3+TOvQ/FF3JjVEHAh4o6OTYZmicS2HejGerOPu6
ROF7vpvWOiJXzbQ8uBoyH/HVjKvnk+6t60ktGhVMEpP1ZUnfvBZtKBiNww1idf53Uvs8/+oV3IP7
+e07d7gfUeyQRA2dIGm41zpsU/eZaq4gNhknrxYwRmeGSwIiLu4aMsh1GhRZCYGRbMyDVQflUklK
L4RhWzpZ7bsamH0x9pTi5rEmIVJbhWvylq4QyNNdGUlvfQBC7HbDW9dgqJNVSHYLmfhGLKjCla2i
VPq4uBOY9/KJaKzMMA1J5qobcGZ5SWbZoqU4nEPTU3g5OHY1bVec/zvFaLpm88eRer29ijAcP8r1
PcETAn35IPS87n19mRSujwqsZ78Rv8PQPmIE5NPYyvUWuAh/Lp8I429tElxXyaeuhjJ6v0MKPpx9
QACkFyrZ5ooM6wYyNEv168mVZLQw7c2J/dcrrf8Cw26KFg6BiE8WCkDGO76NYXYe2BKWpTg+0L/t
W81haqxdPcc2EamB2Q2rsd5sWzXCg60l2f4Vw3QE2YjaIR1H32e0Q+hFFBdYSga+vEPhhw6WfzF2
dPiRvgBwgMACmw0i+zKiRKw1AjHaJdJgcomjvWjFZDLcBbQ7UgYiA9R5M9H+ceiD/TjNXHm2DfP3
kRPoKuSXXVqQJFN++Lz/R1/a4vk5E94sVr+r3ubsbwCHfn7Cc0+j337h+W09oDKG3Vs2myM6kEcz
ZYYl0Jkhkn/ATKCIOaPzBiKUrhJS4/UYiYz/6CoILSw3GxF4j6LqaYJCXV6G3hpZr9S/kg13XQR/
/R8wPA6TZW+lMnj38hP7AR3NbMoMKivpE9TstpT7UR4UWarjl54c+c9DnlUpWFYq6Zzd7ymltbgg
OHAMaW+OvwWD0/xzs/1ikKYbWeOvrAgKPWw8ZBmBJrqU6lAVjfFyrHHRmHLyyP2uGVZ6+NuVqHpJ
8YzVRPFTm5SyXgxxmjuiEflNQzWmQV8evYPf7BKj1rBiRN9i6DgysTcLIoKmUxWrswj/yL842FzZ
ToieOEo5AU6te+n+6jZ30HQiCzPSeROM5vA/83VBIsprUbA2w5D4wg4TjFH0VnSzkMD+uZ+EyZrX
/I16s89zr14eNNPJOGsOidv+XYPpNpZsVYxvevdLuUypUPOzoaQPpPs2WeqyTGA6nvVf98yIEXWm
EoZab002z1ng39z/7AjFQ9oLicwUMKHECmnMSyd403IThrFEJCLk2H8SrgI4qYMb+fPvEEaa2VKF
JIkcmB9ELYfPH74VYzdIOkZpkyvNp5WaGnHZoubOVv4ow2jdTUtK0MfRpBkGvqgTjqSj5Wrn7BDT
djPHRpu0rhOz/Ukpe4iWWm3FpC7keN86N8TlpDdsCv3Xeh4+MMxVVV+WRDraZJNhq9n34ZfYI3Dh
ZS/rdBYLs5OwjhWWMPbkSykhpeOYpxXoJQ/1ybB8kuyVbpRDVctF0n2L/FzqGVcg6QalqV/Xbopn
AiVeNkW/c21o7B9nBUawph4HAbDpy1BBrsTF2zeJ3LGUWcpAq9OTYWL9QgrkCAQBmVI3fW/SMowP
fr/KgulZdJLLGMbYrk3le1Qg8WOBuDrbYeqXYC7kt72I6oUTlUMpunFyt5iajK9/DtTWwOkji1Zi
+tF2A6tVGAL+VCBa5HHxyTt8GxPEFwMcv8+MJ/Uf1SzlnB8i0wiX1C6N6d6lvGF8PztNnO4J+Imn
V1Moao+Syc20PdMXfVPx9gcdeSdJMMDSoUfaosCGQQuy9pKDMXYBMpnwsc9w0+tmyMgHNZ1Feftn
0KRBBtDGU35iYSC+MFCphqCREc+3hqe7kmNpKvrZ9qil7+HFp87wXdH+Ub7AGuE+i9WQyH1aVQEP
PNChOO1xTSkasT2+GvNqLFbMbwmKSdCDiX4/OoRz7Mt7MHQYKY8+n4m7PGX+jHDzXiouyKf2z/12
JXOme0ipN3GJQXx6GFRfdsrPrpbswL7QFxAr9gVzpKAo/R4RJ2a/Fhys3Wp7l4Q+dfH9HDH0gr3o
N25Af7XjKyA/yT7nc2DFREy8jZd+d7f6dUq4hctMfVNR2wNN8vKLLgtxDekxdUcLNeWzF+wieHG8
aPKXqLeiAZ5+tp8BGdcydjUNpeCi7E93ZG6OTzDGgT0Uk5RxGRbb6C8ghnEv4/Pgj7KwXFEivYIX
Y66T91G6OVkUA8Tat7Ih6MIv//gBYAAax+WoIdguPbTEM1Ff8z6wFMVk6aJCGn4ZbCAEo8UNFJQj
NSXkkbDu531QSwNgjhfLVOAOh0r/uVK04H656E+p2RxkbrSNBiE9JsYqTrsuzLcfNShy+8So2qHs
pV2IE1qdvZaxCobv2fgx9sm60fRmv4wkSXkrDx/Qcm9S9y190yESKcXgr/IoC2fcm/IM23xwcQ+j
HCoZ3JIfW9Z8wNi6A0TXAnKcWGJVrzWWvMtDHmwr15hJndN/1T4+mXrne/gik0D5mpRQUNwAL7vh
Cy0IpzCAD7sNNp0ZPOcG735q1+1fNVasU3+2XjSzr+20w+azC74gl3GXOfVB2UStbXNDr9FhUJLN
qsuVtfO9G3wTR1k089hqdjwt21lr+hzfYDu71o9nMmqTuN67KO2L/FvQKncvf7sb2zHIhV7ajGV/
Hpe/t8FtjiG0l5WopzMkpO+jcgnBgQO9jk8e7HA7OHvsTElNJMSn4T29rLyAkCONlkBZXoRDMrHC
y1wbYUEtvXaOHCyDd70osnwstd7o0HeDHSyVt1PXFWOa4Gm+iyaoUwUm9GVNuijAvnGdMPrG9Gwa
idQtm68RfS6aZLJPXrK5sRBwrV5mpJaZzOrO+18MR/GXkReSAA53liFm6OXug+XIZOrATo56Kktj
EmWGM2Jcz6pFLg9Z+VbGLVcBV7OCn2VXPwli/R5+QGeBGTN0KbD8kLKOjtfdCZRaD3AKAGnqfMgn
SJ973TvXvXdG/9sMga1DDOPzjY666LTaf4hup9mFRyRQsCXIv2NXWbpVN9Y20CP8PrujVxnKxFju
el7w0Im/kospVOhmn3GfjgM3ShUyrCeNnJ62+mSYF+6Ri/yboq1x3jjN501cspwePMtSoeQOUb/R
TS2p0v2bbW2brYvQOa8bYnq0HyHSb7HDJti65zB8j1nbLcWPSPzPHceh1Db9X5yRqjK4EcjvFQM+
bPEtMwEAE9AWl4vupNCIG3vWVfk56hiOHJG2RPByNNk2qg1n54iAPjDVZS1CvqRSG5A0BNrn19dH
Cpe44MOJoq5HUhQWUn+in5+HpPgBa+zf03rSWMe3JrtO8ZPaN0hyysBLMcg+CMK8kQwn0cia6fHh
7Abb8s72to4VN3UcwpJ2diT9MReiogLTmQqCFxJcV87sIQQ+2R7fiE6TBceZ2Lajr93O81illNvG
QHaoitZwLRHrkuU995itKNjANcZsbOJXqL6VNHr2CF/MbzzH9MUVJEc1WU2pLu7p17r8AEfH9rpm
7cRsfJGyvSlB5Tw1un13pRVo2Lv2G4KXe9o5OWwUXAcSkSdoBXKaLn7oLRhBG7DqyaSpD5QxwmXx
5eQBtZIzh6oXVRE05tenvnBD/RcVnICp0CPovmzmVQ6qlnVqFqst937C6OC1t2+1dRcIralaXYbL
pDi4Yu2OOEqsz54u+ze8N/isyK6cRJ5r3/zlDtEkQAw4TqzUksmwu/fkjf+9PmDITtYx2k6qe+Rr
9TXyoxpdcT1GwtTLxskZWcB7P02d/TQFE0rC7vsL1a0CplmTYAHamfHJVAIPaROAg8LcXtKFtJQ+
sBcCIcICK5uXfb6R17ozfJ6H/eR2Z3J7EF5k/JCjTiGoboVcKkBAarkAAhf+vjrHrOYy9CDEODB6
buWPtrPfJIDDDeLQWV0qMp9wk6DVcqTlex6bE6cMrJYYngko7cTLFI9ozgH/fWiX8DDFT7qNDYVx
5/otWPAwZ0wadgtdSjaUCGrmS7xpWH3+CpGgCtf/7LbP85zyvCE2QZCWswbpOV47NKgFLgxsdbQi
wW3yMzcfURlNAR6Le4ZabgXIOn67KHxctO6ROLySgZU4c0gEucA/WRjeNBadro8k/IpWEossszco
fhuCGEvwxzV8i8M/KIivmNpeqMHLtDutO2BRIo66td/zqZ/6X/uFY3jQVghc/dhqpM0ZvjODjnyj
ghdIRx5WLRXRUhhomLrbChLMmWh45+jmPLCY1QTMZTt/69XcXG4ANDeGru+A0zrPwJ32pqEnoYSY
29UGndGvB5X26oH1WxfVGuv8r3Sb6sIjc9YdzC+C2YaV6e5Nu/Hcr92sT2+pZ/CY3Mz9d8RWnETD
AaUnPo2LfXxCnpCfSZUGLmkDc8vfqZK2kNd42A/JQx99O1MeieFQgv8BbFz6nrHTfm820XmLREc3
nteVcoBrx1nfBzHMVxX3C5LYebND5BBMRNq3ZdB037FyWijzNxM48NiU1JayMtHGUu/fTnAjCdcI
BMequaMSgV02ZfE2k4ycNPU9wD/qeGXXcqNG4d3eqablhSf5JsUr6AfXbk9mDF01CV6tIQW+hg7T
ByuxJXOlZXopDUK/WiwfXfxPQfdoi5JbdWd9etiF1tuHrvH+BoLQvMA9+d1WtSGBftHUAQe4flPZ
IR8YB9JXOfoy2fM/szkAsmyP0cApti6CyJihpj4XijKupHB036/hVXZIcsmKnG/iedzDS5rg686K
534GTkm8UECBF6d0UjlVrXYohGZIM8JAes1EYbn/dcnXP8PDByPCl5oX1p+6zfjQ3G/gpvWcEhir
Eiek8oKnoPoYRJH8GfHPwe4Z7CU5dKaDR0NO82btldmqHMvJkAOAyjP1h2JuaOBtx8gT9TJc5uz/
bWbkbVhzfpg25/jvQafXlQcs9n3HoZ90eL5nQV1Aq4XmLDgxHXiiskvOnVLJ53MX4SYRJUYAvw7L
rA//ZGPhl1TtFVTF8E1LEBgX9BNe/p2aw/b1/Qpe9i4ik9VyemaQlsTFrlIkxPrGBltUFoeoZvsX
PzrrGKUztm0KQiwR03+ErVNHTDZhH3PR63K57pCs1NB+JsEFsOVew5uDGrDmQZgpsGFmmm1s7vH0
755UXfgJQYy9EFTCowFhdLo2B80nHYF5qouV1hA3G9h2bpstFGcPYDaukc/ReW0+ABRM2ODGjHDE
+4bpNeowCcPA/bxd4IdVvTkTyoGmddkscFMeTVrIJcX7W5VXyWT8PHB4vM+7D0DQe9H89Qo0tCKM
XvRAAZqjnA1qDFtEiw/HyQTtMgxy/88+t33NlnMrQ35rl9B3BJ/dEKguxTiIAjZqmSwrRH3swJdV
DAy8QynreKv+iL9AS+lj3ogBgbkCa6SNgF5HbJ8lSedDcpIpsTovn5nTqrlTXFr4cqipZFDR3U+A
mCa3BYTghZaSsC4pJJrXfcWnokYm1WQYBPu5ns9pYAF7mMdDeVVRovXa4nSXVSnoHpjtEV/MKqvP
mlaMXWrGu4q4vws40bDHaYeek/uvBp2YXjpV7eEf8I8AziI4WwO4sGB7oidUlvOXL7U7p3cQFjH3
+FG/URKd7Iac66D9F46gbEbUkmuSV1xJDeAUmnV+earXhJoGowCPrKnhHEKcxPUc+NhpX85ZxYbq
CFQoWGgs8T8OFgAa1SbnGgbGxgiyXGWf9qgDBJIhEab8H9zxUtVit1CzDDSFXewtqaqKLqHQAYIl
UXgFPaE6AbsNHJthtD/tfj4+MhTXAI/CGTamLIADnl0YDzLHU2/Y6ZzAT2Ie0qAItlkMkH93kGza
DAPLbgRqejiwAcDN+ZGwKr6zJPf8rYoiOO93mvpYhNE63lxDRZnGB4qqdhATBO5YJ6Pa/+O3WS99
en1JJ9RDUKBqzKd7w78DIsHRMQu3c01mBEsK5CB5pa+j3siAOzx9PTMsekXQym9qQzpwSPcD7qow
CHCfdwILI6t1Rr+Qb8M27eGTsJqnfWyVZclLHAzGVaPWYVx/mBYbzolv+IJkJZWU7cJ5nbYZ7hnp
PE7CmYyztpKo/XYDJjz26h2txL5w//cbydO9s9It3nQaSJ2VX1elZ6wBxaIF6h+6UYJa7sBXOzsJ
fkqnqWHwJ+TfIb/WwdtMuftBsOgvwkcJn8sIiyYbnGBqdDMyQA0vh3FgkkuhnoVNUhZkflEkhQAF
T8FBwkFF5I/AjhWQJrbGi3NjDZ0v6hffI/yRNbgkOl1a2rdFWgvNVVSNX6Zv1sbu7F54RIbGyQ7L
GC25EtkzRazbenxehafd/QBd00EX1z09ppRxV0oSkT8Ehbqzz0IgNFZRDesqbVtskTVhcstK8Rk6
9E8OStfBuA+TTj9MPsVkl8KZE8AN8JRkUBrMIo2VIJBrNnD6GInPDhYn2c4qis3aYHQHLZodxt1w
zDvufL76hyeW440ZXKVD5PvcFd+eBzY2yvo91/I4uWWybBYjUYq7sXdkMqLMbA1G9EnKy12nFo7A
glotqcGhBvk+8pOSfgBI46SDtpLdjYwOcyNoiO0UqgnV5SLOtkCA/qCg1YcQMPFuXa/EidG61pQG
6W0klfeqYWA2I1MnRBY1b+8tRJIyK2qsak7DApegknqoZhu53uDPtZ1xghjbyvYckarMTyHyWmxw
qWHwHcW6+RRKzCTFXKAVPsMPN3JgzcL8/3W5xuulLYvEl05Y5O3qHu7KeuR6S4EgCqG4Bd8jsbs/
AZ+fmEg67YS9P4UlRWafNPIdlKpx9MqPj9KdZAiXN2ZDuab5f2tSQuoIh3UlONCCdBgFMsbcq72E
nDmBAZhESilP3IkvxmbWwsvDt91fVmsY3RusTyhv2gZV/qwF774k6TJtBdhX2ao3jg2N6xgseuc3
eRHfOe67ZYntg/aMfsxjcd0mgU98RNfp+S60w4wAsHqPY0/hvJ/e5SdayA+jNpmi+AqhIBt2NehA
qcZtfx4NTOsOb3DJdVlEUsNBzl8n0xAwpH68dTm397z8wy2I1fvlowvG0+rTml7A5BQnZWyL4Nji
OUNa1NP/itwSubfHaxenbQVpo86ciXoBW1b3vAtcszzshWZDtvp4Jt/SK2HalEeOQ4/ts4Lnj2Td
heaVA91t6cYUepevnGC3ZhVtfOYtzF6PZeyDjlLUpsSW1towO9LMRZuK+V0FOddB4hzbIVlAB68J
6NvKU/8BTeWfvA0qbfHW9FB70aEdOyxt8YjpUOIlhV4hMPjwX58dMP5fm3xlUfkC1JsYZCSZfiRx
160jAy6inr6nBb40GhPv3s/K1OFyqK57ifgG55VXYzY/Y5ACpRPiZ8VBMXxFQj3Oyg5SfNURkp2/
bnMQODCT0piFLPtWeTkgO6hhyZPv8jOUJpNFzweMJdYXhzS3Mv22fm4CbmpqyvkttmtCvcTYL6/j
9kuGvirp76Cu9YWXFAMC2hg15ys/ZwveCwoenOS4cNqlxBnhVkcFVeUvfCmO3sKMQTBbQwG9fb/e
tAT8uf4cSjeUJYZtToIzlSZaUBHhDhXNBYfF6o0t2lRBPQzArL15EiHgc/YPpEI4hbGY58apKaqo
ym4nm/jXIe9hFCdc7DzLROQ7QvSsGftrHOylHUzHuLrdB9Qdn++QJ0qg1y9yyhyifCgqj8YhU66y
/13uMvlp6N8WVoaNTouliAjRRjyLw676JGRpAYKJd19sodi3QYKqgZn3tom7C0Yg1oNs9n7orFPg
R862TGPJDffyUeGGQzjNkHy91VxyO+SI7g6c4twdmtyLbL2NGO+zGbTMmpADjjHA+xJAguw/0hI8
qtmrMQC7PkJNUj/As+yD3e5fReQcPkQwaO3rRow0ts4sY75JVOyJ+f7cxb1+Yo9CgJYxEr4AZjcg
+VGGittlVJRx5b7Vqg+picRw4w0yLPL9gGiLu6f0I5enzq/KjX1tWSf9Vl/zmitmXYyVZ369Blru
sAfKaqRKhlGjxX6/NqEx9k6rBVDrGFmjkuXmpG0IkAErQKiQ4IEqOgq82dkuNhyV06Wc2rKlKulF
5kUhY6IpWLQNWoCi54vJDv8mFodN1cf/c8L0eU0nb9jXhGNnwz32oKdjH823RaCLeNDhpSF+K9GL
cyh1y6v1nFmZ270QVjO/of1yDj5t7Yqahz4eG57F/VWgS6D69p3rR8PyWem04dBRQ8ywFDsmGO8O
nmE3gC6XuMN7xURV98n3ST23qrkpfLpbM3jsTToZvtlu0AcN8GbyomyVH36HclHJWE0Q6FkNcaJS
m1hb+ZkOabZePslbsjc3xr8yWmYvdWkDfg7Ybn2+fDZnZyiHwviZ0eOwI843rbaPY7YQMmG8iVVd
/reX13L6/75fH3ZSQfeJ11nnupm/bqixG7Steyh39NZC5lLEUSRAzEF/fIA3Js1HWthtVpqOvGCu
wT337IybRhZaCr1Mq+WzrZqIAOiv7lxXtV+cT9IKRWVH9PVKZBWQ3SxJbGFea89w1XWifen41kFw
cPgzoChGS/W+mQMmMNcdcoPN9403KvZ/kf8gtQRXXLb9oBp19HB0gqaMAmNjQ5CzRHrcdiSLFa3H
pg5gS9evpGp0Dh1nm/F0hwyeuGB7SL3fBpcRAbNyWl3GprBDqDFQ+hl6PpoNJ8+uDRsEY4ctl5/o
PadLqCvFWpZ8hi8R/+98fiWVnxeKno8jeYWhgKavNC4yoJ1qukA1IYiiMzNYPHJG+PEoWm1oBRvJ
3nepXtpVWUOkKYCiPD0+WAAsS2iad/BhaSeJoodHnJN4mTDqBpQ9iDxlWMF9UhcduosT49oEL1K7
Kmeqs7pqGd+8ivr6ueMFEme6g9+Zqq7GUBP41iIQ3lqEzEOO6C+0CWWGVePGIAgQGn29/MjWqkHG
aAUtDu0TnhV5skQlzQkTo+mgzRDwgKYS6sCgizIYfsX6UEEDRybQGsELTA7pjeZQtjvx5LpMPYSO
aOSuf3jBUw7TkBpFmcb2vSw4rBgY2ahEQG1LWUkwA/R5RRMSK9mwSTMt9y+CtR7kp+ZWzjJpEcmT
hliY5TXaqm5OSjOZ6HOSrRlDi+OU8xvLzXoe0S+I0PU5WaMv/0JTc1ZqzqILhv0CU8LptUKZLmht
yweGZCydZztV8UCA8L7zTplipJdhQRVjb7eKSsgEq+IeayKbmGoJ8tcRVyrm6Hn/AZ90mfX2jJf6
mMerkkIw8bSunMUyjiHXwUlZ0Mfmb3AoygFyLUV2Pb+WOXBSfVz0cly4Ogg5ShIIsBLnIhdnBDY+
LX1wwgg1zlefPMp8VZfzPvD2/lEjMAxVH+Zosv9BTyEHpeC0QziqitcDbeR0aKgrfNRDHJWWwEw9
GAVQN9gNpqbu7opd0vP9PDi7tHF4856jp1ZWYQdxjPNc6xgnyOyPcvRqjt4D1CtoVf8sP/1acBBC
MaROn/dxl+qvgouwfpN2bAy76EjCxOjCIGQN04F2cjA1PB3XkJyS5bj4ynGuZZEfcIwrYNqf9nFe
VUuX92SQKrAS93R0kWEgURseFsnpisuPAU9rgXxESTWgPrcRdm6BbdmvekOblcoYSwYIRVGuAigI
cZ6JKPsNXBthZchhEi9tj0oD8MwxL1Nmp+yvd4Sn7sRGDwgiK2N4ruAasy2ZYLdmfhj4l4y8JBuN
YL4o0ds0pe6jXCjKKxHS3Ft/ClqTADWUbjqsRUp+HqomdERRQ1p4dk8F3z/2R+yUGGnIog8ii82e
+urWRlphx/C1otqq7hM/2BkCubPDvyNcu7IVg2tFdQFgnQ5YToiwrHvzFIphSO+P5q+8H3NoQYqF
SVzo21B+zgQqEQqTRBBqiqwpa9m7BudBhvsRK+/iz/L9kKXCWYXFLv+ED8SZJYKNkkVg9i71Ack8
CJpK3XcrV4QiUtya/f/ACGoTAiwvbnwFk4hkFtfkzc15VZGBUAj71vbxAvki01E5X7zuoUp+6xU/
uUvCP6vnH6nMRTk83rfcJfL0HT17jERtxBjkjLlMjLPE89lQK6jWbhjX3LZW5pKGahjn3JDq2Goz
kyGz8fKjrxbBb+sKDNNgjaNBZmaQDde/fHdk4CX1szfcoPJTh+SjPCpe+MFjoU3zI1O+BRwNaf+r
Irr6hD7GHheXaexAnHGdjZufTmVG//sOxy6Lnx3GTazC/Lmvlxk9VHs2Q/tauNzV5coX5zQunYVB
3kQa6wtOunnCeNaoEdxe/PBcRIdbEH1oFRu41eiEglKBzAfQW5BXJq2o9C9HwpLFdp2HTcM9mmjc
ts0rECbvEbqtFir4PHs2NsAmyKHoaa/olMYs51ctqpD5mAZTpAsxQ0mWThEJt1Nn/9vLLW1KRikE
plCmGGhpyQE2ee92KNlWwEFsPoNTRAaDSnwnFDoqMVDHzHugPXd4KRpVVEYMZYPwasc+9SC0hWWI
SaIrXX6V/BcFDWAfhgBtmg5crmfDt0GqAUJa7yf4NQTHABa4L4AejzCt7OM/RtJ7484xt3dHKr7c
deTFGIoiK6hEDf16IA2wZUgplHDrAWVGzZRpYv9WQLGyIZH8zqq8I3N8SlzE45oDuQvjRYtX8E4d
yPiTdenQPl5YDVXgduz8d3AO9SDoWV3D5rVffqCV+FsG6YSNLOZvQ3N0amIB3yXIVf2jFC+cn1dP
xOPr8YX0wC8x9dRnsHt4gU1Ae6xBQjWu/qfM7XFV/+q5q2C9O+6pPgbMZcAkkxcTOs/xJtxAQRR6
1FkelcHD8J0o2jSNG+DiiHBt9A8q2ZMM6RdaEc8ajoNclCFGb+5EGeMqPzeAiU8wXF+hvLh5EEBi
n77MH1V7l64cYep8zGAS1GdiI8/518k+xjUmnuWGR1QFCuBZJSd73cxPDwUAcNpED0udgOF9KlyX
BNhYiv5O0TJDFjL50I8kblFMFuegRAEVjCejrSZUXdv7AoJICMrRQVqP/PnEHrfRJTivvzZrTMPU
FxWY4SAoQvrgqndvC6pLcsNWeJDMlYfrralNi/QwfgvihPiQhyCIq82Pwqe46t8f2B1znNSVNMce
izlFhYgC08iGVDMkKM+tG8LqDX/6sgwFZNyum2U8G1VRsbWzyNf8L2QmVl4UFiPzI9ypjkZ38i8S
JQQ+WY+uH45x6G32vh9+TYE5e3o06ra6TAwPbexa0U7TMm23JGlYkOYcl/b0t+fTHN3+jCpb73xQ
ZnAAOeExPLI1vbZ3HMA25Gd40IghYp2ZI4BCejxxbmQE9vO14SCnoyvWENCB+hER52n1QFWJFDCb
UnDkhqcupA3y0js0E1WB1qzxJjhHbDFoqqYnv+9Zb6WtQDFXe/3OoR0KOFEJe9zuHY097KSvxdYx
Pamop5BhhyrhQYEOtwlm4+CRIjhgTSa8S0B9Q0qEeiSMylU8I7We8ZdyAmjfLYxdXGkL6qXCLk7z
6L4ZO5pmAOGS20BWidktV59xO4wiGkt/o99sJIMRWzdTX+Ezq5c5fhxGQbo2BYjAzrnr5ESn1Ese
+ELEezndIT742Ctk5Q/jU30WWTzIHfH8Pa2ZYxmmPFgTVBVGMrt95j7qr19i9uSS2Dfm+iRgwNF2
a+QDTC1fjMzKddY7vMtlqAdvtoOBAMqah2jXdXZF93pnsrgbIngPhmfR10WWBE312KsSbsCpAFYc
4JPQvZB8T0nGGBBsSXO9AQjAAoJtlLRAt2pmi0O6ZgnTYmfa2QKvl4Ak6YrtjRc3ezSIXjYJm7xP
bkuyHyy3a1N5j31vKupxuyjYr0iNO1TtbXoDfKRIIVQBye8mc+6HgMBKG2iZr7/rPlSKrRceppZi
HLJJcRQSOussSQW4UWCP4X+3C3G/PCcTxBNSbDKGkPY4EVQVIZ4Lae02IAUbJQO5Wj7sCcyAsvIf
rmXcYn+gcFzzl4bRc/qq/nlAcJ45hcH7C7Naqlm89KFDDpOE0wNq168hZvHXbc/ps5k5jCrk55Lq
+dvgpMpqG2vlef+aJel+4C3Afr0fj4q5E69YIFSojx7JuhEFr15o9aJHNFMJt/yr3+hItJOTi1TX
izOEUgnb1dAXKjrRPzMOuNszbKPraE9MCPze2psIUkvOcq4ZjtlCQ0cWsQP1o9ViONdMJvS8bUxF
ubtbww1t6ALASQKFCDDaKIpC9rKJ9Qxyk6ynfrk2wshUoza30xUEbT9NDLLrMEph6jLtQZ4cVI2Y
OFVGj4gUFQ6NENReQ2BDxdd7BdbQOA4YThUIowoLfhGs5o1iLzwFbu8+1ajfhBkIJsYtDWyVwJed
oBUZKYAr3ugubwwTZfnz/QcHNlR1QhmAvuKr3mSs8SVWvqh7Tv/BqyUYZRMWOi5xoazvmr5izVWr
/TM0VAAVTgeb8TXeRAMrjfqWj76x5/k39tD4oDhWe29pgNhP/Hc8nK4TWN6fYm34g37Z0wqJBXtk
Y9vpK6kHMg/lcm1baWsu1IMxRvPkBitEjzjP12tZNtHVKPVNjPRIau8QJK/QCpeeg6ToQaAqa4d8
85DNPJOESttyZaHrkUH1vb0ihDNLBWQmrLczbt+ffd9zimge9h8VaZ8g39D+DdL7qN/OX3WjhGWC
4t+4r8zXe12xDtTXKbIAX96yBwMNSjsn1e+cmbVzTenLEzeLaydQhQtWjT8QZhc+aCAJmSxhtVpY
tEg7nptwKWYo0rjBLOirLvFCymxMQpjPimqi89SNlHJ3fa00wUGF9X4HrMo59aFcuEYmYd47XS4l
dqnE3pmzbfrGKKOkZdaU2A2jsVK3MuB2TA0w/LaQBZ04FSV9iJVLz7VOnEfcPLGwkMWmBVJwIaRm
IGGJAlP0VxUoBCG9WCFYlRgwAewig5mVVt6gzikEvrEGckBLZvywSyvSkoP1Gc3+P5AjNgF8WK2n
48vvtspaw0vtEjbeg1woko7OeMd72G9zHPFHBo9eeMNCy2X1qzfj0Vx8gNMS9831Qrpyl3eul3d0
uSdAyjlDdsnzzOwYu/EmMYKff0eaX4HoZ90XNyZUEAzKbdP+kj7kh5yAy7siuvXUrUzqELpVPDkM
CB01qEjneNndkN9Ddl+O0igjL/U9H3U9tiF7OzAsfNKl2oQ8TdSsXIge+n9YILum3TxeuPPrcUDC
MFT9oj2PfofkuKUUTM0OZELyTetFNBp4oLcK1mdrZRL99UmDvIy0TBOdmOj8TwK0AeToLskwlqWz
H1dPQySr8mp+uyfz6k2TfVi6C0zGp8bWfgcVYEzwDOLTGzFFobf8cO33VG45tZ/W5zcYDiWre7ry
1ME4XWA+dErFctHF1tckRwZ8Dnpm4whF1pc+CdTGSnurzLHuiZiDFM1Ov7MTbAp+g+fgRoLCWlbx
KMk8c9f400aVDYMmDUaWbKNDkUpLWtlyzQk77n/KwuFqKiFifxH9r1ur1sebh/eMTLL6HKBjN5ea
Ui68yK2Kb0oPLqhwmPNCOmWfUB8/H3x20wmrvDv4WUPmALzyG864mm2epdCKsJOBVZrR8xnNT73n
g9wBlspKJfGhqeXVComxMJJjNGbsFsEO8x4hQ3LvrB8STwhWqFJnX3n/BM80ycMhJuTYHjVG+7jM
n31F9Fd1qbWqbBCZ69DTnOhBxgaGBBqx5fpBFEhVbKDlbV//V1tNwVzyOa1FNG0zVGU60rLUumfs
I4IzAHarhCtHjoaCEXdhAcoZDb7gkj+3eWFLXNSy+WU8JKlmgwexHhmZxJHVhpw3t/VsMB1GWMUm
w70wCMvI5adoYuVGtFAvCatBMiQ9osUNWtXylLyVtUyKi4HzImWtVFn1cx02nYJj9UCFtdcOOBkM
N+jk08MjHVF6jU4JFclyXkC1gVUiKx6FpDaPFruDOsmen4xT0JeD2jUj3Sso4xyUNES3yYMk02aE
f3bKmYYsxaMhD+m/7HKeC5ZnWB/eUBhmJb/2yrBZn/XTpcbBBK4HcOCEXfjpJLZqNAyGSfJAL1kl
KlKutwWnPbB9HSm3mxS/96JBJ15OfIRJENhriKUPQGvp95tAiS3wBFNv0A2gx5XETqQoxp/pyqZY
Uiy/v3CMx4cmloOHIYaJSEMDpgbnEVu6QKIrK1C89D6DFa3xce5buyZz4squWIPNJPevsQSUjOtK
IZE4O7lAxaIXSsXuobppG0qnXtmkjRMu3FzYkk7h1/0JLlPhpI601DuijWr4z9iMvVlDKz71BVNW
C9K6k/ndZFjdqssEZse2vtJZwPKBjovGMAXP8Skj8BPz6JPMOZQgmHIR2filGeMUsVQlegQbuYXf
B35oXqj+hwPjrCBNWNgo5YfDMKBwAdkiJzYoM/cS9S8CwQT59HikIwSKoBMPU2yejraMmrnkUC4H
IFK9eMnwbrk8UcOrRcYS1pSU4A1iGtHq+yIec7pgu8BGMOOzyr72jEgXvu0nKG0xTPTNZdl8Jpxc
a+6JPfBmWZGjcKoeeIq9sd1g96nsCcSrm1AaSf3OGbNpE7TWhLbaEGQ6kazo3R8iWzYjvZjeZFJ1
D3BUjUOygnAM3e/N/umU0aAdbjIBwe3L7h0rLFToJcWryr+R9ma+eXmwH21aOFu76zsM8tRhTzqj
Wok0BUXHx4JuG2hvqNHNxq8bt2q1vC/H/5jt9jbRWg5P5mriFUdMiigpXTjiZLGB0ENtJwCSCTb8
zXAshjS7EwSmIn+I9rY9j5M0QxDHVYxMmoPE5jOZdxm/JyR8YwqQ07S/MrHM7lp/jhNqTMqepZSf
gqpDmFuE+fRT82GyAVuT8f/U+anua4hTKrHMq2yCCwHwGuTcHEwJWOSpBYKUcJyN2pUo0kPysC3c
IOh3HDEEB+D4qDFi6puOe7GukJiDjX0R87w0RoOwwaC1UBfuFX1NEbpbJhq4Erwukn/oL3dYNGQj
qvAKXhdHd8tpm2CxKbzl4fkQWKRGSxoie7toChSzCUBXZXgQMRoYaPH7uUY/DDlbvAxIed3/z3LA
38BJ2RUjInMzlRjXZKmIfwd7DTxOEijFcTi3VF4W2aAJLj0qwDUUGNhy3cnQyaWF4U3Y1daMveY3
5LGT5C0LnnTmv951P1vYi0RON9N0t++Y3L509xOKAywpe91/Vc9PlQM0fnDtXUg2zucC7OVjFB7n
W04DiPuv+1zUZCqBtyYQGG2OMMsLq99apwWfcPqX+hx8e+LCbMRM8qJGC9DjMgwtFjPAjMWngLbw
6HG389+nyFtiWctutswjelbwrclGXWB28yIZne7HUn07FTLftngJpCNah8pCHspQO4YbO3+O2nDg
w2xMqEjgQ+g3zKhlaKRXZVTf0I9YOeLvn12GZfM7UIzgPujjwQBZ0+ChTaCzB73hbcNeFPMKUz+Z
awoInh3xSgFlfgVRoW73N5VPec7W9MCXGxJqR8fd0HgcQM94ibE7YZCno1XUNUBkDbbCZWoW/+J8
Znay7fW1Img2PgKbMS+KAY1kSam+qOjnco3i4Yfk5h2Rfr9Zy0UhoSbpwX6Slb1mDeuQvJyWK60E
Zb8ZejPdQK9Grlv3Gs4bxcnXlrUpfUjuOoaG9y7Q2LO30OcAF0Xmdbo2s+sWiWhu2PoNkkrHkifg
LRlqxFVLdv7jhq5Jx+MpB5ya6KT6QAlU5KU6ZEjFZmiUmsJ2xSo072Smmor4uOT6gSeujbgxgTZw
QCIOqSdDI2uS3dK2uTyiRHCn8c52+oE29YFGfC+08WveGFpD5bGKcw2TUV5Nnv+3j3YQ6ZACBSw8
k7RBFNFTwo5stAvhgQ43qlbgRc9ckqDdLq3Ya6nJg8FKtTJGlp9JH3SJjYwig7MN6az/awo+MiEc
xtGOPar0puFtRtN4FroTm4QgYoSXQ9YDDx2Frr0r4XPXizxX1T9evujPJ5ROtFFFnOvnJwgK+190
hOpInjcMIzLhQ1fxqdMrjjYfzHaTfiSjYw8daeg5e8p8e7qEsUoBiMRWAfKaq3THyciUldIbH+XN
780wNjWxQXsGhsGOFv19/zuD31mjVStQGt62h5CHfCoQLZD2ahnkwmqBApG3zpNmN43keFj7hJP/
/kzCBDBr/6BR7teTZOPWKyYooT2ARz2Vx+ilPYbsoFUlCMutJ0vbCOh4g1qoYY8IqJq8uGN6i3a5
6o+/Kg4WGN5EcN6BAi+TUTZo1WJBDfOHX0GND/zGUbFo+gURnuisz0XrObhfBmAKwkK7I2qnp98a
Edl+8GNLyFTWzgVagO//0MJ9Cb8cRl3raZgvfU0bliYH3iFaf9RRE82uMvxTyO/tsP9EWXPgsjIw
gEQFLml9N4VlETzSytJw873kONVctKdjqZ3eBSYA/Y9Vh1xPo0Bf5T7dNhTjyQ4T3QuIZz8KPZQF
sa8jclso7tklUYENDrqN82F9+YY0aZT/7eqkUbUwC9oFtQqwLvqWgkSfm34TjA3IUJol4i5Ae3wO
ROaxPxkpivEETMkkj4hmKpLw+5qOF88BFuP6aQvCvDYL2G2hfSk0GrvxVRJsAFaRc9ixOKcQKptn
nnvzEvKeL9sL4qPOvhcGnfPYn70l1B3+D4+p00+UAOZLaMMWdVnBl4KzT0QSbH1937mPh+oKo/ok
AMBzPjUW7SOFkqSVeidB4w4CxLA+la6JxAaSqNhGSsO3V92CFiUOP2nq2cz5WBjvnX5lYjOXplBb
6lTj6EQdBbv2RzIPYFXKqPeIDtPDB1tvF5JZMYEOeQaP9lNQCtdexUNlkv9nGMvu+30jD+pv8a2i
+EWwb362f4b6FPHkgp4HgpvZuy4IeAIf2HKmPjKkJr1to8B1QYwjVwash0RV6QGlme2/XK2nvAX3
YzEUX48NiuCZV08WiTMEwYHaJcrH9EjNuD40AJRg0Ljdxg8rMvsiObTqH3k8BXx2vM2npd8pfzQz
hnGlt6s1RH16bEW8DbmGiaPHVmTSz21jyKLuBgGU1kR2axuYkRo6ikrJEiCsh/s9VFl4VulIx1Qi
h0aZuaL6OnmuU/e0itkjq2M2K/uahSrnUQFiL/stMoXvYr0sMz1qUCwywjtBXLCS4nTYrRPKeLJU
MAHrLA1UE0FRw5Rwa5zeFc9spIWADSH5LyXQTk5gU5kLBaY6Ycmtnwoa+LO5Y+7H4DhUbWPcwZv4
XiMEyooY6SjX6PWcd0OjRHldV3Gy/Pvmh07FmYNb+SsoM1miLWKeMlkn9TizNlAs4BOBks9ZUdFE
4MqBmb1Nz2T+WJFdKQLh70KzKOtG9Z8KIqtk58pL70DF5B83wbRxhzrccjXRDh6GWcROkKWJz6Ju
/xgwQxXnJleDXdaeJiVgy0AV/eEFiTr64+IaGkxAkmw+2Sp9mOKytYCeHGAhVyuc2K02wYLvRmAg
p4DhGJVE2Yec6eBAokDOvvMB4UOutepUDWSY9KY1GZgJJYczkRVoFc6upg7DzAa18GK9vBRasYAE
fKA7OVM0OzrjmsHaEdAG8AMf7CJ9gVwYXMxRj4sTanAOoxZU1cthN0MkeOZOq60Wmw9Jcaibst4s
XWrJoJdxZ2/hGssjnvaSqjAWPWs0p84X9NlEnOcF8sSuAwuA2UEF8JL15wO/Z3QK0TUemIJ4d0QC
IHEYn3pGXDX6z5DWAyv72aPss72OTUyxNfXFhIhDW4nmGpS9M3NNs1MX5TJjsTVEtuCoRc+P//mt
nuPOvpMXEH1WZ/Xg3zJcz6xjE0FewzsK6YZpacADm2C1N+VpmydAADZOjM5Obrg5cu8GkjItW8x7
dhlY2070aAE0wUAleKMzf5JhJdcZzvTNf4IQ4NC2jCJpGMinZ/kjOmqyLzGmsTSzhcb+/r+yC8pD
V/JZ452RY3B9GsU4wskKT5xuRNLMy8D6SdKGOYigvVMTssMaOmz/LJaw99dZX3lvh5RRoF2L2cbE
NK5dTWRoxAZHCYrCWGv0oprfTL16LTgFmwnqImwLu6leFBntWi3j4OG++JLt8kIwiArIYpzTV/o/
hFrri62z+XMUG023oE5uxo/RRPFdNQ/cRCvXmMiy9xhXBQFqz/QWDwXTB62aIB3K/vms0+7Yfg81
1jjjawNi0m/qdVEz51LGjwdI2uGe5inZJvewITs2xQSLFyQThEa/WbymxcJVeeJI1L9IB0CPNil1
qRBDNDswtrkqcmkxsYb/gVOcqinxUw4jF8d1Nc1iub13NbCHMcPdmdfaVQeHwEGYmCmprgmh/rfB
8yXqICBzbchk/VcpMB+siFHGFRi7HgvhS69SbzmuL27MY/Bnn8TrVRJC7p2Ha9+kK/lU6V8w6rMX
dE/fb7i/QX37KRB9ydItfttjeys66PaSTexV/9d+ln7YM8JTv5/8hCopb6r27oX6tdsXz2niOJbj
JCS0FUcdM5SZMuLAWpT23+18S+Nqfd/pP0LRizTk7hyB118k/z2AEY2No1Y+/JPiQ3egi30GJokv
iwulPpYg68EKnh4FefAoPe6+6192IQjSlhZvbnZ3Yz0csPI1nieSDVVkyPUe+O8faop3AXpvfE8i
kKNxGbaq3EfOB+nC9C1/4fzHGXrowk3WuczhghjmqXVPk9HMjroVcFBI49nzHasFXm0cF4zKVPNs
HhvrrnxVqweph9IlTVlq8woD6dXB1doJzaJNVsBZ746gXiKvr7mRcGYhHhDm+JUlXLLCyxfi99NW
0HDhQdNKzV8kpwpP8FPOZAs2uLCU3WUJyJ6NVSUe6LtsP9xvoVJv2e4/occRlCdPyX+8EW9xZnir
ls4Z0zssTraTUqjFuYcK1R5l9kDVe3+P/7Cg5tHWxUrebRxf6Evy0Lj/u7qppTuOF91FHQqi57g1
andA8l4OZC53dKKRRg1cP++zsu0oxOS8MEoMQYUuRUgv76VlylmfCyDssTD2CpE3qKy37Oc0iyTH
5zCu0jpqtcLKnb8nju+lf4qqieidNuHgxJVmiFr2UGCQ1ShPl3qlSL0bVL5+UxjJl8adP895tTIA
IPwtCdIju4l/XFaTkKUwAlZJZ62InIAeTMsSBc6o513MO3FJfw5Vd0hwfgdG8B9Gi92j5liurNFj
pB+gCHXz9iixQXUbQnMm7828YbVU69oW4d36HAUg2UT12aZU8JE1sCDVVC3u8VQ5ySQxujm2gt4s
IPUbVqS8CdNBrGfif3MK40S3HJABfAGRVe21uhP4jQxfZ3z0k2hm8oH76sT8yHsLxhLCReXa0ttn
lGAHiyCHlQPt2A5P4p/glcO3ni+WuxF73syArTUBk9hsPcYEI+MJqeBbSI1+igesM0EEUPyM8zgU
vh206OgvJCV0JMw7MM+4tjXX5zsCpnLne+xxAsTeykoYu8Bd/q6rPgtigWO0UvEnMtrDyxo7egJD
fwzPhkPKT7QHXK4h1yYfbRuxgr4JpgoTbsbwLt49GQVqluPF3d/x15fjS0BsHLC1WOi9LpOinGkN
MPTSo7HZ49vNIohVuTCy9rYgYc4gv94j/geyB8pLgpFasm5HBFj0h2wk4PrFlEB2zyBamRcMagBP
wSZWG0auCbJYwusBHMUvJfPLguVvuLq72QdFTiW2zWZ6HZnrZemQ8pT3qUmGG6s+f7CBkDuJTspv
QmeL92tDPqyQfjiRCwl89VzTcU63c6hn1I1d7EwFG6X2eFASl99XQ8zbJgsGPplq5gUp9ULzI1I9
dOlCYDmVWAKsFrTgHtXGETRacZd1CVlS7rupCpnkfU13HKCJtMTV++9wD9HUkd6tAD/EWxwz+x3n
/CxWDDb5oFNkOjGLx7F0s8RMJgQ0QsuiKoBSeqrrCDl4W7GkNVeZbCJb8cCsy0gvU+T/dSBzRvFO
ibKd4scTiGzWfe1FBA9PSiis2yARjN6OCK/DVJIwAdwXpVi7nBjOCrVvvhaBGVNhDhLusKhGoVQE
XQNhfIR9l5BXr9tyKYrk262qo3693x2uHmSHrMIVzVL7FcQTwddUCWQWtdRFTIWFSPg/j5nBkrM5
LEgyGt4SoARgVSEwrwPR3W4bKbCp/mzrnItBaOITQcq93PePhdwzvfj+uq9AnkgCcc3Q3qb3sfKH
bs8ophgLar99Z1pn6D4/mwL9k8dMM5j/bK/AB1JXdc/6gNKs5ZXnrHSSGSJWmygrmSM2ezOsoFMQ
mbN4Kg3VPjSylRs9WQBrLbf0I7nt2f60H4EiX8AhuDWxkEV1iDx2tTTg5V+9GL7/3IA6Zl495Uvq
ZF7KmUanBCFs8WJXJ3e+4Az6jKNIGXNEUfGuEPXtJ/tyi79wGasjaxC7bvnhE3x1QIlwoO9761g/
3cYXEUze8PR/ZKfQ47L7NHJCcEb+4Da4c3J3qazwJnXXM3fmzD/eUBRM22Cl8r+sxbsNraD5MIHF
BQJOpyGy242XDqHhochr0oAMDXvr/wVh1NI3Mg/0XUgcY8qRdQuhZH3lHVEBAia7RvIeJWAKsBWz
7Se2YSUeHllvK7Ajmvptp6gn3lVrDe3St23IdM6vK5iT3zxaUfJmftGFboKCJDktlErC1xwWBaGH
3iAWK8XBePTmelvxPu8RK7N1RRBkZ2XeUembE0uQYmOzwrDowEtVw8Xso6adNOQG2geRfIXkggYJ
iHrP/AELtNZYT7yVEPtSQkf0mYrUSH/Zy4WvKt27dW+S5DTRJBxUObisMfHUKVZWxgvWcYD7vrvz
NGBXfoZ+C8eyGczamgGBRT68S2o8PIWEMJHNzctQkAAYjXSq5QTgk7iIBTm2cniqV9oM7AcCeYs7
KDY9nncnaQo1RWE1WxiJbZsjUMLFbfCfzmGRmr1uyWR1rs0LjJhKhIPueM6UaIXHu2+OzriKMIRN
WeFhLcCIj+/jn8MPjVDSRbON5xNksyWMxR1DSZ4qsc+UWeI7D7ZCHue4AjTqIXJO9Vix1QrpGHFO
Ov2lgt+urxdJthT1ln+PyUH+XuZh4zeO0y+KTZ+4MyKfmCc9lbvBra2SZJR/Rs+jHRXy3mvTD/5+
QYE5oAF69uDJi1t86nslW/HERgSmbiAn3HqUUGJJZxoMxTTm2eMKnmZjRgIPmZl18nklosUcJo3c
m6BCFbXui9K//K7j8G7YJC72D2JIOynUxODDSyTwucY0PKXn1MVbm/HeZaMAe6I4DZfEkds6472I
Hl0dCHR+BS2r7NmHoo+z6KqGhz7nHSwWL2GoE24g35N8OsS1Nwbe2YIIZ+ou1J+Om7gHDk70VVtA
oyM+sOxR7AJAF+cRO1gJJ3VmzZLV76j7OqjixcyVs/GXdc2ic+08QNl+kwvTeeiPXTJ4kIZVyiOp
u3MweyMuT3XQp4eqiYdfFwn/q8YgG1OUwAqqexFtTTYS85LjTuMWuZmm6sXAXG+p9BZvh1r96DBK
bb1Z5r2iVVQFD1hPEvB7cjbUXkpNHQyITnMzLiSz9fSE8IHrpaAmLXURTONtgby31bxL8v0dZ1TA
Tfgm95KLimHWyGpaA/hrh4ZXpfsTj763/3B5ekYDLR4UP/gfHR7f9bmhabJ+2plKYACDIUouGHc2
5plOTcQvJWfAlgo4m+Q5ZQVcE4DFjp3Uavk3zYsc/xUoBZhXsugBqX0gUB7x50oFj8tZ2Gjt9Y9f
Sjwz0SnppH17a3DNC6DQUtEzi0mgbWAuZB6z2anzwjk90fb1EfStI4djSVUcLK8xIbl0wJrLYrG8
Rl5IneYlhjm3AF/o0DwgOYBTiubeogVtvSTF9ZTjXuQ8hb095PfkaRg2bE8nZf7+j86B3gALTeIG
zOehNKIb9nMye4D5CouyJs22H86z+ITrK/YgJdd9oFRu3nEJ9LlrXLl/JLJEZuq0yusd1eZ15ra+
WDx99/SB4kSQ+rHP7KL0B7ApW+Ef+jSq6X6tg/JQQiznStt5R2dTOHLP8zV9V4UY4ugAIKuGvy2W
kORrxW9nt04QJLZnTXuv+1Np/Z5wgmFYrfjCGK9wAey4ezZRJiOaKi7zMPAbcI3EXS4LLDiEvMJS
jjo/OkZarIphJstI7QQ/A7Yh3BGCjYrYxKNRiaxNzAzn0nx8/wt75asJIj1yd7+EaQ4sT0qDSnL/
Kj7sn1AYFFeGW45n6ZHVAkaiNpeen35e/bwEHhed48JnZSfLFTklI+wNtnnj6eeXGCZVWErVgL29
8arsWcy0MmYj19cXfTkcTw6rDjnGBQIzAD6M9Gjg4v7BLwMXNfUjKAvcDbnm2ip3yjtQm07iHfAV
5ZnNgKIciW6DpYd6s/5DEM8DvGz8/y+NIH5R1SQ3hg2RPm0ZCmwUZVnDsEXkCQ0axdMYwSBaqOHk
Zfgui/zMAPQmh6R+jlvMIEWQsXAjoyRoRicHa34bOR0WjWnB/SdIkEi4DbJJcwoSkSw0RLVi6aIM
FNWHD6woAA3FeVUg9TumnfY63W8tjcxS6dG7UnE7J0u0/m9PXUwvzE8eOdHD4y4BnUGUc6CWJC+O
cRuBW7akkflzRLVI9Yy4JpzAJp1QUwEQtVmTCEFLATvGeDDcKJKab68UDROm16lGwSj9f64v3EW5
Cp8c5Bdt42VX+Fm5KdMuUvyZpj+T+cQCly3fKcnEfcr+e9TFrthWngA0xLjGEqqtVVg5TvJ3q7Xb
/E9zD+p7bGwRTqimFpbvXe0VWCWjO0iE7B9XP9l3MMuv0ekw/3i9mEr6iuL3nIr22qLDxX9eJIOp
TqbfFlk1I9VbUi5P4J1FUXuM8b6PiLqZDUfLtatcSik9QfltTPvagt8XMuW9N6bYS4v06ULykH4s
q/O9sYBo6kXUj8YDI82WJKxkYIodiKfWCn82eBRliHWrVd4ufu99tSufmkmfUalAiLa+zpLw1Ru1
FSVShVbodMK4aBheJkcrBe/OuXoGOJDhrsAXlbaFunRq8AdQ2O3QdGTYMGu7+tTaJ5BCM+7Dro+5
a9i4R5vd9Www0vVY6rpTJiJnp/mGdmA0ZVFr/6eU+ijAQ7lSgNXgs79TEmT0lH2Q31d+Uugrj7CE
k4ZIn0OFqWQH5SuT91Hl2rTi6/glcrLb2HDT/6NyIaxA4CmEnqnvmQClPj1w3bEfBGeFijgoNPrp
TxAQT1OVNkj+Xb9Ihrcj/jnC9IJdgGdXG37o/cC0ijT1EyJSdkoQselh0DpjLGY9aDsx/8igaMjb
o069+i0kRIRMZJ0mayevehETsPHPRxMFbt/uIsVZucHZxqa1yUAHLGjBul8Z7N19J/z6aWc4Bic0
WN7WFK4C8aOjTdJKivr00jgbhpye4Yxg0MBOvU5TwW0MN3jn8bH6zSzQWDq4xgwCYQ5pe/bhCxWZ
YbXJWn4Zqiji8YdFV8k5AvKILous6nKIO9YXzjjsjZ065uQP+eLbgJ11IJsZTCVsCPXU5aL1gEVd
vjyB8yNUaFr6H04zA8IW4BxetNJICkgHw1WDAasH6azYFMujgFjHu6Pq1HnZGbypbB+n1otlqJPg
IaL2qVfR37sEx+YUtTmpXGmGoYLUC7bSNgR6m7GGP/yNSsITKaciBoc61oERsZGfAoIhBaCfDYJ2
/4aEnu7QpFCn4Ja0VtvT+QfBr5rW0FuB7JnzDNDiNx1MCXE7WDOqJZ4d+BaRDkNPmiAPPpan6TLY
9XTkUmnSqTKaW3IuEXrtOlWk+6DmybkAiCD8P9s6PPuf4Xb1MbIg/fc4JparwISVrr9kQsFBTHND
7qbyKGW3xnMkw3ZRy01FsbIQuFUfdlfDlVocmxeh3WDaA7hnpMot8nU60AX6x8g4AqaT+t2kVlMe
oi+Ca8gViafoF5dzzrdAml8rQmf8wZRxzsUFkm8HEOQ/bCY3tw+sFUwZh7XTN90h2uu5CoryV/4N
ovNiJHG768U+MSTLISzIoM8z8TF2neFl9cyooXIa91F/X+KlEcymEq/Qqq8+/oJEfUv3TI89QGtj
yZbA7KrKFxpRHyCSQ318P/ZVW9QDyu4gZMLHhZ3HhWELAmbiXPxU2JizoZv6hjX4ZK2TntIKoRjR
RZ4uRbI5Vqw7fbfX+4fJ7pcWLqMS4yuXhDJeGVOQrn7R7XsTYSNNNA2chLs9p9bv6bRuiVC5vvho
xCOfFKfZX0w945256sPT3DlXXKvOY9GEqm3bYkYylmuZ2WaeSJVC6wId6RWE7qly24z12Ugi1+Zq
diUZjKelPai7MS6yCiciEYFel62AJ1cUC6NXW1dsFRWJei28OBigAxzLRoBWOqvZOVnJI6hBQv2F
iyRUTVYyJmjxpgHZLN3ngIKGV1LwC+cOatHn24TdS2etb5r571gp0C2xhgC1kzdpvWUdlTFgtOxE
skHjdwO4Xau6SScxdg8VxodpfhJpYqSeBlyzrsKJRauTZb0U/VSq/8hvFuAmj+oKd+666ZM93Alr
VuhmzFfDKQXSQkZWnuSUFEWukjreqbdiZy1Mn3zVk2QPLVcUJwh6t3phx3y7SEFfZVu7Gmuw0iK2
7pJoEse2eg4ID3PwmuJ5aNzLNfBb7h2xdMnWUTab3SpN+H+3UQDIUAXvsBE/M1+ZFKzkkoywVUY1
HDXpnqTC80IQuBy6pXDFoRX1qz5eVxQ6Zm42vGiMrUccM0PqSNa1jzgqzRquSsOvtUgc2tb9Ld+F
lu4cBsZbixWnGNN8yC9PrapoeLcRwj705F3mQGDDt4dATqJ8rCXeIMIzZZ2Apd4WNcHFiwPaQ5Sx
NvY7ow0huFgZwuyk/nl2880YVg69/yidU2dFcR1q8sVmpU3JRZ98RMNO9edJj+ph7GbMNVBmq9d2
KYmuy9DoxNlO/Udkb/9KwKK5k/KZ6eolapLcy9nlW4aRCpRKeLcXMVHHMEvwHtFkhCgwu1mHCAaV
c4PwqBPOf7e6oQlLLAVbtuKwu4qws2o9k4Eg68cayeKgXK5+MPTNP3ei7hpwAguRB/YZHlSYkhy7
c933gV0hDAtKrNqqXUE7shPToq4fPbrlaGO4RBMVEyarft14wVqrany2jBmjG3fmYUQrteaEIwEv
LHIPcpGn8u/iuYUZn5wiHubCs6LMTZ/gDTZgmgE8bGY2mvCXGXxeh2OWK0RDSi/huePDdKCgHNFO
JeLx7n04D1VJ2Pjl+nCEJTn9ros6Lpkf+3FAKj95wqlmiEZw4MgMwYvIm8qkPt2gbUYG8WLLBs+J
roPLRJE7zpODNEkTze/3NLiSrLH8WltO1WxhtmMF0R9KrHpo+QAEO5v/9afy6/kXU89yoiMLleKt
plDuVe8nAVmPrjoWB1YCDxMzmL+pCNKdxvIYEI9KUoywUbcEneFXznAAa5UNfErJHGB+UqXYxQib
btv5fQ9k7KfNUt05kdG8BdJooApaCBmNyuDKETlkfczUr1rXPj86inxLuhuDyiT+5oCxH+ZxzHu2
nX6E4/cvZr6KuGofmi/ONoCBskyCR5xM7vuq1iYADq7VZAezSWf+pUxTL/J2UHAShte6DqKw+dDl
o5IG6C6W2O5u9QJYK3Z30wxrRmQExSGlpVxwxdAGip3vRxZwbr5cTZNmNJxOQ+3z060t1ELV0/9Y
TqJ8B6WY9NuYCbxnZXbSNsk9TzJ+vYBPv1KvAOLcAyWwRG8/28C2FBJ1/JWzBXWVyJK9AAmPRAH3
ts0F9fXYRaO7oapfsyBS+tzhLtxTtelY/pMufs9w+P4Rt6nDMCFVzgjkBkqlFRdCFI/zhc5hexIJ
vPoi30rsiMcac8UkX8nJfUAjQWFKwBWIgMuw0iiKdCTMw5pFXIVleh8yraDdjWDqq3p9LpMdiTP8
3xML7zaT/fgziZBVOu0E1lbqcTnse6pYN36t3ADc7y8JPQ8KWw4KkiSX4HpXFbMymUBu6kHUwSIw
Ns6mRrHjOtunqWzHa5v5jhAssxdwah00F1aGXBaiAH03FdXiGZ17J7CXPsL0s+DrHCowDh70Qw6S
wug9Jeno7rvaLd8+vN5I0HKsSzkUwfxv5WnCk6x7AWX9C4xn1IrVcW0oJeP+heojNzcKLhhpugPi
NL9LcVY0gpjzpAWG3o6rbmWEg9wOYM2lnNXy66qyK51JW2zEolsd6AMZEhzrFqI8skT4qzAhK5kE
SuM5Pz3r7DRdFkqs8BAYUyp6f5+sGRze1yM1VI9XRtj2j+2gnTNo2wmPw8ocGFC48tbvEBfi+2F+
Szf4ebIS8r2Es+pmm5WrZzDecZXu8OteX1KuLSMnG8hFAYD0itTnwYBZ49Mh0XdQc5ngX97crlsb
uImZYbLw3ewjjQ7aTCRje1LD5i7xpviWAluqDIzrucjiQVgLpzQm+kmIDJSATq40jeYTma5Mh5sm
957Za+3ee19OydViX8Gp3idwfcN5ui/cufl4nJJXsFq9DwipMAhrDSDMESNPBYb5NCpc56S5rTgM
A7CnOqk7VcT3h/srNxSFkkRzjL/vp01vx25aKROKWk65r//eVxx6c4m62amgehBBqMmugsZGa0C9
facQyzi6QCDmCMXfvWqQ2gbVFUqhQ50lpzLVz1cXmxaAbqqBn2pFE02xT/JrxhQF9tBgplSP6Is0
IIOrWxkdDwl9JX9QBH79BJVIscpmcG1TGN4MgWUTCncKex3IDJGNGWBEpYFQDgwcZkD0fe90YoDV
LtaMC9Z9fx26uZ8Lo7ylvpIPoVuR+Nr8lmiU2/9NUmJ1QDfQ44Q38ARv/X0NrlxkZhk+iyjzWYId
y4Q5EOq164DJv8uQxdh3NEiZJmjhe5DrfX0zxpc3wKkRsZLrOJBORnEy1y5qhIF7horfK0waPdfo
fesGj8WAEELFtQ2BzhqkD+Tf5QkvMvnnY2iOLs/wXgDZb78YWhMpmUFYVMcQeQbjBKQk7AEdSuwv
VIgUfbqPlkKb1bK4Rvx4wNGqznRlwbayqxPH2NP7/fB4ZYQMM8ev2pTTEUwvbqxoCB2wHWJbgwkA
AGM7hHZx2B0WcscdByFTRz4cADW0kJLFi4R75Gxm5zjto+aQXPET2cIemFAjUy/gxi//yzqtVL6p
Wc4uj+yrChHp8Gs1lDwg0AE5+U7BbLkAyZXBMxihlH3cjoMNGY4JYk5hM3d0Yvb9pRnIaYpSSr7V
rwveUQa8k5WM0Il8dpKuAhyBOaL+ySMcf0y8lAQyX2gmkVDQp302i2DRs2QJpxanqbSOlqPoK/2W
OXgeSfiW3PgoGjgUYGaoHhF8tHynFuIhePqUxb3xW2FbZqD0J7uNpfqy2hHyfE5m/ruvZX2zYEk4
1h9uGkHP23XQtH3aed5yc8McofPVBXOsnSyzGOC2VOZLLL0kPor9ls7W0xZieLITBi5KXOlGAfjQ
XxLND/MIwMGMsa8sDQVmuZoNxFc+R1oAepM++kufRXZKrZaeqDZ2I9rZo5qD9l23BEHTYOrQ7rqU
bKCHJDenxkjrzg2M0IVkMVqn7kbCiUxWNpeDOvzEh9YHz1hpsFsPJNbkwmOhdvdUB1uAs3+Ql2bD
jg1K+3mlmr/ibg3v6sEWPt6kj61H0wQJsYWcn1VxtW+drUAnRW1+jlzZSJ98FJO9DaQrFJ0EZdVp
TdnaiAl9kF0ALX8VAmKMBegKgdUjXbZDTq+JPMnFMrVRVQ6bGqJUXZwe5gKy0naboHKLWl9QtOR7
LAviDbkuS9b+7mB5IBS7JJefbJyrDbdvxoqYCkjm1wNZqfQ5AQTZoOg1iHTFKZstgHsRnaPOkkiq
nNxgC0DQqYDsqG8LIMJJQ2bav+BeuAFZDZbJC7T8ChI4n9TGQ0L+QU5pZro1XzWameZcpVl93T9K
Z9/l1uzxeumfoDffvhYF8W8t3QxLi9ErnNXUghei9HxPHjxiI2BSi1ZQ+qH+RoY4h8U6S08xZjZy
THz26iXTupi/xRbQ/z5F7OkYctR2nn5u+b2zmms1Wsi3upD42OLTo4YpHrCqvdU4rklzTki5JJ2g
r53CB7lLos8s6DFzuuVFnS3I3sO/SdXNaiyK5PXmKimYIeeUtPvlEBz4WaZlmIfRP0BblKdxGBou
PirqkyaBB6moZdoMSBgyKipFHeeXyP02iesTlNfWMLw0eACmwsV9slYvrp8Ulq1sqHo5QrEDhHiB
ETjaWuJdCxSPAH8YvYt8PihOoQt8TMGAEGAK9jOGryMoqVUlkUT0REqqX3aKm4Cej7FS1dyIwddv
3BuO7zl4vXANvUAjr56bvqxo1iPbETaNCz54oNqoQY6mwYBSgUQxtcU7B1Z1CRZwfUQx/ZrxStc9
aSPvRC1invvV40AWeb2adi5VPfTKf0nErD/IcBPbs+0PEOhhqj816k7Agcr/uQ0/aTJaX/lUoRDg
RooXMEiH4AO+czh1bc/0R0ozwktft7c1WOIGzM1Z1sLFw+dqcZXWHKNP8gTAl6KCMa7A9p/j5Uo2
IL63bNAx4bwc9uaOwLUZQlgJCpZo9spD0zUjnRQ8Vz60z6jO1aZhL4ZSvSLh730AzrzfgTWKXc0p
VF1ufVwqm18u7PT6kYGEZG0WAnZbenKtsnPZLnGDJo4mDzA26mIOTdI6x6zz0GJnMN1hIbIZYX0M
GsurrKGSxvOmf8q00/JBc21pk59vMt5YfX19nrPUKSSfr81lGzLFqhvKx9sNz9c4T6gdguaZettZ
WJBh9BtIWQvdeMcA1MLaIgUa0EPy1jHH5RQbeCTsmHhuYHhD7fCtnl8uq5YVUjqM0V2W73hPv7Iz
o4NhY+hF+TJ9unM/Uykog9kuz4zRVyx2lOeHGICNg6wj8VvD10Rf8iswN+EZUia92Q3ZOqgbJe5i
fxIr7exkINI/GYixvLTPT3PeCkwraHLPUDRvKIJQffVyyoup1h7+d2vTEEbTouMppJ6s+nezKkgL
RZYocWWGT0Fo5tgmCckfG5Jh+bgufqOw/CEVyfrpbN54NGB8pXj8M5fvIobdtkzkbyo19uDVStrr
onUJuCGkfGkebPOvZI6WC2SyzlK6rAvezKUb8l4N00d4XLxZFouimXCGTyynbVRtBSekRVjzeWps
GCgudHo5TpF+H+Nuc4WNJeoHG4lT73EImMoI0p8JHqC2X2NAW9UgEdCK5XzORK1C55KavEOrhmd+
L/CrcFAGG1aGZ+lRNNiNO2qm00c/5KK3AUwqBXjFUgjvtUsRgM2IPDj1RSTupWRpCQmStYqQIDUj
tBmViTppIhZ4sAFxQa7ciqssRBKjJQhN72749BuLz/vejEBYci9Ppwhujul8WgN7wRCp/dy70RA/
5dryv6/zPTYfQIb8bH+yThfD/9wbeXT2miX9uzoYpCNGeWvD3fBSEcwqB6J4CmqzjHGDcKFqMvzd
4Wq+rNzyPvwXu4hOcgDnVpoDNt927mR7+99cq9hH1DaKhKgK40IoEMzpgrkUSSwaL3vQrFQVPmkE
gDrcPfcOL7/xjheg+Z7Yzh62NS5SquBDWY5JoH2xQFbpGpuPyxJcQ1lEV6TlC/DKvmIW6RZEFgxj
C2HsQAdpnHL+VJFpJ2wCPGi3gqaGmdhj4FxZTnXoHsiRV6HOI2sfQO9gfTaIPYrU3kh3ltzMmzBc
3VefXcXbfLpKpZMHrcK3TCyygf43BAgLmUndbyVXxs49B3Pguqo5G7lVmSQZ+lMZLS/CktnAoKc0
M/VnLXYhNGcSlzzObdYivGqM6sWEj9gR3O0OuRs/aOmwxdY48AtGN6VssD0m3UkKNInVdVdw6WCm
YlsEowcSQfhIGvGhxGrG1l9YPDvgZxI6Uu6WHCdPTOAYkNMm/ynhwptbcAJR4o5aylAQCnb0oUda
woAkdqu7CldloYxzAxLcdjIGZRhDfqi6FTZ1vA5Jz3keqTVPc+pNdnRtMzfVST7bAaA0cpn8fBJP
gD6n06MLxSdaHyUMcENHJvOt3Lrurq+JfTW5wiOhcBcM7On3HrdRFOVFflTAAcnTTcsvSNjFEPmh
HOf5PVHV49f56w//7xo1n2kZ7nWGwGw0AfepLFzYHE7yuOtLM3ZO6wsQ1WdM0JmS5Wa/kq3tkKDr
qfq9Wm+gX9CUL3s0oWWNhUWkmgE7+j+gy6Ix2xGgMKy0SToRGEltEELe5Eg2x3VTif+R0cKJyv8r
4Zpq914HXT72YaCkw5Mz/WfoYNIF/hun83PvpyB8PZqCvePkr6j9rS8SY+e0aqNJ24eY0vd+zP/L
ecfqNzmBbHvmN9RGSARjX7jaD3UPqlh4nOrg0YGz1jje3iVcQZzk8Jh4p9trwmpjI7tASQ+lTCH5
ulG75eUxYWRIvJrrh1g2c+AMvmuOgXoYKJ/0mP4ByTR7EQN2AEOcQX53wdToXviiF4KKxXze0kTi
q8YhOudFrRRsbQHMT4UWdy+fXta18OIunprs33aT4f8yawjSvS+cvppAM7NOK+OkN9qyt+eG4tdh
KMr4MdVrrv5+VeR2ltHPzuzLDRf3bUALYRWzTxT6nz4847Q11g/5jdwGUCbBSQIxmWkVzjDl/vaY
cX72+PfV9WIP5lEF9kzFYpIN148hFQY+AJpg4ve+L52BiVLLrmw0qMkxRpgcgiXnUlhAvL8EbRyD
E5r3bIN6TKABdAHCj11Yb8dYOJwNe/j4OtTyRf5xEBiWzlo7ZJ+ey7mMUtcaG2HsbHO5D9ZNmLkb
hxfu3zFef+ET4bWC1J+8vME4UQyXL5fZf/BnmD3wZxJ2PPZu+42OHiaTRwDkwPQjqms7XxDxY3D8
Gdnk7CheSdVhqoADA+uAAm0Fbh0SGWM3B7uT384sS+nU1n+aj749Rij2rndpH6p1EQjPL2KfTPg5
paVx8tvBuwcUs+m8OiOcTEvM0JxsbXr1R+pz5mKDkRAgzR0Ybo4OiS2ZOfz136za5ao54YeaRkn/
w2jmUM0lX/KiyaqXE4tbmPGzJQXwt8MHkBkNFoC0Nhg/Q5VhVx3wQWJahgUMA4TJDe1m9oqYqqHJ
XVUqCE7PQB1dad5OqR4iBapt7NBTzDxsYXIhNtBMgsIw9wzZplM5rxgGxytfImkM4WLytii4liZ2
cExUFcJC3kTBZ8QHVfGqZkaBKqGmXAAkcYahoJ4qbNNxYbhRpYoJHz527G2EvNdPiUNfsqe2AQxz
7os81QRO7ft3BDnwL6ienNTybQxZk//A5dTfScCUchW9/MQLw+wSO3IjLE9hLi1eQs2o6LzjV/oc
OW6wSAiJxWv8OjAeC9L/PgsbubWTaXWxXvodZgM4Rqwqs6G/mVFotVmLQE7oLiD0ccHvwuTT/k1q
QLkUj8K0xo+2H2JH6Jzsos/cIFJByrfse/C9Np8C6pQjgELIU5+iNtSkgYMHcYrtIlygtua51f4w
K17QbsaygHTAx6i5wGWUmpmtB5x/j0Dnem4rV4vTweixmR88Tl5tfx4ojb1xwbNUeLLj66/ByzmQ
Moph3i3yO5UQI5PllOk+27Fqx0pt3jtZ/1xFwTcygJ5ns51PX3rhyi5Ii63b8hMtGsGs/K2kdx8T
uAzoyfruETDzWLUEh3uvatoCspXbcpHeSTVCmKTd3LWYkfYQpQ4uPh5qgQ2YOjrMs+cMoJz8IrVc
/XJRhKgZF4mXMc3h9ka+ONNnVP25hWd7Xgzedf9q6WAwwpK6uyvdrLQMT5nPz+tbDXm/out+Yhp0
ntpbF6G3You4JIrWsC/czMPcd5ltdG3TPn4GWdDW9JWeu4Oryl7kxVtCEocd/TCWVVKljVs1n8hF
GvbYf+W+T05A67WWenvEgMGQZmO4d/4/OHaFj81At4lIf5Ey27MieZjxML9KZP7oKceNxGEDyrZl
BW1A3jdqehdWAVe5eWLIbbDPABa+tX3g+CsxLW1vJ+Wmf+3vUgb2A9ICCYZTnoXuc//hoe8yPPJ2
pd0mYeJbFxpSlTz4t45AoNST9G9BaDG3zW0eWpjl0icJIGSUhj16LETovIwLHV1fgVoLIFooaE2O
bSuNp3XIuOGXsIdjn7lkcTJqkEuH71qZgWw5wUFBBcUorJYpVizSCOhKnDFiCq2cUOXzQEmkbSNu
MpcU9od0HHDiC1fi3559a8wIPXa7hRR11coTDCSGZn2UrlwC28pC5Q/tsrlyiDdB+bdr5uKZhbQl
t/6exZgqE1x0JXdxFTvlMuK9dVHkAiuvMM2jAl1ZrsNCPvSpFp5FN7dVuwyiFJpPypKMmpXs5lap
JT6lNyf5q8qesjwKRX1VjIuD1wlikf0ipz2c0MuoqHtFsHb4qB7zbE5AsivMVcuqEeCpOo9mZvv2
WgerLjUNKsj/gvnpbZU/24dLOMdo3ICksY5OqaXdnr9DBasae/UQ6+T243NBj17aJ0Gk/3nDwps3
hL2otXt4k8t8cMtb4TZki0Rs5Qy0vt8KuJ4bV06VVg+WFCOgNuRIJpOuHcL82xu9V1hgWxe7KGDL
f1PfyrGZJPRb4PVGtKNRFabvCypTJU0cALN3r91+lDO2FxTbZKgTHlpUFemV85FZkVpi1XLvON+1
mEHr/keAHiFk9QacQCYM7bvYU14rC9p6DtIZKg4vTQXa2MbenMoEDRXyeBf2caZ0bH16GX1aIVbO
pFkm8IlntuLjc9SW/wOITooCtT5I0N5KMNNUzYfVQ28MTrdY5xjsAR/shy+wW2LmStD8yIsYIJxR
iwhvsMcOLcFaPvKDdKQnt/P3kMETuDkDv0kGFwrSmGaTz7+7b67DuFfV/by8MfU/VTIbt7sg0OWn
PUh+0IrmIlPGI1limd7hqROCSWtu7LEnPx3CN3s0sWj1mh6z6n5OX2lVYJa35nCxOngwEgd0AGaf
n79c3kLNilQM97/wJRN9Fbt4PT9Q6RbPgw5q5oghyTfvJ9z/2taidFacEGEl2VbBukp7pefAS0DS
g/uNl8jib/tRrIz0t9YoiuIIVe0AwolgFLxbdFRyHhXCtPEzQyU0H6bphj877f5CSX5fuIek34Di
1NTGLJXg12Adhz3eIFOCjT2l3+HI23+wtth4jhdtcMBrg/fA3nzIKkAsukejxVdeXnNJsJYM2wYL
lCzy2k6Y3vO1TxWMyRRz/IFRx8/aHOVXm0VbIh2DSTTvMkjMpC9hbzz3kHWnoU9Pgtqu6fF19CA1
SJjd/BLiqUFwBH5kX6IhHkkV6zysUXXkMMRG8dAJIpD6VjEjnLt0YHiXkvTiH/TsccicpQKW5y6b
D7TNqbL4Wrv+B3fDCwkM52AHyT/IQP8NKyW1OIGJbvWnCxmliCXg6V1BVCXk5lQEDeVKEDXqeMvG
i7qrCJIUuW3ZV2zDixwMtZfE/ZfXal+f/F+1EwtB5b5dXKW1nOHiRpgjrMX3nszMMpA5OoMXHvVL
k/c/qiyMH/im2NljbmiYs0SVB4ltI8uk1meeS7ieSAGtK3a3sn1UNwBy1FmTQ2DwEOH1FfVjJQ5v
GUtzWGFzN9kmCtOAO2BsJ1RtQod1NsLb+5RWdF2pHp8j8aQMeTsyH+JEyp/QqL9mNl7/XjVvDf6t
TwwUfA50Jbfc+JEkkL93rbcDqm1vPfYkbaRt8uLkOT1UlH3NIXucCfIJdujhsJ2trfFNg/7BQL8M
Ao6AggtcT/SeR5sZf0jpfDs16c2Jef8CooUurWhS7v3eN3knph5k8Ta/jQ/B5FJFeGCpNqneMYPw
g3P0W5bH7otseYuPlQXWWsfmtk/1Hkcrh7lK2of7nT9u0pGnEnDTiyqeyGxwZGuOi9Wh76WImxDv
oI63ifKKoPzckdfyjqT3dRFd43Hkgy+iZ0cKLOxg6WTkEyK1sfjgJPWIn/lRhwW+8VPgGYNEJ8ee
cVU/u7LML2a0V75s8TAFwbF3RcQDULkavNzvu/sA+o9IdBmSyFyac2PkjCPiGID0axJ/IooHJiyZ
On86VRhigRIEs5MA9972y8AlmbpUOniWtrMxddZCS2JWApERCR+qc9urMRpWJH4vo+F14SYxrKmA
YWMEGtUIPJ5UewA77b49ltF6qDb2EhO9PBMsTo9BAv/CsIOdrPXdOvUmK+huoLrHIHjpL0mhbv5+
6pHJjyT7IuVof60v+g4NVBeG2VHVV8VTW2Xhp0eva8oZrdmSI7K5QSr/5BNbDuRyqjBQV7FQouB0
jst9+TImqlDOx+QPdfMu+bWEzWnbcjpuBP/LGmPR18dHO01Gs0zqDaMTm9/MnS3BzyUxxG1I+Bgf
tpjIr4CY0PUcC+HESyluZyjHMK6nX8ub30AuiZLRtkvyqv7wdEJCqoqTgc9Y2N4XWS78ZSinfOH2
908Zv6qFTLiYEaOtqE+Ykoxk/OU42TXfV3L0zSWYGeD6xZm8sdbgjHieAvGk/gYZ0Z30TT+mXD0Z
pLGYpER1rbhaxiIulXP3Il3wwG9I3Fi0FHZsIIqRyx2TFSt0Lr0DhXtir/sMwPJi1IHLm0U0Tjl4
8wMHPjzek9rrwpa8HR2uf2RPA/i4nLEUEq6AzeHjjby5zmAio2jofcv+Il0L2ZqXT6P9aTyodEGd
rbXdVd66Nm1YVYPjGwCn8hTa+CsZl85Mf60U5wX1SxegB/thJ506+XigUW4dU7CXAy9d66slgFh1
HUSutKRhkfoLgxAcGy8W6OFGUnUOlEvKJv76OJAKn2ZutfNcfT40UzDgt56Zz0AX9uEsRI9g0LZX
45ZIZcRsPjrPStboRro5LQ85An0sT5QXsklpN7l9ChiRTLL5FATXDBzlCarn/ROGDc06Zaqx4FiX
5SXXVFDZDxWlRS670uQLSg/ee3pY/SqGtm5NVtJ2ukvqgkK7IIPamL40oxIryKeDxzvXkVuM2L4k
fD0NdXD97HgkV+55qvIQGRG7AG4IaCec4AlHLbdFIkPxa2kj2kQ8aK+RJeh6b+v7tW9MadRWOs2c
PWhJ1QUEsULnsqO+S9kWGJue9dY6TzyAh15ZMGBdSNdJGDAcnNPr68ro2XQ460szwpviuZKdy2il
wTF6Skt2H0EP/EoVOXXLMV7n1VasJk4m/5myAKwxxq9KtLGxJeP9unJodyIcENvIPgOJBeF3rZuN
v+Os4GYhdnLdaTK/DS6+HBb74cgSnRZd2rj1PE7HOleT/4C9c+iiBnVaqTOi15LgrfQ6PicM46iu
9eP64GiCI7C9wlpFcM5Egph5vLepHz6ruDxN1cZnWDD/aIT/cmF9790J3YHQrNuMTvLov6nZBdyl
/BVR42omyWZslUjSlso6OrsPkKUOAMJ5tXw9Z7QuDJpPW+j2hSlULZRU9KtCNPlp0KMcgHcfanP6
fiJgpn4ZjTMXzO93ydTR4EO7V8W40RWIrEmlCy0VrC4QYQet7pg89WRVyzT8w7jgrBk6VwGHm/3F
rl0AFuPKRCkV6Dh9BQItRXw09rGXotZxki6+5nYfxwoaMq1QPDJSFLBc/eWxcXPpqwaxa5gp0LGw
1NxZOX71jeFoj9aTRCa3o7uhqFTU9mhxjESNr/abEtUfSnjIOSj9b9K1xrO1VP9Px4MGSjsTip+V
S9jfoe9Mfm3IrDVbeyxK59hHkgTfOLkfP4dXYwbBdvfj+8aiPMrLOV+BHMhVX9RSGw0TFJDmb3d7
Q8L8VgS/CDGKC3In1TMWFW4qKio3BdwdMPmhD9mr5qaNonH2q3HnpWRei7kbyUL3SAqCxXDA5jdK
OWGagZxetQv0EaTItpmMY5onW09zhBTx9FSBi0ksCmFQbxjWQS/Th6EPpn1+Kq+Xzgra6EBK4sal
wFqT3clQ4LmGMvVAT/2tpZAatIcBTg1yk18TV+AP+09nUqvHkY+qG8L500UuLHof+Zgo9tWAqDI+
8QHJAJxQkx9L6JrBuK4CXArfXjDq0v22Z7ota2B0aP0Xj/iI68h0ypkP/NOsqWiiVujxXnhfuny3
XmiFahInfRERnOvSmgBLijpgXFV3COHx6KQH9JTNrRDV77NdkxnVE7GleuOZKWJIYPYrd821uDKi
IfyVAVGQZ+hY+hXY7litYpGW8W86i3cfmMoTt8Rp7Vt1RZGHsbuSGe/2AjZJwsTVpNMAyeE9IJq3
JwhBGEwO7NFB7M3ihp1jBpEIjdmkIM+snkUBXnDzxQGys5gOPvDN8Z7qFFGXWoqmBbEe/+Sbp3Pj
bhWgtQlsIiFSZDKwzWOFWGa/KziRVZ83wRFBn6QyTCElWb0wEBzSjzbDJrncKl1zVpYXJgUcpzKF
lMt95OGFyPzKNsCmJ9ONHDcKDI5WXFUDensgxkOG+JeFTzaGadGzqnXa8ZJN+YQKFHFAI1hrFNjZ
BvkAEwrGCOdaeyyxEsBDsbKmy0Qjd/GqWiFTB7FEcEZ9/ZCph57Riv80iiVyo10hFMM+gz3aUEjZ
4OUqipP5BPIbHkhz3PVjb8TSGyz3aDmBzcSXqR9ho9tEl01hIaLnyQr6dzMmfYOWmAH35pDcV9pb
fLixwRt2tCxAa8JsHlEM7grB397urAFT24Cy+a75xtYmTSBBc89garYXmu6GFHuU7UNBOp1t/l67
kodIQSb4w+n9e+fYMczhSKp3H9rjU3AxKpFeNaMCtEKTJjBtvKWg4oNYSBPea816p6+IwTbftTlA
mN6+/apntQ8aKXa3BAwbnIaVgrCJrM+9rRTqsWdx4UOnteyHja3lZWcRvCLK5ts+o27Bhg3g8q1f
+bi0oLt0nJBv4hrRokbpCdl/y7uSAN4cZ+VarC8aoZ174nIDRgtx+0T7ZOx/P0Lxh0GckFmckwpm
ZAl9poPJE2PkOl45npeqKJyltgmXsptd1FLREg01zG6XLLmZJud2B1ETKKmu1pPpklcZZQ/UgYUr
gWJs0rjoH1RuytrH7VAuqSg+VuREj86A3JoovSx4oc4SZjAZkV4CivbBe5z9HYwikEdFUwHju+MC
PIHWS5T3TqED9OZ3TgbDE9BfyD7hAbnZSBJQ2jy3DG5LzSFKamOKt5hgewPJX5X42lbopdlL2jZf
+Zi1QKDtPNPrDpsqd+jnRqtRm+ktX+h8cooJJSAL2EseL+qStf2lAO3q6k5ohGlfCtOovxaotMLR
m/jvae4gavlTGUaytj+US4C4RgLq10NPClEwU4MwEU7WR71LCSqIKROdu5pXNSe1a/T12YR6U19E
03GjwKqE8i937Qv9WPytJ6YM9cfKIcMdoU7hFLRUyU5ZYLuHLfkeCTU9txl9jJNCX2VOAuU9+kz/
E0gAqsOi2CYlwuIV8SF0VLJJng3SPsQFkabUpNVq6aF2/GxQHmw1oS//TffbGyLqFd+xX0Y8eJPz
cp1MuuSa35FmsZmRwCpx01lBvoV9LhG9EIUNdlilkyFIq86dMiwR9GYtD0DVYsmnmX0NZKquFs74
z814xloKutovKGgHer7qqVtgov+BRQTjpzWYoyk6+xKuZMPXb3bfonemM+LaySOsiMpqeju3Xznm
Iu0PsOeFrsiHff2pzAmK9sJw6iB3X/Lai0d6lxLAF3ozPVovI7V9F/jfe+r3QbCoK0KMGfRTv8B+
U9O3VK9DynU+QkloM+yroh+IFKckU9ySGo8CA59sLQ/ypP2mMBN8AykVuP9gUTDFcePO2ruU7s8T
iaUQJO8Ju4+PVoHLSW1dgkZVTOv+8onvFd9CZeCX25PIAweXB4hP6B6FUlyna5dcG9hufs9Hul+F
RuY2Sx1C/jGrXrUBG5trxR6mff/fYuTEBgbODDfIHazD+lVPeXiMrtxvyDB4A93tAto4r8AbZsCX
tjgEwJY44SSRmrnG5SS8/Is3j8C7t4JJxwKy+qDMG0j7woQ+iQ+fY4/eu5wE3j2FJHSn9zNG54AI
iNiHqG2sk9pduhcSvs/isxo4inhyAA/tOSDhmFCf2KtVTS3ylygR1lTMZlZw6VfUjrCBz9/EN7mr
BrP0/TimkwbsAP88nU5TyYMYGF+tSAOI/QOhHji3EfFzDKibCZkNQ3kDaT3knIvEYeV/uYi9Epaq
JRjBWGuLMXavuQscP1qOBP5C0+K2a9i2nZ8COv7SiW6ochWfjcCWqG+iee0EfRmTdjryx0mUVOeJ
yz+FKSfRoLeLHENmQQA3p3tov0XQtIyttEYN/Y7ReE0c3Cs8J2MaxfTX2f5oCPHS3CKrrwPOzBc1
5Qrpl2LOx65LXborPo1Be158nRLfMhomvVW/+LfApL2OcEfQ1Fu419nK+c5GrAAkbhE+zShUpJIt
5VPxBN6qMuxkR15uPURCdDLNl+OjkjDAqJMSZ6nLLg6M3d1AtLyfFQAbsKAzhRCYc7uJ5KoS+dLw
d6/WaGfXF5ct3A0rJyW2zkWLcnHZvYzTqUhBfc6gN+3n/abqH8RSEsR+4YqgoxhsE+hahjSAFmeR
205/VDl/pXYwgyXM3aoeJg3qaw909a01GdkN3kIUe5pTIKSLBpnCwIkJ7BOdddZZUU3xZ0GF9K0P
uke4CgX5y8RT6vI9jn2k+yh+7hc8T2rvCp4vhFwxc995aaz/tfBiktI3uUp61qE26ZK/bAJ8sHVr
SVp181FgpKTIZGDci0ngkew95qImC+EDV3ggMOQC8es+o222f7AsU8tdmUK5uW1FqAxwlDfK5uJq
Kh+4mRzrT9BaXCr2vmrrFi0lA5iYxCPQNifj9Zm+FEU+UK9i4VN+neOOeadbLy/HBQkdH6MtO5O2
jBpHlpvEgjZoFi1BBQN9+Le+aBKq2s99zkH9URrqom+s6JJiTFKi+PH2L10X5ZRn0UdXr6+C1b7Y
9C9Eq/FK4imdDE21eYiHLwxjYk6NXSwHmyZMOzc5obT2/j+2fugyXDYweI/twihM68NDN13JZlip
EXVwas9O0SPfC3af4f3wZhePFhvd17F5qXzyiAobAYQJ9pFLm0RlU3wnBh7Z/SmTC4ElxAgh61QN
WqxP1U+2A1kaQ2LImKkGDoG684B4EdL5zu+9XE4mhmv2qh48cCydg9ltTFPcPQEVz2jYKd5drxiF
XxbFr8TpLn2PJGA+emFu3qbESE8yuRg+sijgp8Z4sLS+WOb2/lAMfDSJIr2hbvwTxU0zVea5GKoh
qIf3qWBRDBX/+WUyZ9YqNj81MfRBuCJnFK4b4i1v+5DQVDIgs1UoQ9nOjraiVtYW2t8X/kftaURx
wZNhA7XxXDX8CWi+2liK709pv2CZxSbP5CwIXiPG09AP33kCz6JXMsbpIPGweFq4tN64s2FEoTea
W5iWwVgkeHJqQ1Y7D86Ro8WevXGjuNHw6Nv1qEelTbvq9ZI4cmFsT5wdV3T4G5GBWIRE4wzUpdYT
fOiPJxHTd3fMfgRmNoMFvU+j9D6ccjvqeFAqF3DS3nWtNbTHbRo0e45pkwWiM+iUNNybjUTBa7ms
JuMho7MVW9h3hXlKfqUBekSPXKEJsdcIAdv+ihGuxyHRrK5fAZD827Xgx0eBpR6Kl1hUpX1JnPsV
WnqSWlgRP/8KNeZ4XmKldZz8C3vlqgoQ9S2OgjWPh2Ite46WRIq6+2HVT+AmSBdOg+UuXLd+xfDv
L5eCUDZd/7tTA6e9e9XN8ipk7M1U2lkWRND9Dzt6B3K+YQabjlNr99dG4k34MgKRIz8Rpv23IC8I
uBH1DSBN/d43Dmq6evZH/SQ+zkkpPgHlMWunv1n9oN+UZjhKpHiDlpYejEo4ugxZR2lvofTFeuff
Y831gSUGkB6vlS6Ewtp92VUR/MiAxXpFN1915BRCUa99lmWfYihDGAH7rSEfFN3XHFryykw5IZmE
RIHHK2RQqajXkc3SRLCHXkWcCI78TANNuhxoKcdzmT9nUaNBiUx+/RDFbcpm2tJOa2memP8zyZ2f
WRHxO+NYS+efvtxXwdl39yk6SK2of/Vm+n196uL5ze16UaU17fmzqnct4M8zssXm3rrq4nYH452/
83tHL0TzD448D9vmMepLXpxG6NPsHJ6rb67N9dobQ+Vzw62LfcrHAjm6BqlKFoV9uJeE6KLrjvSk
sUXfa7IQyoNR2jC6hxERQHkp7kSGTQtIjbq3CxTYtaMT7bda54S11RkdU/tGdu6aDZ4BYjZ544/r
TDXI+qRR7j+SWEkFMeViXDJYFAgjl5fYzcu76HUY8wUTYoNvPZO+LJI4deHrXcVi1p3LB9xaAqy5
c++diOvi33+foAc19wefp7Yxwc+0HtKP1ygAQO7DGYW7ZDkqHOkLD5BYNMn2v21JM61T6RABF2hj
cNeMYM8BtYZOPGg1PJ+woads/Ca0gjxIHRravkBQIxMNjjxt5xxRb4tlKM4NlRzCA2IdiCyyHlYV
sK+B9MNc29WoDchnQrxZFS4sxLvtvWtezAaoHklWIDQ6AeLHRrwwn4/c9dLjWaBi27SYu6Rj7uJJ
gbxMiaCjPyF6s1NJTw522++Wtx/ipAnn1hz9lGvXghhuGQ89jgvIUIK5ajzrY/ruhqIaBxQJIRKB
RzKUxK+N9xe9LuT/jNGR79Q5tAd7y3jYvjPuPNsLjbWMo09pjNnuWGOgisM8jRic+ct1KAv9/LTd
aECTmOY0fibAQZZdVLNwAanGCCRCE/GVI2M4IfjioNL9tGc6GtJpPeExKsNRGwzJLRRVWKN42XZu
EteXBo2KY6l1QyIqCa1Fnaa0JGtFsLucIMYk68ivBOIMU7wj8qcbWdawab48A3r6DZalo0zMlrss
wHDnysBfSwmBtSKGDKs8HkiM1VYmOIimJmgTtnHGJ66YX6sn9WFzh5bnZaoExsR8wJXnvZZCJMtL
14/OQQLzQgnitnhilD0Z8l5v+Mh4yUcMlKHoctEVcUqLGL5UP7EyG+oslXjMqD4/UzoKn5lXLeIF
hqoJmaYffekLOW0ExWKiucxutOk2R9xw5BY9uq/dY9G6N0LxUIHMBlprKOtmMqb+69ApafNaDPOx
N3kT4S4NPzlov1rcL1CQl6FD2eIcxuUvq2uqyVodr118N+hKddC/OI6LTuDFZkncbtbRY1f+GT6A
2gM/yQqnKryDXYVKJcHziS3bg1RCcQ3cydHdtC4gFp/Hfhmd3fIScOWBFiAHnzauh64Tg77BL9UV
r2vw92lrFloNONnFKnyAQK9wGJctZ5fhtggT1arcgnSybYuE/KpSiau6xewoT3/4CtUp5s/nccMY
fUE9xl1vcZp0rEAbjkeELvuxED5fQ/LnNYx0DKpyP4Z/apAL50C/wvskdNQer7h2DLWF+tXqaiGn
480mL/FWa0y2TFXHjkB893cdabWfgnsNYNodEfvvy3BGbnakQqhWK/yQZuf5RQG5Gyf7GaiOtgA9
6VX0xwH1GfKzrIUeGK6YcNX7Jw1bVNTr1ZhTdPk4qnrUys42zf/cfIDXSPumBQNbtxABxZko0NBT
N16X69VRyeZyeAJ8moF+YHHc8iAW4v/fQECX4i3+lbzowJ9+UAvRhRpvVvOAcxtcsm2yilGREu3I
BhCE+gcvrqHJGSpiCOwuDsdbRk83MEQqPjOV+80tVRwTlHX6MSUkABiB3DI8gt2h2sks209KtYc9
Lx9EyJbLIYDSrV+rS68U9w==
`protect end_protected
