-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UBlV8XHc3OwoR58CZpk2Moj215nOpBJsL/4lSc6VOvMywrumUW31RpuOqeO3TXakKCEXhS4arCbm
WT+bs8gHKCCx4PUQGB1mgsryDK2eN/TeNWnRapvI3NrVjHgcfPmXUfqLTewNyTFQyuddp7s+c8cJ
gM8zDAmN74n7cd3p9T8aVOQUFPEPQ5KP2hLgi1y0JKWRmzrJkHt5aCG9GO5Ol+yhSGkqQ+wTQvSl
YlX1mSrewTIrdhXJUkrzp9t7c+5ZS9jA/tJPSAF+C8s3AXWJsGkMmnyzbVNVX0rXaB05p0x3QfqX
+47r5QcDvv+dTQEu9Rfydp577MfvfrA6xbE2XA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
FSR3k4sN4A2yjAMhNlHdDCX9TjYTDFKQb0HyUaegdIPQbpi+ljL+yGFxIQB/6G8IxiNga4quSFRw
Q8+2mwueuC2k4bzIFxIosyyaSb/ouIjhUj49fK6KOt6P8cbFciHxbynHrevxFzkqguP0IpyG6//n
fsXGlcsXgHrLfCtzZy2xf7jpkRdX1aoUYTbKkaBdCU4PxIl75ykwGp+jYy6Lj1X9X+NgjctOjdi3
omAjl7eEA38siULxESb1i/y3RhznchNy19qzDOWh+YVL+S8R6Q1LE2Dy4r1e+7+pYgZHUyniY859
VIK58wPaiLpbUQ3kY1VHbUvTMXwwagTIVGWk9hI5THaAmM6S8Pl3L+Q4a/V5Dc/95XRzEaz2MHVw
UCMyiqSQ20VnkqSVVwgtoFEzdI/UlzWkRqa0qVO3JJuScL9Rc0sXQiC/nYlCzYqJ+chOAgjQ05JA
50ekauum5sfsF3SlaNcnnA2LgG6E6iW01PM28KNG+WjWnBT3OtiaErPBrEbNHwjY2z540ZxIdjSW
AosgpLiFsnKXU9UvTBTrsWB31JwO7KbpOyNXRzPeRvnhDgH/SHGYA7of8Mwksrvhj8uiDvrvClt7
iycr/WyaeP+O62Malt3wsKbiwfTlKffFJkSd3LE0F8YJEcNWkzaCTZlxyl4jRCPVfTTGp1+RPZNx
RJUFU4mxARp9c/f6jemdRhZOE1ECZ+M3x4GOlD0XgpxZYEv1lcI2uoE2QbNkhpfV+MAa9ObnmH6V
3MDwQ3IkjtVZ7NYaShxsHoMrgebIiwhCBMDZzV6rBn/LME78JlUF/mpGyr7+rduPbeSGcQ6TkL2H
ua/yJquztvAIzm7Dbf6rQyU78SeG7xMQOD0/ziCnFUBn1huN8EBkTNcqr78+Xulqn1QRsyUjo9JT
ikZyYOUBwUR/3yepxux39JnLKxx0GS+otSDfnW6Z3lIasrhcXuI6X7brghZ1RdOEvEv2Od/bQYEi
c61BHOc4t3LPCbdangQf+h+9d2szarFWatuao21QV6N1lImJsLyPkHPUx6M4UNcmFNBMtyywlyVP
/avwKbb61c2olV1SGdY5Xcn/OvqFpFfvvfMDdwKf7eW2aMAH+rsUTWt6fHrmlkHd1zovvvKLpKjd
5St2/yd43vBJWy5PtHUNXOPg72n48kbbUmWqUQP9/YV+5wfLQnlGeyaJDJGxMuHo1fuuKaiZs9kT
qYRlpXJ8stpqBcDxno29uS/67BX/TCMmKid7BxT7eKwyXrZCp/nhfeMMhSYe5Lmj7t3lcLE/4J2Y
uRXE1RobeD610YnzawmP1LhmKgMoGzOYH1GUTOUn8VRtGpk6vfqksmTm6PzhxKvOhWtj6yd0jDH9
lzXH6k5KSLLJwYqVn7IhFp+MoGxhpLSM96ScC37oMltE/apLTZgRBpW21Un9ESa9MZpuEaxaHMu8
qKD0V0MF18yAw7Ch6B4BwGaMfzzBNbpvwrV92L+Ii5FxLL9kWYGbaUHvkkFZkQWLOxc1CA3SmSB8
/0nnwB7GWnsmsNkr2i/+5334cf1QHWoTSWZKtHQHGf7FOSI7dVRG6on9GmP4tOdn5jzQcwdmqWx4
dKTtnqp2uAWnu+W9LxLCI4wN5hkXiK3nqbvmcp6yAD34BhCZ+5qvs9veDfQyL9a1V08Tw5fl8ANp
FIaijUbl0Q+ESE7nYa5cq2Odt8unIMlxATE2K3dM7twO6MAlrlX3EA5hgT1hF7LJDGvK6G+doDBS
fn0IkNhl4/Zds1nV5gZgmssxZWbU9TPvN275QtAtAEfQqz7MBRx7kQJYc5NIQFf6EF+2uNOEEq+e
KCleOYgbW6KJZxNedIo7cGVEEL5Z7emcbyHVyfT/MpKzD3weFbX2+Vm97KhS8CRxvE0OG2rMQB4D
o2gMmreh/3EFMOUJcZYZCwe7wmEbtEFvDnL+GGrLzAep1pOi7QjGf3AC0R7TWccm8ScTp86LTjKh
OtIo0OLiZXnYr4UAu0HdtqhvJ6fnM6lsTZgLsplsF9gTBLu7nVB4FrejiBfrPApsN/tcVfl2Bw3t
WIoqLdFPql9UDm/aRuXvCGfDCKjUMIQiAySXTSwvIhu4dC3ItuLE6jdbTW0FRUY+qm5SXBg2+ATb
msKDtV2D4LDhB+PT1hihSfFLRBYJHawfhmaHl0pwiD44nHjlzbowoldsTctJ3y/G0XDZqSQGbvfs
ao2wpapstF6dq7IxWg+1lkuyKWKsJeYx+dvv9c/P1JATWgQe87tycjpjeQsRT0IQ2SrFDelYyM+y
AW1xF/3uEFWGpa6mGimAOV55kDDzEqVL57d1j+VHPCcRAV8WckFQbovJJcwQ1doEOhRd67ySC/2P
RikLLn+qH+33Z5QwHqUtodFaIcIaMm58cUyUge0ArfB3N5k33k4DYhwXb3D03W4JA2Bj1agClGly
b8P2vvHBup2fckqvzILMrp8U7DdG/LNyD4F60KzHWxsi66O3hFW3aZpipjGxMQpbubDIvXkYCU7M
S+luZ9qfqjxheMRq19VYjYaPqFEsbUtzuw0O/3wiR+m38I2flb+2pALJuXBEv9GhklwkxshlbZf6
LvMd8bOcotTk0/C6E/FH7PMaizY25iFIJiy7K3PlOcIcbXf8AaDGzWvRMSBkD7tWcPvx0YVB+ddX
QRja0lr0XDaIeCAqW0iyTQinjRWbCVrDSgMCAnLcJEc09blI+KfvJFvaYZGTWcnJv+AxwGRbz9pk
Y2Nz3L3cLifEZikRzqwnecNSeJCP7r0KGTiceYiXVCxq7BwQaA0sHcakVuwgRzYsdTFzwKiWQvJw
rsMMywKi+WmyXBiGFgr2LxpP76OVFoO3aHlLUDLVaFx+ZrhOuf93c8YeaFB8X76fSkqsD9N+o5zE
HxfZ+BsoUI3bBQQF+CaZOfj1fRQ/8rp6BEl5l8bIRDZ29r5pe9/dGwAC+Dpp7NIOrck3Lo0xClMS
c+VCCIBafZLzc2yxqxl+MZI4RviJj2ewxqciFLb1W3WQTrj3skxwyOuKN5vqLYDPzkUME6pl1ugn
zPg9tf9o3y7fottyw7nFhb6BJeh1WG981E8rMr4h9Akq/iYTQishyrkSerHiGHpoiGgfV0WHtlGH
jau7S28mwKdv1P4zY9vLtib2wlqGuvRzHAw7VWJH4giAEujiOE8uOWQiCirg965xlQr+e/RTrzfD
c6j+8T90HOkDN2288FrlpEw0R84sNaJGEOFn1QOv0hUUMfbn+c5FA1PQyJIkCNIHPnYzkxCabysR
RkeiH/gzaQBttcXwuXIp7YyT2HG3NpLsAEf0xuqOzvxAblZ85RImZGkYKiiQToUrkcFUebR1CkqL
D4OMMJkQkS4Mg8GS4t/cJ4Bs7Fk0c+fMI8MorrUhABKCSHTc8JA+enPWTUWB5inWUm0geL9Fp+xE
lvyiYp+c/D8F+UtDinW8TEQM666YtwGl31gS+MtwC+4jKDndxbZJwjC8Sq7rhXjr3xrVMs24Wo4b
hAD4pDfPd5OBHMq8wQCZaoSP1NxdEipJzqNzKx+/CJSKSg41i0oikhQVcuYNkBB5bKHDcxtehj45
VrgE9yXIhxe0s8DH4GzbsYulhn70J7vpNqJ+hJYO1rsbmuxPOBOrwUCU2tQ/nhypltBWo6AOC1bZ
DfGjjDFf6TAQzbsinjgcOKgzq5gceUSRzHoujVUgbToSwq1SWeKuHRCBdGqE3YoZIQfqdo3UynzG
JbgOMhOFOExofIRohAW7SId4z1Q8Bmx0awCBRHsMtdNYCtyNfnCwzeZjzPE9vtyfYN9FFOAfdK40
7342fWhER28vmPsYhC1Ho+1dAgx1oAwe15GJpX8BB/I4ubcghL5ZJMMB9p7y3e4N3If7YcED+HcW
oeS23DjjEz/q9mhbDxz31nB9haaMqGSdMIT30A0GK+WrmYbqRXQhLAwP5HQ1ehbapOQ6U74wiRED
NdpijsO46s1tC89FL7MbNBfohciuCUEHlTrDAo7fgWh3rta5cDUTUJEj8ooWEQ23/zR+vtPvtM5e
MHb4nwXuq0n8MPksM0REoi3Im+EvmBQvKwgKB4cxgvfSsuBTpvg0+K+cVCJPoyIlXHcURFXMKy0l
JKMUsZPA2MIOM3ruoP0ZLd/YWOQfaUc0tGFnhQ/Qy419jOaYfq6Va5YHQNrH6Hz6ptyYsf+q4EMo
zs+vCf3NLdqlycE10vt3H4rrDdXmFPBNP1w3BbJhQsh9hgRHZKnlAzXHnelNwGot/kjC5rmm9qka
0T+A8x8RlLJKeVfNUOvQtgCcMXJtU1EVpd4Fl0qNCikXb3wChnFyzoebsjmLgfPWWWArZZX7uXPn
dOocqHFR56/RJhYvjYIMeMjORmglkU/j40eDilpbDw807o+Mc3WWkbXh4nWb5kmBxDPecvxNcDf2
nAv1WRzPYZY3TR6SadwEFFjYVo19iE9mefc7bA+vV41+QBIlUT9BHeIrjA9TjQztRTET4Wz9aL+S
jzDdOv5INm7GSPLHayvDRKVF/znx/pHp5EXK8dbL1P3ODYus7/x7oPWmn85Szr8qRxT/WCO8w6PG
xo/rhgOCUn/VLyOLG6vDNWQ6vK/20jAd4+SiYcDCxZdl3kO3yla1UVtP38nmj+VMA0y+w9TKoztk
ggTzTMeJAVkl95FTk9kAijo349qy0tAa+0YpTUzFjC/EKb7LPEGv7JWg43UvfJE4ltLrDmZRxrc3
AYTZlnL/I2Aow56vUBk2jz0g6Trh/NDOGzB4g3pP7BF+uWTIHm0JRmA1KdQOQQKDTLy3hfhb+SAG
avhDQthIKjJVYTEpV2r5h//WHRG+iK7P9Hz2xqhWZN8ETJWt3etPr4FYQJ0L7AjN8FuvjAMUsh/z
aqTNnAKSfiR4i+6UAeUwNJVxZYComy7/oqVFGPu28yZm/qm3vnPg6ti/lRj+Gxbn5cfkG6Jqy/5Q
8O1vH9aaNegNhqnW5shY0Jf6j5rXKkEB2vyhVlfF/ea7ifS88hGBVjPjPa4PNpDsdbd8xHJK8hBP
tn8ql6b3mepCOsBIqFywtXP+tAiY02Rhai44VVsV0nyZYSETdZoIS61DVvjaRQf0iAdYFA/CGg52
uRcp3h4io4Z8RtgN0bbcgn+ySgawC8p8+lQYQ//DTm9V5L6qt0MGa291RSrEbDSnl79u03GQp/Aq
pzsnm0NwZTGfBzo7fUNfezmQEofbsurME0Ch8iEijVpROIpLoVZLujJcP9XDk89L2xP3oRbfjeGr
853os3RjvjorbQIRjuaNrqCq4y14sIAn7MUVanSDLbWkqR9lFe21IAJahFx7RDFMkKIJJBNuA1BU
eXWVPQTdhOuTB0HHKRNCKs66yc251NWuIVEkqgwhOSqMQhzUs/3vpkgDHj+4mb4GnGdnmNJ0jQRw
wG9IQWUp4KHr24vcaHL3q9XnRXow0dZJhYW3W9IcVNeIYIv+YCXojf/IdSwtc19j7xXm9Vy108h4
29j3POjBFnO3O+ncJac+VgG5OPec9jubG0BIsvwqMjVmaYwGrZFd3JusqgCYw0RMesZ67Y6anHEM
dk3c7fLe0bbBa8BhE/rrZcrDvMIu4CWSP6Vt6WDm3Efq29Xzwd/AygzifOx/X22lqU5i3tLVSYc/
cA1c+5o4Aa/hM359mGoItZDftCJCEaiFkosVaRJjJTCbPYmSaIecjzdQq9QnZsJlWUJk7xnThY1w
D3JgVpQL7RL+qeuahsjcRz2wE5N4hNUEOcnWXpSFFZeqTxTcEiB3U6W4QGroeSAokdnfSS8MQGfq
GU2dfsYKE9N5deqK62U4uEz4bsiCRBq1+1Hpjao7iBSpKJ0Y+NL2S1vZ60O6laEJ8Z/0Kh+dHFk2
G20NtREKNkkWeVj2aG1CB2H1QzKbcZmvaJ65zbMrUSNv4UXgrQrBIXbxsWOgc7+isCDrxw4n5Whw
91XFgHfW5T4UCmF9hlnJcqbscaCrVVWQWyiLcvZETOf0+T5PceNd2An5VTm4VRG5tBpEYdWD4BIM
I3sAPvhBENV3gZ24qxfFp+pDW7YtrAdSLIHMrN3P8r11YQVbf7wtO5CiCIdfMRgdo93pjCVhREle
5mkYg/xTHp1bWAkEc8n6BveEJ0gB7VkJ/BEP/Ks/QcaRLs69cywFLm7mJBHv6wAjuN6rQDz0lBTr
8ne+zcO2VT+LMLEcUuijuVTEUCKkr+xnzo+yJRmLRt+WsBIY9UCrd/rrIdGf6VWYUAEShbRfOpKg
RVidNX9z09R7NR7S1dktcJqZkzXzsOVyT2MGQNhPdBnpM2f1G0wAab3MJSaRMRU0fqxUxJHcqrTQ
Vuc37l8PQP49dpzExqAuOmv3FIhzrBj2pNaakZd8wdtDVtLfkIA6poOOATARoRgEg/6plyptVcEN
kaYriaNUK73jqAZWMnlyUsBvVRd2hyidMhTisKproCVXWY7jkyn6VcG6GX7lQOUZ0SV0vkwsYBMH
tOx8rD4cf8FuQ3nGmFjMV+Ff5b9jVf360Xemr7vmRBQa+dDLFWCKuvipeU4tm/QF27Y3O7DGHBBR
g0mGgHjL1rE/S3ScxVmP+IVrIIKZnih7mjy2aaJXIblz+IECdMLtiI+uEdrTiVmj2ua1fRMxUlkw
GlAZQkr9XHEzqvwaxL87DMxfwmGnvnijgjShDO5Yy93Y4KM5+Aa23WpT0eO7EnKd+H2Ajljn8bM5
9LIS97gYY6fdDUUNhiquqZCQQuJ/jrCLpeSrGKCOrqFQ//prvm1TzNGVfbdLOWmJeNetHPMhg+Jx
m3hRSh4u3lHiykrEipFCw94HOCO7Dh9JjqAwWfORMCPXI0eW1JLnseFY/lhbqGSH3BgbpvcTuHFi
f6Bv+7JL3Hdre/OKog9WGRX4nSrxp6ui5xPHuFvUYGoqKISQEr20Q4IYKm+U0xhx471+Y92+2mm4
QibxoOrBB6C3uOcK6LUOR+O1A+mljr2S2k6c4fd+wJbS2xZzw05v5vfHZWAGQW/qXjBZBTEpSfV/
OZDMEo4dTKjAFD94YnFvf1bqz/etyn0stysX3ZZQOs/8t3ptWf+9FK1go6HOlraO9A27r5Doyuvr
IEiVzD1l1hkeRNtEnFfeReHaJpmuphF4LE8r/CRl9Ab3XRL7d/ma/oa6mgpQSIQHbMWXJv1xi6Bc
sWQ4dE4UfzGTco5m6JtMacmmBMWOYICLRrJcc4LxtBqONMKzhazRP984CFeAdg137Lhcc7dlEt1j
6ItjPI9xJtIYeNMMktc1y8UtFIaOFBj99WUMZs8LcuOv0xS3Wy/Rx5pjKMEq4Bjdrsedotcmd9JA
4APMALQYbk7yjTKrKhKz8TO/iXyUQCXpsk/0VYJuH7C9g+umSGD+/sLogwMXcnxAmZkgbLR4V9n7
4JufB1Ex0LNmeSSrmkrmc+cDYeiUCcjpYJIa2w7azcveUKPDSR/VJNBValyeBQZHuWH6XDxMVf7b
bDrY7UkPNBlrDnTz4bQQLlAzrFL3crhTBC3rDEHE6d9l7DrG3JvVxXbZQiFXBsYrHvw8Sctt3Go6
GyE5Lxob3yVx17Dzr6dWBeoonuwvjxoHYEg++p2bOBCLrwM6TA1Ds9PsbTad5ppz5UNpEG7i26xn
Cu0Nkv4lTgx6HkKB5lADUapiXRC4g1mzlrwLvbl7DXHWnF98KIJiL+W4s+Ozk8go+v/vij4WwUTR
yHB8Yc7KfikuNPFSCIv/aAhqVxF9pQkiJxBSZSeJaXyJUTYDhe5xC0dlwBKNMGpKbkuq4BHrJFBJ
HP5V7hSET1noweqHyG+7U+MWgaZ0wemKC6D/WsJ+S0+uE0mjaxQuhv4HEE1nMXrIrm2Q2GBZ4aB3
ZXwA4M0jZpNWSV8ZF74sZguRnxsu3BSDuVgoJ3TusY0vGGb/O7aStMga7mELwv/zv8ixpUm3aLcO
nplumOg8SacFbWL+rDtLJF4Ijzmn5BvdMUrzSqLhhGoadSvMSzDJkKefromM3dFeY/B+XagdORiY
IYj0L30V2cgQbdFMXQMSP9cYP4KhzQ1an9MR4EcUuNVOExVHAY8dyRJQb4zEbktNEzaPiqI43OVL
TRdgmkA52J9P9fEc4xSN9AhSk4wvawYL2Lqah8EZuO2Xb4lDIs269I8we4p2G/Ddp9yfqOZOuTxM
itvnen5HqNc+SzQeJy0t9QswkhF1fGNPpqhyJ1DX8uA0LsC8wOXFYkNr8kZiQr/S96YLjqgMQILD
ndSDZ5H8qsu7Dk3j6Uxq2K46X+MdB3BC/bhVXVrUqK+rMydcY6uTm+Yt/PSLlO8XBytfON7XocUA
parewwpxAPyIlNJEVMqgZHBrc6ka8CUF1EsHd9ZR3FF4RcEdsYIgGxofOMxkZPlCifvopjpVSLwn
UqcosrH+5sfCRsx+P3AqxCXE7UyqQiPNQBQdAXTDu8pWPweUWOK4WUn8tSYkMgWXgL6nUtky+dEY
DooGyERO0arovU26yWf84+QwuzGrTX78otc2AguPuXiQbVWE1kanwv+SGiB1ke7mYj4mQc7YXlmR
7cXOLPHkuPuXxb/667sq12ahilxg2YVULKUObrat4KWThWDLHZsQqWX94lBYt4QKIeOHcCRoMniF
INAbK1Rlj7bG0VMuRTvekD/WCFoC5IAgoLmMbOgm7eGG1Em412y/aI2bfH6mOIHSR7ypoT+ro2Re
/ZRZYWC4lIMgobqSoBJ6UZ88ROg1KbNRVGQo1IxpxgMN7ZJmSP3GTHsmwjgc0aOoXIOVbaGd5FxY
kGJ9YzN3td9oz1Sjz0sMZ3PF82w6q7OgeXcux9yNuC8mqEcrThJuLuKujHYfklhUG5wAFGjaspwj
BBqCQ7XITJg3oXbe6PX6o0GyG0Ono+/XnXZkJx8mD+iDx+XBKOOgtlOM4sKHKXXVgq/lfaZVaEwS
qlpCbdEk6kacWOybCVWujVovP4q/8jD1VHrLKlUkBtKNtxkJB7+0tBmrm+r441tl1n2X0e9xvfUW
0qan18c5Pb/+LkpXJtFfnc023TUZFkukfM4VODqGFgBbL1ew6AuB1aZoeLg6srtw4qBaeZJoMjig
V8d+/RCtJ6FSeOckGTJGiCoMI/rXbocxMKBSsYO+vNeFnedD8OWKd9IA4JLH00uCHGhaZumTeVlL
MvMFsJVUq/5+yiQuWsKSBojji6DUf6I35TLyen1t/VkEAABOUZUmrCE79AiM8FuID+lVaGG9HnIA
tKAubcjMzU9U5QnJpQmiK9207HWu7ggCtscT9aodkbckbBDQwf9YSTJiBtlE8oAxzRQVlpUf7G0U
TwM9EUdi0HCEfCHt73PHrTmACBdtuJUD6rG8SYpPkSIe9+Vp1rBOHi8KIQH/XAy/rOAPbG4pt27k
+1Ehg1hNhGLcFbziW5NscoaJct7hAxiJ9IDDzmhsLWQVCUtMYHnjuy7EYkjSA9gXpqfNGNPPbt5h
tXhqeX8unbywuqCXC7chTUOlVrV7vKeOwEDJZ0K9vvBOGdCdnBhIpTF4r5hi1hDojh1J0HTiPVJ2
MfRMqKUC7i+pIxhZ/T+BP8pGPPMTmeBE3u5xkZRP8FciF3kW8KUbQGFAniIaGdBeBjQXrYjJ39b4
SaYE/GFM9K9rdnG52Vuaz9FaBksPdxxJSrAdrr15bDf3yV2xsajIshdm8UrvRMmZqenSQ/bAzE7N
1cIfHOH4KgC61Eyh3VASIQvgf0p49akNg1DrlAc5wfcOHMjtX5iLOajcYhClWrpuqDK1cjJDJ0da
xID25q+ypUjPpMs7918I9DtCLbRAhJDwDmTTlSapRpBHBqA1DyI+Gm6Wf230kSzMMheiW0DuynIJ
pU0D3XEA2s2JAdJtEDl3vMNTWrZ1uGTwM6QjaC+z2YcWI17Zhrl1gMlmNOemGBDi2JhuYuZqhhgF
nlqIhiZ3EapLOyd2kye5GSqH2Vz0uIiH6gQKE8fzMTz/RnFe9c061kc0mx5BXatlZyMQj0topQT+
5zELWhmGwR9GU3fRYt7yh/Y3KiQHN/BR/WAAo9sXo2xh3D6FuFMnd+bO26hiDaqxl+j2kjqMKO6u
LVpZDGs2Pzq4aaPXgQa5A5EywZ2DkVymkk/5IbpygmuqYnxfW2nB4rYpsF9LY/t9C7o1R6WpGBEg
P0pSVfF1VDXZmtMWy1rbD0utwmJc+bAl2zDjgGqoWKykLT+R/22iQNvcrAmgY+aUCgcuxt7Kw4CV
X4q0OozDK4Ld4CwXHlmIb1im3qlvG1mFzm5YXT8AlZ0LOKsiJR/ReTCNZg43RqLoYfklPHWcgtW/
QO52ZqlKON9/OoBttrLiGGwifdG7g7tGp3fQAKyzhJYOpA/IDrGLF0OH0BeoahFhCK6g+HbZVz0D
7Mj5fRgtEIbp9jIbecutgnyBaY/XHutJRvsVyinLmeLy361uLKWpnGMWfRHNQxVTTb9u9zXnnhm6
XqIUXzpqz4zw1SiZi6ipuZMcYZk2W7UTwSREpTbINpa0+SY2mwxlxMuL7CpeqCL+qw/oFmQ3u8OZ
MVhY+c2h1/SwlxXg4znW5AG++d0/atFymT/ZJje/Cu61h/UKJoeMDfpf27zlN3In48dtAl9jRbK5
xy6eaBGOI+e8xLDFH0eB1UyF6WSBK/GQRXq2MK2w7HRtWfYfJ2V47fIhQlop95q145OJCocKEzbG
RjCRj1ElAOa7zruZfXZDHgbT5/Jqwh+Oja3eCtIv6VeRx3KSfT9sY0fp+r9J2lfrYVCDas4KwHAg
8rnJCZLwY6lzxZACS8ePC4Bwco3yEXSnDFRvqcoYlfLUwit3CpuCccDG9kJ6FDuCzB/nYF0xex/e
xyucNvZLNVXjz7bj8pIy9xVD5NOsPmoanBHvGCPbZxz/z67jmPtx8kv4zhnoWOg3d2SA1KuFqbg0
U8zelQY/nEspUY+pbW4UoHUVVHT7iImxTGcaVLe9UoMr8jjI1+7tonaB43NgB5lPJbUlUEW7syEc
oFeMvX+M01jLEbjCpKe2ISzEMn/IDhw8Rq/m1H1JBe0RxFiLB29zFkbmpG6iRZbuW10zQkus8JGe
lRrRUCd3h+xC/Vm2Blml3VR8x2VWGP7SAW/JhjgyNUj25SK54betOGPjC/uKAh5fW7BHlkHwAX3z
Iuevfxb25eFl2v1bqDgmTWVhfS6NOdxTw7DDzKXOmE9yIFVjsVSadyZz4Vfi9225ayqI5Xf7HyOk
9fxr9Z/G8bmgc2GrXwoKyxiCH26mEHFfd3m0CZJMWbPH+toXOVK8fwmpxeKL+Ttu9jIIdwwbxhle
qOhw2CYUPB0K35DG9qsary2cK5dpa5iKpAxfBM2JZstic/zk7A2VX8hkyjyuImuzLDStXxyCeoXj
gRPKhNMa1JVEmQaxjckRDvL6b2EjaxhWD67En06V5RIamDAq0wNvAcayonaIgCcpenwM+FJoaGDR
oeuFxONiY7MhNUWNmBf3wk0IbnZgPdHavX48zFIG1jAmSvioVH8vUNQ/mxbIXExDZ6UmRuVNI5W2
A8VpknNeS2/Ggo+dGA+Mfrp+Ve3z5pIkUz/pD1tfuvIXYxr2qg/3w1SzUGFkJ4I/zSUCka259kCI
kFEIXAPyPoU8Vqdk/uqbtLOOk4o6g4WbJOFBLd2mhpWGisPkVew4uHlO16d98zGaBK4CfM0OCNEZ
9SjohiuXUqW9rxismRf5bDyxYlyGGfUsvy3efeQqMgheBpYNeuvtQ/qMTCp1P4x56haOwepB1Mpr
d1wn5r3ZZB/yJe42FWYG/OUPYnrPs7KYV5+Rmlx2LCA0XVSnvpYtLy0j8NH+dRihtsNmjALTeJTi
kUXmS2krZj+9HDv32pR9It1PfA3igeoqh22fkaVV627RJtmxdD5dN6Lv7hYzdZcfN1cAVqOt5fGR
E7m54oU+/kYhouUbpZSSvnJa7RyjM6qfbvRhsQapRD3bdWWCE1/hdbSAwwr/CZCZ6AhC854pfOsu
HAEYyrsAkKlIiBAeQqZ8mrVdqi6YueWcJCa+6TLObOUGFhPyB/DGJvdsRBacQEsNsAvjBcnPTimQ
T4qnpdpOqjLoUhjRC8QF7xJZHbu1BZDqAA6ad3si79MahzSM+wmkTRGKWRm2poykN1FWfEPJg7D8
WuEzv+vvQB7DtznmIE61MuvxDezaVKvKCTzbJQWnElqSfphGyM/GJe03oQnSaWRFKXCHLB/HnzYz
0e0rHnUBxaVM64J4Q9ibZCyUA2YFvPIMjM3Lm2mFbpmbjqmNnGh3h6+OB1oNQJWbp62rrTb3YSKy
GrfV6rl6VjRItBpuQ89X4PW5AbrElcb62Co/E6IfiuWH0T+qO+DLVglI+O5S5JFV9ZX2GZDx3aOq
f/zpQ479rwJnKBvA+Wgm6yoECxxzRR8y5cyBTub0VSUlFuBeQdWZtYYMrJ0oqOgJzrvectzEwrOh
WYmnQJIiz8NhzZiSAvk0PKEbCIXmPdD/VpIjBi3LqZx6Eh/M4uZ+B2IsK3+GHXw0zrmATObZ/lWk
L6hW88w91DEvNB/Nh1sAFgJqrhB3ftFy6IfQgW/MLDbb3JDK4p5EkibiwigZ0iMMEI0WB5fKCwoS
7yLbfViMS00NwddpItnNx4m5jiCnttvhLXYLaG2n6ljumiWahUm22NbnCixQULaH3trKN8687ZJQ
tpkEFMWzRlBxpdZMMJJBD6hg5WNKp5SFse9GuO1J+yDJ2WSrEXcwpCYGWG/ygeS6Q5pd09cOzfx4
ROzhpZFiKPVszcIvxY0a1DTcGlEB+39Dr4Rgkm4HRLclO0PP9NW0dC1TpV10PZNKxkFIymyocWv8
ORZ4MIIkjIw/V8U/NGhe2/gzaLXPRb0vVPAaPdiO+Wwhi7ejReKY+lxU4uSDjPJmCFDEW97xx4XD
TeqlsVPBo1IJy3t+CtRzTE2G+NHEjwSRQzUxCdYUrIYn7Kr7ZO/pHyqUWEhixpiLf83ZpFVtDvKM
GdbO48oe2MxqSjzzWcf+6LVOOVl6xxSUghR98y8WTHRjzOhyrZiwQKLQDiB0sTIVNZ1aDs+nTb9l
QBXpnhi1psda0KcRKFgoozfZe5OXlK5bK4JtmGW+3mtCl5BAyShSXQ6VC67rhzleAIYUXzuw+w+o
pUfSlO7WlFkbHgL1RT6cA5FiDCZlpm7cW04I5llp5499SGO8IGh3xt0wxE6rdwBLMWmVvYSMP2OE
gSkU7dZXQB97KqbvQlP7a3jemf9B0126rU18NJZnHmrR+/LskZ/9EHVR6xlFIXGNtaOatKmEnCzb
2RmSztaiiOgPKs4oG/X9mRfmzoQFbM3SffUG1/eLs1h4g8VKL3439G163Oo6P3Ay8CVpNticq1uV
OaWDpNWi9brR5kTGBpnp9NYVd/L76KV9hZWr0DBsSTmMc111zEmNmIwUaljrxYdJsRtvPsVvR7N4
Isv2te/emC4wtQHuhaniYBhqIurGuYkyqgrJi4mnGNYT9VzvVT/xHWaIHFUymlu+kWvf7Akgyoos
U0brNZH39xVBaVExKfXJXtauQOesc7R0Fq1RXw1MFJ+lLBGNHVBzYJIV+FOCYOA/ufKyL5gURnnw
fjbrIjYX0sqbwsaMVhKWESgkJYERsxJtsC5Sy2hnAj3WAdURmTuzapoh0uqN+RoVU2NLPy+iFGkw
pJFKb0GHpGLEihcxBWJPe+75ROskGi2hhOh+TJY8JVsQeSHJSh2jcWlJM85DMWaOmhDI4GpFBR3t
YxvtSNOVq438kPM0CCbOma1NG6dR61JfR6lUzAhtr7jlr8nPT9JbpjrHqIUBmQas1yQ+qvt4yR3i
d1V+dSkJtRjavyzunYNxT0fC0aZxGz+8+19bT+N2JZ3yQVyE+4XqljcJg7WrZFxLtY0ZPslF0FTt
crN9EFQmStYkX+RUpg5BZEjDjVMTJdJYCT20CNxQlGqU9rXRII0AVoQU22x87u1OHGbj4XWWADrW
BomGH0K3Jzw/GrHMmlvGwChnRC79NHC53qZPToTS+PF/X/+gZBc9LXDcVQ/ovJb7Ob7Yr8LABNFy
2zTdEtLLdHdV5yS8/ZPFtbS6i0zrd7RPmfbXy5UkjLeELMJ/q7gPpWsmXAX+fZ0oEmygFEB6Aynk
msnGfe57Pdo9RDsOMm0y1PBnWHiX+qikCn88M8/JaxPzte+XLMhnFVvsK1CdnDpI/uiPZMpa4wEd
hXUbSsaXDGLmwMyX2RytJekXwc4dyJMx43CiocA+kXsmHqPEnFiQIVAW8A5adhPOfFKOptHOIAbH
0DkkqChFFeqls0E3XZG1Zocke/ksFheLtczd+dRT0L1PoVpgcBQt9e9+vQtY3EQssIJuFk03TGp+
dhIHlUP0nyDsmfD3mdPwV0wqZVx/zzHdXfbhyZ/jm7A4fgSIvAdKBJlTYQw4lzh2d6Pzwg5eYis0
4RZbutbTirDcW1wGVAqD+TVtMndmTPwX2580WzKeBYgUbXnxLgfWZ+z5IzOJ5a+54LeMMQEAPmJI
+eflCJD2R+Eu0HpdTmRTdqdqmSqNkz6bgU0GC3M5KEHWbx/BOgSIDiUx9ZvsSTGkHbcJNUP7Oz+8
/5SsQx3BvS9ph1bMD5pLPweEVeR6Vgi/IwL58lH3o3H/LXfJ4zeV777p9EgVW0flNlrVxeNz8U5D
6Sb5ZCh/RkoiV9IhzttGoztmRRyVpQo2RrPOxabnR1aoG9inXmYanpmHQ1k0yG4eHPWV5xf9sG/F
UIoGjDtC3SczrQDRp9v2qjBXQElUOj0D7vgp3fpGUVriiBcCFcy/+F/7HwLVmqlRdUg1kBpJWTed
dXgRK9cTpHfa5DG4NjhIhRxpKkLk+1ox/SBhCbaPpzZRYs4w7YtJ42RlKrNvujmBDIZ51ebVsZWP
LDeeYeQaHOzQCVKFE2mK8o66CPbalzDoTiPe01nwg7kvs8wQmoWjE8Zm4OwzrXHLSxgca2E+rUjz
yE2RsAw3tR+535Md13KIeuc0KLP8upH8NpH0ZNYKAIsKxjh2ht1X16Sg3bvoiU4aSYYrFDN5Ye/N
qH/6vS6/C97Z0vVn05qXqTUlMK8532rSCjfu6IlNOdxdXZOhVCl/DAFvw11PNTyBzYOvcyvLfFEp
LqbEGpuyidc9ikdF5dvJ5ONaiHKh2Rrnq+SyayyZJya1+xOTcZRxR8l21K9Q+21o1bjCb5SwedPC
RCWpFdDVsUwfKBQ169/IzwXOWonbzGSDjQoS9ksrqkD3fZBBI326B9dVapzfEtimS3sQO7+G/QKe
fUj/jq2Siu2OqMiogmv8ChwUz3YLRcsNmJGDhkyy98AlebcyT7T4x+TCR8+wE/3xRNmUEDr1ieql
C2ztSHoVbRT7jf+NHi6Z3aDxtUZn6nDxD4wh1C26qheDlv1qPvf/qQdeRwbhBrAlfJ+aIbK5ruik
OpIrFqcL1g8vUgp2HTsw9xBY8ubG+C3r/YVU2s+BY9QMqNjt4pBHov7elmfrJs0fJUCAbpNbHsc9
1iMCK7Z/bVaE39K/ooRYTItaqaPYhn0DEYBPV2svMUdqAiT7vhnSS3AaFT6/bCRjDV+TeoOQvsZV
DENrjm5GJ2pan5TkQZvGw9iLht7+kLNVcrKstRDMCq27mg8bcBH2mhaLU5elFYd9OIjA2YO+ensx
aioMinop2lRXsBqsRGU1JVBgtmzqWwaZsQsAPFhAaw1yt6kL5nNFCQAhsd41a70xnmf816jgyOQk
78BIIC09fEpu1/gAL821h3esZ82cCyTrADFCn5a0YeZd4IkVQJ0Vn0TuTASc5vcOl7hq2+cPDVaH
E3pOvErJ+N/53FYT2SHAh9Uhxo9HtKMa2ZmrykEW8LviEmjnC7ExI5dOLQDqxIRGhwGIJlJHYH7n
v+dcDjc0C88zErpVpP50vAy2hj2vNNIDPwAT1e/sci+CMzXU/dAEfOb2rd7pbXiBpLJmPQ6S+yUq
K18myjoMQCHaPYwU9bfEIUdWmUYWbWuimiJaqLpXtLkZGl867o48eKWJqTMjd8OelfgHJV2Oplop
uU6E8dk54upgKb/fKd4avIQzzGjq2S53Au5v+1oBsSKVW4HCT+XfQCDralyDmHk+CT4TcA/yA6Ie
lUz3enTYvXf6N+VjFnJDnuPDK7L1fOs2rvDt7nzRYIlm+Po52pRIo2PfY+cEOYnjt0J3QepuFr/v
iekSCxgB02u4Hd4kWmekXu/In/7rOS1ZPXDHyPXc3cZtpyccjc2/8b23zMQT83bP3MLfZ3tumFEM
a5l8RPqOArWH8gS2Kl/r7POIiLR8gUWuMDGaXUowAEiibaroMzdSD8mtq21Xt/PawfsliWClpVMU
NeQww3tdto8Gpb0FaKhCdsOuUl90x8T2SQKFsC0Oqs3AyaEyJXXGrPEqhs4N8/MqIeG63PTX71EJ
oMts8E22rTlKG2yvgABw3wV82ZnYYhRuAJTZMlY/WuAYlAXmeIrHEBQpffQ2WAMJ6UUSwkx2EnlW
5f0NIAp+/3DLYyJKNLfr9JiuCziaUvPbf7mByhqK0NZI0K3loxITs4AJWyZdtPcLAqznqNpqGvlP
/aVEU7MbqrtK/B8t3NcsZz0rb9gWAX54qpr6rjdNXQw7bg2D8AUG6htG1LEcfQowAU8yGifz3LBA
j+WzR/pCLnR5LU6XjCXuFTDrXxcGi7gke7VNU1qYKGZbFYeLsTP3oDHh8oxvE2O7KRRMMAIYogeC
zk8+QWwgBkOfx4oBmw/KZ5MGUEfREtvAyT80wuihuPXALzNWTgOhI0QyE7xtKwLO9WyKO8nApBUI
C1PiVckMzQZMkfXB9lbxjSd09zGUG8VsV8ezmGB1UB4mWn4MlFImCGgWtwMbK59lK9H+OjlDTdNQ
VJBvvuj+lDR+cKhRIeK1jE5D3mt9A1bUHOlEFLGCM5jeqyBXlxVpYDzFzA7RbhlSItL3fE+at/Uj
FRui6vobaSm1ycsFkLxQq8UbHC1xq7WSQdYei2bwyBwdJsOO226n/VbQmLzCCdgo7fgl5wXUIrIc
Vnik/8e2omTJbZlywWObV6cR8RypejtjL002+l2tFKJolRJ8JfxPyepzATFrXiqnUQJhd1VGTAcQ
Liz8L5/fFRIBw2/qEC4xn46Tzxra2tjhGFDjtTADjBlZwc872OGDGucldw9E7zZQKxBBSBuOaQC7
EhnkU6dzfChupFFviT+fKR4BfCTHtI9NvhzdCjUMDczRB/Nbff3RoFLNXabQUHrI0y6evUfSFdJj
3TnskEMCt7yFrQMSqPj+DuusLMFnGcSVAYC1S4DVP9i0YtnTAz/gWPQJ9umaPEfuJpR3TyrO83g+
hh023d+C5/xMn6oHvfgusseO4sVcmdbQ8OlKUQqIDNnZ51YjxKQkELyv/xeF5WJPbUrxo9sA3HBk
QYA7rcMF+TymcGpBtHsis5N/8TzAWvvxHlsQUHFFx3BzohAN1nqt+xZzBLISQyT0h0VTvVBvmds5
3N9uswgyCk3CV1I7NCh35ohc66c6ouAOB22sZF+CcZX7G5zcP1+CdZSjl9VGdPoDzRXtUpkaHWlV
Dzo0l32TOp3gYVGISAyDU+jmkos6352WrU730Gg0/G3rDWAT+2wTIuy/x9iNGkjVRub0MR8++aRU
WnQ645BpPbqS8MnO3ybYGDnh/p04skf70febi5XellWer7PiFwgPvQ2qFeTwWZqseTo8vnGiVI2+
6R+dz2AKj/0DBiZ+PaSAWVdUFVwYE9zU0tCFZvLm+y0q/aKyFF/8IVaysXMkm9ECcUeFsYLXRxFy
R7f3/1tk22Kx8Gm7rvcx7oc2u+68rEvViLcTOztrMsk46DnQ1L7/nu0RoG4CfLJT7yErG+MdC7sa
2r13/8mpSkQzEj2OzhtJUlBxc/gXMxgTEFdAupMwnDZSBCmjeO4WWcAbwidtP1SuEZ/3grtc/WKh
CK6Qf9jo4Cxdb96FcH0i2ouD6OAEyTw5Lm8hmM51yYIlvueo9sSmdsCTnfMfmA+4eQc1qs3onN3+
CGbka6zHwXl/XFyyTNNWjru7Daa0QL6aNbmo7j+IlPet5Sp2/W3XReD6czyeBkhdliiPPmY7DKK0
MuPHqh12P3ZdzkzKYbRP/bkdmE6F+TDk6V8widfbP8pphUEYlLB6kdmE8xIr1Kw1cDLphBz+sCoG
R5A+e02zbAJ03pRI9qOzC24Xt61wsgW71wAFiag9myILbrjAUrR3ZBrIKt0/bB0wwYyQaB6e1w7u
sWdWDYfNqX7IjvRAf42ydtwrwmQ5iEgJiI0OpwhPl95zSCzuW4LKrtxZ+Xy0W7MofkKmJPs9ycTT
9uMq1qHm9UExD6cun8/ryZkvtcGRyZAOqKxRuN8mfx98xlef3Q/3e5PodHsVpKHh6UMbdnUFpwpI
ZjzpmUmkpn0Mdj0DUzfQH6HiEwsAfIodjJVpf9+DgaQ72uvhI+pSdDy8aTwVQtPwJdMizSg4E94J
dmN2/Dw/PsOKd4JujbhnuWrmGIeURxAxC+BQKyDnSxjTeAWrCrejBbRiqffpg+jd8PWJlkzf05wF
/dRHhuuix1j39AlQRDukUSJx7epqnnL/fDheY0m7trOAWQ3khZTyyp3n4FYpvqre1Cv2rZ0oHxDP
ynPHwc+rE/7+wagcDdXNGNZQkpdAD7e5FGa4XBqaZUoqwN4vfg6kLl0Q/MDP8K4ChECr0fzeMEvS
WKkq7+az8KiGZXvnqB5kUGsdnSxonFEthVpZJezYi68D3zI4mqewWxr9aWn0EzYW0j+fQLWbXbR1
81bsUOsiIu7xil5o6ApWWXBEOiTOsOF18mU6ryxQZQtPBHnAx4GxY7gZEcCH7Ipf5xlf+GDOv8lt
aSL9SP6tpsO1jvp4vKptUid96ROrMKeTYxyjs+Dr+9CFnw4MIjMYaqn4EXilaR4kaRZ9BFFZGa5H
vFN13IYaFTWERUIppbtCizgCKtDThtZnGN12bkxhGs5BUc6SYyznw3n9X9793enxdTh8tdePJYu2
wjYEBJ/NrjLS33Yr5+AE1RLr3Tj0CG0BnbheblWqXtpMQuPDzdcadJ+lVVGNPNrzAd+nExgANI5o
yZVqsgWj2ZjI8lJl4+XnvnV+bY8M3L5pLJAvtwIue8btZOt0NcxRYMFKv6AjqMqp9qMXZStboUBf
Jlib11Uge/iFo+xSf1cb9jIUGQ4Cvxg9pCWNnxulZjH76FuvTrW9m+y8vgV4iPvn7W+FLMzbOfzP
q/w5VXIyFzqiCzm2Lu9RXcTWsne+gXD5d/sWcOsXC54OGivHBRhzK1mg+GN7woiQ7IzUCvb8M5gz
XqEa7/srWjzx+2yTrhtTe/0jX9je7bM5jQ9OlIOFJZHIKDxeCUOzsk48EfmXg4UYSYsvjC1qXYM1
Qn/EZuXrSQ7TBYwLMzsydZ1heQ6u7K1MMWHF+Ytdoy+NX9GDEc1dpb/kt8bhoDW14sSHPOAR0gNZ
ar/Jgu+zctAkO9ogy1dkqpIJrIJw1MgnGX3h4UMokrC6XTFELuyQdNQ1eFrsAFAr+vHlHSf4TEed
NMM3d5kqm0n/hsEphuhIQX0j68ObJ+31Di6Q2PGTdhhTgzvQLTyLwbrC9WtRiQgyDNcVUvxutLF3
OXuWlUPUIJlyyPjUnEUQXZT/8lAh7j6ugN1YIjdvzTUXfl0LWR2aiSuw5Lv46RSjw0CMpFPKIzSy
JANTrlRys66UiNtMg+dM9pj94SV5tkOsiSoiGFH7J7OtDdnlqOC1yevb0Dr71SUTGZ3pYtS/iSHg
T8SikkK7rQandtU8w0P0HUPdqpP6fMz7Vy3ZC1dXf+Zt1VoYUij5wWtijlcKTQNkrbQe9dElK/74
UN521aIzh5jkPF44XyKjphvUlZogOz9sStvsZA5Cj+Wmef4xchUBB20bh4FZvExWcPP5/uwejrZI
T57/Yk+FfyJ3L3vvCUeZojFO9M+JTIIulJC2Nk9R/nWrmSu5vEez4Yh13iN34dvSm/5Opho9aCQo
j/i+2/8m/PG6wBflDke83flrM+7ug8y2ElckzLjc/7R7/TX9Wikc9SvPLVsgQtqyUc7j4sTIkQ7Z
roKy3w+9Nt8ogkpztmH+3aP8zV44yJbXGUzCmv62ihEwN0PY0VXIKpjsOxA0h28iaWLMqz0W3+8T
h4jbjLw7BhDagdjcpw1mDdB9BKDrpdu87j4CcDPr6aOVwA6xdRqG+Uab35xS/+7xKsRCF1LDR+FT
qiKFR36UcL3RyF1/w777N4/g67Cr14NjUWkyc5IOghau2LMi7TBSaHORFi9M4B91Hnar4mckPCgO
nlxv4/H+Viikp/638hF1KAtj1UadmyAPAkGfMo/7OgvKqguj4ep8CGgY9wenSFX9skVzBR3qJ6k2
tVpW1iLtqK3KWg6NAX1P8uHz70XU/Ct8rWSvJBqYiG240kcGGIzdjDRQK7t6K/DJKtTf4R30DZHi
XOsBBLZDIALyikoeiWHt+NyMrclBRcDEiUi/cwUuXEEsb5MgJYuXeZG61V4z3BMqDpBShvOL/0bv
jW5i49AFEi8lzZHcY3OoRcX0X/dqOU347N7uLb5N/ctfFVxMcKHKwExA0GV48CdaQkQj425MBUUs
l51aTsWd8JKG+I7+mW7qqwKKanknUz8pawW+c8zvDxMEoFKYNMlK4DFeMcHy44xjoRyGUtUh8Opv
zX2ADUDLLRNzzHKdJuSHLIAQNs8QgjCbpi8o4I1F6egy+FZ2f4UXZqlbOVF1Cn9pY2u0BsHSBKQV
zn16jGTS2fCQdOMhwWBUmu/pWaj4ax8ldW7x1QVmUMIBey3ggE5JBRvMEzc0OKCyt6h5eLty2gO5
xlhY74F2XboDmEBfplldPHdcr88fOpIuINxg5L7qRyEwzjR/nA2HkPPNkauOCqP+0/Bhh8cd0T6V
gEYRlcmrC3lbSXhd2mn3by7HGBw9zUuGQ1j6H1jmA1ng6PkTOHyWjyo17yfxlB/ik2xshWWygeiv
8SrH5RI2biGgH9lXboCFnGLuKEM9VJ+kYnEPmKeDv5Rxdqaw11lk79c+FWwNv+z5IOb66Vk91jvq
GDkL3XpinIGwxJCAtIq7MFKCrBT5vwsv8WlwOm9h4GIvurfoYpOR33F1ZmjbyJJAV1aonxR2SGQ/
xbPXhG/fMF2CVs56yJ+IHpqKAcpxWlXlk0ZGH1+/6D05TZ9sSHKRKoPOu48i0Aw5rue8C6urA3/q
hQNPgmBeyUnXVhxZleiujEj7BL0lDHToBc27M4slAfM5fbRvtUQDQVyjKN33Hy1assPZOiYAQHf/
DWaGARGdBZfoS/nFajKmmFC1bpPcd4OgUtVMirI2JoirlYxcqJ1+rKr/2w0bkGC0J6DchLb5rsTH
r1EbgdRNT7GXn/PWOgdTeM6VQ4VVvQDbx1EwvtRr/RyKV7z+ec89eMBI23IK1+hNN+/tKqsPY0OW
kMmmeYbGbHoqy8Y+WQM46Odkxzodiea/uK2hwJ5545HZPQr+GJw4OqrfLTWxpfahvbw21j5pWGiJ
cbXa/MMbgtY5O8KTyxd3Swa0xXeT/mLojArfgfnBHwFrtr6zk7zMpisy/321IU7+tX+nRJ4wtfKh
tAwehIvExcU9YIPB2ZNAdiM9uyHRuaO3RWoERSRAmBU27AS6HhNJQ7go2nDxfICl8hoMxwwX5SZS
YohAMm6FY3c6HgNdUB0lte3ZPUXonHKOxQ9yICS8ZX47D+eDrfTBbmWtA6v7LE6YBH2KtDJRXj3h
S6q68MyPa9/YiEtexvJ+euTkaKwxmtAa09YYGLdKyf7vZWjdfii3Qfk97djkCIy9AjQ2PzEHrCDm
OelJXrY5fJMQoahp5bz3y0wAlYJV5aczBGas43GSpoCWMx4JC8QXWZ+/cdFiIHKki85rXGwWP8v6
XO24AeJl7dV4QfXZhI+KjhmhS9s1qXyk4p+SfiyuAcZHJs5adxuDixGpr12p52k/6YwN+HEvLaOq
PIvnDIhd4ltcuSI4x12YTyq4V/fXcP1/gBPKOqDE9uMv4BFBHnBO2mrnjTCawQ9MhMYBaVraKXQj
1jHKk4WkvbLPB4eOnIs4EnPL4YRQcfGNtdA3bIsI4TXf9DYYS1KRnM8DrgjxOtpcscJowdayufkN
2sKZ+VxFo9Q9QJQSX7LAW2WTPR8A2Jq3EY6nIfSc2/UHY8kOJKEuAFA7YD0sCa69WKtg1JuCJ27S
HVZIR4McQYj9IKbZEsGn+R3ipqCZQiPbka3yCP35JITvXqWLifGVp7GPWpETF5GceZF5OlUMshaS
sLYfdhG6rlJMBv3/vYM1xD6AEUZASP0O37Tqv9YYBV4yZhavCa+tsglS3kbSf2DM4ayQdaDZ84Yo
wWVqoy6Ciq3zn4t8Blt3EeFs6XiUbwB8JVaiYjdiiSoasr2ZqKdsO9sqikzbvDLD8TQh7Zt8K927
W+OUasEbRuNCnjLsXTI0CU3FGjWnHlBGXYLDdUSqLpfqYUsv8yGwrLcdI97uMWomGY+Bcb+mx4vE
723DX0Nelufrq9ep/Z44ekzYtX5/iodU3dwcwlXPcMaO/qdMDiUum/FRMare/sR37LFA0AetZNXC
2X1IEfWrqy8r6TCO+pMB1OQsnMp6IHd8cNTGY5/H6smDK0U7R/YJqKVmkJsXZUS0zhuzYvCZQh/k
xMsmgwvWPO0XlmKliwmHIIJoXfLqA5I/6eQ9WurkcqGt43uMobrnOXy6AFlbrBsq0wkETetuhkqC
Z7cXz5XJjyI2XTDb47vUeTiw67EBRs3ATjSUvTMBHpWHQ/XOYX84LsGb21gDsdEgr/TfSyxwjzi+
f9sETUt5LVJlWpdrR8ySVaAFmNvtvKLghRI36/Utb7e9v+a9pnVZ13Tf6Xk8rauoFiSHFxBz0KnG
Zx/gfyI1IMZhqmBUTaoGQilrd0N/XNxsmJ9BcceyjGBHA6mEsY0kVearvO9CsqgQf/sOSkbedCbA
pDBx7iEwH/xFWw1CBXmxJ9ND7Nbf67HlgL6BMuTYxo3XwiZ5Qtyvmp39paYk6jyO5z/FG38vQuja
T0os+5QTBHsSyq+UVXQQictF9geUhbrBziqV49XuIyVz4/9AQfo+tfmTa5RprDfHZGnDIKu+/B6e
LV0D8Akkhgi2rd5lBrtx8aFcvVfjs/jUutFh0AnLVqrsUfY9KqMC6lSGCU19uFYb7Xjy7gtZaxlj
tXbmKtKcKNHWVBZkroQkY6XuosPMWXqZ2w+aSmJIcANtkpW/jU12HlDfyyYMFXtGCokectgq7Cgv
iJli67aRRQwdk8QA4u4/+s0eY19HdKSK/KJ9MRHkO6OrySRnir6PsTIKSdmvFPHYkqP6x1FXvsWY
Z9hP1ERl1YHC7c7BvxofCSAp9QHE4+lwK3MM3OFqVOtYEPA0HNBFg/vEBv3DkYq6S/DxSyqSE/Ex
A6kHgHG8ySYga1uPI19wTys5BFpqxzvZMTbIsiXsXJVwn+E2/QHLwjY5AY2Rr4HiYe/8aVc4qz9d
foLRHzHskBT2Fim3p2t4auKjBXU7CfZy4XIrFa13j2PXHWhEmzg1tJ5O8YHsMie4F/Kb1ccI/urq
jVKarnh+LrxASBeNVt8N3rxFFdSsIQrzzmnUDhcRITcoor6Hn/BAZ+4XZLiJmq5HO5i89f1zESKz
fxcTcWIGBY9qmUrfV2re1hgmBPgX4Fk/J+vJsXLfccZBcSt/bA/8g3ecEapTepzBXX2XIKv0/eqB
Ds+sFsDp2lRkPTNk5qxrsqLgpHb/Vw3Tzx6eGzDDqvdXu0j0AAaXXKMZ6I6QlTKirQ9sYIGzaYf5
M20RBEkV0ndAdYyqeWaT2b6bo2Q8wgg1yx6/gwquYo8eHYatGi3ehJfmaq1fDsIitZ0GKiJO0OY4
2LwevwVkOgbyLukWJKhHjy+2W6kEWdt0Dmm9HxZXepav9jX0k8+CLnTP2UPrSN5C/MdB4D0WZP/H
dJrmYqs4WnZ/LeAXFIvI3SvNxMy8ixLDq0mCz91Peub9AuBk9hLTgIfuvrRJ0EaadAdjqKJ79cbQ
hkggogx7DLBY3T67x/WDF5T4JiuwXULqfY7vKvfqIo5DmdCcMAKLu0Vu/6bhMA4jDZGMkyYuCeXc
JR2TFZR2AV444j0XQi5/P2JusSH/4eSZ1tv2Yg7iUL1ZuhzntkwaYV5iXAERFICxH128GIt3ncNV
Qa6uYVdfI/Ssy58sPYJQbGMvxUDK9VeNeUBXJJLDZZHLNIM9JTUh3vE14f4V0yHhH0SxdN6IlCny
riZ7A9m6/CbxXTdUPUfb/OyJy83BNSavwsl5xkTdR//LjQq5H3EfmSFLcmIFsOyV6Xi5G1rpnyR+
l3OcudWv2qfVi++efGZg45O72NbdkpNZeCgPlViYz5re+fQ5ODyJnmFZPLrA1jdER7xK4AOZKSFA
Lr/joOSYs4aamch2o1Ok2/BY+UGpd2l0uKJYMn32Smdk7dh6WMbm1/S5NHMsI9OZSFnxUbFYR45z
AndS+HGFFk1uxjS4oNPhWOxbUI127Nh8WPvNaOZJl/l6E23ldKoxfTvxZdc7JAftDQL6XjkMcHkh
9o5O50G8h2+Vpccm2kB1Y/80UBCWb4koLaC5jWKH4b4mpa3RCV/VYvGqmxfP2QTWHpUKo3b7CGRm
anW/BO+37/E9qZcX8NRbRutSDWxpMxYCfUWjQg42pnSuuaYPvIDAuNxsNapHJExZY8/3bCxLoQka
EeYdB6DHSfScAZhjwz9k2b4UoMrzuKfICuVPR0nqbRHyCvDRzQ4OLKHNIeaYOp0nI2QwiAISpiIc
a6msd/Gdi03a6zAk1WtTSnZBx3l7b+XSN+HIFhueR61XVeksbPwlG97uvxO2qB0qy0v1Z0O4ojbE
Zvil0GkkqMxJ13+B2Nczs5G+3rKv0I0fmihLb9TQybVU/rbYais2CWmhxjL7dElPSw6xC3kjQbGs
bHKNduaBn3DA8pN7KdtrCLV18uABsI15sa1lKgpkVlS3E+sal42BTakvJtGeTw1Aqa+OjtEICd30
n+dG7i3wIBfaRWzCUzXwShUKwkpBnB+ma7Gw/7CoSHyUqf+01wYpe/AA1anufhWqL43Ui81JV6Hb
a42KC13R7cgm0uriOiJvigC6bYdzhqjL4LT759lC4BWG9YUg06VXRhz7oMjo9tfeu+OfeVVTNuJ2
b0pJPBJxRYBDVtkNUo2U+m76WbvemrPR/0iwnsOHeJ9hShdDl4GEtyYY1yTt/ftg4WqhbdOzUeVB
bBv7OtRsBu6x+N2QN3DLaGpY4Fv6/AZ4pOrCZ0gX0UyxV0kI6AkMUa5LgsMHkfhYSbbNGxi5Bzum
7I14M5nQUBu7E7NYVBM07RnuWa45lhX+u7fWztz6trNPGU/nX8jJ4DlXEyAWEQz+cIrYcYe3fAWI
BDFAQXS7wzCjPcU01klJz9ldqzvBqw/onZ3SwKwv5kmE4mjAWTDgVmfUD9XCUQqbajw8ZKkdEXLp
jVYciTuEzB1Pp9CMjpe8bWiXTAACkxJkj5i5BRmafPMyEprnMymU70q9x+bf2xXmeeDLXE5DAhgM
QRssyghunrZcZfbvAi2hRxFBb3u1yDqDEaAIkcOxkeDu6cN6SPbv6PZoi1cv7HcgGJG4kuS2lZJf
bL2uc2p7QoLU1+RsoTgT3MYfvGjT8hOQddmi3wSQN+15b8VKvFZqClW0qK1bxeM5htnYNFYc//9d
YbAuBghmWIGNSKejK1q8aTX+IwZuhyUf8Kzm6RBGhI3jGioHHeiLkqwmSRjfgddbgd+lXeRhm4WC
iQczFAcOWKlFOqtDSGSz1nrudV3Yq/Nz/hoReSyHdMMNthl8043aobpuZTycAM7EzKx/4NUhZNhh
KolUoiyZM4HAEh7IG+dDu/AeO1aHSm7E5XRAREb/Bq8LFPP+b36BPhRd5uqGzqWKXGQlOH7VAk5T
UlgrUTUXDcuf3nrt1zRZaKCxDij5MTZuqKQRRfstTDJCIKqeEERbspMtUdtjgj6pQkRCgldsIbb2
iERLGxIc6u7DMgJxZEojwbj/U9s8aAQ6XraFcQyOr9pIWBheXkvXl0LwDS10ZS+WcNIyeW5kQq+F
Y7jJ+XJuretoNxOVj6sKAxD0/m7B2jSCDZa0IME0jD9Z/OVSDh3ypvV6Om1qyajsModDDfRXphgb
0A10PCnzjxem84bulFr8i6gLVpRvMaW+YyDTxxCJQSFFrnR5MmJJCnuhEjXKIKxsoGVaDH1AkAjT
+/GjmGHREbUzxgL66Y6J8GD7t3K7MY+bp1HxUzkov4W6LE1UXlqz1N6/qiIP1PKNlCJusT+NQCBL
vbAYogThD2w6QG1leluJ7FQgD1JSmy38uGbOC0fjwZS1e8mpKkg+PdBqKeY/DWYAoW6Q5FJw52Ic
ZJ7fQakOKFuS3+kyHssy4uUdCuG3jV+TYqxHeOON4882ycv2gfoYdxYLsY7pPxMTjwO8OYC+D1H7
L7PLNKRGEx6yjJZgj0BkxQg4bSUdqpfimW0pusszAaov984Ifz/5xPVZwACJDKWYV7IAQUbyL05T
4pfrcPr5X/3EJJH2XMlV4lPYnp7JNyCfNy8nXe6h3vl68ZhaQ5gQVR06AU/AlHE2tvu5H4s0czEY
ZnxGAW06E11EII8nU7zQRISpCvs7W72aihN31ul6oZTbIJMLdudRfPk5A8h7TDAMlQJHYW1dkber
331GFLqwTIOI6vLGgQueYIh/SpwsrfMuXPVmSH5zVDivdMM7qMWvOwzjx6U3YbaVicz/eJC/gPy+
B+u61OKW3NIuRKHt7WvWt63NpY3LGVy0nu9Fc6kwSbYHfXZO8XvZNN6qnC2ZKvmkRvSO7IulwSds
t5dY6NCCeXRPd03vJ0JLUbIj5SvD5Lz3Xog2MsR+6iU92U3eeit1kuNjM+0tPpJeYcP/aVLkd6Lc
4Gei1fOREyRa8piWBfgV+HxtDC0fDUehh3s/whQB10Rr0woKeVut3ckkX0pb4/SUs+h1MDtkfD5Y
aFUv71pKZEsBs+j+8l/TNd1RJN/lC0pB1iPEdwO5SNqMV46OhihKt9tt/UQwqAMoFpgaeyyn86Hs
j7o71zqo+y+5hmVNvTBJnSofX3njZ1cG0YUz9Zk/upynhPuEyFyBUcNzGlmMAhA8P2T46LZ9uTcR
GdV1hqLNJVP9XQTfAmDspSMkeUg77Z6CwE6PI7Wou9CaOXDPl8lvkpdu2KNx06D7aUh6jqRFXhVE
L9+uRpXJXp7ITeSgjC+l6SM37F+B2qm0t7uc+CbcKYB51chDZ1aEqAo1SH/b7BdX/y/0p9vyxHNj
ALsNFyvvs/Dt+8+JFYjUS03b9JChiNltiITyYJ+H3vp47Ig4RDT0hxR0GptRfJk987BB3pJII/eW
zrCRfZIJGyF9/Rb+k0ZixbaqQbTJ981NdodKB8O7oM7Rwcsl3avY0KZts/okedFrtI4mvys6B0k4
AVqVEhVwMK37kScFomoyy/hSIlCQ/DST
`protect end_protected
