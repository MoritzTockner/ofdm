-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rhUDL/I/6BBm7Uec2r/aFEHsLQkCmybG19KR9OEHJdjr4evmLZkb0TFobbDoQxDGdlHoANfGAAmv
6A1vxHwcUsAytDkp4OLVHbveB+dsaih9ytEO2nE+hXMEtNbYFk4w0GylsrjNz+xH8RIMUn1Mp4fs
EDzPFkUut3ffEXQBVutyd/5LcTOqGJ+8KyYVGJ2lekMTEkZl2uovZUVwr17l5l8BcHDjr2gXEVkm
G3+m/c92aRKrxaxWDT/vBwCxHmeAHz6NJDJKNQSZpLjdAyFgHTgHvOjmaOdpEgNsAWRrNPC5+y+h
NHQpSf80Fcct7E6INAMGTv9QwYf/pd6rRauFFA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
E2BsRai8Z4TGI5lxNzzIhoj27FKRIMDBDasDk3E2Kqr/cGrVPFMlt8pREi//S30PFvki2S39j75N
5lkCnzMKGGCVcEGDiy1TER6F+uv4Re/KcayDfPQGEZvdQpVjLgd3iLu1ePUhNNplTE/WO+yCNyau
wxTWhSO0brLwUeba88MmuJo6X+iXNOqabdaN/vZ6esSjbzz6ADRVrQn6pxJnztR6yPdgr+7WotSO
eZFO1omIjy4bPRQFDNsUeMgB5QAs0b8fvFTomsmKnGxHuBLy9vO6WBKDfLzCpqX435vssCIqiKKl
PPskEXUgRmTl5cN+NLKL11Wf396EI04GtJev9Voa4ub7sg4wSxwXFdaZW+IvGtQZNaKWdHQvqRmh
P7GiNk6JZQZ6295/S+C9DBgEZgmdvLUWguEVE5A0UhAZVmvJhX6AotwY1EfZz+L+bw0fgt3J7xJh
RcUkXNyGny4v9IIZM+kWgj0ItJrttY/L/0VGdao4Sa7//Xes8mseJvZSwJhBSOeqqMd8CYeKuORk
OHUtNlwEsFy5hnsgHdz8kchNx9F0GZJR8ywi+nfx8tUImYnphdDgWJBLhDn7bf3ikz3+PYLjXLHp
Lg4FFxXTP4IZqbUTs0CJ2whomdCAOC/HVe7pQZ9qoJbIJlNRr0YTHnNP4bsMRJskHiR81KGh7Nlp
pzInmgcYXUkCGXejaI2AO5bFz7BCbolkIR6QgSkbsvAZJ0t7XQuW2gM9FH6Mc35gVkKlBGmMglft
JNRwBZgdjaGoqAHY1xqBEnWfWb/6pQDAfnaKWb3JpVyn6n/AJN4j7J2hiEqUQjbBDng+egU6kem8
tLMUEuOoRYJNSrjlGP7VLL04l5a4QJ6eLkOnLUKsenHf6GNQb6/4+Y11d9ZDBZEcgrRWH5lVUl6M
LfjvIc8wN9AEXD4y5bnf1MbGsHWrGJxgI9xVeiemS4EA7DcfeaT11r0kWn4KaJ6aNOLDEKvgJ2NP
5uNxOHUqXSL+HHqQ32T2eeQkmoqADWXDX6sdFfQgwXEG2GBL1h8YEsKr6lvZvwjniR9tHlmbbl1+
Uf0da8suKwHid2y7xrigfhtiRq4T/excRpaZsV5pJGJTRnJbSGDfPmiTsSlgPPqTjcHqqGGLcC1+
bkxOd+FKN4mPXAANA0RuiHCW2MSpznuLmgUW5ZWd6cO4Zu1T3V9eqUJEa6TcPgO/1BrKGrypN/Tz
cXbIJTW1sRV0UuYsB6UPVoprTijI4BspjPT2VatHyMa42HNX0dS6hGpQNDgwid09UVggzhoHRwCw
+ZUBnpcJSx6KHNEq73m3j8BlKgXrsrmcf6MvsntEXqfWDkhM05koXqyetvg39t5HyceLbHRgED2y
U6hwJVWwN2HSL6NN8MWvlpm0S1IaRK+lM617uR9ZJsY0gudklCm8voJGgBa09mOKhYonbQJDu06x
yoWREI+TBy5k7Oe93vqBm2GA1DPndTMk/8DRFwP9+VgPdZHbQdtDkwKWin2b8I/F7oWJ12D3PUXf
+JsN+hVO6um9Hjk+ws7eM9J7SmDKUaTi8/9CnlSKx9MtZcm92vBO7TiUPLHrQoImdpCIMlmnzeyn
/yhx2fn0PKhO4W9zOEVdazFnoYgt+H+tqz7UaV+QIHPQFBLB6E1l0Pu/RGNtohp/N5heQBLQzV4G
lVQGbyCL4onDVzy9T8Lq/aIbj51bERf3hs1AoWqLzlFOkstds+kx8slFj46oXVY5m6bon8jyj8MH
Jc/PSqFG2eYat2tde+MfC6mgQkOzlkhwkwc6xApgf6DnbHx9nRmGXZxeIBs9k+t10GQl0fxf1nTI
VcuzuGs17GQwtSi3ktGxMwRcwYcTH2Rb8vWfmdp6V6kLr4sMSJdilZG0lH16fCA9gQiDTRJswWnT
bux8yBzz+4KNbIcBEnIt4s7VZVebmaVe0MoA8iFpSuHTxoU6CCQw+/YdTeJWfgfl2PDzgZQNCIxT
Tkao5+Q8XP4AiLj0rVMUh05OqUrHtHuRwNAY1NPP496lBWDSZA1y9dnrsn6UIFV9jJiIYRcHLoaJ
d7PI6P5neAHWixxgsT7L+46vEVuvJ3YK6vyc0IYO9ckOmx8uIS8EluiYWuu5Xwl/at/HSNNYE9by
RMtSWaA6MaC2m8mhp1NrNpM6cWpAMuWqnMok3GeyHBXP/d3CFoXTIW8RXWG0ZA24BhuDIR6TXjUW
LGuURN3qlW6AS/TWXjqUlqlKCSi251ho+PrtLUZUQD3AaOlXtdqx0qgpFN9cjhAKcgCw2+/xxGEA
hJaSYp79OeiVhRTpmfzjyN9kI7a/jG0vb+tZNUx+GDbFUvKfhuXyCvUxwjUDocp29X2unzYtf41W
3tiXLvDE+0/w1TqfQIXmQHgzPCy/JF3F/Zcxn/ZOmTLwF395VLc1149SN3BlacNBoUT4gRMampJQ
2bVKn4/cic//7QpSR/nqJfjmQwcAlsp/1ntU80cNd335KOdttJEtTR7vaDykw4MVtKz+8qKukQ73
uDMKm8qqAQjXwoK3trmpM9J966TWFDn0u+R6SXRKdJQqkKBVfOWZ8yISs7SxZYY8pnVsB+adbPMK
X/0cktG975omr5zrIqm/6yVsp0vlBTZsdMBN5JN6bhlwkcjsCtHBFjJJsJWeyv7jk7lgSxvcr5p8
7oRiijPc/1VGx55QD+ydXnEhr8gluDztTp8eOoJcy62Li47Bt/kPAIdClye+pS4k3N9N7qR5LWb/
a4FlPVNkhugGWn2fvZUrTjI3oK84l89wroyqZR89nsupBAtSOnM9mpG5D+ovfWXzI/N+/em9dAh1
z6CFRAty5LT5GDItfCpR5ewnZiN/O7rCAQtj1gQDXcZhiUE556w7rWICxDFf5KJT/uXdmtsQc4T7
Y3plLHnbWaymzPMxy5rLmIcqt85pLfimXkHnbnCU0tm9UnnVQI7VXpRO3Pz7/nFJF9MwdaYiASmC
0WxKFO1TVBNkQ6n2FohW5IaWOfsr3K7fDZo/5UcrAlngdMFoiVSeaVipva9vB3X0sxN6FpWh9UED
zsp+DLZQUI1Tg0G0OH7EOgrhbvOb3Ykha3gRSVwmbnA22pjbPe73+NLyX7aV+oCpxXRkCtzem1wQ
LPjd1qLgGnl5ZT2WcWSX++CjftRVITOnX4KbdDWmZWSyhPI+2FHKDLhOD8Ily5qDeP7iKonrVOfW
nDSiBH9ew/vbnfiU/xb4Mgyhzzn0CdP6zRCBsMJypXq+7YgtyzwnuqvD2EL35ILMOYsTJa+KIzmT
0Wlv4zm/Bh3c2g2uuKKuHKdnMIpbghQETA0gSv4daq6nj1yruOavsF7Zh8YnfuWHDk1PgndhUTFL
4Y1uAx5+qFG9juW9iU6ta8QzlhH1/7cTiJmanQ1V/YEjV0PFypVPsqLcD5US24nupSjs2zmmz6yJ
OrhPcpoXmoScywa4fWC+c5KYHA3F4Ot6gS9UK2S71Ht7zCQF+1oSdG6Ef+K3STDxPuNs2J6CmZGG
nQeICCvwxCMnRMwJyEyKf/doFTALIuc51yBr778DGUWgzOQJeKmoWxCy+a2K/mV/FZGU/7lTAL6Z
iLxYWIkgaczfti2XTxg/sDoMkN6PmsktJQA70TikmUoviFVSVMy6Xj9mwfIRWITpLEgmnkYepMxX
9BsIgDLASHxlqcf4Oai2ksPx7pFW7B/i6op8HaIQb4XA5NNsWuTFGbkot1ckZ88V5Zbfw0mgkwZs
0QTTob10Ydj3lN8uPs+J6Fyr3WJVPtyQtfRRDLI6niCEfvyro7FDwi6xtiswAm0y0AGYOdgtSGpo
NOqFmMlqavKzy0l48MWE/Mop4Y7sp5m+RLt8V+n9gyBdFmfUA8bTHyXaZMnf7eOH9zf46MbeVzCq
nrSwbKWEMHb4Gt1T54gAhZKSLVsbXs4IxDTKL1jF8lu8kR5PGgyPWG3tJSeRhWo3A8oq3jBaocmh
UyyVMsyXCl8by7N8BScw9//keEiIQ9OxQphC5Yc2OqYDXmd++K++0yJdPdeTLMoHkQlX2jQVMqCu
9iGEBJV8YwcDUlfLPFxZo6yid9pIclj5VrooBdDTLuPHHCa5GQ22rHHuBPUhpzQ4FEzw1D4CU+95
r9AYJKgEzV7HD69cxfpD8anHOpmhCSEZeA1VoAJVt8iym+qVCyn6beKZ0ZyFNn/hGjXCQqWtWnwM
plbSEHxc9+2fowDBNADqZ4+vzFZa1XYBXU2kJaa95EkSvtZl+qcnlWph28NNF1zzblWDBihtjzNd
BqkEIAq7QBU9kleu4KzwyLLy8gIVN6xIOvpG1IW8oAhJqN7pd2SMlnfK0PJTfKt/rnruu11Pee2R
CuD4Kv9p541R8ZtffrrT3cPM/X2m0FSPghqP+5IXBCwylMWtGsqD9EFX5PTOyFw5vC2rMp/eYlqS
0jt9YX4MbF4RLsCvNBajbU7B7Hc+n6NHCfm9xKcTmj0+4EqfKlJ2YaTTGLiwD2h4jL/yFR9NWYwv
ZufEcvfnsgSAnslfuWN+vG09GgkTRNoMDiaHztcyi7p29stSP71SjMme0cG38OA6BjLuBImwiYVe
Ikha0OCl9nrhfIh9YVidsHFZa1yBpxUAq5n2wzd/zH2x2sYLPQ8oRNAVOI5vnLjkHtYBy9R2hOn9
qgdHeGlmp5z+/oLyC7T86xLlaKRssMH9BcGgBUmBhQNBz0QkkGuDgGEHCp0QOFZQP/jNNTDTUCVP
0xLuE+icHeBWgoVXjZGNnXY9EtdvBwsI/bHRD58Ks897vvj4bGEFUOK3Yehfm8xQFrKrYP1/Wjoy
yrlimAtUyuXblddG+BLK/rU3g6tIKWmDnK9OHBoadQImpREXORI2fpPj1/SqQufst0eEm9qCPVYP
8RiSzUIkY4CJKyHY1c7TgbIZSIf5i/vTpwMmwp5IIqfIawPgMuzQmJ00uzJK9jJ3Xf9Zvd8nS8TR
EOnoa74+gDgRG6w8p58uvNp/J0fGmXamVaF2EGAwqlEJFcqVBaznNrwxXUBLGqdLAGwzCSVLFJ0+
iumy7FJ0Ruq04m0G2Awjm7W44H00BGcrsRgnBZJk0i8t61+23IXWto+cfEuIj5/ZtNdTf8SgWU19
5r0ZMqjmW/qEca5h80t4mtPhx8XJmKkJuWomLNVLwYtZXXo/ZfLiNUhMhrP7hyC4Uvbw2afYBgqt
h4UrfaK/M+mxgfRgB3vZykqfIC9IWYvTQ9Q2QpnB8vXKuXSqpfC0fnLDQHZjs+rpqxcB9t1f7h2L
BD3m9xOaDYrBmLHSSCuBPSuzaCbpT+8SdjZDSSGyK01EK448onFeKBfEvF3JCTegaVd0+2PjUeGU
8//AWqvaZteVbls1vq16i08opk3niqHB8OuspECDJBjpRGrfyF5xh7lAUBGC8ebrj1Iftxl7XJig
YesRr/eM03lAiMpX+NtJ9IS9Vzuxey7YCX5PYgZEGoLLoLEs4bCRaQyr5ofDl9Sjciu5MKv/JVc2
pmFCtVguBs8c+2di5lJLj/GbKH2ei/rOFBUtdKqKisd65COBqOC2wyIWXOxtcnsWXuTwkH8gWA0w
lyuZAEC0Su1NDRwHo7PAet8bg73nX7QJT8IYTHZ4N7aNVskL7zIRK2NHvxMLw4U67i2Zf+Ud65pn
0W0ke3/Jsc7Upwuj6I5fVCxJZKQQaE4X4H+0QzipTz+veviWUGvDR4OWs3c/l5DKniPdIki43QK6
NrqF7WFZKypN6kdAKJr+d1OerH2uVV4fjEVbZ5FwFhpUV/hSRZzv6/C/JUiilfn6mBvg7k0GWqHt
qDHbyj+dOadQjAkSiWoZVec1ZESO2xkWxTaRklcDFkT/gOIjHOOsij6nm/g5prPYxGEN421Rg8Mw
D8zBeEgRt2GtbdJGVlSJR+8LKBI13XMRtyw0xbTtJNuoXCZ3A2IGkMG71cJjJS0/8kJXIy95SBRC
Yk94qDbL3g2nEgacW4UrW8CciEbZJ4CdH2qa5n1Np3scxDYZvjFSs2kMa7ozeND+yF3hwK+Mk24q
mIQYPSjTtEPor0hTuTztVNbbSJPdZnkieQQixTVe8fqAsPb2xBIYoW9dbtERQkx8kDGd55Rr4sDh
e5PCeOkaqqilwdw4ffQh70USB5J2U3BD5pl21zbDj+Y2KgMBMEd/3x+1cbiymQJE99EiFcHqbXPR
nvf9k+PUDPvoO/J5ksK45qLhamz9dD6PUd3uXLJlgv/jgkj2Mp+H+8NpdHyyBV9+1ag/+EVGhz0G
jb40in1RS59ZkKenGSBqjp9YcFddHnV3+c669iaGj/gGtkplFaupkMewbXvUCHpo4cBCkQoSY9BK
0ds/WCE6UIHqbKFLoDs3hdknC03vEJ45q8RhM1UNQG4khJ9LyoYH4QHDHsfaXPojuyBJ6bgdS2SG
JIgxSyivfwrVgEaOKU4ukbm/zq32ErFUDlrE9oXulTmfz85NDo1/MVFIrAg4JohfIHudPsrxJZne
JATfUPEUzLfJYXiq1ZXf8GWPXzmmyE8t65Zz2I9xaOT4si2jRSMjzJermUaOOTtQrP9rLw4uEFVp
EXZkcFkqiVVf5O9vFD7WaH+LdnQiIG4sTCzNP7fnXFh2tMDENQGWVSU9u6f3QOIxZPw/D4xMdnLX
XkvhaTigGvWpNRhnr1t8rob8yotYzEyjisQGc8BiYFY4mlVz7UdnvAWOqtWB8W91RdFnDLyF7KX9
AkigXlgZwKjrB789BK9fZDAqKzkdi8vIzSToyDbwRxMrzwK3yGUhPQjs3oAV+UOvELwnqVlqhdMo
h2IPzmLW3Swd26jM0SePL9534byc+hSaD5UFqaAGz6sSszho3MmZS6BSsKgN7jr/ptxnCbnBubt0
PEEc7HaPnnAxemkEE/q45fz5TBxU0Bad2Sw7LDM2rehtbOJwGuzwKpGXaWS049stdEJ+mj6RveNi
Jt27z3WEIssgBZ97a3CJ+HvI3CVSvUYdT/j9AjM7RsT3Jne8QN/eY5EZfHgI5LzQpsnFdq7xo4cF
epoPD0Nl8WuuQpJFehPFc88RIDa0fXc/xpgz6ToKGUf5Oq/n9o3tZlCgs8knEUYr2G3qfEdCkAoB
XG1tJQ366mh69pUTxFDRZIgV4Pqj6VEzr5cq7lmpWriNxOzBqLoN/f1U5IgkiSClnV+1uHyGcIZn
0jTCDHKyo2DSrtisramk2+Sr4S9tBFb7lsezVGr9QhGGFtRgIKGtpti3q7FF+/vnkOPmSCZm+mCE
viP1OEInPaPaLlCjMgcRg3Q1PaQhrqkfLnOv2DmURaoqVEanY6WCi9sjcDt4RXrq6e7fH8ghRDPC
oeYrd2wraxHnq2WO8/W4NhQx+iJk4uAn1gV504rq4mCQd5p/Me4ZQLOwXDBXOBCDXIthZXKodvOZ
+FcoCl7e9PU8rkNWDwZ/LQsFjC9McYIIDCkvX+8yqwD7ZulLfdm9RB3aECJ+ElmAbBGYkpP8x3Ab
gaq33pUxP71upJptBegmMhpWRfxZ0XoNK8Npd4XejaVNiKfPHisxWkhYcSgI5IOjwVEncXUFPTUJ
Dzd+irJFU90qsyKCiafDufab4hAHPYxPNL1smehKcHBjLmMZCPPCbJ0trLqC5br2Jij/afknUjiG
82ALV2Gc7n4eHpLk+hMX6tj2b9J9AmQLSsckGB1NyJxD5QJt2/RQ8IzGpvEAU7tgZG/fnLegLMS5
o3Dwg0ItqLFZgwidtkdcxCTNn0lcE8e4Il/2+izgTR1IKy88CG9X0L62jGtRbvDQ6Sro0amb0B+0
okO3Dcfu8Wr59Q==
`protect end_protected
