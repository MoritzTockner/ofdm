-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K8l2uDBL/WH0yqq/PCO+ktZ9sJwuX8iqrtVlbvg9c6bcUba2IzmdC3sRHB/8wh+PRFsyOwd+kuOb
A6J/anoXE4TaPHuq79XMNW6xkfo+b+0ZxMt13hV73EExsYCQVLw+xWSrbZdnkILGVA3pGyb/IAYQ
oepBqcMExCOUF+MZPzMBElKdRP/tf86r/e46L+K9JHfnJiDmCSdIekiFoElcSdBN4aLerBI3dnMJ
B4t4E3SoLVoSuy/t1OvkyqggSgqe0hv9OxvHjENINNJL2iZwauVqPUpSuhDh166xrrTJyPS7B20a
wLDzW53Rair3254/jjTOMruEmGct1Hj88Ow+nQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124960)
`protect data_block
OYUOvwUjFYcLio70nBPRqk34s46o0Qin9A1IsAJYFqlolU4q//PHRuRsp0eMBU1mGDtZaP4FjRZ7
CMPGIklcfUkKf6HPvcYjJoyhGaFUomvhTEG4OSKx4qwxd/143w9dKknoeqgswur7sQEw44ra3bce
oq+jM8vg/pLmQ62Kd3qhmbhdy1c1WnXqNe0TfuzMsLFSivv9ZtHRTMKr9iS++osjUsfmHfevOLZb
5YNVoxzniTh4hcGAJm/rAxjJt3QOUDKHw5fCNl/CFfHsGgSGU3mZLy33rErSBwRGJOGEm8V/K2dQ
Cq3Q0RcvBfkBzGilNN6agIt+smBGPeBESKBllpuXxMo8QN0cqGNzjB9+eoIh1Rk4Coa3tzT2rBnd
C3+o515+onyg0ju23Sg4fNfNC5ZlU4gh9iqg+OJDi3qbUadgWq2MBFqOnUYHJDvEUxAEf4xPngGf
XZk6XKT2FJXHbfJrPtBjSKAUGgnGYi0NJFAGYgCku42ZXJOpHVDPuhRf+X9Y+QwYGbl+gPVaQRqV
MZ4aHWdW2x7u4BJV7KzyKAYpLepEFMlgw2XP45pgcS0/7lR/DVdjNK55hcm8fn0NLWtyBoQW7+an
V8NG7RwX0BilEF8WhWS3BTja3PGe5HT5pDZ6cpuQRaMWsTN13okc61ZwpgB6dkxq+xhUW8z4sAjI
vQmtNVm2XS/gG+iGCzmhITIpK+ODK11hjS2bb1t25zx8N2EItGE526PzkAr/Tcsj3iGLZru70RAz
L4uzUqacyCg3DPSbh3gZeCeaFs4qa7I+9nF2wkY96wvVPuxVdihO8mgkIm8xzIinJdCF8e6PhMgn
t4ElnB1P1melDS7kqBOWo+8d+AmiTEVjIyM+gFBOQGgLfUAuS4/CUrFEn160W99Il6ITb1Nw3U8h
1t7kQXRc7nGMX/BiFOo6A/ifGh/Us6DaRODgJJLIX+1mkhWx7w1k2RPEHHtpWmLywh4IVMOVcB2B
qWiP1yZcFSGgdqTmgyU4DgD26xi2QQnPDUmzI2tEJpzsToTKiOzOkaF6bD6sAM7T4+LTIwJ2Fm+i
aDDZHt263pU9xcJv+8yVD9g2Ie65qfd1ToTxyMBQteyjRPqYSQ2P3VeX6DGoFeaQVgKYuDQhytmF
/m/3vOxi5aLfwdAgTDgjcHCCRwBLjB6mEJzdOmRVH+5N7jTPletjEWhnblTccGbJY8by4MKM8M9m
ucWFWsAI17006pl51cF/QzcW7+2NXLY3l8eTMcLaWj050sJSr0Nk/4YERzt1V8FnK3LuPOmTQYMh
Z6QFJHAkihYa1wRGOyw4a50jGrVavPzpU2LCSUg7eWOFPKVfaOXuwXI4Wdg1gv9CfL7L+RM6eZ6t
P5WsBhais7humvCFbGMhmXC7G6x616LMCtZpseu7eqYr6b9FacXzc14dTCoCzagKtiAs6FnDJae2
IIP22iDrxHFDRabKftFE0azHz6LIYRkGuzl47qNGj5ceL/qryNlYr4NJHTDQu0QDYgrE4y+IfhqM
wXwgfIrc+QyGSYVi7u+q4CxoCe8EYRgirbk8gJ2S/cP4tET4cq8t3y2CHW/s+PIUnfdmcg3pxy6I
dVPo8LuaBx2/nnMJ7p9lNqdXD1FbzEfRjf7ipNSmKzYx8Pt1c0lnaHRmzAgR1ZI92B0FQh28KOdu
cpOcGMczuZDPSsa2JYRfu8Y51aoWN5YZJh9EIQ6vY7KyUie4joo6yXuGSr+xaU5JJAp926u95+/f
SZldF3f+83FECb1v+txg9KsoTZzGkTbbAvxQMoUKnx3sV8S/ddBvPgrhA/n9JP12Q+2GmfMKqocx
SSmo9q2EppZhqjWSF0MZNt55CMDCY18W4Vj+u/8mYvkbjeUPt970jhKGLnfSyBibo+7wZIkHqo9+
LQEbmYOu03SU0F8VF2stG95ViGYIiW1Jz8QH4vvutQRXXtxwG/wrLwOc/XtJUS4JHrgIv49P6Yo2
LGTxR4hh0iMAx2xv+IeOip1IHgTlffsNrtxO0d1h7auSwuneSiZEaBnsyOCu2jIqVKMIKGJhbuHC
rKEsvcJtbDH6eJqIUBuQX0L2DN+KT99ZFaKU1PF62TaXPo9DCzK2gmJMrHYlrII1WotP9geZV14m
Tp/QBQpn+/FSaEvuuEdAwUsAiCbgiNCnBx8QFcqSfGGzXevfwLAhSebbE/bYlzvp/jkXS6Ot1x/H
7qAZl1Asp9VWCZDfhILTDckfFkf5u+IhEKGGzyh1Ugn+UQhUtSpOVJ928liBlzA5AasYFE1nzlxs
YsJXCDN6ppxZftBZpjdXaqb10zaHHIoXXAT3V0cCc6sHiWViJFALvJVpoWSsAhrGisikFYVES/kt
SLu6VwmteRRzAlG3aJ9tN1aAMl83LCVpgJAyWsfin7UzaDIc4BjJ5563y4MmUH7PZsDJmSszC6St
tydjBKH0Gu2kkFH/cp6WgJt9Zbl4qXkN8IE1G2TRNgoHgjv7KRF1elvz/bgAuevJsxqbMsWBBcl0
sqITMMI8a3tXoHPSoUpRs+aqEQpSgnk0hpX9nN7fJw4Q3Flo7bHcz9wqamSxIlCWSL6NM2HoYqLZ
6btPh0aVmXG2Xm1EHZLGIR2rynWa2fbrsK0sv9G14c1uOJSkqFRAZXs+4ZeaJAw3jL+E1O7t6L90
10jfZM7iLOyv5e6pMtUlfoCPdk3Anzx5IsVtnEN+NSx9hJIPStMCWkC1TvF08KQw4TUYYGQh111C
6C4N1/rVwsDyW1wbiOq3uOr35xtK3l7/dN2F5oLJDKlPt6TeADeUf3d8ZejMSyLQD0hzv6SIscBD
2S7NYGXy1zMy/qUhuQua5fU5C8538Bblx7cNsv5hXZ38Nn0ijXwxxumrZKeprz5SxjbNK3oLN8Sj
uVrxBC//GkaOSTduUk+vWEZ4W3enSX6W3lA4l4GLo+pTD25dWo0X9XQIqG5G2eLnb5AqxYx87BDy
F4BlqIcTjZMgYa47TD9fpth502OzPXl0dhKAkImRy4k/9dRcqWZNe9ynoq+yZh9CIsP3k5huURZA
jOqtBaZu6ZXSiFEMaQtWGMxrVc6fTyJkb5/WjeidsL6Ixs3f7rCUHmqbvnE495+sKwYjM0ScnlVa
ZjoBa8h7M9VRSBcoH8SPP7DqIwJTUe01Xpsmw92tv6otr4zwzuoZFT4R0tZ1UC8EZBtoRWgegoHv
ss7ey53DkScvAIGi3CoRLGSGthjVGTXEfwuvNTKCF5p12bSaPgOnHD66SSHfjiiKOijXwcoHLkty
wH6M4+X5YkoIcFNYRFVLZGGjPxXKLP/pk7RXDHR4QuSrPEHR5ytCyHxrcS01WCQt2nibj57iO1Rl
Ejqj9Uc2cBdKRyFjvOXo69/OHnkVErniWb8w1/UdUE2wEEr+Gg9xKvCHRO9vfz14kiTkDJj5gYLt
2+hOYXebluMZ8G5uG8Swju1f7lKB90dBOSZ+cUiRRx6wzt79hNxOZbQPfWXc83+gRfx3ILY+lmJE
MAWv/wO6yluNobQSUC5zUiCvmKdqMny4UR6TWbcdknz84XlzSlfiXVH2qJc5lLNc+bg0HZXpoh/4
fMyHJhOqsCHI2aTrmuVj6ltBT8Kc+t5jk9CdDOIeC7L6CEUUm3qe7L2IFxFErY0Hl0otRkT2bu4Y
W/OW9gnSCHe+gPYyaCf7LlwDzTX3Rw5Zotq0qyboHOlXAoeXcrtoQa4LicSDV1R3i1Cfn0NCMiap
O4xX0gEksR8kIrF8kJadH4CYleaKv3L3kRxOZxOFPWEjoiyx4JL/wd8S5LpFj1vhozf5I/ATYQ59
7HsbDBwnZ7noIJtfkI+Zk21cAo9UJKIokqqC2hhsmXXSRVCxYStFLToFZK6TCcpo0+Z4PYPW63zc
NkZVGSd6BH+H78QqMvOXEAJiLWYSzGNNbx5wuQuwu/2z3XlayOdbV0tBdGKHC4PCgHhMJd7zlRTI
XUEmyBjGWwOVKfxGUTeOH9FTuwWqO+SZ1N8rlcNXwOn/34pN96ykEUoPBcF5qWbDuqrUVgQCMXzW
gEk4H4Ahunja1+Btvjbj0mTb7GdRbduBr+8c5UYHD4Jb76ZQoy5PFDF+5WS7lf+3u14cVjOtjKRL
Y8X5COstCHski9obrzL2NUXh5cPtW7nqQF9mz+dt37l2Lyamf67wcfCQzZ1wMKGZvcKjAKHPKUs5
GHueUF6+TROEt4+BLb49L1YbQiIe/632w8j4Uee/iUH2ETBjZSdGN91ZIxQuAXAHmej62FL2grr0
n3hnvmvBraYVENne6DLI6JGiOTg3VBsC3lDg8CrergGRQDpv5NxBcUo92nCRw2QF/6GaefYRIgEc
FRIGOEy2ayE9Po/cUeazPtDFsHS3htRB3ViTYb/y1VilLH+wQv7x/nxibVcuzRbY0XstWj1LOhZe
tt4t73c+lG42dhX6HejtWaz5tu+bf3Cxk+8iQ2r2tD/q8lmZGlTXiz6dAIDuhg1d+/y89chfBwzb
K7EqcUhEmMdhLOsxlt4GGBmqgv9VGKhf2oP4VlvSlRW2tbdKJyZOaDy1fxeYnX30q3U5VBBGBrzh
znq2zFIR8fdo0gdy7bug+qwfwDSqX31GI1gtqWYLgn2x4lImv0sPi7eyA3Mh46eoW891KGShcc7m
NWRvymi8TBCV418F1BfXHHKxyJddulDH7/Fe17EGDuR0M/YUIv5Vryr5DZGC/2oiKyCzkkG8+BWI
o19syc40seDDpUBVuaqwzIqcaFGyxQ+Fao2YmESqrj4gzIgwRZCfCmcILJy5OOJXPzeyegiVR9Wn
WlwCXnT1TQtiXsFT0eRzcvOQs7RVjFSYyJ/dNn6B+KODSPUOUDhDo/2mdquPL8HFDEQYGlJyZHcV
dq1mkwpwMZgbdc7qJZGcMmV0sf0QvDsyTAllulHEWKWGA7NH9URFEmnXAsJGNEvbULLVQ1fnw6VE
MMlfOLkH4rHmiN/+NbWfWjPu8k8yTGc087P6gWxWMX443kBIKkOF1BBITireQae0K86aLNKqMqXD
SFw5W6drdzLWTbQqeZCCS/IYtpKDni83cPz07WsWl+5wYEZzjjnBFQKSyokc5pzMcywSB0A/KNMK
ib1HG3HnvVKbrCoa9TJDYtIjneCYTghdlQoJKDdC4AZAEGHYw8ly9z4eFXEmZeUPBfPHVwzynRh3
cSZIrJxCGI/fJZhJUaZFnOq08c0ZKUbfdda8OHFDtSAT2XMEyVVl4DsN85TnC5l5maPzIVdHXiwc
ZZRk/c4mIM390pXM+iKoKFsUChhdL25vtFHy3xCRgzl5kc59ddGk3nrawChfPXySoHdY7n9YMdN+
Lbh64e7rwXBL6sfBvvkZXws6xv97tqjczGCxGne6+IzFMjRNq4FGRIXX53FTd9GN1rt6GpkPlAwk
M02j6MnASj7yTYIss/cFJ8PUG1fXuEFvqsNeqnnJ9/UfV1jwNTxqgVCJ41nlux4w/6iE74ZvFFOT
bwtPuqg648KAwTGCXfhVT/lwC77zkLTcQIQObqIrJ6HAohWnveSrj8+0LtSnXXESBlfbsojx/rtG
D3pNxddGn/pMAHXR9mhcvNIZNfpyk9m9CLVkYem8nc9lhgpWn5W8fMoC/eXsATpNl/saRec1GFU1
2dewXNnedbO9CF73Gasvec8XA6xQmn//KSiI9Wcj6m+57fHNlqtPtlbXxCe8XP2PTbQ8jFy06kMr
jj/ZfUmBHD/8vwf7mJGr9kcvajLKeXoIbW9vy3I8OFjYm8qFlS4xjWDJjTtvMcdeMqiQc81X3wTG
C2J/fpdaqtBCrmncMCRFINSCxGP3pAs/+via7ftI1qwqpYhxX8KOxhWOjAR1OX1KDDc6rl0qlfdt
uOsAA/ya/d0ji7hPqFDwl6M3l1x/WC6DaAu30IdO6lyoCP1TddNNbdbG99wu53K5X0YxACFxZ10L
D13Ysuw/Yqj+HjRqU3Akl+QDN1gbhiXsGqMYBMbBq0efpITvdbbJ5SAwWqu60FaUbQD+AE7r/6ml
20mJv4bmbOuVVpxZUd0ECnPDcZX+CNRqqfyDhNY0a9F/lnlQEKaHUXIUpRwvbN/aTqe2GuV/i/V9
j1XFk9Jh+5J3VeN+fzbZxEdnAPK/GmN5B+lcke9tzYHKcF1+UCLNENEAMQm3U3eTeRo+k+AjPw6G
t9FZSA14GyTEGsevR8h8iUpCnyGeyoic4t153z5xY+aXrDPuwCGjCSj7tH97GnmlHB9YH01lNbV9
6J2W+zp2YwMP1AOLoFk1fwB25uNHlMxE4RpvHgw7YaMTvEwk3J8FhUmkWm+R2kw6d782C3sW2F/P
ibiHNOQXTsQZnz2p0q8CMI8oWwKPTAL2dvbyNwF6U5QGBhyKBLLTRHD8kU1k1l6ZpOXxL1QRLGJT
hpmt0qM7oOzqHFL+qByZ+5exFvBd6FI83wICsLF8sIF4i3/jLxZ/Ot+Tl+fMa8x+aVFDlPgH+axy
vDQuF0ULi4DIxl8qtpPT6IS7UbUhOu2ITcN7pAEiXyeLOQPaCA9Zd1PjW/PaZtLpvt6b9Mh9MPYv
yARwc57Hd58ZCPBMfeFmmTDTEeshBKwKo0BbGTN1TnWL2sfkDXjQ4pMnGGuhH/z+w0ZOS96hQ0Og
lFEMW8df7gIvarDeOmwO1BJm0jI2I85TN0Bl0XOL+zenlqnDxLwLbJiJuzW/jyhGc0VqFCZrtIku
3JccPAGl61RxgmKjPYxnkxRw1puLuDTbzSNpt8+IwslNkwcqRHkg8UMzanckgQw6H9fthh9zAvLC
0RxZap8Iguw3FqiY8zQ8q0x2mBw2WJxmtzZ4UhgiVaC9eIup6U3oj5w8aw5eK/GJWjZ7gBlr/ocZ
lull8su6HQbqu+8TUALQo38hFdd9epHORkjOqhwnhuDH6hKByb5m6G/yPrqT9j5byMg5N3/xHo9+
4OLkEpY79LHI7bhFksDnR9xVQMNRmed5udZBwjsBOqJCCvc2UoW301NlolCrUmbUoEqpjIjIMF2e
PKPYKucjj2CdB3yglIEnPXOIqZZR5A+ejwGE2nXnPgZErhLFVSOm5/z+Eiu5aAmbezD+/RoCcYEg
IdOLZCCcG+zL3zBsZuHuUYMxZ5MaLgJhdnW3O6SUk52A4M/9W0iEzb1oomAKtgk20JXmxLVFATJh
+OqyZiB1M6uyZD9XfIgIBtAguWtRBx2nWjd8zocUTceKMvGNpIZmduxIcXHd6WpzNsJVgmoQp19O
1Gg1qv4p34u2Lw9lK9xTVt3OVExRGY9RRc0OoYSxuBSOmgauiDw/cntHfYj/ca3HZ3igKgBSF2wy
UmfUNnKEZJ1aFU2dUx9PSiurBuHrcyMgmWiAI2WRQje01HLzuPevSgFc4J1rGnKUkHvx3tXlq/M9
cGMFUSCXgVaWAI2fKrvoEMsCrG5rvllPIe1PKI6Ay6VQyvHk1uBAIgG1mrpDXeVl9h9i8JiBRn19
u9Z+Lnshgh0Y8CBeWJE7+OPKplPkAZUu4k8XkI8NndEmJg26CU94a9//6DPb2eSLTtLmE4HUf6ih
ldAwXb7MM7E/COrqywmJpBOSAa49G+3CaT1MgqithX4MqJzFwH4eHuX4YVs59HKPq/Dm3HakuRh6
tWiKVy73VlEmgrhflN00gbnwyC5lSawOZ0Iuznn0+mXshwnrUjH/XEHp9OMbyqKWEx0zftgveThQ
9f+eXmj2Q85ZOlGrWaXjRPPy+pRvPFb0MY6SQyXRJLOPTvyh1a+CUJSTYN2ycniboyTkpP/arUkn
/XENj3s6W52RChlwFIVGBcd1HdAaqOK/+68JHmvxl2qYN3CJ3Qo3NLH8CH0XekE+JncA7EpsT5OZ
wPTp9qjnuxgISX9O7RU0vyJJ1SHRBpYbSWTebQCIy+TXDWGfVo7aqDOoZSQZ/UkRo/bAwyIXDnPE
0H4Vi9ZO2IBRqv0xXfHrBP3ivSlrTa4FvMzR0kFVyxzd8TyMG/m6IVxRDxHCkZ/oSwebTErZWXRY
X8REaAU1N2Y6pAijDFC9s8Xz7IeJieYNVf/MQEjCK5C/gha9O3lLBB4cMo6mOmO5xLWhgaxrFVwX
4li8MEtabQqzuG9bsFTtMJ3G2EGIQOsboKF9tnIA7S51DhhZeN+Um0pGlAHQcniSHGwgekX+bGoM
RZ1CbFLkUqyK5VzawOFHd7YVoAzqyXplk36Q9kMuaNRVPRaBRm+Mv0Tr0Ug+QIUkwQCP19NeW7ZG
jzYAgRF7oO3bLEF4Bx/pRdJRLUNK+YCm819ch2Th3ZE+Fu9LH5XFaVb2IxCm0vKLJQYr0GcIpFrs
h6RZxzl73fh2RnL8pGhfF0+SvxTKWe/0eVRDAUedivRquFYzfnFMSWvfBk5+BU3edudEclaRrFMq
fvq6TLZw8pcJns4tL/wTXu7VM8gUNa0NKuuZCEejB+bLL2pSXK02OiIvDYMzFNci1NKeFAqQZMeg
d51RZKD3JdvExY0sUdIlyvl+vsFVmmTtZCMZHNoAMrIHRsvc3Q4AqEmXMcsj/Mb77QTtqgf+RMtY
/2i6yVqHsTN/tM5xWTxAHl3EhGlw+geKKRTSMMoh7D3tKpZLrVS240DRdHuwFGVeh+CrnnYGui7M
OKB+QvbLQWI+fRUCH6V5JEDAmwzY+eefWKRrBWwvt+QiMVduG/DOtDpOQGp+VNjT1z0m6z+qjxTG
i//4jma6qjfSZf4/tcTATa33Iuh6m/2CJpvTpDUxh4hk5NoZqk8vNZN8J6t4K0OuzfN38J14Z9wi
elUTJK3HUAHZv+MkYNFImc0qisbBy9NzD+ODJ7d2JClfE78LWO5A2/oyR6dZzya5KFchrxLUnXvm
UJfiBHz7Wx/yVBa8fcoF1/+aEO+fQ0InH8a3gCUPLimuxQ3OQqMqq9NrrctC0ixyXO7uciYxPRA9
en0V8Sr36Z5DA9x188a+BK4lZgXS8390yDNF/xsKgkPZp7Vsev+YuJnISH4R6YBi6uYWZFnkxt+C
Bk9k8iYJLFes9IKxSETiTJbtQCeYYvPWLe2eVevVq5DqYrLy0p2k9LYbGvU+STDqxlAhR35dbZN4
o9r7T0vSmLUxp5jQsl248wz+Nr256xkXfKm6viDWDAC3HikELl2xSw71tunoRN9bziYempfjyg1A
YZzYX6wPMeF4iUxmRhHXzuIwEdIejLuAqVGdcQZkaWiEJatTLtxD2+Gt1qIsawfmJtq9y0F6xRAo
PrvejnaX6ZiTYc13BBmGDA4QnX33EplmPkr9SrpaDHoJBWpxDgWOctLnoru/cfZoZEusxoya60ec
oZ09eMwaCnHhIfduSC8sWlzcuBDDuyJS8fxu1LALKgC34W7gw7rIMKHBecRdxYlPiidELzJtfoKG
GYDROvXenvOEEnXejcIr+D1afbMSacDU74l/XPDtVGulpxULWaOGpmXj03AKSvk1kwCy+BCvaPOP
yMdZNyvJiRXYhhm3rtKv0CQU2Wduy9ZoWzKUv5i0+4W/eJ1AVE81Nb0dmn0hDdD/DTnLL4yUBmSb
9oE6O1eoEw8A3kNl9Xp4VOryiSH5r2P89fNQmiCY2H0bbH9tliyGvPR6U4vRgbK7n1pahDhTiAF9
RWWGJonG0Xob4khDhEDf+dBTJiM94kBwRy6XZahTFMwAy9rqbd5yqV/zKmnrScCX0iaEQRgEbjzV
A0kfZLdQfsHL9uxZI7cb99Jj1GQJEuQQKDPAQJTKxwnQpAVvbUq9gY5U/vvwouhafT7ihCuZs19f
HCITVTIMceAjKRmMR9leazY6ZBC4SA1xoqiNq7hZR19rvwvg4DJYyYpDEH8VhhismfCy4jO8asOl
7PPKB1ONu/QyLKv/53cUwbCPacMMHzrk+ApnHN28bFTJrwpIqtN39m2FfM8DiQ1/FeIbzTe3x8e4
M2ptMKlB9B8oUdacERUU7qoGCupbO1WSUYiy84tLXqIJsK3I7hxiFDSF6dqm35BvcvudL6gTpV/Q
LNH1+E6qgGXRUsxYOS/+Wxtj0/MgO+gi79cDZD310Rm2GdzLktK1S9Pq0cKTbAZIocE5gSwc5u1I
qwenyrG7ycrHoGESSK8MNrGmOYLoDcmCisINntJ8XxTyZrg6DZAdpWUZUmOD0eC7nHsd7CBhgG61
ToR5ol0QQ2iiJM+UM5uhFy/3o1XmS+c1CDrPSQIXE01oI1RZhWsYmBHrVhmjEbWcgWUQoKQOSV7y
a7TRkx4olNekZYinv8Jdo0xiGVy4eCqdf7vtrnpJSFKb/JaZu5G8skRqMdg8IYIHK4QCTOKCkVjl
iGTyo5r99HaBKg0x9+66nJJFqXZCkuKenCwPFXIHPheZmE2amBnzrr2LuhgEEjfOWKXd94dhbIR6
9EJPMTuclBCmRSEDfurzMV+DH1XHhfLxMIx63wHRBhavtiOxUmLNHsBKVraPqEYj8RXsl1biBlQt
h60g49k7QAadpG3lvbqxgHewqNpOGukOCc74Qwnx9+D3TK/rlruU67bzMFtDkL90SWDYUhU66eQZ
gBh1pzLGWgghq5x/y1O8whZo75gP7i8DK+tX6hs/O0qAW6QeG8nL7azEXyR8YN0NKdqwcs6NSTTj
PcrY/oiWOkPfShQ+lFdqjA8yxGbhvUyoYaAG7dn8hFf/vZZoACjrOOT3VS+iZSHQpOfUqYn8w2MT
ggdVVk6zn6ZG7+MzAIUQOVoBqReXanzFqFVarUoVDSWH5gazRiEnr1meOdwZRUc1sJmNExrd8HCZ
2qXRCBB7g9E5V+UcD/oZO1GWJURJaFlJhK1iJv7zjM4zSE1NTQl+XQXriSSDMZQl14d2G0RoUHRy
4FXXqt+B0WhD/MccWgPfBzKCrSN0cRIqpQM3KMKvaD9om3TQtmDcgy6XQismBhrN/LPIbr0IUc0E
DS6XUA10tXmV/bKfi+8mFOdt3Jg1fKyJ18lXJeQ7vkgs9/oZwMocc+SRjnMkUgUUxOzFrSBtA+J9
852Ju+sqfr6+1h1oQRDKyTcOttsuQYEsGH1YwdAxSXrzYMBVW7OQpCX2RGrL+StR4b7QYwbEXqdb
lAJrfjsCJ09qm/X14ErJPGAsV17HTfb6Mk+ABPo+6b1+UiRZo5ijJ4/XuZYyduMQipwqt5pVvke1
r1tWnI3+IYkwS0dNYWwvzdy52hIZ+IC/iyYWysQNDG9DtKgl1ycTSmZrt6PHmL1JD+W6K92qxHyg
pcgO3VoJrmVCmzzve8dESkaB1VuobZBRXYjgPOCMwJmHMLVFms/4B6kGjBZ+EmhJcb7JHQLnWTjM
EYbab7Yeu03WLWHGjFdwMHegWoIzluARCKhzwjGV9418zwmt87wQHLLrECkM1UpaOgFxoBVdqbW+
aAdnmorD59kBHi2ofCnLTk0t8Kk/3dhrNDAfrXUL+8QI8NfT3GD7LE+cdcwX32XT3ZCpOk6o+4qP
FV5J3ZDtSRvfRppgUhrTvEaXNlCgN9DgV/coJ/JFvgbGczcDx9TYqMYZUjZpdQ/WNhmW+6UDDPsX
XmYsKmAwzh1EW9EktKIaJeuTNgQL0RwTv5xIDrZyMf/3uR+3yjbiQSRIgpplbFRFL3k/qj9KuUTc
7FcbCWxH9tHjl4wmcGWGEzABv850YL9zYnluNjmqE1Cz2rAkNkkFbF12mU9fAQN51l+nXkZIyxZD
uPDvSrXH+MYKQc45f7UqVbI0hOAB3hKvkois2x3WnwIKf9R2q29fUpj2JBJ0Vfzz88oiWahLQvE2
tn3VkkjwqIuGLbc1PBnFkj5JTTgXEjhn/VpPiwCHRcXFpetC6H5GD75mgoou0CseWwwmeqE3+8iD
eNfxhrAUGLX78ckcUdo9TBFoqI26WJrInemOTRhyz9uLJYsO3ED1aMlpSxZCNC5n80hHye7kmedG
Mfr9OUmpN68f7h+Jb/ylag2cBHxIVhYZdaLSNn55Y4dOaMi0a17ox6xnDpg8lagD2E6f4aMQXrCh
5cF6mrelzAQc0/e3M0kYQtzr69Ied8qMvoPiIAeHgOQ2TERU6bPIJzUbZeVfrgDDumEf349cXU2S
Ztq+Fstj+gFELiTwresBOq40UeuyT/wELdeZgKufdhfJFynr0DlQ8xL5FSN8h8yaulBajuwh6V9R
o9EF3M2K7TJ1U15vTjeGwaan6ebouPazMprVVzbhqbHOkT5gJ+YdVeALzIz+zhq7Wj+TWYLA1tuc
KYM6Dcsqt06HG9vqtFlfvrHtKrvpbxLQOPmI65Ay3MayiNBU28kv8bJpNQvLu9yMHJN90iW9S+WP
69SbVRnjAe+HhmtGnZ4eM90+AuhVQjBbOpa9a8xVehQsJ/wqMEVG75JiFe5DH8w1kv3AwTe6KoOM
7Z498Sf/Zd/v8h9uwzhfD36n7+6GCSngoD2A5sK+PuXnJhxfyz3oLrONmJkklZHrXJsdEIfqf6NQ
/dFe8edrTTKPdzb2bJQ3SiOA/DWCrRBWJTr+Cd2ZhXYuPzlLVq6Q0HzsIlVkNzq5+YkUx5GR1KwL
M7PoFPT2CmkXUtFpQGD4RPtg2vqj5p0QrqCFtIVEj85SxsrtMKFE+YY2RIcMx9nosWJgBuiny0+M
Xpch9emVt3OI98LP+1DUuA3wni3XHILtnX+ZgAGfyS6/fEMM4zIP0Gn0B+z3rHhJdj3fq/Q8Aead
AFhLzc/wNGA6GKns902A980Pj6CoN0Q94A3EV+xVudhCZ7gUaTrAN5G1+BjUAZvnegHR88jXqXqp
bDFbpM6hVlBj5t34xGyVmik/69b4zTVzKdGwbWmMIpeORkxX3BeQCRUrDQIJiyjfDIrwB4nEnkqz
K9QfajzWSu1RSqOMyY8v+I2gGEMSaWsekBJVOUwbi08TYyKo11U5IgMYYeLLIPFu3futk95dQQV2
XkddeZDdviDG8ZQDAsvsw9mhPZYEoRwRkURPsrzbIzDB5hX+dEZgkYmNI97KZb3c3vejAQYixW6B
yu4BHsU/ubz7ZRIhIo3eYKaZcD2KccQJM16sUHly5/Qvm7LB3ws3M5gU9f9ptuLtVH27ZhOi/l/o
o7ndREilJVog9o755XU9YodBFRekg82++jb1yUdq1uUAZoqA1310J5zc9GCdlUnGtZKX2B8JSRWQ
q+s5HcMAofOVomB0jKvbZi3YFPHsCwzQydYiFYxCMt4vvi04E4ejmAY8kIzo34eYFc4JkmtH7Boh
Jx5AmJhiNBurzZ0OIK6//3djKBoaTFk2PJsJUvkP3uIv93TqhDmeVhmu8cl36QGfMqYUL0oLVJC4
OQfddmmhH3RM8oGdjxkG0aeZSP+vJaf5D0+mxKRu1weHobWpkvd6U9e3K6zoTaNVxkgzyhluVOEG
eeZsk4p0rKO03oSvP3+H8hByr1ZcFN1XOM6x/I9eTdkB4JaR2b4TOjHHIBBRPnfP+yk2L4YowHUf
uktTngC9m7JlNI02dvSHZBqQoEA68WrOCaZU8eibmQ//osZxwRG6GzgVyrKojn6QEbHI7XeWqlXM
wa6bI/SxmBVYcCDetLq5xikjqPJdW8n4mDHVXztO/Jb/bamuV+lJMjxGBnPAo7CYm+5ntNXmiDuj
XoEWNsc/HygmTX5gT+2ytbnTSllMzz2xZWKGEpjhhXElvihf05EWCUAKW8VNE7NzmOXfydM01s7L
sVzrZivAPcmTKWjRzbfeIO33/GMOTi8G5eUHAZDEHQlw0Ggy49bmKMYL8LKT38Ux3Mat96SoKrSh
Bmmq3G/sPFvKramipsnsr9Ku1bf/sNGjXLZQ3fYA3zmVHiOpIv1H0iOVS5VTRGGQs+B25xtZMbT7
m1dX5n646w9PcUbC/m3o54jr9/+alZ1ELEZPmCTzPUYDTnm2+s8zpY+oNPzm+l7RooVIDrT5qv1U
by8akHKn4HGXTMcE2pwZZyPhWNzE5MRQ1mdBfg7yuN/Tcbau1zWK4drRqy3GRWOw9+L81BRn+Obb
4rsFRkrxaS0WhO+wKpr/af7VkeCnqza2Y0s9mkizxqJinjMYGmhh7lH9WaQkZ4V0/LbUlbqlj3e3
wnCKpdFnMFtZPfCocU5fqD3OSKSOuenV/3FWjrcqmrEW+Su/d4VsDNzimDLHc5jU2YwSE+C1P4D+
wNLtVazIBxKBR9IGCD5HeH1C4CwmZxeVu2UtexsNDi1cjQMIpqfUHe4hIhuO7NtQbmrB3iEgzBq0
ELndTWAFmo86Vyp4+/RqFBpfi3Cm8DAHuWNsXjB8BpTkSoxsg/G6OzI4A9vF0oiIM+VcKh0T4MTt
R4e7iXYORbi0j180jwpzzO09CMNKQBN6VNnygPS4K2YGsWatPOaglR4qJLC6uCZTlf/YI3rvfhU0
kf58Gpz2SAOqMc1CcNDYwcEymPbcRnL0yRtZINxw5jzMi+p7B7cQBY5yT0M/tl4HbkdsbwGoYn+p
fy5XuFg1lSwrLcUbz88tltgmk/tOpOBy5ZyTirw9bp+nYwX9/7bgQZheAUCybTkszs6hUDl5JS8P
Ej1fYOqkH3RrAD6QiHg0q8bRBWBSKmkKqEIsvveTPz235UaV0p2hvT+uq0dS0BzqXX/lpcLav1d8
zNc3BFGkoTONbaM7ZPDS8Ii4UEKNr0Nt03l4t1wH4PPUOGrEV43ujH8kJO9KPv9w/E3oCwg8Nynm
EiAU7Tb5esP2f+QhrTWPc3fVGEtNXr84kJoRdNeFg3dfjqb4F1zuHIJvTtFJuG8szFvNWiIPqQGX
tXWEXyuAsgj6/Ezk9cbnrCtFTNj1GfgeOnyy8fFfSRnXH8vJNWrglddbhf6qv1qwixNVV6TJcwuO
KOQV1MtbU8fFQQiJGfLGYOiPuSzA+4H4n5nGdEWUigYTveQB6IrZmRMiUsOFtQK6pamKzhHdIOZq
lWmneuT3e3QS/YVF3rAR2/5VG1V0aKKyOiqUMzwaOFPTunc+A4TxCSmaUZbUDcTFXyDDMM8Wrjba
08bzmOuuK0xP621lMKV00M6k904U39LB1iH9DvLvg1iuVtLItxrzFZN81k7F0wBwQuftEHtumxER
WYQyCT6K7f+OO9GXEPD3ujANEt7lWunU7JbaDPqCnIm51YDzpYZdgAxoMBuGrpjo/Cql4nuW2WYA
RI0t0/3ccJp6GFz700QDOA+E0JZFU9+Sj0ogmC/h4wyVvOdz81cYXRD2l2fLiEcL0UNK02JNjs8g
efCgVUL5cOfi0llArMj8OVmMCPjYj1mFsHx/dY+9cbE3TvfKPRv3ssxCIDKMrQbOY8xX7wn9zkCt
6v/Xse4wxCUP/mWIx9M4gib2nHhyBix9mSjLLZReqiICoQeMLhbENMMCr6sRKIlSB16aw4Tgm5yN
AC+27N0UBPAZB2zi9FcwL/JoRz+QaS5j7e5sudymM7a7ElWuJk1Yfi505uoRcIXMAgTvWPAviiCy
4Yvs12rjjxeWrm7cOKZNlUHTmldlkiGy2u/zDb9WKUy7d73ZgCs6ygUprgH8x4ejbHEcDuVoI0TU
BqzfSmUdm26DxiR8xLGfO2sdvtJ6rgC4C4vN6J9PqLr4ZFbhBNhm8EwIuxq2VsEKzqe+S9Qih6e0
3ZyHK0p3Ib2S/OHdGnFJ5lR8rNZpT42ZlTvLhFcMEoxFtt6ePegNTqBV/uqzbYEw9AMz6fMRvfon
THdveeA2G5GeONiRNYGCOFaq4UqDjIAdIrqZL0leEFfOmk6BxjRTGj2qStRWnLFooUHbNfnVLk1I
cEXqPuCE8Z4uRqmo98KMl9+iqCkx9pilgrvlm6BZNduYRkWsXXgRE5JZOnuK0IPeKQykIyK43Kry
JvE0JpdFiUx5+zVJn/yDN+6vspLj6s9+AeNVhG42YMKDEXyonIC7cI0zHi1Uqtnz67A2xAJaytZA
1UwXydm8vOyirzdFxc7uq9n+Aw//02G/WheDjKntuCB36u++aQW9fIFVCpEdZeTVl72dObizM1uK
lmOWJbkZ5/rWoPYLITemIlKgrha3x1aNO4Q+HyS0yh8L7OFp86kAGY6dPRz6vD66whWpPNd1Fb0Z
VriL8BkAF532/NjCE0axPbzK+TgNY7sQ0/pmepxwilfKvAauZNYr/Pd3yIY0nZv+PcyX8nRvXxjH
6LeFEjFz9GTYUcGkE5+M2QC8DUV7N5+m72V4lLqy+wrelWhK3/MFrGOVH68VT70AKLONwHwaxf+r
ucJw1YpHfWpO+EOQ6Ypqj9w4kpfLnSAkGW9MaZONyGMkpoRidHa91HG/axRzlxtJhkP/ClZukM2e
fCMhzelfoAaLAtYFqdZY8N2swNieHKnr97YvFLfAAX0ZpGo6FTV0F7gLt8DmeDPyHRCCQ/s9K2BK
RR3ZuI8q+EklVitr/qCpc/71wL0ngZW/vQl78JnMV9SyHDMFq4SGxL9a24nIyoH5inn8qFGf4vog
+AJQCubbs4sfcraVROWanAxi9HKIDEqkCUzjHVRnuRo60aTd++f6OB6yEJgDp1NYJY6rRHt93+5k
lz7QPhPgTfLx3MpLV/7Ef+D/O1AxR9qE/VKIcFooKik9Xwc6b2kyo/ZL7cDu7uCFGFDbxCadZnyy
Kfs87TU9Z1eTkNF7Hew+zJyQl3KDTl5aJ+lUlyFcUoj2HTmJagwTSsIgtay2U8WixH6VaN7kGV2t
uVRGhGxziMG2bSzzJjGecFmFvYsRbUz6jUv1oIBw8oQrZecNnD6VJ3D62lZF1h2jXC47/AMBnpxq
1kcejAjbO+a7odTKare6kvKGlC3OnYdHfc41X8/jiojuc0GxlfDpJrKRaHBEGCjGFPlX9T6Azx40
ue3qWrHyFzXAu+R9pojt0UqLd32OWB5J6rzqACNbc1uzyFA2LKOTA6q79oz1bFvBrbeatKVHZ7nU
ebKY7cuse2VsdRW9IM+aQGAyF5CX52Q1J+TVFGbc+fSSY7vqz3SXAwKpKZTl6Jxa41tDUyMZToYE
qUWNgwjlbxSQ7wZNDWXuyGfRre63ISt3BmctonMtLrI5Lre9AUjete9BGzQIA0YbikOjDc79ReaT
y04IOBX5WAP4A7kUx3BTIfKX6WF2B+7ZwEny70+8c0U5HLoQ6sLbTY9sSUfXLj5eyAnLFCeVoH3h
iRkAUAq7fCKY6gbW49BAiKpi0bgEgnAvNJ+At4ztIryRqw847HHFmXmPVss65ewSD6CeabdqxYUL
zzqEbDdC42KIR2yITGK9sZAyNlRs1IF1iu5QtEZFHG1KQfxr3K7u2/+zUXtDxDx0xL+rV0eXKUcJ
/rfMLAF0PH1O5ZZGtk3X2qJ6uRDNm664j6UThqB1FvwlFVMqJj2zoKDAsoyskgJ8R3WnWcpzbDIK
wUzdfiUdMqVJqdZAm9pGRrB9uApzPdBmdClyyaD4I4Da2lpJ1dlNX3bspC9QSPV+dPWJN9D8EOxR
DenNbbRZIV/ehtKfZrJQTyViFSZ6eH057X1h/xF8did495qA1VEkJ8bKT0c+Ox/3xDsWzqvhyOFh
ZP0Bt3XCsjJLbmVUClN3flpmsw94BjQ7QRDNrBeAt8twelHTxBHdAH6kyYFRNiINr9bynCXIov53
PqxIt2B7XocKuUWZrddE5FgUm4wAsdsBYjq8pIuul4WQDvEtWK5qNaCpoRHU3unDC++R7i0RIqaz
CLWoIySspEwPKFfXsykryA46ijoswthsJE1mFFxOJ6G2UhdgTQjE957ar7u9TqpGtH+Re4VHKiHP
16jKnxgn0FsLnXIp6ECwMQL/Zv+a02/rvHObkdc8ZCNshleS78nwkfxpMsES+1mRTNNsIyCohxVJ
fzYMjd+7oTTNxeZeS/JYBrFyEq0o3it79grlToIbd3diLFiIr26jdiHysOI1JkQX18lTKq2kzwY+
jSJVC1WcpvGUGqzp6ybSLB399vIwQzNb9QKMypAMsoZgGx0LqCSSNoOYJHEpDW8i7jBALwIhIsWd
1k2rY21n40AQ60MkOvItqQk/ksMp967U0g7DSFeatIIMmbe2BNZZi4ZPnY5nuqx+FCv94UjMkcsw
ge/XLtJoYyigMRr8It5HE3/Tm6X+13GIBprNqiodBhELbe3iuvA76/PePa0MHyB0l+k3QFjeBWX0
HfvFEqPZaMq4K98XhLpExSSDlG0xkU8Wu554/59L1B/X+nDhLMRZ2yeB2TuXw33tqIs2JPK0sZu/
OJL0Sv+5/1uw9M1iV/yuHCXpLc9k6PPtNLTnlm7BJfSsjrqde2otdNwj83xHJop+MPrzPtILz7DM
EtkmInYYyGpnfpYecr3OTqa6r5PiNScy2nyQFPRcWtdlXrc2KexnkLgpxocQhBxM5viSaCKrbiGx
6hBuL4ndUJDtazKGcQmtq/Ed3wjoMuBO0HvEKGTmdj9mNiFhhzqZgi7JzSZmFeaNAxAO6ckJJfhw
NdUKKQM1ktFgFzsmhfJLUZNlvtOz+aPQrhymqBIl9MJd/vB2Kf1bJXbRgecXd15J2i5IQqdjh9w1
JNZ5zmTyWZbwaHQiAa7zPQSfBhkpmLxyOZMDrXAK0MSe58CFWJ7S8SibgBsb6H8kASHixmanzhfX
em3ffVwZOLi0EKDXMgudq42WYVZgdcDap03B8lYI3F7ejqJikFdRQpihyIlhXdBNSz3VOXhndsPf
4DvVEd97yxYC0+G5d5HB0Y+8AuWrtMtaIfxSq+4GFhLItsn2KYWkgYs+hyD9i4TmnlNOiqJ7Ewo6
2mZJAmmEVkMfHw57vT7/p7Q9QdNnrToYJQi2EtQQV410gs0jNkO9SWCohJ3uuNfwogeFNIJHnqgk
4nDIfv8Zk+dvjL+B7DbVxGIs8l5Utui0rfeuMXeWzdmveoH+RRjDJGv/vjZixnU2zJFe+5VG1dmo
sy1y6J0X99eIHr7xcj5UfUBrlM0Hnir2S4B0w1pFWrBKt1PGwUHi2R7BpdiLBAJ2e4nyaN7hFurY
6TS9WaJa9VwXVduOcLmNVBrhoZm88CUs/7NTW12m3ZLFbeMiLVAcp+qQ77wKphGF8D7H/WswgNhN
aGVoIJC0ueS+MyIrtsDlHLJ2tuv4xRH46oc7V9EVhzdS3ON8MapPx+X5xA1JOaAm51sVp5aggc8R
iB7vzQGYrdiJBFi/tYIAlASJwp0QUEbEMaSA8iCicuWNMe43qdnk2WNKsCh+beULroR8qIacbv80
J/018oe/varVxnuV/gI3UHz6+dkEEZDijSRkpaTI/aONW91nLTGIuhBSQDStAhWNxP4pCU1skv/1
CgpoIHiHm8HUqRY5yt7h5k+Uh13YtK3A7mxfq8CwWDMQYwAv2Hb4AKdUeihxg7Y2cQAmLgG9U9au
b/x7ekAjs3fhEAatmyVUz+kf/QytTWdL3xu2kH0Zbf/WI0QQ2PHnAq1w9YP0rS4rFVR7Lnq2ykyx
6N2hAtH4Ww7FUs/amNgVSwMDnWtlarxM9FRmPNby9wvxuyNvZpvO3LDSp4u9DX9nkLnT//UbnPzU
9TJq4FoRSRjqYM8iFJX50lpMA+Xen/NB0mEg/dqtwrwo1US6AzrDwy4pCW0HONOs7vayLygcRrtj
Wnoo9wE8hmmxdizB3cNM9xGtoh0CiuvBptT0PdOu/r4qK7KTcAiJS+clf8JL9oR2+Eh6EOZNYvRa
fuoKItkqZgeP8+vuP6zidErka2DIxos6lIMKH06ggMe3ct0aRRjzAbj3uWoccn19+BkDiUEo4lrb
QFktr8eMMIj9NJccWsb8WRRKZbzPPrPKA31FJtY9iGnOMbcieJMznQ/k1mTj/hOp8YClRipzA8lJ
Zin82cN+uLVwTo5d/WUGfhp3O1dhtFQSnb3lzcDjwwRofJvXxgeN0r7L3ISBVex/ATh50uR3rN2a
x2JLGHr/THC56s2cubuWTik31y6z4YoJPii3qTA+oh/jCUcIxUkHSPnEb0ifPHX4VR/qq7wOhTuq
WHktwWebWArsb9KAIUHVprShimzuQ2pY6TWhwhDv86HDL/WUGCEAv/E4fgdu1FvBgXlL2dP5eU5w
rTKnNfgbZ2y1zQJrshQ2K3buBJxuymYYj3IDKWKfuk3Vbs2lO8AXMFZi3Zl/DGWk7EUrqkPlcdnI
5RY8W3x2LYZBtMxw/E+4JjaG4b7pb5p2B9KVGQWWADco4urBwu4sOf6d29mkyRrnhjUHfZBkgyrD
zdHMYaiAWwRoCQ+yePFOLyEdwu/VpTMiI1/EwOyrdrGr9IXiKrJswteUuqzNDwwCIHnk7vYQH3Mj
XjwZ7W+8tmF6GfbUAHexGegxpGwEndvAzG9RHIm0y/3tHdI4uTn+2yj3hSB03MckzOrqQmBip+xE
VtsUOhBOeYFicYaxYCoUWymK7KL23yUC/eG/3inQn+a/xEKnWcozAOEcs/oTekjZHbd45gADb4N1
nq2K+dApv7jjObQb5ZRf9ZbRPlQqWqOpAwv7egbI1ypkNNwnMvFUCLqRzNOp3lkUt5dbo1KBncgz
WV2qpeDHvsrhzfFj6FInFUsJ/MGXHAI8sYtKKRqHzPm5blTxvJXUotqQFcJqB4XIjCYfWe7gohJd
WjMebs8X1lKi0yf3SKCItpuPUKaPOFId8cIfYNBA1yHJzkYo2E9UwLS2FvYXEVcMG2QdrfHD+aG7
y85r07PGX4Cb7lUfDzvleXOlJNESNiQzURxvWwxA+UgyFfmZKghuDkW0eEdDsAa4DxXeLOshpMya
JVXXoca0IyM4f49ttpKVyyThuiOqp6xpQAqCzKkG6exVRoqqK2RQOvfumebjzlMOY3JVSW6Cqn1D
geSDVBVS8SZxzporxO1OOBFePFgJ50oUFOARfVBwKsKrW0MjJ+zGOtlVeXIu+t44fJINDfYLsxYe
Ipq2J7oqgTdKBi4hH81pyPJipn5Elt8e8Pc2XKn04jfVL01tYd+eCg1mMUtO2Rw0c9LoeIdsU/SF
/+P0RYquPc7FFIuA7wPx9S1wgRygApbNjQZtUdj6ldPtyXHKbCH0yGBur1QbOuWK5KymtxrwrzkP
dmaI7RERt93ogYXO0L9OqHq3XxSEnWNCN0HNDQtXPNXcYAh3DNNv7SJFp+oU6ieD0oGYuq6QJjGB
b9cJ+yCRlatE8ci/YCUWhjx86WVzwz19QY7nZC8YN2fVuclkESLYm6aY8AqF6WLhX3DAYX5b0+Az
Dmoky9dD/5ddOO+L9Cc6JRiM1iDZMfAQBm2aSYYgLubqQfEoESx30ZGAINWD9BVwEd42swuJPmrK
dexfXeuS+YTSXva5RAOHPFp9s8h7S8BL71MMayu7M7yR0wkuS2IHXSvaPjqPVcny6epCqM/jr+eN
3WrPTEnncyMjeIhX45LKZERbuVDP9W8qKl4oxvoyeS4Cq8r2qSn5T1w2lPZ1cenOarGA51PmKHp4
m3ESJGWASDmeK3y2hOe56GQdvJz56Dqc0mO3pqItM0eijkpqI0o/jEoBusKPbdchLGtIe7S5En1o
sc7LQdcIWTHyts+Q0/ZLp2yRfwZKg6xK8IQ2yYTAH8ezuafbcFt4XmvL4DsmCLCI/JFvZ9XWRRaE
MORVGBvZUp/IjnGzC2u907XM4EARaLYQ+p4ecd1m/HtNfQlHStQyd+v3juw37rHCFw9s7VME9SRO
khPMGBmh6UD0gxm2kmFe6hqdx87z8SFKl61GPrGBLIT+8T9XHmPfy6ARHoxUkluoK1Z5udVygS9w
39KFJqW4h0eQIXP3rMgZrwKA9PXSFz7C7yaIwcRstv84Cz8gNo/bH1wYwTbPS7SUsPKbdfGk4P63
UmGMqv7TFzuzZpQo9cxH2HvfpZp1PNWC8uXSolRGaZk+vydtLMH63eWrAf/U5tkb1wXTy329EP0g
4+aZMeyapIvDLGZNHVqzhoJsONBzGT20A/rQMrGoaxlJtgF0/B4QUZzpO3NCG3GoHlyEsbDNbw9D
+LFPCLN/JKD8zHeEAW6Mf0DwofRLc6YCkcEWr+q7tZKdlw4P02nwoYN8Q6mRyguus5SMQaUtpLGc
NCx7VeaDBX774Pi0Yf7hEWeYTJ4jm+mp4q5y6ghyLTYnlHiS8jjWO6geVabTLJ6+EyrafZqDnB5z
4/t0pGUgDZuRZMcT20VLggZevPLaOhTu5xcsezQcaDF2l0Q0oKpMNbiwO+3DNnymPVbYMAVY6lCq
/oNmC3Bzuvzh7Dkmh4+9+ZX00arZ9zGWbieqpbOjU03efj6nHMl7V2OmwpCBNDxMsB/MvdoA99PN
IFallCNv9YlZa7Y1ZApgGMGC9CQ8EtfjBj8j+OSsgLZnH07DeMlU5CS1hIpeoly+qS47N40LN+OF
243BQ8fmfge2ss9Bo3UOgj+/PI3EcSnbwe8DJxWhcMn+mYoJHkk82WlRUWtJCNwTmwtzqp9r+qWx
npPZYwuPUax87dTdQAP+jBgkd20I8u/CWVCL6Fx31xT9PiBHUQSPAreVffMQkbWJQQ5+qQd5SgeS
co03umwOsp3KytnjTFIqEAzXxggSt3ZmBWqJmcDcPu8/AxQ3nmDMgZm80z4oFCj3py4MZvoQ0s8m
Cc3knQ9T4YfGbI5cb7v7jKAM8UPTn5ejLTnIUm/Z4MG2KUis7wxQYWXc247lvDJ2PNjAbNY7s/Ss
yvIcvn/Y3io0M6rmZTnPbXfz7kdfAz3R/zKUyCr5x3MVD4u8Rodqe2wv8vxTvplmyV3j1bhgcAhU
H08jpL6JyxhRlWMlga+kBfKI9bPJ1hu3KT00gq04agHpabCp/Ycj9KhY/Akv5A0FBo6HOqS3eMy8
hmDvb55Ik2EARRiV7P/ynwxxroMHK9tO6rGhge8qcn1ni8Sl381K2pgBcZhZN3V7zkQdGvNp3jHx
JyRstkSu7TJJ8M3TZVC6TbMu2RsHqclpOMxxJIurvokE/xUjKDbzDDYMbrCEM3nr3CWcIEdUshTw
nmykSptfWU9sLOKWEgplL3NDZ6adk0CVbw97N9hT2h2KUHOq16nb4wQ4IHSUcgXxApbPqhbhem1C
K64AanzGcXnhJBNnwlbNQkisnsxAFiscyfShqefiw9zQ9mvLwrDLboqhT2ADrg5zP9JMeNeFtqT7
omWAWCKFrtqNKvDbXvRI3kAvNJxDJPFc3WE5XK0fQ6RZns7wnyrQMKuOdeS/tRaVgPO4TrvSyab2
mIm9dOF1uqhM28bauKv4jlV6R1H0LUqcF0IRSsh07Ws64UWHh1kSykYQPwLZJWh1M0xmV9axXF3K
MOD0qqbwYQxCPMkXmsXplCfrY/V0PFFNqfAqd+Myfz+DarkfxlqA7E4QFkKN/7wZTENBToN3vbMJ
L9KCfl7NbFGRYftyDaVFucGrqv9Pzzk3N79wz5Nb4E4ONYaQPEOEWFyS9IQdYHqcAYFcwWIoBxWK
eqkK7JdZ5pc8/xdTa9rh4UQ1mI6ZfHXrnETRDwqWC8PlYiKBfCbz1g6+s8QDAPM2B4QtoG2yH6yB
t8OBscz8tCN9EzqCUXpaK/aVFAcEypR1BzNkPvGWDULiLpvvKN0/itsvJspJSNqVu3YCBHeiNRJv
Rt1xbHpunt3gYJPNFGuFgI+BeUpO1QTIsCgF5Vlf5Q6z11XLGa0UfOTIa0WRFo1qFd7g4VHhSMoq
Ggrd0mw0lugRoYfF9gAwac6nCXggzslXndK4pBw4frp0Vfh+6xWGQIzy4TcWvZP4aISSR78eijwk
7bnfh65XGCIdfuwgbe5bEnbkI0ML8Xh1X2ySySq3LPI8q99SXsw5aPUQ1n1TTvoFUy4t1HLX1eGy
8bgv0IQggELNjeYTkwzLkZ37c2y004MaLEz4qCBFTVMsLOfSYIF3G1fCfeMsVhHGYD9egI2ZbqXq
dg7nW3inhHdOHDGJGPEvqY2lJEFXzjPMElYxZ1ZQy09GBhA7Fbik0JVCCiw2a9hBrBnyQIbNjDp0
0mg+Kv6/aKt+a8SogJT6UBP5RTm67fuv1O+c7iBrPyTFWva9E98q6c+Fb7LvgYV6L1BgCvTxvj2s
qaA47sTZzYCoVu1JstC3EGG9FbF4NX43mvVaEPPKqAM4NgYDC/UBrbY4Pl2Caxy+FP5As5Q0WWw2
yC/fgRFin4zRbZrkKP0lWxPcGgo1tLe226nJs6sGKKnI40aGwe5dNHonvQ7vJ21Rrv3CmTVlFRqM
Wrm3STuRiB1r1+l+ycfOTIGqwYtjxtFYn8wmrjA/gCOKT8jc4ghTsj+/ok7lgztOALcUBr4+J+70
93cT6HNZAA0bFhi5gI5s4s7BbuN1reRGZiaO+srSWtwPlSG3ziAXuWoTrh2msxmCPSNbYoSIoSM5
2WSToQU+FiEA1SkjTsJuqNIWa0Qy9KSTzcMXLCvYt03JLuRQNc/A45aceGPSpeHisojKiI3h18cA
69GJzoTnssi/EC1A4gbWMTUzN7CSwla4SRstmp4yHOfi+2xs5MgWBF4NggU5HJjQDpXdSNl2+4eG
Sb3i/d1dAmMa2f35FjoXN6P/TwiH/ul8jqcl3fMcQ312tbZgDH+3uEnyFUVjXdLeAjd/B6/6oJda
m/89vQ3aVp7uwtNs1xpMh/uxJJarpDusRZ87k05bmqKB6B3Rnk+EQJjjP+Ep2MRdzUvZWxzSLZIt
uw6oRCx73Hp8Ov8l3uZXWgxxjBzsBaMfm3F3nDUGTrrpn7dDS8y3UWgB4FeHQDZbpeuzN3DX25xI
pq55pB9SbS5kjsAAP5QEHauHuvcPzHCJdu04oKoeuiCAU+/mIBeC9aXqR24hUk/VYX2LRZv+qFym
0W0FJrWAsIMDfWP1pmN104wjbqjbT429zPoRl6iyTIVH3Cqqz5jjxthzTx3uRHSw3JFN4V6RAVPw
TM5iFyeYwPeEID2rf2jFoKH+0utLoOljIYFLv57poaIHkym9D/ewg2BL3YRPpXs5Vs7XAHtvxwdg
kohD2fOSkA3imzBpOwog/URxR12VYh+FmEEtNFJsXxLGnzomySHajNEQdE75u19lnyvMO3fgUUNW
PMwLEom8bK6kAoThVxpeRDGOUASng94QKcu6b/beYo6uDfP9l3pyiy4EmyW1NPXiA8gl9E0siAQh
/GyTivfcBUbtwnLUZbBZ0w7a5tVWD5/IDPDpqGHR06TdOEwoSJydkW3YabTtSWmzeCQrzK61xTl+
M5Xpp61164lZp8PFaO6u6pmd+JLiyxnhXYabcABqaXl0kRd6uRYv60ZpgKggGGpkkOn+GkztvyqI
9SieuJur8wonlWctYWAo3yKl3PlUF0MX7UNLlByzPUqMteZP2Wq/qDDRgf2h2j8PzBLcfK60grqX
74JddljR9y5+0zDuZTNIRvXhYGd8CCQhARilcEJHgfJQ1j95UuslcKXRse+W/l2HByPoQ+QTRLBK
ETTWXDVpebdiMqkWeaZ81C87bhWR2ft5uYuv87i4HWt42TvIgILqK+4+gs446cUudT06Dn2+Wldn
bTTZGOSXeYk7MkryGOn8Kd878xGgcPfVyOyNFmJMCaSTUIW/vNPvidgopIiApXriS2Qv88tH/c2M
w5TAhoNire17owPJMuFua8GGfFTBsdy1Bhf0fdYCYQu2x0rKoR/fNTLEnOxMDBsLreRD5gfOmJ60
3JCrIRkvgUgYn2P/ZQtIKvFcszOcJ2cgNy+WRkM2Ut7cKH3/DcY+S/N2YmSfv0U1XbpLqE6V00m/
RcsKJZgtdDs0RyXUOqtbj3psBdO5qaHH2UKX5Pqx1HStHnyj/0jf5ZWkLb8ZeTza7JE4flLd7480
FSVeAxkoDQ5XSbgtUhMK8UlaTDUeV47yEOKRdkQGnAdFLHNV8whPnnVawrbiAZtEPsP4FNRmx535
xK0F583frPjbGldE+6iXKM5xw9ocaAjAuJRI8dd8i7XVLe27R5pnrgcnC60EjRgL3QG9zneL0Gn2
wULZrqTCYmjU7jBhD2BZnDczFXthRshgzDZ9wlQF2dK+dThUxHzrM9y/OLWzeiF/LYsBSyS7j+1s
pXfJGTTsFJkNK5VfQaLdRgBKwp78G2Jjz4gj0zk6IwGi+FfahU655s3qKpUGNMbxKQUHQhnDtxuD
DMNYybvZ4xANZOCFdWRRxLWkgdW2UpWdc2ygNibc9agqw0qjC7UVBjYUicd8+DKZHoutCbsBcJtJ
WwuKFqA0G8Quj6cp6uTMBcbXztYPfhMejX+yOXWGuDnMCq6cegLaiGKMoBUwPwtObGGnFBXJ2Upx
ck2K2Eeq6zjyaXKbEHmqkiriqMkYNCoJQj3mDKpKs/Vx4lJ/HeE13/Xlo8DR3yu6zDLpEyqzgeX5
P95UGw/1Z9ipFF8Y1A9R4TNG0uNlJaRQ/bFdmW3UWtr3G7akkJvezMmITOb2MD0k8XAHuzU+shhA
VIF7iWQFtcfqKqX5kW/GZh7LIMlQdKWG7NWPn0gGvqcUM6GDQzESMhpZnsN54UZZPlsQ3Zw43p9P
1aIwFAvxtD2q2voFXvLdKbMWIXSoOnPIiOxxGXZ4dM+teHWEex/oWrYEvF/q+G2zZa2Skfw6/pNl
5Z2KI/yKWtjRKZ2InJT1g1wFg3ZYc2aIm1ma8G9R/WKrBwyPpHmRG3MsRntDkVlADnIalxY8slQU
0O2L05bPS/B4G163M4wjMlPafTLxMX91VoM889RJ/tOBFWiM4wVH1puoo5HiGy4y2a8v37W9yeWC
h0yiJWbhsCr7TScauQ9xvIgcxBLAjhOsUme5NSFaixuyBS6L0IN2LaQRN3ZLUc7xmU+DEx5NmIT6
vbYUG3rLzA5fEWzHbU3zkU1g9FxdpWNb+ctOQmKttWpVaGCYGS4urscGrHmZQBnEGq5qK2wKunqk
EY5V3Mzkk/gMBAV1T3sSKQRbB9UM+njb0UzsgtNe4aUvRwRQVLRIk8RZ7eomasJjC54tRyQLZ83e
RxAFA2+hOBCeB1vtRuznOiA0nGNvBFR7EoEjL/yQ+V9acuNLaaBCKGcW4TMtmwDGYaCboUiKZ6CI
a2RuUGPKe3DKrCUB50dUF2hMLq4z2zTc1r04d+RHIohD9obnxBir4iQ0Lwl64qp0JtdL+z4wJ9Z+
kgmvcUJy2WITPjqHYANN7kPD5ZZ9DP1BLr7cmARbF+bwcu4JLPsrKYF21OgPO+z9iI5sUFFLGN4S
0sm3AswgE6Mcbcx6IaHWgAG+pfE4Eke8Jqz7hqPi86nuU4nLtwq3qZW7WXDbY8PjmjgLTnOx8KoW
PXXBVZbkmA7jTlFim4qv5QCPCbueQt89vo4jQ93hKeujgQyu0ErYkvpYiokpVTecDDMKSWnQtip7
5C5dRO7tAmbLRximvOFM8s7LUp5FXEtLm93+vvM93ShM2inoGypM8EPOH7jqW+CBQQ9AsyfaQ3XT
+ksUnatJzlqsO4XW6K5EkhI8FVgZGA+9fJ2R7jdsz/NWZmMdY+yXRUkLlbM/jUw9+uUtHI6Cqo5d
UO7fRGrQ1K1n/1bnA7bI/IHN5CwqamxYSJ6Mw/cK4LVpjjnA+2H7JQ9Hc64yeXtxAyB9GD7bcF8q
gOkK4/ZslTHeE2eCioVREk1tuAx6cpJqZCrzBpZDOPI+3rpXECadJEupE5hmeUbc7F6WHxZzb1Uu
dLqbU2BLPFukPqUwQpTda9on7j4gxBziuPf+RtbfGjySuNzJk6A2mSM7KjGMjd04MskqfbtZvaFd
nFZl59WU7dm3mqMf6w7sTLEAX2m4zPtJFnUtiXa6Sm4vXMBNb2+6Lzb/itdNj3t8wMpUt3+yr6LZ
IaRhY8+pnsfO0r10cuBv4nrj0BSzWnWlX9NFMlVIhC8e72hKnjx/YGA9RmsO6hGIgiJenKNeO/9j
mUGbnsuUu1UpSnrOirFXEK0jV4Qt60DqUTjJTwinTV40UyPiua6AB8IHglQhvrywKvGnKGXWj9bx
eNF4m5lhEGSYEl76a6XcUSku4UtniuQFqXU7Epc952umIVT3pRLUWWX5/wD+adzhdHr8+nkf3Ybc
lXNfcC1KGKfQukOKi4l0jpV0Zrzwlou4DqzuCuhpGWaWthKi8uKTiSIhKyADWs+T9YTFfVO1j2OO
uZAZ8DyI5bNZO13shEJEAWaPKRpWpHbxWdzIh+p491FWTVcq45MBDtqCeyvE6ajIQZtvDpTd2r+c
A8IW9cBJeN5FwWqF+Mu1Fn9R957jKUmLvQcOBox4UekztKi90VBrqkpG3IOnSlnwGQs7gxvlxBQj
vQ+imJ8RGMCRDPzwEzYuUosQBdgF4DFlOwL8JfzQdxQvLjiuStTukmtL+5vbqHNJmg3HCWGQNR1t
s4Yfn+DBZTszh3rWlzPQkh9cPJlRAwWOxZ1ERLh+N2312El2LeetFa083avVipOGR7gHhko6sgIW
6QcPMX13rgIx3EtNvMemx/0LNXlv6L11/NQVB1EIExuGlzvxixJV3LGrGBh57XdlpiCIirWCm7dG
lUkhIV/Whq6GbZwv3GDwfArwTABXozAJvYPYJOewpAsDK0Lfg4qvoa7AMyDDw/FrzivqSpyx4UO3
fLhqWl6a+D3Pi4uKfco/AbgenrTtPiXc2lx2QP+2Rwh9ASvM2XEQwWMiuUO13UZWD+W9h6pc8K5J
yfJ4yiXxD/BN708s65p1HRx3zF5HH1RKqjMIRcpojJoI0N5wX/I8I7mmvvqJJvYURf5VK3clEnnH
4tbm0bBNcUN8Vh+nri92ax6KfWTOruJk0JGxot5/OJKh2JtUJqLdc4PGKkWZE8SEoTMsqTHV8XVX
BHpowkZeUAPHliu28BJfiK+b9SDmIveLcKT2yfSCmL63GcDcH+9HZ+wbDwdVkfGtzU8h9L3PlUFx
he8FCI9I3/7cirRaGS/nw1ytCHF3OPMbBUesB/MRJHDtpV50sFtmysASgapGAE+QP19/oiftsQfv
UDZMhGV+WnGQki4fENaminJBpq8TPe559nedmOUyCuDAEhwGrnerD26aBl7Qmrnl1FNu5IBR6Ani
GPA9Mol/S/gp6Cf0hzbaPAoX7EVqXyjpJ99QadFJlLb7c4bt7lD3fyBNpir6MubS1ZvbNcd7sV9Z
ansGH88N9/Ag2EByWA/L5y8zK+gdL2k0Of/u66O1rUGMRdmXDb6U5R3YJXOF92AQmZlAZvciWAyG
nQ1uUexos2S0USw954Cn580izrufhGpH6KMgO0oskMdSjEgZAnr4ueTkdD4kAlLCFCyDOyMxIj78
KfbM7OKOCPx72FzlHr3XozO4THsFfUpFKkqzXeU83dpcjg5b8M9Kf0rbnFmAqY/mn4AS/vsoFKTh
qpNWLWv/nzJoUBYYn9UXcYeLBsw+nh01aX+us4cR/j07ifSHVwSFQvpBA3WsQHdWbt0vQ6+Ui/0u
hrkeTx3YHJ7wxzgo0tBcRQKyf0rDuOUkcbDIKMj8iQp1RAuEbz5CSBbH/57f1FlQkxE1J1f/xMwu
hCm325VnKxuPFB1zEUoZsIpbJW46WDzprl4pJMK1Gy0bTgJSdp/MPWiDdPMGgMFvqYZD3MmjLDKq
ecmqMq0qUVvNSAGnavY9xrSM0EU53HTAQ3FjyLBprdPzwKIQd2vomeNcmxOPY8aZZ62OkcCmWyVj
GPPZxjb0AL9TkKDdxXsqe6BpCUqylS1M/5gdHbPgn3BqgizY5tO39YMJCIZsV5fAQeheavxfE20c
zG0oZXy5hITjxCcS82MpHGIG1pbp7A1rPGKeWWl+pCfUySkI3sdiGuSzeLrmzsVQ0zJjaAEVK7Xr
hWsP7HkjkacIjPQn3+D1AMhlX322meTpWx2wKzSXet5rd5G8DILPKKblrQJIqcMTgezxmt/sWW0/
fwKf9SJoCLcAaLMBIWvJk6uAMPLrZnIpvVSqHYh1unRIvlboadKEeL1fQS6iA1E0pbQXvw4UBJGK
DNC0op+i+88NQH/OmSPitytJgnbXtBlhM9TuPu2zDMx88UIZBrwSo+iPmVQMgWBbpekuOuI61jE2
xP324uMimkQ+NVTUHgOt62cZn42GBMxe2560KSC0B6AsrE7A6tI7/rQY2rGjvcvNI/dzpZmmxlmy
Za9cj0rhymGLN+G9l3874QZACmbCR9nNtkrcSlHEZdcenJekyjPwNy5QdS7x95DI/BnKv7PJJmZ9
LzBN3NGMbJwYP//uVQNRJkXbuvx4oS22O9mnDUzVlZ7XwaB3+cR4XnCI4RrRa8gORng2erdaNg6S
zGMhjvy3y4oYfVO1aFNArHO6D9JV6rQ+8qhj5n5zIyDrpkMLQ1krE4t1/qDtcr9YJYF4iQCZHNwl
QVC0IdTkJFVgPbCJAU5sDtyftqSGd1OMCuvVsHPgAavQT80+QKDohMxkBdl+ekaipToz1+gRDzmN
/KCkuDk/u2KHvlK0hptiBZmh8Cy8WO2YASQG1TtDBjPT7kG1zE8aYP3CyUPE9kPya+8aZtEtZsrO
lKdgw7isFvfC3vWWA0fVeL1C+iex53FMqbaKNONyL53Mwe41d3Y+7mLHWWSqMvut8erPbETOrto/
tiIufpX/MsFzVLknmPW0Ao3utn/wWepnWR9nmTXNYPgR2XlCpFiUHtDH/kc/eByD84DBsFy8gPt/
lLVmn54+FrTaLlB9bsGuN219lROb5gMLP6x0nk1wBu/3lESU90x9yrFYqVJG7Z4uZ+EpMDqTOSoK
ZPiZXTcOuqWxrR9pHjP5nBxnIoIwUzBxWpgjiR4kiTxFw6suG9S5q9p//TCEwchK5wFbEptMKMri
K/HYwF+0HIM8J/fz3AJ0eetCHGl0LegpkiJ4dSF/6rFTZyGq5sdpd1JMtGptUSPQ0xGXjOEJaDZp
ah224rTw5WBTQb2YlMc7wsbDyh9OjYZ0ywpWBEfh6xt71OLQKk+Qk2TSGsYI3R4bnijhgRiHs/dg
R8bLm5Y5x2XzAwTiFlXp8eit8JYn3flO7NfA1Ip1emK+EmfC7WX6KRtdqz7rbnpN9XGSZuC7+D0Y
irguTbtTxk5UqFEJWAGepVNR6ztP7dlOYa+laaOJ2G6k30fOR7L0Jabs7fYQ1aB4s3d+FTXFfunZ
Poa2GM9B4/kYbd5gVS2SGp1ERuVxfmxCxs2H7lTV+2jK5vcMScAgz8gT7NLyCFdhrbQW3Li5Bnwb
NyPnxBJsmvV4EvXqC2GYvo5PHhFs/gae+bG9ingXWhQXdQPPFn47aeukwXbecdWNtnL12sc/kHl4
lNqbMkEq616mf+Dq6BAbtgXKcuvGhS48lkudWDSojI00z0w8eNFLuCIy8z/6PFevrUcvaKdz72Z9
kQurvXWv4xnLXvByfc6CrcJjqCJGtDLiC6k3eYZJMJrmswFrJ6aV68zDx3nnKuA0mnMFXuWghobk
gwBTEjXS0OHZJgP3bw6dxlrET1rpUdRFSH55B0h+hfLj2P9J6ECVwhEywP629oVxBgMS/6cOjXSZ
q+ZNtOn34sbZCmUo7bqeuCtnMJ4SB/JH0uoTDkB9xTw5w9sPg77+ZrYrYnmOTXIHOFTQ3I2DAgEB
MQ2cYbyIT2jbhcvrFdKuQdhZg5hAYcDqaR3p61FUBVBOWiWCuqnR8/s1KB8PM8G8nN6+YIG2e/7h
aD++a7g0yUVyFoMxyaVYUzSrpu0aEwxSgQvlptEYLMH088OWbyFAZ+fYalc/wK9gc1S3DjEfqyRI
jgNDI9KMg3Qc39XuPe91NZ3FF0ePWpJ6sttE3yz0vI/fUtsFv/uviY+Mbr3EWxMOLLCA0/kbOJuI
Hju9bIWqEfgsutZxo/gV5hfuOHW7DNM1eWl4ahp0vLDj7qJRFa81OTsA4YwYckutv6pgEg1EAIH9
7/L53tSz2ObnuQZvk5IYrlYaYL94G0FLRBJI88SfrwbJQJzAwRIhucTAAOq0sOwM+04M42yCCOpX
UAMVRuUBlvkoIEPo3lfhBY5B0lXmxSRs7embHijzHCxCQPf2EF3mzlFIuqxoYyatek+9y/cluxU1
SxpxWA4RbiONK4Ge02aXnzjz3/80bmmX3sWnZIvgc1fGYYdb0Qm28qwEfru+6HTd2bLOiBbCqFbt
3Li3IENFkmn1/5WlxlRnMQ56bohIuJOcr6TujJdnpxQJ/J6106tojuFpvvbb/lwBA7ei7IB3in97
mgHOC98/ePSgMj3Vm3NRKlDT04EloCpFg1gCfJuc2wrFUaIBth4fa5HkEQaGQG0WHSEoYrcbs37A
qDfTmx3uE6DZMYgLH5Tsww/yag3MMFx6nMzB5NNgPYrguHjKX3dUvLTu5BhH/jpBrPi8StSSQTqq
wQcAkxnOYmwMyHSnxLC2yFvnVfaMGTY9Sn90q9fFM0JpozPBWWB3x9va7n62Rb5mMlSPirb0Fxlt
2HORugEBkSe/XULBzahWOUwvZ/L3KfYhj76ZnykxqQoZUIuK89v0lM09UYUcOJiA1Th8rvPznGPv
iUC/UDsORK/R73qYouMUzAuX0sUwVIZC+cvwgAXdikgvCQ0FTD6/PY1hKy26SiVUcjqbGMvIS2uZ
Y3Ya99nYDjtffIl9d3iC7GBHNYh3N9ZbCT9rBKaE+whMRhNp52yqaVGJbS0M383lylcRIqWVPfZW
XrcrtgSdZvOGVe8ZNlNbDKb3XoVarzVA9aqG3CJ9PjtAwPgQECzoArRSi43kLe/x4dWRM+vDSB8A
kjH5X8yJf2Nt9djFE5Z69rcMuu37Udm3t1SZsWXQeiF9CTkSi5cmXSezjtsop3VQZ3s2oiYQpjk1
0D8pR0hrd5E0qlexeF/w2V2FbJZpWfQhF+e2q9C4rUqtwN6bwGqta+ot99XuULlkg8IpO2LemfRq
+0lN6AEkMjS1bMQZ4iNb6pccBvl3yupBuIJXBK70nw4WbjEdTeGRUSCJVWFCwE8CQz95x2fiO8a1
Wlas9dIABB4X61DakRZFbGi/XRSXxh2a5JSAH2U6smOI/SbSvxEQ/0teVOaYwnwfaTyou7po3zQ1
TooiMjkbzuU804BUlg9DxQ5cIJiXHiu4WbW9iEZRTsj9JFW4VjEAWw+unpTrqYSWyOT/bOAO8qYx
+BCYMIz9b4Wa224CIBdGtYFcFl92i7sQCVUklvNZC7N0txkxtXDogZIssoej4880HjEz4X41EtFA
tezW5CMXLUYEP5/9ZQFMk1gwA43X5641eq2slOx2ZBiXMdkLjQ4CDkMjVNz+khpV4VbBSDeEbPJs
smthfJE8gBtZyd5mg9YCmVoLWshyCXs11DT11w9DNcFwMIrq/i2XfrSTVEi5lxKME81RD+Wpu1+K
F5BYUZ+mqNUCmSpU3/nBYhnCJ848elN1NkxbN+umzEahm048yG9Cy7S06/uFhnicrhQBQQVzt3hb
wTHylVdMvyEbYPrFh5Sopvpg+jtInjCFlz1ZCzPliG14sn0Akw8oUlQIPYyPQO99r4/XbEvElyWj
riohDc1VXXdopPxawysdc3YDi8NRxbt8UwqI2Xuub2A1P7wc7WpEzjXWvHlVqXcQU1hQd1LUYR4b
8oLdG2LQJISCQkkLBe4x/yt7GMgucjFsV4KExSUBEgLZAOba1UOErcLdOwrNC/4No8ctq5xaYxd0
47KIAdPokM5K7o2+kKXgXjhvSPIKjhbYsfu4Kdl6GYtBVrrxaCGqHozF/sVYy1T+yvrFpVksc7Rt
+rpvX3Ne/BTOWgsUh0j5aVwhCCda4EepiU8tedw/2g5cjugmZarwusrKBI0C7+LW/r/CblTCechk
SJ66MzpmCbJX3I6TdW1uBpSP38PPTDqW5oq1Sks+MjXeHh4ETo9tDS03dTxn5KoGkL4Jj5e8p4ja
AZfe8iIRD7H+d0D5xcQyXTTNb7YI385LcKTuRHrZcnfFilwrLgGGA+sxFg42vTDx889C5gsm/Sfs
isMuAYD4igKiQOYkxgOCP5w+dsnHvlJ+0z+ksbYySKr9XsU6NtczA7o7Hzr1ng5vagh8UwvGrRtl
arIW0+DpIg1lBOzVB4YrC6CXOS/YxHOON+fBuEHrWUk0GogQw4QnPRB4WK1sfArf+gtIfMSPgemp
ouciTYHmff74Q5lLb/sUn28Kwwzwiabic1TQKU6hP0A7COwWq56xF2TrKIReIAsQqtS0pKlqd2yb
2b02jlZNqZGHgzrK6ydU10JrdDZpSl9i3wqlBVGknsjh4bHRw23ZwTTaDMKAZeQP9i6OeHyGZvVM
8GcMgu5/cKysvPTSkQE/JXrX7pYJ7MFpicdBbynf8F25yMfti8v/dxwqO3SBCvNe2c0O4CewW2Rx
maj/DBNfXWr4nCV+4ps4bclRTuGxfZnUPttcoGU/TYhK2F6RQ9mM/ytD7mETQtpbeR3VCUCKh5vv
PCAaFuOJWJnvyfkN7L60ykLUfkrcSk3Lmx53TL2HwOVKeB+e48b75rA9396SZvWdiWOCwMtpWxf4
uP2lHQXz8lqSA07kclPkpWw7QYXu8pnWXEmW5b2tFrxOYxLbpyZvwu8mWguHdyh4nZacM8+TiO/S
+c4Nn6voLInNrliUkp1KlKa72Lv6cJ/5o38YOwm6ro6Z9S7KV3ODGuch88Dfsw5HRXIkmivnu8/f
N5JviPy3vyE0hKRpLq2C1ykZE2UQdELDwFjw6k1V/enQsePcxsbz07tUbrj2BJ4NgIR9JxdET1oX
nLkZPB0g/pZCkM6KJlFcOacUBbuL8eZoU1kIQTBw63Mpst6bVGOt/5O6IutGoWk0ZZJRYOMKFUew
u1Sh1ctMjcmaySu0UfK6s+CMfzHITthU6OrFoPIVCSG23pR9gdk7dzjJkeIcI7iVa0ok6lie+1c+
S3n+R7V0M6usXphHIGGecNN4tHOsD3zwZV8+oFP7qL6DB72d/yjl0VHtVJ50xAR6uTobHtzIN/zD
cBMmF+cyVdSSTK0tc9KMjHbSaCUE7DNrmH12hJ2mKFFoXJY4mYG8zCzEd8sOdgSK/v9Sgtso9381
juqRZJeibCEPKJVcvfLNSxKeI8G3N9tjz2/Ct/ele0cGUScIQSuEMKa92SYUfe92RyPFtXgVXwLl
p7pGzyf1JDhZPN61IzxIkUdDUG4KnncLs1z2KkkK7bWqTLM7OX7qvZeu0Hnk6E1tfze49x40HR75
o+4H+fyWD8HHXa/s6jrEGsq8o9IP96SnCKZapsMHxtSrF/5Yn1Qc1OqWbGulmRELotn84U6LWoKz
iUJN2NZQZBdN5KIiWtpWsQOK2FbL2A6VYku/L8id+bl9n4OVQ1ebRuroFTT9aZHVMuMqJjQL596e
nfQX+8nn71GHbsBSvmWIfryLvB9hNRDbBq8g1WsaEy2872v/C/fAWYFox6nXb9NCLFI9aCnquq3q
Z0Z4o9Vqg9u4/TFTqC3yp633+CaSUKA0COWblpgSSnRL41Uf4mm7euu47EdD8APzOz/tmEMYZ3ux
F+oXurY2r9SXpg+6QUBrIZlmTlvMA2ty73dJfIa5dAUGBeOsjtHtmMaQm3ppipw3uNI0ZIk023wV
7kAAm+6MjlJu1uzp7gED+MhpFJ3pt0zhdSwi5pY9vzLqeNnzEDKmRiw7OQzUclCkpfy8qmXXiog+
qDvP/M/pSYyAYLqvtU+xvXnjuKkSSkq94tQdK2vMM4JE0/Yi2xuZ6BBQWFAB9knYXN3SuUpVZR8d
02d3nVhX4m/x6pV8gksO4U+7ucxbAg55dSvKg4LfwuzyD5wHQt73GY5Sl9kiEpMKHu9uQxsZHVlE
6PwqoWKc55X0FHi81X/bpMLrrDcRuEHejf65V7VklJEXqmkD0JEdEa2yUlrY7XuJtyyl79aF3OU/
3mfcz4ajk6Pf1xC+qG3PJjeKab70QJSSui/uwMEQiwlMQ1t6IQdntKW3NnidSTsvs48Zj84Mv5oT
d97/1+3MvSiN9/3jxwblob1G0M8IHnENNJlk//QzAOE6oF+PXJnJzY5VtCQ+q/ZGQcy2qdV5O5/J
tRdjgAHmnMIqKE4sEAiGD7/czbBsGOj8MntlxQ/x6woT5oER/RTE5pbVcfT3xjBSBL/bni8DzEwd
LwiENAuyKc4ppThhFK7+9bcCt1s5/LQ3JDA0Qmok6t4ra+GLVn0sT4AlAXDpWNG1immrbnmJ0ope
+GRDp6r1Ch2JjLl0BsRsjcKXhlW0tYPklBHnJTIekEMQbE8jxoDoEvSGn3x7c/52TIXRPGJGu1Za
/YQmi+GVEa4+sNg4RLDa2Fu0JP8NLkooWm1Cxt5JLjwVvfxoxQ3yA0+Nz3R93JLWwMU73Dkr77N7
642rbV5njQY6yTaRnZg8p99eEAzRmOpp1pBn4uBp2UAuf4IAy50Z7ixLcKjhkT+Gj2aqkDmEnPji
GhmAcQ43n9ndPM80h14PKCjwhScYju5MF6ybZFFQWdPRdorGZwFXaSMnQXwFnFFdZoMZ6UNEa/y7
TzfoCDNxhHvMgKzWLXbbr+TMIOEp3qNr1yazp5BTNuH0C+mfYq0HgdqEuOnjagyDcnbgoEbXONnM
C+NV20b0kapkEh/KnyKruM09Hfr8ZyJ8HXP26YsmKgc86a8osxly5bLJCMp7szcqk43/gdt898EC
bvMou3AoiOgYF5ZIzZYlveboekKdDjdjUNquCR69486ZZHHlT/FbRcyqh+KtKY+fS1bAMm7v8HBG
xT2ts3kflD2pR8rg8KntwIkeb/aTapZRX417UwklH8hUlTVXOD0+ZGeDXZ3iSiRHVyMEXF6oveYA
iO7WC+jWnNzaJHEpmcIYrLQerM8Yqeevks/3cwVCWUEj5Pc8lBVXlYTANVfCXW70Dpzs7i1HPGaR
Qi9rD9O+oXFLwLmPOvrdYO1OSDzKFh0MAPBWo4u0xzsWKDEhJt6LIAKxwAqCsBsAVxeZPxqSGFNG
hgKI67ndbSB9LSL+M0QOYe8mhJWMERjTh0VOqvFx/CpIH+xtqroLwst0z9KkbUpXUsQlBN64iwvy
aeZ4rQn4ryKuicQR96y+SCMoSaJQGhRvbPOCWodcGjFruSqiPuNVa87tN8Sl2XpypydPlL2rCucM
x5x8vAHWJFapLs9KrA80GLVo8HKWP6fMI5Z82MmCFawDOfRcoOnxdOH9tjR22yA6MFZAJx7SfQEK
EXDrBJTFnSLuJYE5nh0VbFd0JMhtmgaCjYZdOdiq4nh9YLNMXNbYjtAz1vuyxlZ60jcwrffX6oqS
YtzgSgq6MO9m31Ltw0a7CQTg6lCYbLv3gV7sIUGwvqt4e/rhjyzretXTNAdaRdhBcG7x+YBZX7tu
2xHfzhdlo03I57nBQVyIRltBdFsWIwiqZ4PKihTqdrl87scpBdoZ/KZeGap53Xmf/VEgde9GI16N
hx/qlTaDSxUCFjnGcX9w0LemHmDCwuaU+ylvFVpFUFiohhVB0IlNBK1GT2/l7WyiWzvRcCbHx2ug
e1ZJJfDZIlm+Q4AjjJczfYBNb4WX+UAN1s802HbePPTkHI2oHPtG3zdpSFHOp031ygzGEWuNnWP3
DMVsErd8SnXLSM9ttkCTfbnqEofjqK26fwnAxnVePEH6Hr++Ye8zUuN4or64nC4zSs7qxjxkbFw0
Www28Q7PD2tx1C6W6HHDDC4cKoSCswFKZ8ISglboCxaCDs95nHAjR60hhdViyi2Z2YUEgNrn8Zaa
d/NvlV43deDvbF/ZredwyzKr4PxbdEx1/1q+9wsj3mAyqYtwAJVzKn6gWwnpBtSl0sgf7nAIKqeC
UZj3f+BtVfrAEo6G3VSkOippb2+Xm/3TPH6X22T5yreDLue02GrzMry2FWaeR/uoTIN7w4SlWlHe
q6F0vd1S4AyUuANAP+685VrUkAkPWHC+6EG/zdAq0DKHNFjs0NfcyDPH9NUH2d5BezbdTRX9JU+l
Nq1LpeCzsQe2wLF3b6xKZaezS3v1+4KlD7qqM3YxegW0yuD49O6+Mf/gYsWzzqOtrBuTZKxbLTfd
RgM872S9R0vU2KMsVpJrIxo/R2ON/U2OK2+PW34WCYH9PpCuB7M8GvC3omHn2riGopsofuF0+WaT
Qu/E7FhAo1unI9FHPAQYRQexRUsdYsyI9j/PeoNSMUbFQ0ceV/EtKSFBThrXaqA5w3gbq4HJ+V3O
OxcfLpaPH95tMqya7hwT4ztdfeA7OO7Rpc8lYfG3X4SptNRIB3ZXAUQOvc9ro7lwSyF9NBo8suYd
vzdrsxaqvRlVXVrRQPtdX6ev+OUSNUxwq/UIcDUKeMFowkwV8lV2AN+SVaLU6KCAQkvPsCdniiex
zD+wVY/1xZ0eHgXMGudiH9EGD02i+ojIZDX4kWT/EQgJmWThPvP0DRWCpmi2QbCwW6IGPrKBVwCi
Yflti7CVVYYhSxa/nB4EFJaTaZ9EpZEw+a2muetxIjT83Id8YP/Fir9vZQqO/J0PNqCOnBhOMui3
6dmPUjvZWwlOQ0th6AbOKDn4g/AnMj6xOcLT1Ty4LJENafruRrqrtYtWnA4fgT5fRtl13NqOad71
8OBdG5Uz9UNQvNg38GAEte7US3T3g9UDR5IDu60yvMfPfUN7q/OyljPMTc2gcWSzGtKB2jrseLGS
wIAlZxiUSpv3J1TqG3/Yz4x8sDkAdoRRAY1xYhGo8xCoaTdY9H+TPTjQwY+e9zRHYrK3RdrhixLR
uL4FdXhDFsjg5sqk3Y926Z/+hfTUX4w7FQe6kd570JKdwRckA7A8mE1iOgsEARMq3hD0ozlL4iOk
Ha87MOZE41q+bQj/qQi/Y47LS4gYLkA1fZ8p41n5/7bO0aTttVwgnpR63+2utgdj5G2DP70ole+Z
rQY9LhVu2lsUkbNpHh8rJJkiYBzAJ87N0yK92oYrBVasc7VELIssFgbiGPOoUJFnCJAIxihMgZ3B
nxZnRtJq5mgSrjfcpfLxVs+k+XbhnrpIicIvqrGaK3ejqmLJwo8zkCdmWmOECENTfs1IZeof+R0R
DJwSGt404Wq1kAoybtPLmMa3RGm7lqZMUHoAZtUOm/NNoe6O3kzjJrlRelO1PusgAEgsW0IvUt2U
xAdHwCecSrGEgsLQ8LoMbudK0iXa+VF7Xsyj3gBkjXr8KIykG6gp8xfvfgqIwr9heLOPFjoscHz5
RkEIZHNTJ3P+1OsK2wej0tQ5wTswaemsi5Z86QOelIq68e5AvUHaXZaBw6YTYflXgaGs4GaY14/j
s41FNACXewdyrNE8XUzyZBBpCP2VHop5gU3HJ2JaMdEsDKr0mGrA6D2mgy27yDd1/aWaiy/gsz/Q
BdHbpXeY2zsVm8TafBp0pB/Fsk5jdeHyc8Yaqu+i440271Rv5idkzs2yJAx11QSUr+Wfa6NTPf+W
AvFwZCkDCeYZq+Ox0+UZK3Cz0NwwxPe14vsF86wK7nIQZU1B/skjVXM1KQR0cQNGd8kHzFni4KKz
dS58cXUlDtHbAAigEtKP4ae1yHbaC4YoKq/Eod2B3xQAGofDKgwGrytx7D1EzYhcUkZLBdUC2NGN
W7sgvIrmkTo2mF3Iscp65jsuBG0+um8oK1sFB5cdBvpmTKBZCslG14rL+UC2PCbU0qfS60b5mhx6
MYuj2hUX2Z9Al61I25BUKqbM3MRiiMUQDDXbQtOmouAdYCaLRjf+nQxN7s9zuMSFlXpZ8spFrq+A
/+EQEnp5B+tlgkLUL3bRbwtUEXFN+OgZGlrVmnZetnVvmBr+EQWUEe3sIB2elo/HEd3Z8RXSSAFa
CVcYbXI8qtgO0c1PY03MpA8NDTv5D4ALH/ahBt1kKV0EO9kSoATlaNqLWlcQfI1f9fvKlc62Pm9n
GCGpqRqqBa786VSvfcVN6JcMZTCWIYZmIPlqwXB35VSbiguu0USdslG4FJXFaPzM88Wn/CRrTdVF
vl8UtbFogxtan7eDk2ysbF/GX/FRLIbTjxWdRtRjdKW9m8zAMyE4SG6xMWYvFC/3yYtO2YFbqplX
awT7bd3NetIxpanJncSehPMqL2T/lqxm96NXKc26JFSI220qhXoC5AM8dK+QidmyTNWP0FNieyB7
bs6FTRHQrjVW6TaPmOMZOkw6K+9/4V41OE+TZgvVwDBl969A7hYwaVC4cDlf4Nr5lfSdXBOwBM1t
ie5v8MBvRxcTrJrm9CtPpwLQU1e+GG+K8D34IqpssT2nKv2/VWNbFa8EEv0446RWZf/10noDCPyF
voe7olNdb8K1mpRMMgH+2LYjQKkc3L1Cv2R2xJFEJhq+FK/xFe0i7MqAtai2T0Cb45HBV2PKY3Lh
m7HFWvi3+Nvhjfr5MAAIK1dTcl3A6Czn+yT9QbMyPh2vP8eRu0dZGlxoeWQREKI5tlKwlrWfdvge
z9fENYFazfYpnuEZAToz08o4gzSj0agdMe6NXykCWEayVNT6x99d1Wl0ET6tUe7zpeZqfr07jTrU
4LnS9/joYkqtPXE+K0SmA2g9AVCiDNGS2A/+1zkmUrrx8qD4HpodpfVzFpnFu8yFjECXuw7efC9g
ue0Fo0R9Sv1kvXJYRSHOBaSuXnQDW5XwdlaAVz5TI6GEmSlel29HazdpfzuKVAD5sMh7PobTQmzq
YzVHRhc4ENPhhOtowWqUC5ygBqN2exY4DGxXKbcDdQ4wOxFlfDisrE1I53wbO41Ftw1XUhHoXCdB
zzsyA0LSnqgLMC+cmWr/T8yAmJMYLqOdNJtc8ewwI9RjO9JtKgMqH1liGfeUFjQSuvhvRBttozo6
VGGHHSL/Suypkf0tkg5nxnorBiRGaz12NVOgo/sY9XtobTZcJlpqQMnev7Tn8gYIlsNwfIdfRT0j
HwQz9PGpyp3U4HHK3UZRR5sDG1cVUQAfIwuXaZ/O1FPtq8JPqtSiPJeWjzNywjReAq9E66pT4rhC
Ol7Xhx49wO/2IF23irDLL0lerKg0f9djt5HqBm8OkVDuLKKcmgTjCoJPuvRqNIFfQ8k/N1wcX/zI
zzMj09CNyBWsjIoFRCdNSyKO5RLrCOZ+hX2g84Oz7UESmkYPup8X0XBshDEdjUoJSNBUxFmC3kgj
Lg4KhCoLsMANGP9pE+NRTZRVSkmAGdWJYxXQqsZsU1teGzBtfQVH13iJgZ7pp21mKMG5HnLFrCMy
/pYtn+g9i/6Gk+B16nhJBnBEtPNsRR+wdLt+AfXh8dfQvbLrEllKD414hr57VFR2lzb2ri483zg/
ZfwDicsFKwwzJ7e5jrXs8qlYayMLhRKGAyek/srw6khC3tM4p0+uHioS+8S8RnpSNk9Q/j1pIL6A
BZ3J/uC1EKvF0m4YGPpDKSEetHgJY7Al9y2NRHUfcsbsId3+ui7CQgLRheTEY5g/QVCXlGwBsYJz
wKf603rqCFVJL9jCi0cC0ZAlK4DpdUesoNRF0e4dl3v47dqxwaVZ14Ardb4XODYetiw4FL95fcqu
dGLbPqnDezsanTozuwmZl8xpq85+Ymw4J3Z75sS8pEFU1p6APEkuyR0gvTGv/rgWyX5aABVsjBp2
u5V5zyRIxFb/RBhlbfdPC8JcOJo62iOBB/P6aXTJ+bNMgkgzSfruYxrKEN4BAmcFOPoOLAT58znD
gb96k2DyNXqd0JIQBM/ONghfo2WNDfb0RIJtga7pAp5p0J25nGeMiQ/wz1XH4YcHrJFlvy4amhmu
lkHe+UD5SqTowyxDCW1jS/r1Vdq6LCojhBGN+X0V3cs3lWdJQle+NST6WwlxYVh2a6FWVAYVG0X3
bOI7AGQd/uTd/5QuNqnAEB9WbPLg/8bii54QcoIpFjcI7Pn0ew6GL6tugN+hhXLx3WbzRdPXCiXX
Muz6VjVSTNYXrhKYs0lGjtPyo5L0ZXEtVN3xAky+FTk8BkIt3UlqvH8CecUHOSJFJMSwm1JLAuiM
AbYt0ypy3KIFjldL1pjRlMVVzHKH/xiU5z8awTYlMJUDeO4DlXUgRFJLgXJNPSq4j3pVJl3jvBal
fccxpIUk/5N+qAgBhgnfIrIJp9fJxcmhahw4fuA8o9RdixZ0+Ly/IlBatbjrlwJzgfyuSzT9iolc
NxV38wYjyxqNL3bgkrOi7fqXL3LbyS2RA8jChHYxKjfAZXdIn2mOEum0NC7mJZW9LQolepM7XxQA
U5ocCe5iYiXhpHebIp+y5SQmJlfcYZG30wOFGxsFTDA2bGVpXZZ2MPklyle2Lj7rgnyTBKW+/K5J
Z2Iy7w7GeaP//FXmoGE7o/mwAdKMD74gDhj6xla5lNrbmJLeJHlJibFX4mHBhd+XJ9S0jlCud1Nq
yWphRNmuHVLWpYGDlQv8Vmt1BAzqFdiCJ+r+3/2AXZXXqF8dIhGbQvfQ7xe2tvspjuz3wz6RXXen
1JQ89OZ+Jmpks6qK7E2K1eVRa16c13tuad7D9eAll6isvC35CCpBEh8PTIr/lRCkWX2gxbsCsQ78
euyvqvEuiju3DaqeBmM+V7xHWpZLdd0Zek9nW6W+xTFDBDqm22v5KIjJZ9cysp3ypoeSu6x3Q2PS
inDnhvn9Aa4rg4o5f8R8PmtOqLayZJTVCP/pLJLCKparQTC83PBdBaXupuL95ESQxfqtAK43z3qe
mAcJMeQ7uyf4coFis2NQNetkyGagHvQS2cj4/t6hDnGbSGX0R7lGYMDbd7ZFsKtWFo3e7Bs0SSC5
WbrS0kT4SzWF5b/xihW3AmUO1YC9facQoOd7MAcZ5SCN4DHXsUGtR3LXxC7GHzaLz8SSeH7tY/2S
VEAyEy1Bf3Uq5IwO2Oy+uGTzdjDNi7SidjDEWiYqmGv2Tn/2VX0hBH0vVOaB4eUaRRp4WAXxoVWO
BufmDzT4R+xjFbH4NK+5wfgKO+dEDwxRt2SXs+eoyps1L4KRvb6HA5snmzaeO25Jivdux5g7C3aE
w74fhX2EztpYmnHXRfMcKwH2+4fwOgGQvnXohrpoDMKybxOzOpJRMQH7GQr12kg3L7MGpsSJXBUz
2oG0Ui23gW0lKSFInpIVz3XbNd4QC5+y/wz2gB5i2H/Rap0UUlX/tg6Oae01yNBSC63K1WldqE1q
yYcLAaKlMBAzRTTQIIUR+R9ea43iebZB3JvmSaG86H8hCtLOjd2U7B2nlBDx//62hFDy7Yp7+SMd
avuIbVkpUIbq4ZqnhiQN1xfN1wu0553Bw0LXsfr42FO79iaqvTo5OhyE4Ihv0uscrLWm0tW42419
Lcj8958145wKXYBnCkOoLE0di5Wg8IJPl7jO/e7G0w3zsXwBjMtxSYDf4Y4VYkmVjHMSvBRf8EEa
WVN7U7wS2yalvcwMsuc7jT9ET7eaFvlmJ0U8ycdy4cVz3U4ou9OerBx4Qxz/N9M4nw5SdsdZclxS
8+3vkeo/U3mmdBt0yr2wkxy0oOsGZwTlW0TJkrftTWQ0+2cTZf1BVl7sAHx4vpTHPdL1/SGzx9/T
8BBvZvfinF5lRXCLyOEMEnQHEKWpzuEVgbDvzNq2Eum35Rk+/+WwO8SX2/Mha17C9N0tLy2eKnQn
0AIGU3EK9ctW744sdTjKOU1KzNGfv4r1wEwa9b6LSica0IX0QrRLdTwEHVPJJlOfAdTY4dcyBFEk
WugPtprMJ07uQdOhSkKjmDyCE2sh4/U8KWzKMQU+y/u/gxMo3cDzW/JRezLK1wNOJYULem+9zwR1
w/uU9N7G3XPTgulfNLLGnPpQkOt06eonvOXFtfNZ3sKIpdrE0bh6DlxC264iQ7aYWXZ2nH1Ue4ty
mi0uvM/8Wyu08cy06sZSGwkhZ1At++18K5/SHQ1HOmFx3IOsr0W3vlbfOGEllqF3Md93WQ29yGQ7
IxsBSWWaeKUl6ha3pVrtH0wb68sTv6Qf725+1v3aATlAsuNPpmOgteE6Yp5uzdBVtTqyJ/uDn07w
KS7kUWZ9oEHIR4Nth0wivCxkYTfpG+eMP98TdlqOZiFYQ7yTj6/z/+BX1pKtf/QsPxiU1h4niiqa
BvGxthtBm8pm9QRK5snDuzyC9sWLSEyAkSCUBbOoDFebuvFzxXnBx7D/c6v8X9g492x0FnF8vdh8
K65AFg2uJFnpP81W7k4lcwf8XACN4LARShMZg7iQUE+X12tDK4Raufv1uDt/C2lh9NIeaczqeBRn
OKP/dF58krwwmeVUDrnp8jvJDvOzUCZyQWSxin2WlZnS0Q0Ev1NfG8vP2s9SoAQa4VUv4FU3tQxS
cCiv6KsQkvip1gafn1AtOZ/owvuSFblEs8eByk3c8NdOi9TQJl1AoiB8xeHfY+NZiYv6XuMVc8aE
L6gpqJESp6pmINxQJSzET9yAF0pv54VYH1ASIncksTnHFH/LFZcXmQ5FOm2kciarV2ZVSCmBKmvr
a6/v44eZVrXb0HE2+eC/uWSW14Zb+L63+/o62Ij3mfnyLDcAjPbPjsZErS1t/aokSp6vuHkhkzQV
XQppl5+nJCN4ZFpm8dAnR72XppNrjXTfQAJLjTfMA0PoBxC4gXA3EjMchvfEBI/2uqy6jw1o9OxA
+xa0aFjh7ntCNHxlT+T4kTakGfKO1H+v8b2tQQ/xxdCTG8NlTIMHHE6KC+1nKK+MjvwNDs3OBB8x
E+jQ5fmtiXHkViGPL4G5bwqpvSbMAKqrrKQ683SW4/ZNwG9r75bweO4t05XqSDLjgfiiLd+QHQRd
pguv6ZHgaBXX4Z+/s9Rj56pjWVh9qSSpFyqIpKUKrn1AjOXu2wEYiAeFxM1W0irU9UnywfZGbMHr
DsUx2e7WY2D77scdc17KpxcbUs0RI5qxN7pCdrBSXO4tH97PJTUSJrOIDVW/NWwdriEO3CmPCEVr
DD/nyujjcJX5GMjYhVWPEc/6lrXWfxgYsoT3AZq1KIhwxE1NVFmH+uRui28cCyFVfTusLouruLB6
tF0P2RNuscmZcC2zhVk9Rxdn5v9zXGcuGdXscRA1OofjC9RDXE4frDgF27mR6U24cY9BKj2AUqKT
+00iHvSy0E4x6vIKxh59qkQbHjgQVdyQMFceQ6Q1CRLHsvQfKiCj2604twSRFWadRvwxTknkiQ2j
5N7Hvsv+LttK3GFol4KrM9ID7TJ0cD3REjQOqfc8USI4Cw8QUIu58coJfJBQlhl/hOdJYaBiAGlM
pW//OrN2/0ZRBXBcMKbhzuKCH/Z8jif3g7yPWsbHl1MfFKf7nExNyw0CZia2fe48MOh4zymusRbP
5DePhFQDXnaLnEFJUE5O3fTgbKiQwSDvh327FxfCjd2yHxA/B7OtrnXigBO8Uzu060ZDSpg2fWyT
5keoQrVKg+3N+PW/0ge1QWuI6aOcoLIk2ZxpYltx+2pqDyM0HF4QcobRGrbUVTWjGp15tAOGKvBH
1BA8BOAm5zpfSAEC8/8KvfsoI+XTkzW6dGm9mqtZkruQZTBaoxwrK8OhpkKnB335XudsQszvaS8H
4rg4C3kRagNHKCPF0cKUX/77/akQYmGVdU+/PZOaXIcuYEILsJnNsWyBhKR0W39VV7FL4ANUhnzu
NTBlmwL1PWffYCBqxsd4yYPBTMfrbpGWdVuipUhglUn8iq2cAy2fqL4fVq0ukXnJmAFfl4EfeNv+
Dxp9gyb40T2kRgqWuS9RUD5aXTxDNAGAjfv5lIBHU2+DNrWr/fZLi0bPNlmcqP7QUkSiHtrDYKPQ
GCINxjkZKsO6tN8Fh5Kr2v5jnn5KoY2S4Klum5MxJgkK/9j/lYMej4sW6wJECbrQJDcuuLLaS6GL
sTS31hUZtg5vHih18q/O7zVY+Ei0X2YPX+2M0azd/h913bjliKXmchJIKz2xxUWtIoiTdLN+gNDh
PzyiEbAyYoy3Kr6wwQspCbQN8tx4VY2owCcbq93KCZ3PAZOlhR53wGfXIZK3e+7Gw3/XbceipbJ7
L12BmsuZH3gIPZo52MXWkpMkarnlENDyFfKckYIe/loQhE5tfmnm2dVT2Are552WpJUdR7IDhUNu
860suKFv5QjkPuWyXjGlb7rbqc0uiglmxkTcNKgDly/YNld9mWjxRRAYGQ0rjEI2g+KkOoyGZg10
0NVPrYQvP1dDlo6FJmJjDMIRea5F753GrfXyyfpzZ71Utx0vIxF+5HjKtFoGTvImm+L7yeE/hIyl
Z7IcQUG0M9FU6LRaBXD/38ULbOb173sA4PqI0Kub3Y3/z4bbuDszxKazedkcqZfzFagoAYCwCErn
hfxHXv7q5jrOFxbRI4ymZt+VcCb8qQgPw6RP6TIXAi6AA+KDZg67Jy+bXj38paf7Ze9JmCiZmOOq
+gKwdv4sK/0Anx5jARtoXh+a5kDIh5CPq/mWs2pNX3B+ALoOLkNDdglVsOrFAx2aRBHRYnZpkLcy
HZH/XELZCVhweaJI9c4KiOL4M6xzes2R7QkOa65cJQMXrP6CIi59MnQwJpElQkrj6ILSqavL1nBQ
Ype+g14RbhrLVOwd/8NT/oWG3OSRwvr7jKKTPZ6Gy5ZfDCKN93LDi3h2MD/eFKSxuv3I+g7UWtRo
EpzZ5T4RsaQN30h+DvXWufHtnEVt+GxEkHlYxBcI2OjZppOZquJiPe/BU4A7WKlxAXOl/93yCRu7
RhqjNlhSgcuSCxNAAGwG+x0tvlpeSL8mn9aUJSDR0y5ZGmtfrlrCGJSOu94rorOsbOC4wDGzijLG
wSY12fz/cOIIx0xaQE7O5cftr+fZ/vkUcgeHCP/u9Mk2XMwydvZeEpll7TfqM6BPc8O5fd+mVw2C
8nUkTfG+WXcWR9hHeTzxVUYUplDatvYwUkhGTGkaB0p3da4YBWq0E2/ECcJOMQ+pAbUhXPFuabm1
V1gVfMwUywFyhZzDuIh31lNZADtQUmLMYOuir0shkR4mT/MNPKvQ377pmgbQeopllHtmck+r7A+1
jU/Cv2Q2gR5c2UDRKCVDSyjrFZMRmt+tlfwvZr9dbz+gKk7+1HW670Cr2aHhKGXxQucwFoYvfX/F
Csv+NAJKHNKO0jHeMdTx9zdEo0A9vk1LLhqM6FwwIfVDR+0OOirwsNbVDVZoB9KvKFCVRMivDEYU
/Ks9mlLQ9tr+J+KDnfNLd6ZQTRfJ757lyLtaNU8gimj7/82BQpi6E7WwZA+00XaFTT4NoydO6bOa
WRZFjA40N738l21jtAHBvsCcKRWDAakr+tXRetb8NbasbdKjdPb74AUK/SaOZudKjyNVW9mVOTa7
Ye0ddtJOpNL3FsqSYrr1OqBlcllk5AlSNUxqdJPTDGbbBpQEKLDSn4in9idgOdxa8qD5ZXgMIGWQ
Hfy33A8wpBe2paOgflW0jK8Og4oDV/pnkpzzD+J5wtRdZ4WfdXiYqioUo2Y1IEcp/ont8aL6fMJs
ADLZafPHLR9Sqh58CH722t9HcIt3lQDRfxGGN8LwR3fV250vRFadCgg6POK9Rue8H93eMdb7xInb
XYtDY1ZeGoQK6lbv/0ZScMhUSd2/04TY2CV5/OQq8cZu16Bz8hzVQCkTuD1p2+Xsoo36dIO5RXOh
WI0l7r8DHv1ftQ4xOd4D2asfaQ1hrnPpDXJ8gOom6DvoXCGGLscE/jK1g7JaDVVM5S+J+gLkxbaC
7tERQ9cmTeN1ZO3VztQX8kTswn4fhfkjD8jTrAN/m3QunDGRQ5ZQ3y/xWDH5WRvTc5dknvlkQobT
yk1GnUnd3Q0nQzMaj1pjwMqP7LMm+E3UOLhZx9ARvTA2fjm16dcTq2kKkxXL4Tt+STbjZl5IRweQ
wKBQ4L9ARNQ9VU9BjX3uhzLz8IYPGDJ9c0qPSbpV82btSWd5YB1aU8o2UQRQelBxI7QQ5yD2G7Du
59SKgUhH+KfRtRn73LiesU5nBnZs5fD26XcweZzewpH59Fu4eo3HsK+34BObrQQl56KWdLVE1WMd
7yq8PfyHoW951NWSj5kmhsdNFNXpiSJhjYtYP4wncBbZq7xOEIYvR86pKit74B5YbYlw8tmV/teX
CZg65YoDD641JzEJ6c2BVuLxKaOrLnnEHILf+3gkhT9Fo7YS9RKyhg7ixwoenhwyfr4I/B/mnL8o
mzdeGSyRnuEAjDfW+YBlhBpubyYeEd49epGoV/fXnKmZoX8YecIuPVlnMp1h2zjKrIgNLjHuaUex
nNOgoDuM9SoP4hdWu4yh0IzkjBzlUf/MPm0EzLe/h553mFr+xeH25A38ZK5KyFSK5y1vqkzcGAaq
Z25AR30RP93c6kms95jn7UmqMvu49+k5+ORVp08NggDabgFSv7by6Jm26J6L26V3yBqrOIxCxaHI
js+rLZb37EIoP0xEj/QiMSb6/oWXkxNN2+4ZQMctoH9kfNQMmo3nCr5Td54OD8o+0Hj3WY0RaBlv
W1aD61+su4mtGbmZEPJqLWjKykonbQei57lL/Zu/6odweYfAafI9GFaf43dAwqj42p+D6UKtueBz
TcPjl3Me1wLosqVhVesBumpeF4FUt84jcjBHmOksia3X8p4EVzp8pz/ygqYNKa8OOcPEgz9kA4T2
krfw64lClvnfC0vvMQnrm4hHrjwiDfqWkXBRvtme6XxklUoAiMm9ryZO4K1JG971Kc0zVXAFigma
vOVoyI5PAqA9xS64kcQYybdE8T4wbzstvlx/Ed18FO2F4+2+jK/QbhWAWUuJe4TBCLdb2aWnWAEh
jWpgqj6Bcpj8hcxkTxltHQBxRsHbNHxjokucbSXr0BbiwgGaYoqDgYYitqaj19NisytvptIy9h+p
nv4ecBe1fNRizNxokAwHktb8UHDXIH+9W0Y8cB1Yl1fDLoPxt2CEsxN5PvfVz+7l2d0ja2pY+V8X
m77/48Gr17588lHsHsmNgSVENRIr6lYEanLBjGZtpzfuIZnOhQGqMj9ZQtELMZIcbt3zl+nSeqpB
JLk18R2V0vG+EVgfCOLfKxn9zVpN+VtKNqnuAVM5qz0DR3OXT25AqrsAmv4fXsNfCzcixSWfgW/h
piaBZNL8tYhkkb2RYmSRpGYRfkOmUVXtVkV2Ggi4ynZ/fwkSdQMnKm0nTqeZ66eyRXE7TGTYX35L
J6CgjLigN6DdaRJbALJz9WLzXM0eA/mKgXOSGZ11dQXDljib1Mk5LrybB4PBPWlI4amBCkRVIpse
SFojKlxYMosgb/pgUVCj5it3jyrSUrK7IHAxUByVw5HMadrku/NNN6SkS1H1rq/1iSE/Z9v1Krse
xQNlMmgN0GkOyRSDtSRDIMbFBJjokTcqTSXEVpWZZd/2umhz7f4vbimPHibHX6lyO5m0o6NW8v/C
P6+OWUXPhI8KeBnt2ubtxYJ3aK/zsquZvax6e6LPLtgRCGsff1emqZRcDakqKbTBOzVY82w4kHvD
PGn5uZ9PCyqXp1G4yLDE7OgGgaruv0vqgb1cD3MwT97ObR/IqlVYr5/jczhN4u+tancEGsN5jqKS
SLlj/3U0M2rXkBkt68joRnGr2EzmZbpCgooXDuEF0rL57Em3hMwwzxlkyyZI3EcmowPbGagmnOFL
fSANv83udd/iFLYI3F5PB43g1ZgWjxOGHUQVVfbk3ffPYAynxKjDwa9bUitYFP8JKlJnMsV2fuAV
H2d0pyIrkQy4AmdnoDxU+BpuPbwwkUBJXWKgdEB0IpkWAnfPsihv6FHBV+E7ZpIHaQqnsP0DBKPt
C8tzPUAWE8K6qzdtKNGkxl+7CKTBVMZeF2KFwQfELPtIO3Fst3qEY7KQ4At8CDmzfovPPsCtSYDD
1h8Hah2nwi4+AxDIqKbjrvYE9ee4J+OCmM0kV8e2BWtSfEuG5JnLpQQ+hNpPceDGkFRGBpvEfLn/
s71RbyEtLcGv+LJaG5zGbcFgNohyd0PoLw7tCdELHdTttELNpdJnEKFU+NlnpJPTeiXFiHz5HdgE
2wbo6VMqwNP2QweNKZ7q1jtLY0oAjRj15uWcLnQSPOdPvUHX0JCGo9/gZ/nqcF3l9+hDV3cpHOqD
kZGhCIgPSExHJgT/F1R3EZbc/vFBDzzTXOaQyfQZ0hbWy9TBhQA1mm/GiwBTthFwnb9Uq97cZxht
iKy0wQvl3Uj8SJqWjzORecqe8PcNbuW+N5/A9DqIPINNi9N11OYtJe2orghPm4blHz8Is7d9wecd
BQVlylV5Dq3zlwdwyalhUxun79472BMlfyQRjgtC3EJ7T7xbPwlBLCoXXeJGekwsIUImrtU0948C
aqizDYT97kUbm8Uznf5WtMk3N1vZF93Cm2hokB+JGnWXM1nw/Mn14CCXZee2Hvbo+Xm0aNUX2ACU
IOk5mLGTP7vV7GtnovtezXfrfkdMXZ8bi6o/k8qsPymQh0cYdIJUny2YLj9xui8D7H6l+rAj07Py
VjAtkRH+/eEEauQuD0TdiRaBGTu3Fy1KX5LUJij1xrR1rEBqf0AUUw8HxOVBu9dSseOdP6pIduNf
rKIuDUhXkG7oNo9UPQ7Db6r+mCuFFQI57edvK/J+zprk25MlmMOKvxKt8P4IKsWy99GlZ/Iescbd
WcD1f9Jv6sTiHUIzhPXXB/3pIxe2Db40sUQHMnd0XkJolFK6azhzH97mjMxSkEo6bRZZPkFRV3hT
DlrCvjA+XUkbDO8qeC1ohu+M0oJozCce6cTIQ/rEcjY5L4GMRf55sYFPjA0hZyFvxxrsX9SBPVE1
6h9hCYdzhrkW6weVO+rtNQyrPVf9YVQ59DSa4ucEl8QQpablGAEHUwrBmHE0n6C1UOWAiTyS64CJ
et92Cta9qu9Lhem2iSfQO1LpY/enSNKQo1DcL8wyldkhKTxyoR56FPPMNzivFhVddrZILwdTfvUQ
ErodlMiuv4L+4grPZDKewuG+mk4UzMBkkVCbLSo6mQ8+4mbOq5Lq0A7R0noIFKFCzoXy/RUJ4RVi
9nK9TY8ZXlAM0pBES4n0YW0r1f4bfmQlyB+ZxcjbAGOK3eZhAQNokSZNDHH6bxtBd7RcpseZSBAJ
eOOQqP347flVxxWapJ07mjWQ9TjEViiCsZzychnfdQ56v49QP4Ctm5YOTadFdXPaFsuu1ae7+nsI
9rAT3Me0KoczER+7po9Rvh9JPIG91REkLZAyXdB/yLz5QWvNUbZfu44b2XogJ95bK/TyHMxB1vMH
tVsbgHsCQaGYrlpYC3J61c4qWWycIEP1uiwdmCI+O4UG2XXaDEd48Pbz3832hHwgkBSW/mohHW8F
qMMoVnIvT7kl8o54q139u05TChW6E26XSYdVT7C7ti1Jl+f4kq/WglEV0Hh9k4m9HhRxKAx3qhSz
8v+8ZltdgjcvNmyBAiubKDhbKTxz6AUAEZDQbXtB7O90OaUfyBDDCTLEz6nDToVYQ2FoVoYXIrne
Lua3YgCgaOU8VLJ+enFLhqu+jQAvK84TX0pDiS+zxrZpyO/JMLjZBuPVC1LYtBuqQL8y+JCquius
wK/BbQ1/c3ViGnXrTEWdOX5Bn9iSPcf5Z0682WgDV4gzoZG2gk0UzdWqo4iL+D9IHWeMUQe+h2DZ
HGNySjGoDt1FOotBvadqdtqwgI9RjkyOUpQB3j+RD3+4Qf88Tt4uCdXgd4EQNxQ/dizpgYht8/kO
AYq5p2yxY31sTP328w6SaIh28aBycEJg2eA8k+0o2ony5DpMXMzzIRGfnj0PiDbbAU9kBmqHEQ+/
K1t8jahxy8dWAm/el9qrS63IVgSY9dxz60LG96kuJbCJf3gEac8UFnxbEVIV+4be/ExovaPFa2Z3
jpykQIJzHiyBUpU19Sx9X5WkFrvqCifANZ2t/RMTsV3raC0z1oURqMt3kQWaMPEinumUXf6NTBA3
YXKFjvNwrdQVdIK/qCf/jLH1pxqdeHy6XVa8U6ZocMiArLv1SIjwUxM49r0e5NQ/KhJIAd47inhb
OUoo6Td6jPi4SfFy3mzPdMUQ8qzAXh2ZvJ/nZl3lX1JGUG8yyLeDEm9tOXlizCwGGaKdYljva8qe
N+8v8u2yBy2vHdSvghma8ZH7VQBYmac0XBJ72GmXpsaR56TmzSluJy4xgSocK1h6WkfX9Kr9Vp89
MwazhrgNptGUGafk9efQZXzzsnQ/RkOqF3JJKbjr9ctXKjUbF2pdqATXjSpYjMwLfDxD+a+nlXYF
J9/gaEio2H5RlDxkPv+yL+KHzzyI0OE87sOHHRB17Cc2RbJmj7p0xL3B2/SMmMI0lMgWLlh/Pz/a
TSfDv4rZj2Q9zFxi1+mlFJixEJ7TNIwrbz2vvv3A5jpnvhOUb/x8ZSt1H1O3uuailzCyAK+KW9gP
wxB7yS+d1uHvamhc5LGXwMO0CLTH28Axlaubbl+SzfwA9RuFgP5N3GQD3vv7V+Jdz0DBkBcfxTld
nT+xbV0lDdP+XI5aTnn9DMZD0v2gdVEue/SzRwIeQlmuvK+k2KUdnVl47p6kjUvHuZWJCzzbvknm
LG9ckF3hJl6kSScc6ZbteSApiQupzJLp/3oFQV077eoPHAAwD1r9D0dbUxBhQsWS2zrdK1fggDyQ
wjAEMOdjKf+ZOqsoy8PRBEr6CjTLb+0mkDS9CIMupnSw691ONMyQGFtW1zEMpGD6m+7ZyEzYTk8u
gXioqiAqFDr9S9lG10G0JjmoCub9KBuHVZ9AiKvge3/GOHCQI6gd/oI2OXOydzLgN/h4ocCXRdu4
j3xPbcSP7HLBBLqi21mVZQMVQoqQ42UIIKKeSOWL4NsWpM/bwvyo+24mtmI9N5gXXffEGS7PCTDv
cynYCOCByua0r0Tozsa/1VXzvXlrUfogWqtMwGjrlLhm7Knw8zitJmW/klGFbBK5QFCOthhBc6ut
zEM7LS8U0N7kFyW25jhu09x8Ewyks/BdYOXGHp10jBvdJEb5THcijFuhwKjWNkxL93LdBtGZZbvS
PsspsOSMMQc2odC2PWcSI9IK3DO0cetGDRO1fUeoTzduwEK5TlCyM7jRvl5Ext4jsu3EsFAG3leO
ByMQl/WS74pheK4Gr0dMvYqWsDkKQ7Od1dzpHDl7+xSVXavq0Zo0msHobJ2e8wwIORFP4QMqPVQm
pAyg8cXuHZT0jP3xuBB8q9bNANVGsfWEK6vKDlutSYvM9Sbf+duFTAh5Dnz7+xlKS1iKR2OkYNNS
XGjpH/xdfeHF+v41NJ5Yb+bhgubORdMO4l6wpNYJnUZ6mrtkQS4Gi4DwDN/vvHtHAP0QTJLWYI6I
9k95/fDifVH0UZBPAktdj9o4P19KDai7pF6u+mRGhRI7+L7yxynO4Ze+uQgxftAw/oakigNZAAgM
9Yn4lOvCJaUOkaYEjeQ8LdkN5BOPvpUWvbvQmzIFbitiFGKr1PZEULRWUAwTx2RfpJqd7m2899XT
pLjQS6jdzziQeRujskiScsEQwp3YhbaZ0pMshFtwjFzoZwCTe8gg9A0DcIZflDbA1aIWs4xIjzjw
mrgzkIgpr3p7JZosy2QYiQb8ym7iQFhriPeJOXs9wR/kIFaPktWSgWIjC6UHJzQJk4DM1P5NverC
PNh0lEjU18CA76nVKvEPXaOFB/kKIa39OwxtygIeZeCRpkb0kJFYLImzQBtWKxAE4mzstgpvnrOe
LFKeBuBbUMZ++ld7JcFO4s29YEgNvCumju7pAfSkcdkJGWen0JdfXr/gH8qxE/e8JyFBkNftOj2N
kRpgNbwsuVY565tYLE4BqaXvbysHIjrBBn/UZONn2URDU+b98E6iCHu2d5q/8fTkh2zWKHbOaJg3
Bwz5Jp7NyveKjk2mLyyH85AHYQt11uSHuHa/I8GLPemBoI94TxkxtOxfanlvH1UcFVn2Z/xfI7VV
KOP4zS3hXtlVy2jRzvzr6TlqyIooJbhBflIQKWX0jsE1D+s+tOO9P4BQ09DCWC0UEA2JXrsEvWIU
93aT8COcXDD+VwbUAYbRgJvn32MiVqCCNnOcFLXaN0rnUJf/h/u3OpEWFhdFOzCyhVKEC1C61omX
NT94naP1xpOZEZWzu3HjogrpojABv/H2z4pTRvCIoXBDEaek+PfEONHIi0PHzELjvtkn5G79JfdM
6awEpudDFXVHWFoGJw2dMREbRJ0CdYbFr3w/BMF96X8/VNP+Vvzd9DuDhe/EdXTUiahvtGsr4vbD
nPq7GkONtlWPluebbu9JkYFLCYca3Tt0V15U5UST1rUzAYQBiZCGpdIPnjWMqZ7+vpEkCIiFlVf1
dWAvR2bly2ZHsSI8JyFYgds1w0//e5FZqm+MyIc1osjXuMvMaYfHC1ohzAN00QFhYoEJIDrm/QYa
C7umMVHhE7w4vgRjftSQfeYb8lPqEy4UAZkL5UgxGW1Fhwn3P9MU3XY3/uocog8hyf5ezlO/E0c8
mEs3rxII15VCOsBmeYDgD75rHRtZDxF+DY1nnOorUkhWZcSX1oNYkDc/DYUaBKjSNJsdYJE/mNBJ
IoigXdGTN1rOcdpzIEKZacIF/u+Sh7GpkmnGYvSJP89vP9tgczgpuHMVYTcFHh1acObAcssQpBYb
oFAyTk5DmFV5YcqO3yULPaM/F7IwJRbiagShtjNry203+s1TqL57kTeBqNdPYBMXtt4EciXsGqNx
OpHhtR2bzn6iJ3yVzmWjkGBwRbwQBMcjqD5cueATssoqlZme+vW9J7wCqj7nnyqHUvwUgnLjAV6S
ClaHxrGqM5n49W+A0c67ROKE+bdhZllZFtiopre3VEXtONimF1AcnrOH15hAowgWUqahGOU1kqZq
2qmpmV7be58YJ+BT/k0c1HVkxmzdQH6tp9xwJf2iLcs+L8tJAyyBuLiv9Y694CLIvxsOBP6vUNif
Up0jhiRr6AmJP8CVk4nInUfnc3kXr2JEBFelASSOkd5EgD7ubzjImz17P9Dkgn0mCius9h/ZiZgq
TD4Gh2/lfyK22/TF4tepQUDnhUh5Tn4vLw2UpReuNw/VawsRcwms8IyH6znRAiTKE+PiD+bEGhIi
x4RCBOofqGEdArdrvOvUqqHFzEKUPTlueUD2RZ7Ns3X1C06jGermEXneN+ffN28YK+0VMeJ86O4Z
dteUHi7UzSVSpTPLNySf7PntXC64pXtCqJP95+rZxifDFuUtaexzIh/nfwdTk7mhrzLUiF5IfJTQ
TDkcAyOz5zik9HL/QMetIloZUx/vqzjVlRixWyIaBZQHT/Q8qF+OYwgFRfhiylQ3kjP/seKKTMj0
VpdS4ZI3BWGMoL2PsHNCrzaSlQ5ATOEy5xV9I5UzQSuTSxNtKzPgJ2TWoqDJXX8t9q1UP6hntXKl
y2xw7ijtzsh08qQGTkJkGZzL2uWEFn+w48ntNWBbvjomItwA9ECn3ep4eoDMi0Ukjw/CjNsLN2Fm
EfD2zxGwCs+ZeLNZ2RkqkwGodY8B06E9Nh/0pGRc7vddtEx007Ua3TH4C74abMA9ptuCetYmdWiq
ZtHmjJocVYMiLRr3nLTtXLDuKmBAqJ233S40mqMcTzc8BgPfzruJDIYP6ixnASCSNbxCxBjwQgoe
vsbCpTiR0rIfZGLVa+sMaI7ai3tyRHcTa2GBf1XbqdvLTBfsubouad1CtJnI4DvFdxxDFh0ryJWP
9LQED1OKYqpmLFW168pPBbfe9UIqyS17wSIqWiH9nqU+e5KgG9SXcyN6KDn4XRPXLOY6puxTArA/
bOyUyNtLeMWP8BUDLLl87MXwUYWNfhDpGhUUYqvX3e0kw3rbuKQG5Z9DT3nqH2aw9njBctORw64E
+2gUIPVW0ItO3WPlviaYI9M5h/bwYjoJMSa2dj60788oimaCQOdU2MZVvH3sEJyzNis950zXjQLc
aADPpk89AyG/OgClkV3owwJgOcGxUm7hkbKEVC2YJsYzL8ZOAehkHIcJuOfz/8/0lnDUhviFyONp
DUQ3OkRyR9fOhPskT42Ev4uifHvKC7jyrb7cj7OkyOn1fJqHT8zS6Q3RS60wGtx8l5mFxTHHrTW0
9kqDc4ph4rbMwmGrLd0qT5bjyqyM7ZuDDNr6DefrbggXWZzKWCA1doRXIx93EkoVLheL/mcM3ccs
pVP7kmvS2q3lzM1pHTvBE3ucah7l/SeaZNiZ7ZKjmiVcEpo9Fx5aEyDn49ccfPSfab5+HymbSR/x
kbTOUasOYQjdDbwLq/SoBWHO/pWuIoBk+XRvbCf92megdbrQZzIveFgxRlsMnDKoCW51u41fkjl8
x1t++4/m1mk0WKxGNRsB6ZqoE/9P7wRNdRa5RHI2t3Y+TXze/wU15Gc725qG9Jg9MGlht8iZ1XXz
CFqMN4BR3eDs8g+0r6A1jwouBDMjuD1j7RbN30wZQNTd4AtwsTMaXV+rXU98WkQhbS2ImRQlWI7u
EoG3j4Vqm1+IsEiAtQHReT/0+XjjFP/yBQ7GMPhfjNNPA8Fps5BUgJ3VVGfFmm3az9Mu2/dRbnfd
jMbTcdBTcwgpX7AsoIPZeSmzpATXgq/dHjPmJ3krXfGoopGdAQ8aqQcH9mpUunbDlX+X0/nWlwPs
qeM7UFwk6dZ4630A0z+VbL3QVhObyPyS9xsoY614Y6Twy18rIP/8pAvaFb6IhopXqmuLvZFEIy13
VdAaJ/Fh/cl8PGeNrvtuUU7w/p1MotRjoKt989ao4a75+Fa2jkrQOXpjt/5b07i84Ce8i8Fg2KD7
j8or11+vkFavFE3NS4EfAPFntoWifCKdiXhfgSBeS4VHKGt7K3CHKhCjEEnkBXcrjOmd9VLg7pje
ER/71R25VZklcT9BkKVyVKxgSRdJOzUUmHi1OvpIl7Aropmxxf3h/fgmLxdsfc1aTaqWZ6B8Z1RE
BmHMoTsOn6qsF7Qpi6uH5p1JC37iQM60y22hyESQpAeNBnsiPDipRkxG8Q5YPSk0V7Z+6qw5B6Ld
XkYAIRS+pYgeV4JTK9EhHyoT63wIzKHrhxKGTFULqWfiuzVf5KY1PmmY9bSMNw0B7/ApldKdXUv3
um7eA4O+HWyhKmfJg8PfusjcXiZHbRtS9DtXMJq/ay7vAqMrwTxYE9P3sl3jArjlNeI0dwQlq77H
L21SU1NllKSvCVGrAf8UO7JVTh7Gl/jMSnoJAcFjV7NLUJpPvQw9lcIaJlXYcIZin5WyqHgvk8r5
q2SFvA5CrjAujJMomRboZSQKln1rJWRpZpq0URu7ZRABWiIn/hKMO3sIk4dKkFrl/l5aTFUQGrXu
n0V05jV3QgGU1wGc2kNHu54JAokkTS6OvP3EfLZwVqVF4Zp3nGV9Sqgqp/qdOg4KKcylXxJbWBTB
nFYT6M2QTNEqsF0H/4LvHYYkNGS7I5zqCfrwUKP8xvZouyCJ2DIkzlTa0ibPid5dlkBNfqszIafK
ty8vS8NFrJqyNgGUQ/WaLiUnfFIh3N8LWH3Y35nfaguVb0jVwqR3zeJvOZe8otkLRHtWESbyfalj
xnBVrcTIEAoawdEnbYM79XDHyBucKttSnf1H39Wd5v4v2z2M0B56QfmCCjRyczyrgzf4nrAVaKO4
cZASjYkQUiLnC/gzuL8EvKn/8JLLv2YGmfVsYYgQalFK+Oj/0uxrfFXZnoEdD1xzbMM4gMkB78bv
PKF90AGozE3jrckQ3v/pw657mAlSeT0MwjUfYBiIU9qjHvdVaSycW/YYS+QcE61z5nXaDT8Nbch/
eyh7n19PDSh7xIx0udY5GDPgdh0Skj6zPmA/yedojWsAU4CaWrBapV/JpWsGTOD7YmAFtdbAsl/I
N8AxYocOkNoljzdBHWUEM6ldt8q7e1SuaaOwZMi8kzz9HRNBJ8X3T2FCLb9gCBG1VqyJPO2zO4rk
Mf+Akur0NuG2yORqoG5VWmJ7MunKZeVzIaFauIoEG+zLWKaTNx8nSl+NcyWw/rnG8TGRVeMqgg0I
fPH21q810s4xk/tIHC92bW04wscAjfMcV8mEVdF3BezKxR7kHWBznna9rWSEBpMezvgA3kYoiQQ9
NALEIKaHicXTt1R53jN2LxGoQgOrKmLRmH4qUUz1TXN1IHDtI0gkhk4XbC744a38aKCfafrj3Na8
1O04vkHPKquLEWsfkqEjYoxf6tt4XijAwkwc425lWuMCjMDrpIyQUlff75qmjabVi1obE9SodiU6
a8/CJZrEtJ1XBiBbmoEtxix1fkTCNKtXzeHHtuK0qJIzDhp1ZhyvTlb5zEW6M1GfSSh+LhO4BlZD
pwOM3VoNMgnnfRB39IXvD+sjCIDkW3yxnc6TIgbABmpFI7Hnp1ZDXzo5mulmI68kOHXi8ls6rcE8
00xXOU/ilCeAcrLNI8DpGw6FhmFyUMq8FCwHroasr+TFhYFoTbuClM3xPmoeZUOAl3xcY2+MPX15
lmNe723PC9T2bNe+Dvg2NZCiHgYhEigIg6QQJycwdwhs8AdV3rCEuAGQLAB4arYNVYZ+fmOZGryU
4yLkt6u8uT7sP0bwYHXKPgcZqms1ZBNiJYVS+pWrvdGUpxseNpgQG/x8+YdnnttGotHZZFGL18os
LnmlK6hzlR6HbQCvFAQZQLC0Q/9pDRvvMsuDAK0bwiZd7K3jQ2aDui0eXrDJmgBVmS4N+WpQ8URi
0e+4O9DDlK0JlTy/Z8I1r4Ovz2mbySO122uqj0Q/Och4LFKqG2kVH8o9tvIj1QSo2JnKiaN/NwWc
bPtf7mq5fuwrTXnZK06QRgr/rF5v/3qU3kivQ9P+zBWyW2QfNrjiWaaeY08H3zE+0XJUrT1byT7m
jW/iY1Jg/Bo1VJ5XrcluYY0p4Rzv3V1LwJf/QXo1Nc1cugxNH0iN3KnG54M+/KSbTTQpr/ndsWFm
Fg8htrq+ZEFJhQAD+baEDuJeE5C/0Ux1gjWrmeIx2xnGzLXj9kyhqUUXXUcWiQgJ5EWu3u/riDQU
UmMdscknzZHER6xDBRK1abcV9s/cUW0Q3v/2YhLujEf+C3bJfVpYbIr35RHqwpSeqGJxY34Mah60
aQUy8fFR9m2FuMfn7757uzSks/eYpD0ioDGsUuhAyDfCjycRcFrCwGfq1EW+7kfMDObetqSkYiSJ
YYSGS/NlYTXSLSg93eLTBBAInj2X+ewUnounQpGUPLmKsxeY66L9X1NiHvIW0/UX4PnN2MqfI70R
zsnSyzFLpglKir5PRHOQztXuJwGdQ8uW0dN7Pk6SMJaTMvBt3NCpXofFpahrK+pPlcMrwI5qVoH3
BrdGLxU21R3ANTupVny+MvGtauUARCtt9eAxZ1VSfRsCmke7BPhPMKHzwR+l8pqepNlCGMd9JWTS
lklC5SFza+r/xHSQFrLVILuF0Y8eInYmmwnQosVviF0FPp/I5SuJjTbbebVCE49VA8CMYTlxaJEA
qFgwbxUYK1we/x0W8aeailY2UxYOl0KAWGrRuIXHhca1sylEqaDv8ujusZoWy1h5nqnI6ksjTAGU
tk/IUVvi4waKQSp5ZYX4PAs+6fsGxoHKv7YPmBJs9h7JwwxyX7ftv8ubz8vYf6VkP6kM2ue89kTL
WUvU8v0yyzTSKEupetKSiiVqAKjz6vCcFtuxaVH1Zec/NBiO+Pp85iIf7Ch3f82CFHssTZWYoG8J
SqJAUgnDuq8uN0TxEZCPk73nz0aJgk6uxU8zWS03KIhGFtKKLIU0x+E+SEDI8JiRkTYiW35ApkCC
YLu3BXWG86Env8MFYgVtUziv+gjrESRj8F5dMDLi1AG6IluHx8xANwW7yAHX3icuSRhvs4Su9AMM
vUYJtSLxYlOfTVabBaIFzN4Xk+4vHKsNNqlHIIFz+UL0FXhwHYrtvR9bCQ5q0cmPp7sJC+irv68c
anL95SqZETlwvNxTR0dwvzGMBpGiaMqHxmHbBAX9JkPlCsn1rEL1si/Ri+MmKcmhsm6Bb/groqIU
1Nlx9b8+sqDboDRUZp/0B8Ph7Uwnu2Bi7+2I9+odmjW4gTTY9LBTYlFa1rt0YPt02SV/hj6HU22B
SWsOE21SK9DhOD/OcYytqEi9aMpINXlmxG3lNyxwQD5GQCYfawvBcE5Bmin5a8EdkUPfBtHXvUl4
k7e32q9d0f3mhzqLr5jK8L0PI1fYtnI+whYsjcbCa3DiMcDHIqjDh5vdD7sYWtdDhDgRr/zFWiKk
ixUOwHmKyc83be99MQ55RnIXTYlwuxLGMjaG1JRpIOBM7XFnNgdj9Vcnzw3clZYy66iL6TUzZGSe
2j3nAMMsqJ4Hr6i0rfU2OMR0Q2A9XHibu/J0BUltk3bW75ycN0puLKnWVWJXBprDiENvwmwzEiT8
AWuhy7Px+mgF2I2XjS8iaZJw1vCHNApymv4ApXXFT/4KpjjkAjeQ8lGWL++btLdkkW1mbzyQQDsL
hjPVKrNrS6fcw/M1q3gNXybm18KEkIvi4kI87H8OBCE5NSYyqEdvCrESynmyNHxlRCQG0gQrqC2E
zL/cIr8XlGZCTtDdh3vgsT3tgdV5OdRNwTVG184wqUbk2nero5Dglr6SbfWWXwasBYJcQ/pow+Ml
KBUPygpLIngHxzftsEOEoOumywTGDx4zoasum2jYFjSSZj6E1HqnlBAQK8Ehfi1w3DviV1qJ7aGf
0WVq/lRkAft9cG4wWbNT9VAFYggmOwFKia9t9a4+Sy7qNfvSye9Ah4Zs/T7R6KEvrKkU45KE8krO
43j33l8PiMNtn+JJn+UhavSZl+eD82jhIEWWB/PTAmpLc0BUfcLNUFEqgjYv/kFay3QEoi298H6X
mwQW7O91nD4w4E3WLl+IYBO7TwEn628XaSra7xQHU7pqwqmRfW77A0Uecj3Zz5HadzAhNIxl+Ra2
PbporEJ7TvSenI7+LQZZJJJRqZQ3lumsox53v/9AXay/sU0Ufkol4xA/+ovwe00BWsF7tNJwlBbx
3tbHBXr9gvH/T24ZevCQIFbfgRsBDVisM/vy5VLMUy8v7nkjKV8Wzz3mFncdLPqNhRBHEZdQvjnj
Fyr205Ilk6I0i8WQMjEHJsb3SC65Zxr3qdNYlgi1Vcz9/W+E5GYHQGuHtk70mYcwHC7vt+OIVqzC
uS8jBv7tcVyF4ugRmWuHsRt59bkrGCl1KS52VbAOLRWm5r8s6aBY1xTujw8ZHuH0p942neafr9bq
zkDi8MNJN60rINh/LgDaTFIoID+zrj+LOFJqzk7GZ3+OQ6qxzQhS6JtED0LWGOzi09SO4TqZeOwH
oqUlT7B7Fqn9Q4QGCjHvn8J/nU0mevYFvt4Swj7EKBfCYc8MZJ02ZJSxmLT23s3cBQBpRCKGqjI3
M8jocPfTj2vnG9DAV1znyZfvjRPIibhuiAzKFj38RsQCYSVpfD+rX3ZBggD6MbrTqv79FbwXPooj
t+OGzKMxj7uxKzz5239pe5jgPPyhjZcnYCcAhli5YtxX55MlDl3zRsuWcXJ4Mya41B611yRL3dJh
4Ch7CLl62Gd2hzE+ijKRdgO+/EGKrLI/sRB3rDMYn7QN4icyJHfKVSAaZ14XubMgge5OnHDf0wR+
NcYlCJe8rh3f5bJzq8VDJqUwH1odRd+GzxitCAw5FwwwE5OGRGiIkqQbkwN5SmIduVS3Q0eiF+BQ
NcfesWWyCsCRNd80trYXC8C/Jpjy1b/k90tbfiVousN9Vpk6wI8rIeRMSd3mBGI5a5bDTkiM3hi2
3nDJBDtkLbySl9RaiHnLuCuWNzVYApipP2KkkN1tyUyvPhUTy948VSWgZMvOUhZ3UtNQ5Ps3GTY3
7uhhe4gCtBCey+V94bFkx1tHdOdFqrWeKUx4leXdPMZ5IcPziJ3a7RvYt1teBDL9MOw+oRU2rVsp
7YvOy4xq95sBDmdaUI594mB6Xh3mHGCFCfUgtBfr1MhYdI8CZC9360d+x0MvTXNuTJ/E9nAQ2Dsj
L/gFyMS9VXaM12JF4YX7G/a99xs+xX5JLyBjByOOYjnKCcwmdleOINnZct42KN/BP+N/Oe/O81RT
5BCuIfUiP3O5qlRsOvs4Ovp91Ac7AZo0RCIEVEw7Sc93Oy7GOHWZdzbEN3Vi/Dbk/ZovhpBd2mCd
SKF4P/DrYbfh1vdVW0TGvFqP4zfpIk+M42oDEpiQlQpU41ah2DwGJLlGzt3LEX60vVYLHiNutV6q
eBz00cyvIup2ZHpa7MuUEGoT0E7TC9fJtl3BKSGREisK7imxiJfEesw3tHTye6IQf669QxAETgz0
TOzaWY7Nl5ardqea5o11+ZkhkladLnYmlwRvS9kIH1aRGAgV50Q+gZnYcmEEJol50fi2R0orOaJK
vYt1fhMUyqZh52I+IBpCCrDWRQayVqgPVzOqBpzl8c5lQh40XGAuYvueB8jOxwQGX+fX2Z+H3Jrq
Dv2iCEiCed1Nu0N8XnwyM8gVBCxJRjVHLPFdQ75lXUuVk/lg530V8xLBGN7zmfh8PJ5dv4b/93+i
IE7db5MwxAcmCGb7t6NIpDy3rWAApDpO3FLI7YrMv6MkfqrLzbNAnRjIZTo59ajqZ2WVpmNYNvde
thY7I0pHq1OIIPxktgR2Zrh47Jlx2yLXBa3IQc1Qekv3h6WnZsddPqlLIg2XGsg46xb9OppSXPO4
SJNJ0MVxI83hjHOpPU5RbhxX4JJHcyv3dgsJzJNUNf/nCWF7UyjHh6YDjehCmbrYYYH8aNCB1pgo
D6vONgQkO1quNvuvFIu8ue856yBjxUx3SnMG06MU6cIKoOjGkeR3DQZqKbL6n2Jxle3fFvk68ii8
ceX0V4jv/H7xmZLF8u63AR8x6bxBZJfR27vA+Rt90DwTnHCSYK/v33NZU7CktPyhRLYA6YzFJm3W
kwB7MTRwtQXinC/MU3zFlm1DCg/uWOnzjn4ogTfGxVR9C3Cw214Fg21Sr1sjtyzzrE1ZxWGsaQBT
msAgbjYc52Y0RnKW4/krY/dyueNLG48dgpDp1JdEJ0VZYYLO/W/FfIgym460FZkZkP+eSKlfzog9
U2tjODOjAAOB7OgKvgkkCP73qcjcReWKu9Q03nPVNVXdQvFrse0YJYGI3mGVFEFrrEBjRVpmahYn
6SQeJQg1JJHDcWH9Z6yO0ROKRCBfqnC9t7dA56ZwrRB89czeB68hUZbPfI2EmfJDYpsjtSlk2Q0E
DaKSn2oSVysDA+qWjtPBp1lysFhC1EyYcX0BPpgS6r6cX3EJXW3dfD4+3kn3AesMMbHwnZc1rI7C
0WJpRfGJPnmxd2xPlM4fYFkNspOmHej72q4jJd4zHnTGA3A/FTKbtrxASVOpiuFI8eHK1+IK+VWM
myDdfwCA5Me/4WwFf+U5PqmURmmCV2nDWD8In2oyJthBZ4y2JQ99blt+e+AkoGZjq7OwWfeqs1JC
sQH0d39ekg8614Zv9o4bdBq1FmmZl7FbuNyDUbMBrfzR1h1gcNSayPfFFQK+G4ZrUoEG7ubmODDq
uBP0JlBj1AvabGMCMO/ld3+aEq9mh050Kbu1Ph8fEgZXicnVb7n3CTsHfw7rlliMtiVO12DgqrdG
zzDgHhJiDBpWPPmvXe4ouLwtWsO9jXXgTjC9D9ZZboqQF1kahVItRQkcfqBbeAdrklFv7vHzSFjW
hB1fUJ+xFaph7Zxk3fPTjCpZY2l0uQCO4UE6a50nUWK9wsX9jrTadauAxVFv6F+amRjT0KA8b735
YaEU59u+qd2PRudZ2dYFJwopUm6QBt1ntKpFvB+KrVurYqiHIkyGSwvfObBNp5IK6/JAbJswlFMI
vjudohvvs5iu19/+ps6SmQSDdWK+OozEFDdYy2Dc2D+lD5D9M2c2y1O4kIPopSy3jJPs9NZLIpSb
B0leslQV8auPx7OklqLjr5f6xmawlFPz67KkxKJ6jV2ST5Je6FpGB03yO5PphrVIRPIsm/oEu7SD
k0JnRPOKNdjZoyDiC4J6xlAoWIg4exTvAwsWW/dT2gwXPk4cODO9QlHi4G9/8IfGNlKy0i6mFe3D
K9kSuFJnD+W0rfRVPcYQMpOe5Cva14XAUwh0uMVRcxmK0PBRLP6kTS+Cg2tTnBVNrNkorqdR4gOR
VD2Wcr9o4NY4n29tKl8F8w6g1WHbB51IaKWeS4DO2V4Sc4/6072Rk2LgYb6uX5f/x0MZ2wOD2Ldp
qQMLB62AD17kXmeYMsvMvcCiAtXU5ZyUNq3E2auJoG9rb55/reejYHGSP9fpdVxaSQBNfRuAKGG5
X2LlWTRAClpbIrsfB9FjvekHkHU5knx9W9wB9KFdmy9+7NYC+qQyLJs9TmTFSZ5x2XqIE242+rX9
yRKHx8ZpJ1uCAppIbxLm9YbJGCgnOlwai7bXDnJQcmFG3sejeu1MLCTbUOuxJPBpCosnAg71RRll
XIU4aIekbicG8l+8pOK8fVBVco0q8EhMmNHh5G3S29D/GH4eVITmaTWBwymiC8px5LPH3XlXCiDJ
XbZte9HHPpLvkpUiBQhVYNzvT6A9Zo0j9n96I83tjYXfjy0v1MIPnXCzkOHMvL1T+CAzzzYD3T36
DXxrJqZmEw4/5EfixU6dYvPDlHJYSHt9cYoN0KKA4kNsE+Y9a0S9YkOJJCOqWZpP+vrM3qbzu0wc
7PeQIxKGVwZeDCrymhv4TboCRy+jU3kURJeHVv3MxILvqH9Px384Z7RGqkdHa1SUZo9aFEKRsj4P
BvwqkIS1+/llJ/R0/NzSDYa6CcfPzk37WKRUZ3RDXPwmWh11X6WxLV+K9v9FjUIpf7mUxlX8ovj3
PUIYNaHYZmtUovhCqBn2ygq4g7fv8gzLy3HpiNuna8VVm1Vi2IfJ7Gg3UtHnxk5LJ5mAEZTsQ4SY
da420uwSzNnT6I6PFd88xcKIsLZGmUiPH/MNRTsGS2bKlhMRCMQ7DAMGwPlTFScxU4W3TTuYL2aw
q0KEowL8etJyZzvbrMVhw6RJngI5aCjvdD5UIZYUJQmNj5urxVnIV9uKt284U/eT95VNX9egPk/e
+viBNsTDBMVTPreuWpodOUSbRReUu0tqOwoVOU4JiQoGYCdxXNqjxjiDYQ6CfQlXh6A5jOcrNdoT
fuhKyWMwsBfybkAWvnyRj7ADPAipDPg3mse7jCHx3db7/OkfNX0A9JUihvj0QhxfZ7JRUQnJZE+a
cLQ/5+IjSfjxv0xe7x4dgGzC9eJ1xXGNOmCocoAyhYojsxkkaP7mGF4CTCgG5pr20IsZVNGXm3cn
K43KF6ezoxzy69d8g1cb+T+StSOnp8MG25RD+XP4pE1nt/W2/6I4CSXkqKuZUIwXeOQb/xOXJJux
yLNL/brfS7vuRsCyu0zJ6EfeKW6q3au7rmeVSJFrz/7v2u/wNY37uHIKwR7ovWYqnz0LEvguiSbw
3Wo50qHXp1STlHw/IvpqSpotdOTSVyI7puLs98WFiwJmKirB0E89pVF39cw9s+D2BL+NnIzQp39L
K/uRRbv7FgVRqYab9hvfTnrnM9p+4Pe+37+GrcRCr3YEDG8aA7Zdj5TE8w7dsm9v1JVzKSGcjcv2
XOzOSvrvEul/mnQRyHI0OWNps1b/8B9jGy5EdJwbMX+EFjmd77iSvlskzcSQRqlTKrElWwMuDlF2
cN9tC3/XtpyNcdAoQRLKhFJQjq6MnNdD+X1BdNDX0vnzqiHwkX2r//UA7MNUf+evfU8ND5voK1qm
kCHUiXZ2K6RlG6cYin4XZW5zU3DVU9MnNFwSAFXCItzSU32ScCIjAY+sLsrmNWZNFnEU5RQ/A+yW
yh6plDy0GxGN3O5mbLiIQ/4GHWh+wY8uKK9grLLhXa/2p7ZLHy5iaDDbVpLxLcdfn13Nrw6G7DzY
0sy8bbyol2Ak36e9ENNEDDmvVkHeRl1XZjfsK9LKEgvAs4wzGQVKeNTnEUSuD313y5evBXN166et
bMSeC76PLSTHIinx3aebrqnMXt9wLqzHPHwdpmgn7gi6fZIa68OpqqDiW1VmtqndwhRuABtOFY46
PGXoOcNcrHjimTpaEMy6XwA6qCgYRJ7pbgShfw7sVflPeN8gzFyDP/ehTzDAZyIMpgSBjqO+ko0h
XqqV6mlAfgnAsK2mNRm71MM9nKGLo2LeVLvjekdLo42+rL6X6MjEgCRrSJBLeBs2PX4j+OUpgpR4
tuq+T5icS9k6Ana0CzSqIPko7A+ajLhDTMZ9OTAmGGTLKV9SSO0nEARQjDLt/DSMtDIG5O/qep8V
b/YBYnsQG4HbIFYU1aEH2QEybMrMGrK3DSu24tAKqso04FMAM8kH7LIItlAxvve1wzDLGOeLATh8
B4Wz9fZBHQmD2MKyH/ag9IMONLikWa1f3MChLsr8k5rasTsffCpdleReL+KrAGHo4/bVmqtZBYlK
h1Szu1hmYfpa2fw304JHnRkaZgjZ5wXqJGCTDi4C8qmJelqgkkaYqksog60vAjQ2QLTotMds6XsP
xVxMAYBBbPPgv9gXVl4mtPQVzO0SycFOQmzS4S+Y/pyOjBfXTUhyI6Wkn7JrS2LzPry8xsbMRcrE
BhOcqyNVTcOE4B4OLWNL12sEKxi02X5YenmPw//nL6S4VOk5GvJ7ECvRHlFnO+C5vOsikO+csb1n
UPkmeLHzDBxfSj2e30Yg+C91/UqatEvj5DHluH3zAC2eV5rCHyVPLilC0iZVBBfIOTOCBODnaI+K
txSObAQ6D+/v2y3SF5M81dS6y6nKU72lQXvNSZbSqaU8CQgbLoIm1bIXLWh05UWP9tiDPbixHfB3
2d5KiV+01Sy1tQsDYM/E1yXnahKohvCTl54iWS2auUDFLrGfN7/OSpQSJPjo00n9Fav0m4rgTUaH
9CWjoR/SaeqggdsHmYe1OSBUNdMoGT1woe5k93AJ1t5gK6gOTIGaiKLp8hzdslaQGEmkBCcAsoDX
WYf2JjzwxdrnI4hnGaihJeiKmlCNwhSDhqCoRFEzUr0uq8khYd9F8JwiwXv03zeb2Gyfxd/Jg5Lh
1aRJFcBSjyss5yUkxVUA7K4h3Ecx6cDlOaPH5cMwv/c7JkhjrBtlTgCSEmWL+QeAXXCabsZKLAfF
jY4bCzHz3R93+oXMesU3JOSNko4VLDjzjpud04EEZtWUxNs/q6pIufIWY7MrlQk3mNKAWR7hu6MO
ptxhKdcrP7WnASAN87ySSOwVbwzdCRXip2UOF8/tPp0Qfiaic6Je2f+Kh4mO8AKoRi/L0ORQOPmn
kxYh3gc4fsdRkRovJ+DJay3vMIFp3IveK61w1aRg+P0TDglKjehQUVOB72sPyEsEdez67k962AvL
BxLpj+oew50Uj3R9uUutlbWlfWNoavT4b/aDxcRKkohec15GP/DyIx+6irGJV7U37/e/KKILhnwZ
tUutpFzsTWYMkqJWoncOtzlxZ2tHk/BiWq5vBIab2tA/Cwf0VDAbUNh3keA9AIrBIUTRO0rSIbSm
ao5bdp4bqHoABL2yPOEA3ULWCP4StR9I/UWWRgujCY/QQK0oFTclyQdVOSpevkG+DvaD3V8yoxIE
/JA6laL1uxNRI1vHheeKPdMkmqZejyq/3Pwy1YomV3ELc4iTecPeAo/BCX70C3yUgLrvhawBGdDN
PlrvIAHsoU48A/gV6DYsqR+ZnFfyqLetfIDdMorde2rcky9lKsC0Db2tJvnLjq6o97nHWFB73rWe
2v75GK0xwcMCts+e7A5ZWtNK35uKgkApfucEdD0jKJwwNuNXgpq+GA+98TvA+/eU16642ZWsEGJg
SVaeG5VF16yDbWGa+IECQMi1J3hxM6EcU57TaxJ+G7/ocpuuI6pczZaVjsS1fs05/GGeupAc5cUE
2h1YblJcjmjPxtqBlBJXaM/snASltnHUp/SrJJSKzhwCsKLjKoCkaYw97dQABXXb4y1AzXNwm/Eg
BKDmPR0EbQPqmk0lNrJpZgolo5R2EXFAnzTw+BfESDOEjnt9ZAjijt6hN8T7b0OMyT1rlhs2wpXT
PY6w/7pLJHF7O4ryG/eV6b/xwEvqwE6YNrY21mn7JjQrIvoC6RL62R47+Ak83HXmfY7JjjxElmIx
Tq0pOu0Zb0j+DBggX9JWK3GrApVH2jrgNSJfggr94Ujc/7MFUF4HD5g7n+wMAK4QOp4axCQJ+30m
BoWo7nevTpzwYAeUmCmqTShHc7n1kc6L6ZoahNRU6fH6M8wGOksLp4w4Jvb3BWdgqW1KZKNyNUSy
BO38b4HbrE0QeFa86c3AimcC7TuOnr3OFmOncLR4xYva7Kzg6JJYS/SS/RfdCCt7hiAv7YPB0vG8
6my6vdVbyGPfk0pbgezHJR6hThfn37KudiZw3HylI7h1+JGf36NqmCbyjegdCiazDdTzgggJLJGm
m75vAOsWFXrviy1I5V7Znx8ROe6M8CcGPHKDIYp/t5eFdRB7FQARsEVXKwqJkdCcrgmewkVpzQnP
UzMxtArscTPnarlPxyDYaGwCPmqpNBl3ClyFFZ3bTzK8/dGru57p/uZPS4mpeRy2wcGqiFA6+sXn
RzmGuVkIgjgW2hCSUkC/1flbeOV0s41vLXdnykTnq40VgyQoYbaKvqaIg/4nz7TXJVZqnxAR08EX
kpobavK0me2fe2aXTZr7C6N/N38z6mSipbdyALKHLiih7pMhzg8tPv3e9XrN1hH064Uh8WoBsC1j
cnSH5lVo5WnBSjbWW5DqA4xgRQQ9eM5LQtdWOlsoTyYUoJw4TfBM7/dE8yd+2t4u92X2SZXlzOo6
P7rhortvFDA+Qo3vo8JI3DM1hIAn9Jrc1mODA9oXQ0OaCi0eu6vSi9gMg5m7hu6G+WXvE2zAtLlW
jZIaWAtKlcSM7ZCtzlDd1q45kxYiIqih5rUZ2FYtqVNkEdeSleGka0MXDfvJLlUUitQqjQnya6zX
IYAux6731ALIhKumjBixzhD5gZakXPVY+tE1XR4U3UK502yXKJDZz0GvvVTn6RVJCvtHp7KeBfYZ
XbrP4MJS5uvV+XTjvTm5ihhNyzSZp/l5TVp5Lmrng02q5D3/k2/CCYE++JDp6DROQ6cd8QIeFPdp
TmFkgfmspxD+mw36LZmmmN6DFm8QxxEO0bKOlLOxRPLUYpdGgw5RtZF4V1vo6/PI2gittph07g6V
LPcgoHmxYOBpBr5Rz1L1TgIthOWmYGeOJfgdqxjN3MkeAbr9P22abmgYYddN0XG1h81v9REFVF5u
H17fTCM1EtveuRf8dTBk9hqTFGJMgbD/1vYmScRo3v7z0DwAgY8+3kIStLYmkayCAmblgmg5Zqca
5reLK67ptXakVKaxeAcK+VaVpjZ4o2G1l1B5lNLeupeyUIG1BVmRyB4J2/HHkhWcAVuAKCrLYJbW
cPC3NknChpFcuMDkvamDq4A2c6EW+d5WSV7kzoVnJjZG58TvYSXHwp/BaO6PjsU6FcFhanOLmpCk
SaANmgElDp9yubma9d2r+Vs4I4miNu6u58znT0shaWRniN8nPahzC/IR4A92cNQtmsJJAdpIIbac
2kE7xeOfPnap2qx0hXNXc5VaJaFOvbdzm1qpuHnLD5Xex3GkeDkOmU3IJ/VzIyuY6KQF3T8c6F4C
qTSu7NajAx/79lHwEzSUhv4pI1lQ+hLMO4akBOWPBQaxEL/FztL2Ra6u8fA/vTAnXN25585axQbF
BLhtngHnnWuJTDfBF+vm3Ppxy3pFdT/QRv1jyNKVxPIGw42zluT3OqQu/ZRoTSrCtO9W8M4fSLJD
EL4GlMyarNmbnltIq8SIPb912KDantbKc0yx65AZBEH3Nz7I+Sf4iFOr7Z5R09MWhRvb8ZOyjG1r
HOUE2UTEZjY6zlOGmbd+ONxbEEfqk95rOgdwA5oKRb9EOndvGzEl1Fjan/WoTl5jWIgqsma0zGpg
/0Yq584BUy69NofNhL83jWSxJk3ORyKNgr6bkkRsBSHQT72xJFjOebV3X3M/PNqSX0WnPHPB8si4
5eU7v60kQP14J727j1rj/fryxw8kjZBq6C55Q49QW4F2ni4DcFN9RLdie60aAbmClc1iCEEp/Jb+
UUkGYNNpeuNcn4S8JGDMlCj/o8KQ6Q/uR9bojPOMYmASXqSLgaakD1Q49CNuB96fyJ/hsFuVG98I
ungYndyIuHdo43yi5qa30XQuQ6zbyi8SzqITLoTF7Shf4qoLt1cOmpSrfRddp1yqwbARUddM8g40
h1dv4SgiwbrzsiHK7iKmLhX7zMgzham4dbcO+UnOILFG+9sc0fDn/Z5ZgURFmsRReshOUh82urnG
6foDAaGGbzJvkhjBl7VSfJfSDUCLCNwV1yf2gtWWmvIt+X80dCi/xjPyuBaqZB6g/0bZn91sk77L
KfszpLKrlbXgQEMHYgyJQk7hijwoO+yJSPwDajxDcecRe/rfmFb3mAoYwatjBTzLTxIk2F2A2v9F
5s1nVXPNVAk5/dCYl6xpxNZw3S1QQG9V+y/keQAASOSqUNXRZeq9C0jY//NlpWmTLCWwNKcC+i/S
dS4WlvZe6f0uLs1+MFXY1xEyh+6L8ga6Erw6NGi8WiHUvAkbyuey+XxzJBIPgROMn2xmLVx1IYjX
c2BkKdHMNapVZc7159sc9Ju4npGSVcAWZg608oWLG3rqW700j5vea2adT5MdxEaw0rSr2y8kE7pn
q0AhhOrdDjpCnoGSXsc2JasLBf/EnpjMSmvVFc5+kKT8FMjUH6BzKdZ4r1Wu6NdJFO1u4CAYvsak
2kQx8MtEv4QHjozTl4lpHRTSElMNkYP3t9I1a6X6gQbcH/WrhYL3B+7x98CoxnsQmlIwF4IgGYHw
jxC0eyLpPl2BizbRE6WKwvfbmp5aovsOB3ZDnhSQTHHpMsMNDUEDULrIEanDk4brctpimvVcSbNu
sOXky2ial7a9J1UGi2RJVV2UgNy9POPAio/QO5E9XXkpe7z47x5su/PMEGhpZ27FsVgWqOr/bzr/
aLDQ1Dhj91j+S8gGScEtKgkJBOLEdXy9e9qMoOTM7Nlr72+3geAZ2N/3/obrQ/T+FkCTpdtdFvup
j15eU0B4gyOptYJIR+MLU/sOrfJfOcqlk58fdvdpCrH7yp+EZSil78UGlkNJYVMLLy423HYyIMhv
wm6GXU8R6sBIyb1ahrQ2xTzvr1MBGiMY+LaGVjkjgoHAXXUxLxjLlYSWoGUATagssSbIR2ovPGGG
eXShriJ+ZRvwF4XWt7eSyq7kLb6oVVFXDzspJp9YDwHJJ72fgitzhUfCUxfWb886Wpxg+lKxYkiz
xVUGWZXL1OS5LNjjBJhQMBqtTMYlPh/pFfQL51rPywxyJHd2F7kfxYoQjOYiRHz2RUfRJJ2uZyx5
UwqZ0xDlztM6uXaUoJ1zhD/rVOsUzooWgoOzHIZGpLZe/zB8tDQZy2yqADJFQ0N3ap19FIk4Fjg9
QYzz81+bWQsra0jtzv+chdcydE3yn17BipmPTA4JS6+EcYnqlZ1XNDhgSMmysqJ1NcB1bLMJJCb8
tiM/eBLfk1/6YH2lay371tTO+kukfYWZnpvzvol5hbPNl45lfW87rwyYnm1Xg9O5UatBDUmcuOs0
uG/a2PC3Gub9nGH3DXqiVukObJ22z7un3tr/tAFTxGF+ufLBIuQdUK6oa5/zd8KYMKpt8VC4FA5t
mZqzcpdG0H9q3a5RP5nUOBdm3eE/ERLMbS4uQd8s/sUkE2dDloIJtolv1TfG2bvPjtuenpz34a1n
Gq4GRZPtS5HPzxOChRUT/SQN6uKQgfpDnJN2K/vUkMlrXpycjntY6OPDMkth9LmoPGfuCkJcytSd
5emQvRoe5aujmLwPGr2LRR4rMy/a7J0MraDkAJZP0MU2ZqgQYdsiuiyihFsdUvjxodzL1a6wF+7q
wtvhnrwcLrCW3aOHT5dGfVrxrSlZO7T9rjpCfyCY4O8jWzF7Rg7gD1jgaU3JgirzaETRyjf1UPzh
fHk4teQqUuEXY3LXDFR7Y5XcdlmnDmljmauIGWlH0wSyadhQYYLwOAcIEWGhcmbP/OUc27CJOL2Y
2nayU0dmi/HJ8RVDczic0n6OtYZRWxNNZGfSEvOYDo7eFcti+zPe7lLs6Cf+H8TZUhl4z2kVqII9
Wze+km+fb858FRerCclh9w1IwJuVgpMdZFfDsFnWcI/J3tE3Yo6kTGQoh90IyGuXS/KToyg1eWrT
4FYfTG4675kDx2ygDnL0DjU/89TsZOuJHUCiuc5tgkOGjm5Hu2dZhzO/gbKsZ0CWrPj/d2UTUbCe
ZMX/KFQpyrAIyyG6FZPfhHZc2Dasu6A75FGVhyB1z8R7u/dblQ4sCEahwKAo4GB7V2dXsnvAcf0m
0Oq9SUDKYsJsfdktwDjh+Ta2UQugzm7EQ8qvkh1H9liWlIE/rhYB3OKMbGndLVG5ZoCaj/fmA/8Y
b+1f+S6jN5O7a5vcW3PkP9vgCr+2ZaJYv5KZj93/7pb15uhmaShWvR3z9bM5Zm4ONZ8eFcOe6Xuq
Ig+1CdwEeeWr8We+ueYEu0pmaGOgL8kRd2/LVRW/nYXVYgP2FaTkYtMBqw/xmhcVBQH+F9Z0V27y
GKSSEe3ByWSCnxtU8X8Ehe6phyZbcfibOnEf7jL1YJnxyjzki1OuExwoZ/nAVquMiCsbJC5jvIhH
ecE9CzFrh7L8mt7hY2RcaDeBjxZNvBCcqgyQsHRGbv2uzy+3k/Nzu5C+Lph0WUDQV5d77Jqv8JXo
lpFVTIiEM2jRbnkfnHj590xjSWgdgfBkWUpTffbtQohMyTZD/lTD7pymsSc8YpQTP6GqJOJK6qdl
JRirQMfuoXnuamNF5ZlXUIyUWUYd4LiUzkBZRUKbHEADIwySFA48x2DGQEQ2XTFvfdmERBq290sp
W2QWGTnDFlCsL7zPC7506egtJ7spPOiib88GVtKdyTDzNkmHAGBI0tJxs1x6lnY6VnZJ1iO/nGsc
u/SR31ANkDIobm4OKAF1+ZBn6UXnNHRq4RduHuGTcjK6c1tyvMFn1LIuz+etj7PmEmLk9cK+w855
SZ1VXWfxShnfjtp8TQeX/FzjTuqkmk+h2mjYE7Q/QGhsAJlp7bLOUVbe49ZEzTDslc/veKaMqmiZ
MMtufFD4NFQd5Gp0C2msgIlOMTtrawA/CjmzlKDXlUrAXsyPWc516zwnU+7rmRYrGqXlQRe9aCkf
DZQP/UIp1oRY/iN1xTnK+bfCtdEYo/nXg7m1rB82UqgyKPiUMUwiP4pIM8X4u3c56Ig75J32pRuE
UOP/t4iiVoDOhtTsRRnBBZivEn2fNugSskoWU5zXeKe/bIL9pUgpWyiSMSI51Z/MhO2gi14zjPfY
Kk/07FbLfsWIEpmv9jaXY4LQ8I5kTJ6Efp8ThQxSA2Ulj6QlSm+udIzOm70iE8QZo2IBZNZM9IdN
tXnQALfcMtk3h34OPRqxsXnziUOzf/9aIi4Nm3m1emzxVcKclNZrKFobAoUV1Trd7LvhzatGHv1o
vjSBIeXl7PoAKFDPnPHqzaoAi2melhDonJaAxKJM1y+fcolFSgLkFaxDYQVRQ499lf+FU7ev0kwv
7nHe384bKffS9U4W3EY/20a8rn52/YtPZIJIwlfn7SilPZ0XuDjWTrFnxg/CVelxvVwUQsgTXiZg
21kSBG/uq6eCqwwdVvjpZYO5t+zWs0617tCoDM37o+7A/FWFSx9SLkmrzY5VE/1PmiV/SMJhPhyC
EdNptLzWsy8KYWmd2jNRoDGvmShAI21fqF/kLOvpAHFApa7umGPBQqTWPA5odWbQ68y9NVLf/ssq
2WDK0CH2hqbTkV/XMDCHk3ohunxs6/3LKaRW2eFuvKgrIyAL5RlEhndZQiGmTsCaA/hkekrrOdQD
n/8PfGt8zudeqbgMLmzBYniCp9kRRmenTNJLZ1vfyzYfiDZ0bHFELQAhxLR+2JpFk1Osl9uCwlQQ
S0pgYMbXAGDctqR6RzpdwzCpV1OTabD8B/okuEZNVmjv1IYrUFJHijUmYfiDflinvKrlfJgqf3Ab
yjVuRZUMN7/CdK6f7vjxVK52z8nVN74/Vk5X70aP8BvuKpwwFXsEfhxnpsvEpdbDsmu7DurMmLFh
oOrDGLg8wK5qonI2w8YBs+/So7pIpOZ8gsfGL+FVSFigbUoFErCSW9t9sFb4u2hxs9e7DSdctZXm
HH1kMIP1pVS9oyv7GUnYfgkO5tRtf8hBTYeRTBOr5wJbq348ZSdq2sdRp3K69fmGgBR+MAUragB0
PwI83/Zvd468GQgg3toiKq7DRpb/TAValhNl/2V6NkdslTFQa7IqeT16srSD0Tq8NceDFVcbWJfC
O3PNy5EVM015vmFbonsd+O2TYnDEtTStHtjI8KR19Bi2gWRHvg5+W+he5OsjAHuK+FKn3xWL94AA
e17l6hnc0MvRxNl/4kUEjo1rcYAUak+/y7jAWjMkj96fp/VBIO1zuC7diJv6IWgjDMDxWe8qwM9h
DiCBI9Ij9wba8rXT6IxYNaU5XmR0TDLFq0IeHExjiQwd754uJrrHk5zFRMFrmoqnKaq2kV0hXU52
mK3qN+PYt1HWvQQ3RYtp2Y/hJINr3oYsVkJZ/skoytxInZ7S4cwt2IjzakSTMEr4dVselkfs/Ox+
7LTk1SIlHuRm0kc99AlhsJCZHQHgEAmzK0eeNtKdYxwBmvMiSqPSTS14UpWL4XSTKmQin3yoZs8Y
K4cxGhXrFA7TX+Ug6C1OGt6JSE+SatvjwqkhYC0N/1SBGqT3GkoR78JOoVamIh/HOze6e9b8WQ+E
nplbTDYytFgX7xjn1VxZEAisU4gjqBLtaREuu2kIcruyV3vEzje1IAl4lJglrd3Svcai2OUZxqDT
8dKorxyaglu2rqM5azdNFspgCSYqnQn7k/jgqLY62/3/XcfO/bnUqbWkaWYe7MfncsIDjlVJZVGb
hCaOlrEw5z+XFhDHG71bUQ2WlB448la7lRJWNMJ+Hk/SDdf0YbXMJu9gsJEtXim/VsUsh1HuqAjM
mM+8mp3RebE1iwx9V9jWtcZPUDxFj47bzMc+aGwmM6OmozAxWcoGlM2f9VNPEYlVsTRvDa7PHCDh
tE8M5o7pzc9yYCozjLCmcSrnz8x9UWYd8vkVAj5lE46kVUspznO6Jm6Ev+Q9re4FgRCoudcwZJWl
FquVM1GahBciBDhjLfGjmezt3z+YNbVhM1ZeZ3Fs8rG4MHe1iOk1yya5oP9bNCuanEQiVq72DNMf
aGnEl0Ul2m6NBDzn0s6u7ISZOx7PrGMktxFJGF7HJxHeW5wVrh4tP1C2b3Y0XNjDWqEMBcSDNkIq
r5DjFOaxf3hvfHe+7jmn5IGcvdJbVI8TElAlaJ633j61Jgj7JGRZRbzau1IpeUqRXvrKJXZAeErZ
6PHIhpE/i1e1NDp81USWOdLF7ur3TYUNKuMbu4AX7FNSVCMI1fl3k0M1HPihBsLZ+Aun+/mayEzk
LFM1Al8i62aAGIyhS6PyL3ICI3YEeOtUwPqwO43FghrkqyJlRB4+DnLCSR7zqaMh8HvejG/z/ZPU
cvn6ngLcvrUVS61MeFcZ3WoReODDbXuLlmQn6QxkJNK8yiJSF9jkxwJFVpz6fe+lpo0UXF4d8fia
cXaWveu6oTNRfDyO2qcsEXUOg5u3M9WPciMhbEs5rBfm86p2qAPxXS2Jlmhy0ViG6iUBtr6Lszc+
hxXLrbYOYy4OHQfjIjaGneDOHYNBq5c10OrUnAn+17f/Vtfld5spq74LMVFSR8WOOdfuCUemSxv2
6NOVPhkQO+RWwn3P/wIHcD+25TD3jsrm7J6BDPzDD95Z8dAM82yXO7SdVJ1CbCqWJ7YNyBZx5fvW
2OhrivYyf7OUquhPM5dJdDGWqkVQ3gJoS7HupkG0bO2C1QT2JMlmCSRLIuV4lnKq9z+Q3uLb/Os5
KbV16a0tLoSpiiH6PTnRq7hvlO8s6FII1+xSKnxzMjwxDVifo3qQJxysgSX8/CXOf8p1b2vdsCNT
CQuaqo+bO0cBYx1eE56yXafEHgptusm1W0R2oP4ViouZa1egOQOk/jaMTdhB3QWoviZ7KGb4/NnH
m1zpelOZwV45W1DKHZBpiyVIVga7wB8Mw0zWff3nUobQJykCNIFq6978DWGT1ykCI1YqKFbnmJ4+
IiQ0zYC6R7IS4Wdy3IxHm5ep7ugU5arU9UFR4mar7mwtRFbJthWSOWfeRRrPsxFvHMCLH4eZbt8R
m91ClibPO/TwQHvAFqPOBJKZwPFNWT/IebnOSTs7BNz/92nZhVv4Fs32Uh/XeGY6wz2cjXfelsi2
cQVKrv+lUn2AhVLMv6R7qw5aazW8akai4YUiaiv8z+BagUGCozgya+/mHYy18MxMklbPOUFYZ14u
aVN3Idt+d3EryYQwYHUU3j9WVqVaTPAXvf2VzQHs5gIIWnvh8Gisb9lr1VFpCFJbyx0gWk+GyD8C
HEQ/1LhMiYZR/z1DGdZsbum5kQKjletAB1nrrPZRNE1ScrEfOTmCiZnPSQFhazVHBTkGD6DNjlH2
79pDdkddPUrLKDUTgyS8hH0MSniq53Z7ZXZ1fvNxY/z8Z5T6IMJLqQvIjRG8tHpb6utCvJmXSk4M
cNfBEofQeABFYGO+crV/NYks/nGAP0Ym5iLoQc3E6V8sSkIhKbYJ7C/MIJojFnIBInK5k4rky3OK
440PM/8MKn5v5oyUnOPNuyxdtSYPHeBMkossKIvA6oCl4wXrsTcruEiaMHr57lDVlj5YtN99viF0
oM2lBjrB4bv+3BFup1GW7IYiZh47HIpA1tEV7crs6Or+6jPodQHunGEI0t9UGGnOJLLxE7H84FHn
hy7npAmibApl0Ud2HBxyNajmcL+DEmXBw94+t3z9pFNXfFgt+6q+VnhQD5yi8aeqTJNDvNks6gDD
ZUhGxr0NL2Cn7BNHhxkYpUSu+aIoSWgNN/f5tkbNz/fO/oVcA74N4JU35Cd0F21VmnldxtE0cRG9
4L6/wIOws3m0Rs59Xb99/fiaXjKI+Hzni/buwFAIGbNae72jayPlqdYdVa/L/pjGDhyv7buobdZM
63UujkDs831cU7I4ttdjusBV07/ZljWpDXy3ofHoVtt11NP1W4ctetVl1ttlBxUrOvjJCCiBboir
Vo6eYW2CqpLYsglGEuwnOBAcjXG37HLHuwLyI60/McdszClm549eW4rUf3Oa9usVLi5qKPLlwxIW
yn5ILKmh/zw/Mpkt5ILJ+4TYc81EU3WmCehV2HEotYgoP6Ubqh24c3/ts2qb/RwlpTQ40ShfemCn
dMv+uB6dscQuWWERQH02BGh5c4hg0SufA1GTjjJsXetHJeqeDwrbG+wFfhFHjkbXoonXAu0WDc+h
GtnpL2oUhLol2QH/zhpDp6U4uNEbUtZx7/eEkWP70XCnV0AC5O0jWT7iDAcFQonU6ZB4KQyt521K
NwctnUUxi7LScge51SvKpRSGmdyQBpBC55R9Lgh7OvcbiWfYPdW6W6xEnQsfaQ7X+fW0migZxSft
QMyvtL2dmwag8mQdpktW3kivedDSKYOWLdmNruFFZVqbV6AgF+JEJfNkvPyZoHS3XuDnGicClfbm
tJ/fM3Ec7EqhapA9z6j7Q7gMFsEjWqS1uj0Nyz/m53pn/s/rZfKTc/zCtarMk0Ms5vSFBulw6Yqg
1mXFIR0/ltArOC6iEfq7wGI8BJiK6mnIJ5j7d6OCNTlTt6GUeMnZGqSNoiq9j/rJMfEkdalzrWYF
ESJ2BNn2USR49XauyyzEhXx8H5+CB6T62b/S6tVrTxvOTs3l3HyUolQZzJ3KuVWLsiqs9zI+Xj7L
EIDQ/x66wIcuCY9CO5WMiUYJKZlpzd+6P2iS5gLmubMo8FwWvi52aO8+pCGiaLzbsqSfTk5k+LoU
EFwFvd/VukqfS87w0Mh+ClurKH8aaa9t0eMTmKLmJExNUtJZy14WkXNXfBGEwx5k31Qk7FC3NFd2
NQ2aQDy0fHffDvrixmQCzFeGtmkZSdRDbDpANo6jlo4WaP0ozuNNJhBsGKdrdlVMZRcsfl4VoSpc
iDAQn1wKSvP5LeAbAqIFwMb9h1cyhvwPzpcGRnLKhAz/7NYSY1lUdGFDLEt+1dyLZ1miEYWBjwuD
UIg/GJELMS9IOLDTIskjLdApcVUy+t4aOLOQ0Fvm5zNlj41Sfx/gvnfMsFBi4bS+2NJGTCr/lEm3
FQPnsTG9Dx9fSyv2v0T4FVAORDTxt5ojQg0jKrSVI3/gFIRsm2BZjnA9rG1d0euPA4vZT9z7Hq1a
yXDIviANapzQKIwPtNVRMUVaB+BcnJxFXvvDpes9iwxxeWrdW0C2LOxGA8QQP8luSHXnZDZfPvEF
P2C5TZi3UKXCuXU2fgYnIzvLMPvo5zf3yjMOs37m2wbnPcRKTM9ebaRNV6087QqLXBTYZs9M20Im
f3Xn83cLiRPHSRymyBKnO9aAYh8Ws0jVsO4n1Bq8tnclltMeELLWZNY1oGCM1sKnZYsTQpyJ31yZ
7Z5WVQtOouYtcEk8M6WEpWyuW0xUINT+Zl5oDuqK1QpuASVp5HLfBonLRj2xs1+tbNO2McuDseCH
oYtME0WbacdrZn+rKqR91hyJbaxOLpT9Y5eJdP80cCzZ/bkd6A+mOpl2ozEbR/0ioCeh/MZEnATW
OeKGTj33HdumNE5ZUzaIBkw1VNs9HQl+3CMAH5XvhTTwKjFdXajZXtGAeu4p/zDEQk8Tu3y9FtfV
8jukdtXpScVYyyxmTKOeKltMftQrd0t3c2DkU4K6M3xj4b3738JFzDw9PLL8lisKUWGM6pa0AiF+
WpI9CMcAtRtda1987Cwsub+Zb+hA0jcJvCayQihcGH2sF7Q0/Yw1mi30kn5LcofEa45ycKHVndoq
Q1RK2BVKfMzNGG/gWn+cJKaQFQ3A+5cfpvndPqfjeM/jreYBABEwZ8WnPUxaHDePRkVSP67JDxkF
75b23/4TrVPpOduSHuUifeyC0hQARkj7zmz8Fqsq7omCoe5g/s5sa+4Ca0t0b5Yza+KWf5sBVpJX
1O42W2FRoztDWDY3N68n+5ugwlCMUQdbiK+v9RBxyPbQQlNKVEs+sMveie84hAlEiR4+y0ULRne7
1FL9ip6AMJzOnKnnjCy5xpPQM/HbbdvZgC2qi0yeOdXuonmz/lbeJjAk0NN3DRyeSw8rnfvvs2EP
FrpdKYxI8MugS61b4NQdxxBrBkYvPX2AkTYHgxrm8km51Tp0wWcZDoAnFFaOUBe6DElIfPrdg7uF
BLVqPgzqRkTiG5w9AIM34gHSfJhd26Mrs/4ElKIwm6JxD7dctjH0SVZxpcLY5yzktvtzdS+HcLJS
t0Jju5zyiykwcF/RC+rz7XPN/UVQamOoyhUyl+/HiPH/BZJgHUww4dxltGKKJI8BdrZBjHuliv8t
bL/Hr2L/CjkeWRCNZj1xyeh8HRnpohaDknXhq3sjDUtkOYFzUBvMrNCKg7UtsGpkNmtgkRz9u+QJ
NNps2FkdQuUA7mWgt/6Ypqgw9QQ5/tURBCqCZcLHtkp6nLAxRE10aSQQ54lrYN12YZ7N/PK6Dz5v
eP/hQdOOy41JzCIMuelPlhtVuD/SO5itypn80GSHLn1SXPQPaa8itzGAdywWf6N/bN7rP86pd92O
UxgBmEZffdXwqUcWqQ+ZRGT36qjtxtgR1OBwkVbl+eoZBEnGtJ7mwaupk4KZknokNMLIhl9DapFn
E+n8nCucJO+JIbZmsUEDLH2LbrO4NPXWees3tgiUQP7LTCoBXjpWKmidkBAXG+rdogqr3YIJZHNw
6s2ziFhTEsn7DIw5t7813ufiRa+GjMuVNcyaEwlra13iVBRFfP7+AZ+P0CQrDVg91MSKM3EyJ/7F
PNi78saBIvYKWLJbs3Vqhuh5+Kp1cz1u4J3we/wMgrHDq8BbCkdYQKy2Y/7acqTVDv+XJba4xqaV
SVBrC+w62UgLyJeIJeimMGTx+yHL9hL1QO2bmZf+9C5A8MzSdiCYI4GKvhoO1RJyBdUIg2dUBAQe
AzeQUVTROeYhevrM+5HUsPh8Cp/fgSUKEM8gn/uDhq57I0L1ewRDJQrEq73T6myj65Ohf3lNdE8C
dxRvqOu8OW2qaTe0kb69YRc15ywp3bPZFi1KfsG119oxvgO/tfZVN2n0lrwIpv5iS9s1kAMIx5nQ
3FOpe3/qr0LSrJublHRieWU1aDtI+GRv9AltvqrSsaMp75KEWLVeQI7Xq65eYIo3LJCvAM/67byu
ec09L4cSvneF/cBRgsShlOFQuiXhkf0RYN4cy7Gpd2rRRPAJKH6/5q1taHdRYTglBr4cQs0UIfqS
c4LgEhQEnF50OE8AYjuLRwfWoRZxCMLkYT6ut+Ylvo9QlTGkK/N4y8xDJ59uF6F+mLg5AxjfTVAV
WIkHlfH3tOWOsmyum8PSo5mU45ZBVvBO4hrZYG981wodp3+7M4PjZ0/X3vbQi89BO6uoRHlRLSGg
CX6Ou3gxMGvl02Q8DeTDDIT+uOuo+yFJhtCYvtwI9asGLev7XOQR1VYnOTekO+fdSRCUR1YCY3jW
Yedt60WSZVxKWOQEb+7IkLdHiNSIVczQYsTE1JW0+nix+tSO+aLd4BGGqigFy9HxipwO+Q6aHT0V
YsAAXwZiYhVT0UQ4YrbgrCXFP/TEdumyqQeganZrHTA5IJaC72Gcysg2Uv++q+KJ+Y/krF2UtAXw
GNRNky07shvCMo5YLCyG47yFjPFBVhjZBT5HaEvDODPbcqh7dSAiHt/vcPnaLFNriXy8200Ht590
fNvjzek25KzpQG0g+Adz5laI53MsTyBGguTcFtrpDn77SNGjf8vZ8zf6zZZcCjJrmfIAogLuTz0j
w4UUHt3O/wSsyBa1g9D4jTDhJIa0td5/rzXIK42uPhY1rMzrJnTI+UFRFz8GS0qPkLSG/41BpFVJ
vWpds8SyehJ2sftO2XXtfREVzscuGIwuvAZ530+LkietyTEXKoPQHXJrIy+AaxnyXsSMxjXs+x2H
+EPQqOeLxbgNChTt/49B8uiVWB/D463p2lQ/8okV2wtVZTG2u5O947N5g04noHp5i6NlFzGHlM0A
poRyTBFsjS1G0WVwdeF3zceB2R2LHEwEg3AUvBbC3xqc9PnoA2adv86WIa3exog4h2grA9F3ZZO+
SOWEDxYdMo6nVfDjJYbVsGde40U+3nna+cQBjO1Z3JoAtNeX6fGNzT3UqPdpixNbSjsTqzJGsY9A
FYL9u6CLw/tzNKVulNtF0ZbOsY2wXMCKjTQIbSIHKLdt8QBtakodoLBRRhFQ8cauSdpTFqcil/1Q
RhqqKHKYwNimbWvP2F4yUHYLBUAB4LLQUZC65ADMPDz+H+HqC+WJ78K0b3e6uBqVMsphZVLCy7/O
m0cF1acLTg3UgL6ErWS2JlIQi6J563khZMqn3LkiaWwGy7k9u5kTSANBOKEMU8HWLR0hUdmvPoZb
ZfTOcmhpgFEu5gtADxCnPQaPFentiGXHDV0BBHReonoFPDY7TKVE0GHfR8ptGg8YOAfPeZMfD2We
+zERenvhSr69CuJlkFeiJt0WFMveTJyKc1+gnbef+DCHeFiCFiycy9NLlsjQoO28vgKU55DO9oRP
n2g5idsS7ZZzWKgbFqNF79TA/jmLwQ/0pE5h8lXFtbokb60oTUclhcc+H4HZcO1B22M3f2MZNlbu
ovpqowNl7ihlOMWwMUUmtotLvOonLhCzrRG0ZGNcBFDCVfgnMpPG3Xxej83LOS/kWGegcepyyZVi
KqkCkjJN01uCmj5a9CMS6kYOLqGOh1BrGux4FhksYPfsh5HkJI7TocANkFLOHKZxO7BEjE2XLcyV
OVPtbApvVZ2pyhKVrhASqyY21XZL4ZuqqfOIwDl1CSJuXMX8CkrfQQniNdBraypp29/+PThzkAPt
2BsR/I/qcmiMBbl3VypJts9ahMTdLhaABYis8e6+E3xxqVcuK58J9VTQuidKUUbNpwIjmWo5AGoh
TX4FFccuGDkLAikm8QgQdXN5F51dvWLh1n00iaqfbpOpkDjFPM264xxB14EFI9wE3ZcOahNfHj4y
GSmtx993+6kr3aDhJ174R3VsSlPtHdvH16VnVgohJud0WpgeWPjlBrsTJ9pkXSJmDRsoqaML6xQJ
fKqbmmo9lC8q0uGc4wUYuQMWFxJxC2l2vZcZG5AFf2/MbXEZyIjh5y0P29dhRPK8nxpldBG5vMKc
JhD5yYB/T+Xql0jBIDYhVrKFfOEe1lqYj+eIs6q4/DZoYqbPhLhqYPKGxKIxbv1/lmP4IB79lbOa
z35t664UFQTVtRuOGSZxrf3l7xkeKOf7+H9FRKFpNDCEIN5bHd34SSN4SRdIU7zp45sINcHKlqkl
TdM+2m1zZQZpzoOg8aobgHkYuG7St9vLyYVWQNUOVSuQ6e7ypYj1rQEaIsk1RItbd5Y2QZJ1lh2Y
X6+RuD+eHI7kOgqCgOw73vXkyhN5lBM0HX/yQQxobZPIKDgl/gIHom23+aacEgUmoyGvYinTtEDk
5559Go1rFz65xkma1kTaNqgnW2P+lveYUuJCTf/ymLXLmOzAv3wXPRoKM5+TRTB7XW0CmJfd4Dm5
pUh8WECIsW6JPV4nvQM2X5HxoYfc6CUJ9rUkCQ80hg5WgfqihJGwKIkb9K8jWFeNfwhDYgIpqUhS
QW0mpMk01tdfnJfPO1hUIxVwWmhBRhKgqhhkOnzdoozRukz6MLBArFdLgV9iqFRVbtGK55d9Jsdf
dQHEyRffFmgrReRdO2hucYjzqV+rAT02ibtne744LWtQx9Rq2+CgRj6MHxGPLJUuousXX5Ktht+r
7NQhWTfxcI9MhdZbuq7sg9B5SR50y90o785YRif++Qa5IS2CiOoS9eWzWLjs+C3ai03DNvXYXgzG
jMc2rQi7b9sN+btrqOHYih7zBPeHOzbsRzL/vMr9P4gFm/Hb3xvICns8Lq7Y2qmxsN7Kf3xJj0AI
7zlMDg+/7AZj+YmGVznmf6U/3gifmD4TwdqgQHEHoYjLcbvwhxqjkyVZbA8dFJz72Hf0Gy06+n9L
thIovDBEV3mj9vv4xHsfyefGcKzeqexij8vPDtS6zwHQBg3LlFcG41H8RegaRk09SeRSC/XYjGgT
aw7dU5vVwGzGORopiVweTZ8Wu9MwUlem2jdr91wfLQ0txx4d19cnw83QK0nsGN4vHdgm9b9UdTUy
xFL1EJrCwxS7vDl4lWPektocQhAXwlIXZwvo3WERQrw5ybO6az2rTDsnB+MOWrRHBTDEyj1sqKJG
dhFbB8QcX0/2ipIhMJX9EIZC7Bf/wgJCTipzHl6dKCUJHt7rsphS8KQYL2fdN4XWphCvYw1M/7J0
zQnKtsWMUxT6y4gA8/XnUIByw2Ji5alxEr+qr3vqgOndvFez2zAL8sAcdgOLLTzOrPoUehLAkYiZ
7CUOPdrgLOjz8Mnw4c/5+4j7CGpVM5RmMW4uEku7FpCX6CeO+gM0GT+Xd5fAjTKTbik3z7JPj6aZ
srPBaxul6ZpAkVAeWpdBdOO39AVYdHpSYFlpaI7maqECf7gFtBIvOf+/EUz8vv7ZHUQaPwZo4l7I
Ex9mw4fslMIwTGHpzyeyf06nj2VxgTXS3bgUsp4BXYWlhI0sKIzSfKde+mZoC3QySHBkDyNJ0kwn
JEw02bL1wOJomtstSHpAndaoXaI/eKRlcAP/ZSxSEDRhy1P8Eg0zzF6yylOzxVlrykVpUEKFQamB
N38qJPolgTEhGkkz82fZ2UpMIdZ7jBhR7oLrqVNc5O4VKpc7O+XnD5HMJNxv+xDqK4kB4dvxcDcC
WWsXW9kQ/9dnGnIe5DUfrHBlgVLg/RW4jl70lK0IVgYjXhGfHKNSNiAtqNpaj4TGZuM0HtDx0hAV
9GFwRkflAAmHi5MQ7oDOM1R/H0X4LbzpJXNhgUEyuFdgvzhzxTuMkjagB9/NLTElJH3epRwOuPl5
VcItpPgXtvCmZP3jg68rzfPnt6zXIqT4ZkbgQr0tbkqByZVssGU/NTDMZX4Rtm9VG1JPrBw0qpJG
KxIIbrZr2rBFMP42xOLXt1NYPU54kCJo5GNWvx669ss1stDkbqVxrnLL/9kDjyQDJqF/4va/s3zl
QmsYErp2WWoGxfbQWWP4vypG4Xvyo4KXi93rEV0/5MzWzE7wt6E+Fd93B6fyyTm3//VZ3pUo9V6n
J/rAgKcp2OXvfjtNaOPWuxBxRpk4cds6D6ezPudSMLjevQ10m0W9ja5wD9mHrXdheDEz4oA4cr+e
i/t2iJqFFSIAYRG+Mti2YO36PFETDJRSsADkW2wn9k7WQs/aFoQLFjnx7l0e4qNPiu8+1382SSxB
gUH0rqlmhp/+VachInb21buYujfGwDVPEmSYunU0gTNQDWMXXaeasaJhRRYaTecABbZGEco3/I2S
fiKSRdrM/5No3LQRNq9+c3/k2SPzSQQ/29dsND8q6AXU2tQrjKJGhn7R1g67Oy6VmpSnIN5VunM+
Hr58xYk+P644Vbz3wmYb7RI9J+ojB+XTKr7r+AiAt+QHSu8AwCEAirIRKLMISYBNM94kzBoVEWf+
B821oJu03dAtBWjGMA+bMXQACndN5OCd59QnfX//YKW2MgommGQJ9KAFnONxD5oaXqCC3HT2BY5X
fQViqqfunrn6sxuYSj5/Rm9V4fJ0VuppJJXwEqAjwnxTh8qSVh9HwDfBlxoSkSyov517fSQNx4sL
i30ktpjd4WLoqG34OYoPTiVc62wQR9pOUcIk6bv8R8GxMzq2LO4QGkkmKrp4P7ta67XxNUer7mug
alVXPICyftmLDCsYrOE++8jZYk/+gS0utAIDaTAAx+OHGRCIQB8MQ89Y8NCLEz0UhmkVHIZX+RUD
kYytTKPgjsxpIDIip3ucljPSC1EtyKHUyKwQUHSbykSz9ujv11R6v3aiLNPJqJ4kJm7UE2LFCEE4
zqv9juf8yYphEsGwLewNPhQVCrVoi2ZQ5tG6hGkfl9tZthJNdRS3zcjYwXu6mn2REZs6/zC5PeYL
Quekt85NUfjjAVMOKG7YUkOcnT++xI+f0VOresnfFG+FiCJGtpkpqnlt47ABcIfiGCceU7cYNQu4
zM5iqqFXvRsq6uMPpn9X8BX/qreRd7eVuf1yrPQ8m70uKNBNkuUEqk29BXNnwCi/dryn4yqPKWCU
kmiMPiXu/X6FtBbC9AiAW+BHbY+SUzpHNZ4gSZexiyrXvY7umCzHokB/sDVoUucS860NbG8zQm3i
EM3ZL3mm7v6MdArNbNP8OqxONq5EfHJ6tvyHsmWH3jAl6FchYnZok0UxD1bdcXhaImbNOSL6DjvH
hLG7bUHDiuJYJJ7mSBcXiddSvfsyR6hSF8rRIO8NXgomrogYyY+k1SKclqvdv6HyAfAs8v6P/KCI
rDSzH6Kzc/DyYLr7exMBo/IdcKPqM5KWv6tPPmh8GSUifXBSndl15y5CqVvOSJdxVaYYF/KOo5CE
k5ZoC0hlVfq5uq5skFfdjiJikU5hgvvkpsgo9X0P4nSu9lHtM8uFAYAuz1K2o3FohfrbkwaV6jRV
/oibXUPlsgeg+ylI4C2lIn6lcLcG0tnlGTjTBOeL0IE/nkQMcMvSVOeu44HmG5ku6juOniPg0Vvz
XYMqwT1/ndoJSYbKN5kELOMSKCyXMTkb0BvxEDzeiMOokIEmpUjQbsL+1Y7J6ZlCjjBTC2h9nTBT
7WjJglPycwb27x7A8j+krqD7WG28+5zcHBoAYt8y2Hg/7wBBZJ3jGFDZcK1ypHTp4q2K9onRo7ss
8kd4d3MszuDrMGSTg+JfnHUg3wB27gWt4js/fqFKx92k/LALbK2FCZzEyMeIPjeni0bsRKFsd8gR
+0SpORvmn6vOFaz8CqROEOMmsDXlfU8H9vfX4LgwA06LHGMzmANz9+OABiM1klg2dc/dWe5vbFTH
CdNQDPyjZEtkPqgPlpC2Ae4TrF0rWQvuIxLttO2hRWjypg/OmasM/F1yKIIIGK5WfkjJBI/LyK32
AKOKDYoQUp+Fn9gpIxaaLmPyfZLs6rqEafvkQNcTwELitANJnhvMcn8jo8+VBFIaWIuzmLItio8F
8vZ9Kd4tx9qIbyMtC4JqI/9LVOb0aNFCntjqM8x5eznf4tcnNaPyXsWu1AU/VWcN0DuWTsNoHilU
h8pdw046hlz8jdXn+M3u9NDc8u8PGBRYU79L/njIiDT7zOhjKwTmFtaqJy/C5HneQ4AyD6+HXAxu
Pf0X0A2B1drQ3zxyhxTBUoDNT4zTakKBx5UTJOw5pBkyEUUgfmIlC2z4QAIeYc6cDnKu4U2Uzb1L
tloJqwcRM8X/528FUHPTsggau0cwLR3lWrqCvXjq6uFCKtIBIjMzBfsLCm4l/CKrTyZzR2LzziLf
yEU+isHsCLiCEG4Ol5fwpttQwftfd11bBgE0Bz2FoRkS2yGSQkKJGR+BWg5ggF8e1S0B+u+rCuMa
f6tutG2e6rM4qkuibFMBQ4DaRv48keWNynkojVgM5MVp27MCUK6Q/RdClSnIOXkpM7ZfJwJHe4xE
mpJciFQstr6p4lYO3j26RZdSN0yVVU9+i2cjGjSuIh/cP144nb5oLNSAkAsaneDWzlUa/YUjQ1Wl
tYmNIPGo04VaL+hjybluFFIw4KnQifdclVG/O3v+zt3jl0JUmFIPY4CQz3c26GsW+qS11LICgwe2
SnRlIY+jeR6JW/Z2pIVf2mWrGe+m7FSvfAXUJJDbi44QzLUtlNaHXThEgePFdrgERnyiVC4YtRMC
GgIrVVSu2g98/vjjS4VySfzIxYkwes5GXbqzbB2wTWENgrELnJnmgk68V/RbPCkYLmLBEmnIWKKr
em0S1XJWBg1Rvrr9C2GdyM4QyKfvpqn30TAjT2oDZobwYXBH1JH+0iPadVjw1V/2B1BXgGZgMMY4
NTCDs2eL2HOyZC+3PGgPiNbrA04Mr5EjRQnU+YFcLdLaprBK+fC/dQSqHfhIzitUqpQc7KlJYkBf
uW27hNf2wYjO3VmtqQTasz77HG5AHlmUrSoYJFurKkEeBq0lgNNefJWSON1h+PJ7jQiaLX4PJWQ4
TYJlCoCT++aVI8tg85m19My34QKkWeA0N8h4RR60To5QkXAETTfQN0MYZEHCDCek4kaOCh99Tcyt
u75zPyDGJjrzBGyBvUIk2vr7r8MfXniKjbxo6k4N6To/7XsX9Fw3oPQnAPai6JMkA4xXEAegEm8D
0+i2JKd566y9SBTViTwwfNxcnsEILnN407PKhAN/O+lgb2PAcMcQDFxyz06E7Jq3ge4rFT+WfTU4
2KRkW0C3tZ/tdSpPuatOr0NSZYIZ1hxj1OQBO0DUQZMAAwfZ4Jk/8yocFHRz9xYddXS2ccPcoG9Y
jhmn1aDR017cQylAUCHM+IK3E8Dbo+tuWLTmwVltS8XzulY5HNuHmvCQBRNxlnOqjqGScnLcP9dg
1oFBbzlyrN2S8ZikeyGBdEQJnBiSpQ//yNp1mJIja4qXZp+WnDqouzKSM06e8hABIEZm3pTvx5zq
MvHUobGzwWcjoJsE6VGGdeKebD9NBZ09jMRbPSbz6MF1XpzI2NNyRgGrbflN8OIDJLQ2+EhOeVvZ
oklVG67hFjPwURwypxRMWjnQg5xs3zGNaaW64Ce6NRqNlo34d38xz2hGB+tDHD7wix0W0p6EFuma
vFt1vJEB2Alc1gc4V7NSuGhER1aQNPceVywh6JW/apeZUhi9ZVE/tRhc5bpeuJxSfIzEmJmE/7T2
JoRHOryPQVIDmfbEKEp+FKQwJEzJ15MD2nCfJlJGOcEkZ349d9bz/dZE2JL1L1ZNPPRMNNCHOkMa
rUDT/3FtdgG54oyBQ6Bm/LPyCYn56J9rABt7A1qjly+Yz0WMO4WUViEW9wGa0sMPrk/wNtI2hZV9
AMlKU+O+XW58RoR0+C+QX2fAdyxtSPxuYZ+iOQs/A5v8HOcNBXHq6t0lSAczDk3A2uHeMxmWu2l5
VFoc+dPviM0lM41jFW/dOQ9fFmGLItuxIrWtNpTFlaN2gyHb5SsBE5XqT6tRjgqF4Zfnvh47g3ne
rJKb94As+R6g100BlYY0Qn7n2kk6fZSGhsfMJ9KwAzYi0z5yVfdig2eyDcdP+v54lPXB//rr8phT
+Dcs+Ajfar3KFhUxThh5y96Knc0eqqdMrp2N0pUznkNKCm40xntWWgHZ9bjU6Q0xDNOxxv546bmd
uZOsdshbQDVjwVXdrSKqBqjgksbSC+cIm6ZBShugN0Ydg025n1nQh+fs5qwSdv4/2bxa7yAJfCR3
QROilTU+DQnXC6CMtUkkRDeMv8fJrghckDVlFdvJEpQclCqAeVw61l2DbiOKi5Fe3MdPgIF5wVw0
5NLdigcuX+9CDRiCIPnFRH9VWKaR5ALyDoU88LQDm2CXSuMPEC9EHsWyXQDb55bEzFJXoQ8qFjuh
1Es9+ZAE5O0EbgEm1+YzpmApSfC1sfZnEzZuVXg3ws8erTikSBTyrndoERhGA2pegaqEuCDOh8UR
jbH7rU/1ufUUrhnHyHkZYKpo3toADPU+7Y9Mo74nPvAvfxKm6u2cKbGjLtezuchLYWQTQslQlM2N
QCFk5bp0P/QgAKPtaD9vKy30RiLZe6FZDLbh76FHi8DPVkXsCmLBItSgNG6SPqdxZpCDsCPR821M
JyzlW00maTFRopPhlJT+SGGgP9tBrUPMHUfCKzb/hsPRcpembOWDLZu7hULSRqzn8U/K1Xi4i5iF
CDyK32Ql4De6phD+dVzkgUK3MKM5ixZ7WP+o9ryPkctbd/zkemr8t6Oo77E05E5yyrpNiSUX7cZz
DNZRup4nuSYfvPd7yAm+tr24ju2trw5XnRXrKhasD0Y1TgIooGuoTmvTl0rAB4X8j+KEw85+XsfR
/N0idgZ2SKe95rkDzen3j50Bf+1D+7ybievUSIoPo1lRiq7Si1lTKfX5fUfhb1Y1iqMU1y/Eggg3
HzWtu8tEVTiU2OXqI/Yar1jynFOt+j5VKkySBgUYy46meUVIljc90oLvsEZIXv80rAczFHT0NSjZ
JmVKAjFwVgRF4oAtQOeVIpo0y8YgO++TMWYlEovxHKlvsGwgzxqQ6TYbQeGuXE92Al+LcDz6sySV
ePqCAf42WWJPKHcJnOPrZJTm20bjJ29HQEx3QUhwFnK7P6e9NzoEZBpfw/jOev0HFJa66ktQTiEY
K/3uDw8rFdF3qhrvcVmHZJ5Bv/r9572sdoumzz81fjqCxMKBWGGp2+Wja/z84NZ4571jt+gud0/H
LMvJcouxgCIQPS005lMRx6n/mUL9WOg1GuvLczZc9IjBkT0MQJ/SI59vNV81iwais1vSlBjGLN3N
XlSsqIWs77FbYa+y60SgLP2y6wqpg2sAEn8hpHHflsk5pqw22DvCzbRpmHflUVZNf83rjy7aESsj
2dCfMuQG467NJpFF/ivd/3NM2c9He8vtP7MA/GM7wIWTkwUovikNE3/avWA6jPZTEZ9iT+LZjT2f
lwhcLxsWfk4TeqozEJJOANwQjENbvJzSBtMGrdsj5+GAra2X+2zrwGb2E+8atIYgoYGtmEMoTBsP
hntmupL+BagV5Uh8Nfwz//ncwNUWzrc+up7Vfjl43kk1htFI5XnQOv/2KL2NVh0p5mpCrWPFE8Gl
5BGXCWWmSJg7PsgvXtPKhJL2m48cUKkuGvmdhXSbKjnrKFzNUf1KR6sX7f8SJcor8Zv4Vj5CJASK
pKxsFeSpZ3D/LQq5Py9WGdeZm8TUrdn7hRFUIAg39qRow7986X+q/2mkjb3RM4KmO+ey48UPSjuo
vHd7jzhpl16k8YavVfK0WZ7AuiD5vpicFazxkQHMVBHw9nql2orqeJx7/15PmhVUCaWv0uqtuyZU
rH+XxlaCeP01XCvVZ3bc8bhYoj7Al5yibbskGVeWpRMH8LoffWXbqn240zC/HrvISuqOIqRkWxPG
gcZJRQcaat6aXTX3NExWfLNzFwTYwkbrAKN9c4H38CIFtQdiAysPVq2AELS877/Fb2b5u1KIXWnG
esFFWsUn+a/5C8BBh9jLuVUNvzmiqyy/Y0g+NyhuPrCX/BvMKwjGEX0b6KDHeYqlqEAvOXwpY45L
TvgcJvEjDC5X5MJqlIdndaeajMS3blHbutRd0DKV0lbBcOeGtst/wfBuXaTuwg+o6JaWMhHq9cr/
gojyyz2AoFBiqij3mFx0b8IidgNqAQTmZQeReKIw/hFjZnDzlBxDTkKLDO/8eSHj+9sdic90vmbz
fH9Wl8m1DPEUMzqcKux+N/eh8yi2/2nwniMXlX3ftFaUKs8884oVQncCdPo3hq51ffhE8QDkRjBz
VsHjvyMBQII8vDAxE0OxdciprBNP+ijfofqpKYccK8u2KYJOp22WTzADITIsflUbc1ocTd7Sl9UD
Pzr7ZbZ0kH1nZgZvJKmT74Rf1igw3Bmc/PfybNJPS/jaCVbALwOHjWvvu/Q3GHWECqphJUV75Eid
muCD1uBNMttxMb6bvOKYth7WiUVjZQes1A2s+9MxEwfv52kBr1dy2oxsLEPEvpOiJyzeQ2uBkiMb
VE/othSB0/2vTMTuoFJAGxC3Js1kaLdwjJna2XVTNsUO+jaVStMNDc8gTpiXONls5T2jFdLwXeJ6
gCakIztiyomHOA7xSmk5x4BK9iijEJjWiXrowMIWpRh9pro91/Pr8gBJDwccN8nc/ICkL8r/DoKL
kGmiGjyDoIkU67CwweFhtF0jLyp9bVwC5tBasT9U2xOIqzEwbO2DkF3JCWikYOdT8LtdVDOJYvjb
gUwInM7RFsrp/659yaCl+8gTzlmco7a9N4ArQs8PRD13nmuthfQ7MAn2EhclbdAuk9UOU9mAE/rQ
Va9kKgirVp6fIhBL/3lP7MeoMmx22DhnirkZAMRXTtA8InuwQW1Vt/IOdBcKapi8pMocYJtU3L3P
EjFIZdHwyG923Vs5xuQ5B2VCsr0IjhJLTig9rrrivFZsTv8E86nThvBlnB3n4k1PL9JE7lQqlVtG
y2ueotcxWwMb/qo++xtknUYd53kxsdjrmiHMEcKfrL77eXHbhKqGOsN0CZA1fRI5IktLNfmdriKD
vHsN3YtLtkfa2sXaWEHiofxIDyjZ3YBje0B6HqWtevBGpSrb+AI9l2hjWLeCfjmh28jw4p9GSQ7d
xX5rTk98yltYH4l+qkVWlSyNkGnBK3a4/nOSMXrskxoGJ/0yYm2WgUIdw2Gb11Pm1GikgLwp326X
3m9CEnmqAIc6L1dKr00hGsdWHNXYo9tqwDvJTukRuV2TShP35x1KQ+mXyTYqv+8E6hZHAFSC6roO
QKlYcM0uWkNN2JjcJOIlNF/Y/6+gNrBI5NhuJzRtBSrywSgyY/22iLpGBVE7AuFiaHdyIFnn7OJG
eTbEOM45NAydWVDAAsgf9uRtTJ06+V54kMYlgn3YW+sq9rkLASoiclOWlsSj6QLFDrrGdnA34Ssj
OryHQaHSYVBmCvHr3NUwLz3qTkH5kklgw5yRiMNRTHDGjhKs3L6HdARLsEzhxwbBJpzIoryB+S7S
gRAhLD5ajsYqUCgHrXKj9XAB6bxi9RLP76ivwS08NKUy6VyK79Ne85HDR/r/B1HsOa9DtuXzj2B3
aokA5OnfPVGUCyeHUD+qJbLlFpqPFo5hdIfddugV15gqaLIGX9VsiPoQA2CjItXyYSEKU4l8PM9e
b8JUEwTpkPjb1M8rRskrwwn8r/fddjqKKN7niVqblfjy9zAe1abiKHG1Ua6C2d+oQqy175zr2CoA
uy8xu9onH5pUgqleGL5utJRDKSwlwXGH0fG3DvzZN8ez3gRxDfsQF6pjdUQZSiN8HfiHgx4kXd+c
+MktJ6NoYrFXhPXIndKWeaOjoXiRX+80ax7U3p7iJyagEk4WGnWkAozGdi/6+mh5FpEx0PxQIlyW
fz9iCbpQ94yf6OwWx9N1nsdawFi7IwMcQid8d9S6QPRiZ4euKyA6jn+0RRUjwb7exA0d1fFS9e/v
jVV7gLn6jrxU/saBoMBymk0Z5RHfKJSYOsrmBHHE8H9b2p2fcBG3C9QHWwCvkeFzPdrNcD0/qX/n
QRagsmqTEfUMX0cmU6OL2EGsg07v8uMGXSjVZPsE9RlgcvtRRpQO0zehYHhXyxIJ6ZI4rkisa0Zg
iPtiNcQ14g9aGXZGpfEITf7dJYOmbLhWeWp4uTtuci7XFM1E+RbbVJPwoDTW5L8Su0C2ZSZAjZ+K
5PuIaWGuK0UL8Z+sVU7A6HSCpvRlfy15lj8fG+9cFLg1zY/kRIE8LFFn99e8oabdp34hqsQtLHof
2zjLzt0MXFX6QZsaNCBYnFpYua+XKnwITRlKUw/CC7s2d4FnQHMLgmGXsViAwzKFSDajds9RlSqt
gtuWbUzDH2N9j2uNGtxRBxSY/86+Ckq33HHMoMC0SKZSsMI2kLsGrknXItLaKjQ+xofswmoItEAp
1dXxyO8KDM4+p//l/r8O0c7p7tINEJUnMYePKdm/njU2MbrnllJzzb357X1Z8jp7Ckoh03DrNMbH
lKKph5TjOX+vxNsEwi9NyQOTBSAwJoM2WJiCHoGHBvt57xZI/vrW3ETBmOf2QjJXu15czFWfaGTL
Iubb3m7Hv+VwoEW34TlBaIAjSUW+Wd824Dme8TP4DUTOGqExkIHbMVl8CTMZZNbT7zpfhBNlMe+X
+rk8foLECt1bGDcCzeCfoho4dTnk5kOBzb23WopLxJAz43pGFAkSP4xtQAmZKsDQCQOkwJj4sODE
QYkKVAzxfOlvlaByTNDp0e8O3U9vKuZIj5MzIGSc7LVgyn6UMzclqOOEqQxUwX11EFuCLmy03C6l
8Ir2caMUVvva7kdjqsNltaO25VBZjTFm9XmoVK3YQ1fKjUdNLFGUoPiHL1EitLdjQGOk28xsEcBg
2Cqm2nMfyLK9gji+NRlmnpAd84/6Blhl1J0hJ1xf7pKyfDqrpFLQ7l0CUVJF/drBc/ZWTPC7Hkt1
wlzhgh+xllWtU/XACNf9L2zv03il1JvHSRXJWOKJnkjgFeazsj1S/Vje16ijGFgoebS8S8lFaPw+
Gy1BCyWgqoHQETZJSM/6bqw4q56VecP3ehIydfMFL+3pBiEVjLzO/JzJ6PrShd9ev7JRDCnW+e1t
SePWDN3dxcYW79NtiAwVd+wNUeIjhkyTIw+BNtmqg+mk5w9B28w5mSE+7er+oXlhZDqtQ5y+kTuQ
cfZeP9n3peiE/EZcoAxEnLYIUaBPMfh3GafASNOY2Q4AocheqfUNu6G2aBfhefuz8h1YFWOUQQ5X
nR0z85mAIMZ9a3JzykbR72dL2m7oCwNzEoK8AvWoxW7ybHPi4s6ktB9veoMyTnmWyn6A8xSMIQTF
Ld0HdaDmshOskFC1jKLyHaDDpIik64zLsI5lJwkoa2t8jPRUQhFx2/vSyQW+IFDvsA3pu5+yymXG
iRgqQgqTy4iypntXP5oTlLSs0/5S++Ir5HZV1EOjCMaq6LFm7ptHiMiv5RdUm2SlHYeGBEqYf4tx
h8wD0cuY7c2nfkARe16Emmo3lju2YhlANn9kNZVjU9HzJde3d7AM4AaYYaUWhOD4/ls/s5Elobi6
yRP1EuACvSconqW6ARcBF93DC0pnYPnu1a96YO1ygEJ56aJR+cJscnsQvEbjeTJTgdVBe9c6OuAK
NZd1q7q4z7rQ4j8POA5vt28ZCZtnJxXYKn+b0XEkUV7CyPdsFej2SZOyFBBN4V90edI5PVwgQBgS
vXhEawURcrZjveq7gwTh2ImSmohR8NbNkkBlp3K1vsEWCzZBUeH2X0Si4g+fN+NQy9jvIPtMHOBO
JGXaV6Jk7nCaN/ctBnvl9mEOYxFsW/DZJikWGsDCjzFPWCezWpZWO6y89bX84kaxZxRVJGqNb6RV
NZgJdwwcH/atEaG44VHIBttBXk7RkAzVwrLCOJn2K2yii29ETEUU6+6j/CBT0QxfS6q7PPmb2NbP
qqwOv64TZibBG0UYyfTfdlR7yE1CLwlnQ8Hwr8hZuWBhS/L3eWkW7ZcxLynqxZvuUVD54jH5uO/a
uwE4rGja4Y8H3fXcnmEcnV0nTA/e5MXDNksuTsY5bwqOyi6PpspiDrftKudfH6ib08ttfDdNt4qS
vxE1oAiV+H2Hq1g1EBegW1xrxkO7EOTdR9b+eGspVlIty+6CbvPYuJsffeGu71q3Qb1aXMRMxkr7
JMHmaaOIJYAeJ8KBKWRwUDO0n7xJI8Ra21ttllN7yvZzhQKar/uWVli0youtwDzmBVszfcVoyAGc
u2oNAmOZlun5c+5iyG+XPyKIaSDNlp1r45oiBnutjwimuXOYoXcCpKOw8n7Zz5tkNuTLp2psklRu
QUozSR36GriZJa/LpkVZ7yFd5P7PyJAWLO9dWylnnr6V7yg38XgKjBA8KDIIEy0x54gRZhQkTSxG
Y8W4rvSUR4I/+fpgjUkUo04hpqgkijDsazo/A9bLeOs80Bbk1zzqmS16WaXlbT1sE6U+kqZx/9pl
4sGBwqRPx1yzwqhTZ5KETnZBV41MLXyPH/1o8b4yMyuBLKxRLa2RBvvEtvTS18ONacOGB7w31lzp
jj+p2O+fmT4tpR1gLtZG1eN5ndS3BCHWgCqGDnLQMrp5MrT78/QliFvqE99htU2OMs19ojyNRora
Xi5qEMcBzhvB4MxxGPnc8tpRimFJ9S3FKoPcg4tglgw++zfT/UOAd82QffWawu0qvY9KX2+MgvPp
TwvIT+g45hN0Hgp4Et1l6Is0+CofK3XZWxBoDb8j7Dtg25SIFPcXfVYgrzD/YkXJQfp7EB0ptAX6
0PYVn5/E3V1wCmrU1gvEDuc0pfmHJg1rafgV/WXFE+nddaSpfX+liA2gMVC9hQxZ8U9TLNLOcLlL
+tQIGK1Dye4Wg3nMqaXfzMOj/dl0djzaEo+V9q6M4MmfiRJ0D/4uymf8wXvs7I8MC7TaFuQl4eSv
QEdyapSWGxsGzlIranDfNBcAfwp2c8LHZJW0FATVcM2FZYhaouSHlZnqEP7ZvkKZhzeEjg4cvz2q
skZXoQ1psREo1vPjNlK9bLVncrOgqFtUg055yCJcxvBKpMw1QGGeeVroyvPJulP/7/E3fSoAuaNr
4adVzdgtWJpQf7kSxi7jGsndMFfBmVVMcJ/YnMBYjJkAz6ogpsGFjWVovRCFYEn0zi3xqw5eE37s
4auVhgPP6FcZLeTsiPSG0GNDaQsXwt0/jhDRVr3AIZdkZuMY3b1BBh+rlwCR7HhTzOX+ifPfURGX
36BFyCi8sSqRQp3Iom988n5grVCFugXfwiRZkyA0ty6jx52ZNGEG5hHbvbbIDMxv//4P/QLjgHHb
RJjONMA0eILSzViFdjL9sOoVYazzBSTVNnImOk7UTFdEOsYknXENDl9opWxOX6GDlyeSVWKKKei2
23fkq99mtIEltlUClpUpw3fvKI8WQ8npmsdaX5hXG2DHfTFRFBw9GMD/WDx9X5nHfecX7VQgI5hT
ai9OhTIoPgHFosxFJ0O0GFtSIwFnQIkfAjroyNOi3csL48XmMKhCf6bewNcQbn4dzkCrwbfx7NGX
uPeExrko3dFNypK5ulYnGN64PCJyjngV2/m4xZARGg9deAB8Og/KIA8mnlLdGLlL3sBV9XzV7CAh
+khqCqeyWkzWycn/E9fpM2KineuwOhoCSpJlQRxIj7oJn7diDgDG0RpdGvD+mq7FD4F/qdfCTXO8
HdQKbT8GQLGfGR8g15UnhcLegW4mIs1DL3oDIJWt4AJxpyRrYfl9QcOxZx+ing3YdoRaZG6sI0e5
nxIt1vVQv7w/gDeGcnXrk8h9/2Z/qF9WcNENS6OXhdQZ2kTYt7KOByogGyMYJNzwOEJqjjq1xPHU
4L70e3m2tZsF+qTh53LNxeJIZcWbclkiFhyothfmhPNDHKNtgpWl0ehJmxQgZK5dtqM+8NHsosoJ
a7ZJjejMTSTeY3xKXh69dAm2waVojB3jpBjtdURNwfJfmZiso7qljro/nW6aEEG1qSHnTTztPev7
CNxFoGF3mCELg7yvDQZXZLFzLUrDpSo7vPEfzlcIFv9qDTrt3Asj5DHfPQwcSpwR7nmobRuUoSob
/g1xlCt9uXHoxzpU9GnW4dASA12zi3VbciGFwmrUs2PMqz+par0zdfVyvLFlwQ5gGqdu9paYxQ0z
oDgU/BHh23F++nBMO7DtBRomdQsbwZv5WKGE2wumoDLbS3xueAYzoN7L+2oyf3laxIpHHOgBTt/J
/HcDwazVIr3SpVpz8b5NYLp4/os0jqRBF88I0imKyCHZM7EQ6x4k3pU8mygcTAvbTZp/4tcUix8e
0TjtT1EffwbBEByBgC+5kkquvNRp8wjbEQ+80SPae5c6zYeLkimOCg/JYbZiymoRVqb25KjZbr44
4R4ciUVulCVd9UTIgfKU1Vf+Ri8kk7Z/6XE0xVbSJg66uoM0/lc8dg/pEE3se86i0gp3vB546wbf
jPeBaUmdpE2om6N9ezItlfAFyepW/fAwTyV0jqHqyhP5+sX50KcM8qZoNzGWRnp0EolqWF/LuIgQ
g0LcxE6+WeuBJKoJSFvXOG5OQz7moeiFlnMBcu08/2TsvzKHhaWFEvg2oA//ehAjhFK0dScrGKea
Xz6SsvFZ48u0A6qD/rEgCN7Rrqb9HY60viC6fO9DZIrI4TO4jeaYFPTQorTR93mMLBo0BUFke83b
A6z/1NKplZJyT9dBJlC6L38sL7RhKJsOWogYHv9tsJhq1UO6EP2QZdut25Y6A0b9EK1bBFTlIQcG
8/kg421fxsmOQL/CHu4llvMKRm9VQvRd+z18UYJhxmZ61rROJqfDt2QJkj/+TdGQHph/WjE0JUuM
hL9h/QFrd5TGn38Okl6DSwkt+e2VNg76wJeEuPTenMs0EXiRJ8Y8lMgPhW2qMCDKFxweKB4i6IQX
hOaVMIDLlWYmlUxDXx5BQV1E4pmmWIJ2158l/dv4cS1bKPauMntKK4JNDRu9SnM4xA8Ynp4FjoaX
VuoKkiJxpRA72vh6X2f+lPIJgO7mLXCD/PFCk3UvnfjTjONwD2tG0kPP+vygZvaAZDo1K9Wc2Lj4
fptkWv3p+4ssNz4QKk7ueGX7QfQ1HpURG5+sZw+sMIKiYLNIJF7qsWDkmL9yWbuBpksYggD6EQNZ
q7qSx5wsqi1YrlUcFPya8cuWzcA23fdjKaKKv6LI7wgU9S6TrkSjpWQBk1P4AhI76uM0asYK/TbW
DfZsid4EIuaR3BFIlXYtv81ZcHe7L5cc4MZCmp6NiaAfatbMT6SSCR9X2ZYMWXw+PfB2H+UjymqQ
HLe53ZjNjOit5iPU+3QseO3UxK3UArH3cPOD5i8cixNqGdO+o/QzlVkT2DKor4Fm8gAVAQtZ5qv6
ONLlGjuM5q5AlUw/arJ88RfLd8h2xRyP9SnnwKxQfAieOiKFj5T63KEwxhe42+0e6rgj+BoNCxww
HTzLwnqx1A4kFmEwzq1EfWth45pmiy6hDGsz/j1qNXY2zljCqXY8TItMpWaqQkNT141IMCJV/pyq
K6dJNXgs2nX8I6B7ecYAVKbZSMi8R08tXV09JUpUsNUc3oie8Zi/QHXxI2uDDYjqzf9bLwbAVJ9Y
oL4D9teuvlp5rsHMBXiFI2x76nQuPSAsPAVusCCgqT9ooTNcDvgRWyPnGCvAey56QC5N4CIm5naV
xrvjCsSMJCmZ12V8DPRZy2NT9Ay0LH+QrTVmPABwkl6smyLBxbNJ9IRlZ5FgfhPNfTbra26uCxP7
vegtMF99xhyhHmf4WGFc0ghsLWXrdAtnI/kZ9+UKo/J550zRiVYOHO184w3YIQJra4I9w1XOdZYE
0glfWn6LcNdOowl1a9ge9HM0BGUO/QylcaUAxv6eQdxh/mx+ZqbcjptLt1zLW0kZTkTGjViQ5aa3
W6it1dZ+YHH5Q0A/SOaNeu7baIcQRuLFzBvAeMxFZ/KolleQkie3OTPK6moyfWFbvOPsIlUdQVl2
H65SDFrX5K1hRltK7XBIcbltjjNK0uWs2qOsR0HafAqdOL+5x+5Bnh3aK1xltHSVaRZ0ijReG6FI
KS37QSolIoDl42JnhadkAFbLBB2UKjUJTW3fY7X+6ZgzIMdr4av895FcvA78se/L+WsjnD10BCHS
l9VBNGdZyWDi4e/r2Q9ZfivPcXI+lu4TYui7jPvSDxT5bNK4gGooxHRghgy+QaHwWEQmmDh8e4nA
CmgyUsQ/+1stem99xSv9JbH0mKI3D+45s+o0szOVj1J2A3hyT2ajfiV7oB0B//3NCFuUJyE6UwAu
rMAKKUsaLEPyUoWLk+dOAkQlj6GUwAaPrSj1CsmpVJsPYlMS4Fw6OSTIwLiPZ7CGxE6/bVzcEzmK
qeKMmJLebC5cKLHcm3P62Tyx5tkia4w3JETdU7iOoaAZn4nJ4MgUC1ilxm8sTFzcC5LoRF93ERtr
lLLWh6GF6D9HmxgOOSkM41djWNUAiRs5w+7Ju39PeuGtlgyM1d0hSWVkPKK4k6SqMu2C0zFij2Aq
rEBjbQAsRSq8UTE2mzALuUG0HCRt/cc97kMDPbqvtXG0fTAn8Tzs9qRyfW2cPk6uNMesf3X9Kdqi
Iow2ITRRuDeFUrnd36HgPMy7L/SfZEsAwOlRibBF7s6o5CuZCjz5ntic9ecDo66douCAzSupUxUt
WOm0HcnWRKpt4oS0dfGt/feZfQ2PrC/y+zXlY5QUXsPZrMyIMyIPOYcimfxfI0dkFH6Qp38uPGbf
gG4961DKe1yughY/giRqteJAheQ7AsFfenWScWmRB5v9ae02+x+mmXQm+mt2aNY4k/XgHhL5eu90
UOX1nJw8mNK/X+D71OmEFyEfjDDMYXX+2713cv7VTTg62DcBlCJo7VOcee5yk4dLjhQ6kcW5VCOB
Ek/fvqVDFFYlLHaRg+4Co1Ff1Adep7jhy4nmxUdMOmwHMMEEF5NA80oX1kn9AqFfd6Xwmrrpv0A5
826jKWDtoORPHAQ/JJgXosUx3qgBxxyDvRGz1URT+qBP6hDX1JubfCCmP7/MMrVWMbrt/vIIfQ5x
KCiQ4fQEYKrZ7Z4uLDOSWG8LsaqgOn+QB23j0OeWEaKle+nomIfQh9K/TqdnGOZySy2tQrke9ytC
sk2AeqSPHBHCAwHLe/bwKslbN/0wQ8oxB9uEyEL+yVrVKksampnEQ6sF7gUlgPBqQ1nXL8WcTn/a
mcGliiEuukofDfGPnIFSWKC2NR34d/ayNbaAHPVy49xEWDvySya8mUH0AVWz0qL+dsO2UKwMIyPk
8f/6PgsfXeyR/S1yuf6PQPWVIb27bHf5Rpx8GTHPQdKAg1OKyQfejetrozKktYy4mENMvJ+Yucmi
zjQZOq6WRLiVvoSg7EROmh3dW7xnxv8nVtg4ZuUUcNpj2UxdedqNz8yxM3RfBeJo7Uyr6ws7wF8E
5B8kfeCQyDg6HOucAWexwkSBZG1PjSIIbynk2C6JjSEoq2KdgE+6LdramFtTMFJVNjvxMvzcgNoY
Fw4yAJk4ptfg6TColy1gDTBtJ7Ilyg7leAV7EcvlvKWkdYHkl/b3xHut0UEkVIKbzBWUyP+TG5JX
fJUO1qAtOpuB0DYA/KZlXJ1LrTg0E19A4beTk3HdNoYzItTbJS0okupv14zj4gwRRs5Zs1LlshGY
XXJJ/rk7M+exjiYhMOSPaWcqB1l4ad+7Qka9V3eqqPP//AJvL7zNA22j0uIk3xMD9AV2oyMnJZX/
4Tm8WB/2N50mFiEZgvY8Pifx8k7avlRtSdISTrEglXUZpIuQmEpHk8QdZmM5Vw4a91mWLojUqTLx
Asf8eMCErsTm6fZb//g7ZeR+1pHXkfMyFX8Ex8dFU6WupsZZ60+eIriU4AQHiPsvtHIp9GM8r2IE
5sww8830jOvmCxhSskVp7Sjlu+tRKh3SBApVjwEmqeDrUlU8rzbc/fg8g0pIpbe1vg7DuAsE3xeI
pLSpYr5dtHAujFzDkXVC1xqQPBzO2q9/3BvLikCaCJSXQR72zBHlrBPclYYdTw1UdGqxCgmeD1V+
bm7aPIlgw4dt/PMm/uMrh5PmYJ90BIhDIvoGWc5U45e0dWfTabHBYVj9C7kiDiZsb8j8P+0PIe4T
hvTSotvCYDw82Nty0XRROjIaBTCi4P9gq/vGSnZwUYVdzZpAcm/HAgH/24QMqO1om2RMfuv0OwjC
voCtgsNr5RcoAQtqiOKkPj/WMz7brHpcWdf4Hj+tUMecwW1ICaxFeUBsjUjwpVMQLnsWhUEA1R9A
/iPeNZF42Ti+L9n0MVK+8Imob9jIMHrCgx38OGIWfEW1FkHMtRwTJkBsuYyrKIs8JEw31YVh3n8S
RnBBtv9jcGNEHzR7SDjelIfSzh+QpHEeyNDRSbkGLVdGa/GAmAwARg3AtIRW9wt+r3V1AjoHt118
Nm84Bl+2YWOzLdD/7GWQhVea++QYnAzJlIEj9/L0/mZM7rcNy9J0OssCSWaL0hz0R2yvorr3UkQc
78xCrKO9/zMV0qKGXvxsBXii+UhzhFuZkTvaZB8Fh0YM0H1Y7R/EpPQlyhHL3wVVBLJ+LoWyMgxH
wFRmAB+QFf/9BX67jzC6XsR/gT8pVBOZDnDJupcl6UgW3m/oRUlnWeZWYmyVibvybXfOC+ZRLgon
ao4cIqTmVB4bsfv+f1cVglGeCj0TrBpk+Sf6FGIpaFMpoetEYdKt6RGR6oSE+xJnewDee94km1QR
4ee7ySHbwsecAYlDrBsSecHCdGKk7PKSZ3f1NdxGfHhmJbRdtwySkneoldK4IU1x/ZG63Cr9l/2E
mqIsEer2RUI1rUMQ2SZINqUpRY73biaw4BZczWpgbyUL+5QakA7XPH38AaTsozFVZ2emsV/+vrpW
22Zz1y9qu7XpEjqwznu+b45+a9K3A2dX3OS0vlusEMd406qT9QJqeQJCpzD7QidvV8bLiXrnjsjr
blMzuXisGw+ZPO4cn2yJEDQu4gMFfbeENeOuZ9mqwHzcvHpbW3X/+HDLDwjN9WumrBffEY6cuy/K
opCZTLMitP9uQtvLEeqy1nP66HWCRFhmwcQOyS0k7MsmiBYglVKI9j8I4317OfnTPVIPrXNBE/2z
7xvLswvGoRnivGHOUQAbbREow9xJzgF65G3PIS8JEh+rRAHXagmVi3YKpaLoUE3axfr23w1zUg/Q
OmSLWvqV5Gmr5ZwmVcJVEJgY9AJOTmRqwa0DiAzpYqESalFflV2wc+yOJ6zPaZrGEj8jF1YVQ4CX
eplUt5tKhMQDk/JNmjzvivABtJW69yn6ijx3rhi5uqtxXkZU6V1GDND5gWK2b3ttYLUNBqXt0AOK
UPOSQ5VikaYq/i/D7izGPVRhfoJq+3wKoYxpXhq7RL/5gIPB6TsRvitOurYY/miOF1GL+Gkrnxlj
RVZmqfkljQPoKf4qJhw8Ms3EBeHzNvgx+49C1aviF+7xg7nSXxNUrxGrC3zNOem2JmuD5JdBmstu
il5xkOV/CpTAlzOc4Z61eCdpyFOYmAmja+BxmvmigNWGYyLE5plU5HB1CUNElXR8QEslaKUclDh4
SYmwq8hv8YFhY7RJzVsi+sIRtNNzpEZMK+ksEikHfKG8lyTn3P3qf/fKOaPvQ384zXaER17cbUZR
Lunc+RW2scHqS5oyrhzD5MW8WgPaMLSX6nd3jRyy2N8HOKdvNF8ejB2nhph4GpXVuqIo4ks6s9/P
XPzSBOskUIVM3qWc7YPRGaXf9InYVVsycg05/NtfZvOewJrJa3ZL7C0ONDoyip8cnm1Xte8w/HzZ
5mXoNN3Q1EbZPs0vDLIuu+XNxlGjIhaSlvvAjuES3n8TwVxSe4UzfrdLKvHZs6MUF8CMN6PZeR0L
6fmMjuea1O68WbZVO8QJWlZDHKvd5Eqn6lB1Bx1aegWoiIW5/Y993NbaDOcpR0pN4o8oaxG6FLO7
2YG0efgmAJek2axR6JdbK+5f3G/AYXTlqC2EvAz7H3SJC25MN3Cra+Yoqi4UYf0kutlKyJDgqPof
NdLZ1B07uFzI4yKlNZtxVB2Lvy2s0k9lXez7kxFX5jjXZNG0cqWwuuTf1qVnX8vC4XuQHUKxzuAD
5k9Q21dHsssFJ8JsGjY+hXh72iPxzVa136dPDn7UtQJMPBGhIxtG9nv6GNFvViLzRHthuZmOjU3F
h6FRH7+HjJfaps1bbNugvk/KeO1BtgihUSz/xgEVCMl2ZNMzDJsUCCk/iwhjJXWuj5PfY9akxEYh
90hrKVHqO5A0JhaVvE67/QKY23XQhmamSM+izz4+upd6Tvj3H4ilPq3h0YPxuzOe8PCbPIRGNglI
Sjqe0f8o1EnnnLuz+ApnRDIGngt8yYXNDdCRiN1Fs4xuYqty/4F842z8SAWaloWV007UWMElp1U4
enQBdtCib77rNomXF2ZD8BpJfzpLRNwotMlyBKhTaQdEXXbDj3tyIcDjYBiu3nq+Z0snI4epzMpK
qGxTzvruIAy6kAz0l3ztvRfe/edXCol+GlJO3jylpIQqol7s1K9oMc+2SnTJJ1k891KCGV+9tenD
vlwa5M+RgyErA7Pef+2U1KOCPCjfDp5A69S/HfTLfQbzfYOn6kEZwpIAUiM60Qqu5Br4MDJmzH/n
beD1Bxymi1PHz/hn1H1IM1NV3jF2rwTxMpg3q7oz9n2uKBW4ofFfTRL61kIKqQkfElUIXjZh/1I0
rF10bLKXaG06zm6VT6y2aLm+idOFwyKvhJjZDhfa4fmmrBhtOIiDrI9RwKOcsPGoaopm0yXbCW/b
0M/ECGihCz+700y/TSW0foRX7mSs/xsdM6xJtKugau257WwAU9H51CHZD6zeCDzez+Mhj4RvZXc9
NWxRG5mYBT/X+ABhwxUB7M9kdUF4IhVj52vmOcDiBmf72xyAJ31mofgJntUUecMASonSCVRiq9EG
Nl5BG6a+sq9wHWkyeWs655P6UlIb2d+VF87mH8XifIHDgbfOTOpJ+bzJc3vz3+5CXJQchT4K/Dzl
TQ5zClWRGUKrw50JAqZKN9FPJ0BYc70NSxrAbHxdRbLpnd61FpeGhyZ+xbdGXDXkOdFYayyYORbs
JNejHy317AtAeL/oZVThSMQ3kUDOMXA0Onlk4I5R+mRAzJulBmG+Jaxi++MjKe245d5FO4HQ3s0J
q8riTnKDLSoXEj03UiX8K785OQUfjvRg3dFWB3KaSCEi4Npmep1w01r5Bnmu7pJXElGj+/zFk5+J
XQznGUFBXQdprJ9SFZUgMm+bhvviBPKDIpqrD5h+nfHFanZoHzUg0sb+NCZ8AjClTWWTFpXEeZ5Z
KAtugCJNQtUlAQppP4Ebx7BUhdog51pvz4zHThNnSH4txqhhtKCtA5H5BIqhGsrCN/k88pRn9ho9
mKFAnQih0Ncwm4SZj82yX6z0G0Dz7//vrGWkBgCndUerZumLa1oGlPmmvF70yW3ZXOTUbmdCaipa
mz36mRMxCEzGXYsXf4KhUzH7iVDJGbpIEIAnMW4GfniAcaNa3XdxA7sEstMXBK1Vh2/KI9YZM9H+
Y9hIGhWDFHIE4Z5YxXuhwSxnO1Z36kH5J2n+G5zJz2QTrl4UjyaszGoVrc3etKYyY4SR1frGzMGP
I/qfDe0z0KYnJKav8Yrbe5MOsF111uAtAVvgH7oJiv2gg8Eic7RvhLXI4k+woxQEIE8QTVxnPSMa
UpLNAflisbP5OjV+XaXskJL+xuveu6eaPwValvrS+A0T3cJEu2qEZ6nJ/3LG61WFSB1li5/9pujx
N531I53/xKQMYASezNXOY1NA55m6mWLaA5DQITkAP4yj3gj1HsJwHdZvTqFFWHpi5o6DlGCmHIzF
aogqSccVAtkD6YRGbC3/A+S2uCunFxBb+dmYEI+UpPwdzY/qA/7YBWUS0ops6NMZ1bsbTMaEtXaU
m72DFrHxcg7Mly4K2B1U2fdSSfiRsNolvz6Y3dIsbgkFFLsjbTSk7CVqbPXA1uhUGPEpPH+NzvQX
q7jLjMogfyk+ERzIux/WxocA9xhVwg9A2LWJqthcTZX7hKNyiKdYJRrDDaxwej4zbeYWbOB6mbhD
FSwPHCVHNIf7jPZZuJrjYCo0zUqZ+s4C2rp3FuocopbxIdbj6qGRrzs1AtNYhTtkxB9p93YbxUrr
VNHckGe9ULKLRmOcby3eps84JxTL0H2u2MpRMg/ti4Ksy2AJ9qTG102FCxS2Lts4WZU2GuqOoXoH
cJSFTQ0gafBKFgQLdD+yJYKhA6nhQJWmxARnyfBM+IZWXQWHS4mIFFn7zUqtD+FcRTFd8mPTWcOz
MShAYtXMoMEySKUXgPuzogM0mAYuEtd8u+h+swskIngYqwySpUarYo2UrGqT5CcQDEWrIu40JEYE
iD1KT9sGw2+F/pwg4fF492LlhYW/bZcI4CsAFLUJZFClGqTBC4Q6zlyW1K+9Yn2PN2srJtiWiz4h
QNXXRRXk+QwFWePRo4Jwtg+E/A6gYa4nv24Kb8pSN66KDc0TPjqLpllHBPKJ+MwoT+hkX/AeGd4o
ctUR2R9+TrsI/hncBlSIl+kWuPbRewqtorLgAqEO0ho6MdQzI+ZzidrTp6Ru92n2mTr9K4sX2IiS
EgKcST0IhunGIHKCxSTet5WRrolXkc/TEl1wyBIJkVovb6doolZOwBrKr2kpKLC/yP5EAniraPaS
w8c+FwIneiLIyIMFBstOWfjtCdyT08pKpjndzIZo11yL8PriH1H6uKueZrcDQ57SJT+LPafzUu9x
sSDP5W2KJhKiDLPo0hsO+s2JA8/qljJcBe6o2lbTfwk/BgU77y4jfgAn0xQ+DJYOXD+4hAObWaWH
MEIMG6nlFNIQpTzPxUEgh3xdTwxBE7Il7u2bEvKW7uc3ogqp8hCGyxgEelHXuzkyXmPpWbNhjv6B
8GZPmIndxtdGBJwfctDKIuRnGg71RCt+Ys6h4mFMm48mAdm4vrbn5QpR66WaISNfCNrV85702y0m
Ir7FywwXo+3Rkq4AJVZry2LfYqa4u6uki3GwmIGMGDoD0648Da1vBdf23N/7Nl9TkdQKS4/ZiRIj
satvkS/8yz8xfdbuWQjlzf+azO0ZzooRmHA4V5YRFkHiTyDP7UhtfAk6O1wYeHacJ1+ujNNQU56U
/P86CcJ+FWgK1SYIXJIZ83IcOHrZFvczOIOR2eZR4ixdDexmMkf8d1t5huOPhlLwFTXPtykoEfPN
J+iKE4XzLYceYAk/AtfhuBZIuQQ9ZODxub/nUUzepG8Ept3AYvvTtFQk3e2kxFMQxsY7VNqgenIx
xxhK5C+RxFtwhTzipmuJm64Frp9Ife3K/U0Wvv584t+MmsrhJyM80St21K90vUgGo/rKA0Aefbr0
MecZqvpm/gykFxvxzCCCJcsf7J1pIFdUgJG0rT9ODWdUKSuUrdok0Nz2Cz+n0+JVRwbsaJK3tzX+
kdzo+51D7ssrOWaiDivfJuCHuVRXrXZboVnwpWy5qX0yOIKQNRmsZIr/H9Bifi2q/5P4qeJjTrRP
k4l+QAz1EswCYI18agH2Uipm40Io+Wro7Tws37ERhEsVvVDOnca6v+XHqDMwKjlzMiONNmOMrUx0
RLmMBaoLoeebDj+IHOBDhM2RMrixrRdbIN6xghGsTeD3VdKT44p8METETBnu0KfD3Rm90YMSIXvs
koAwwH41+R4AAZ7wZ5a68RzHP+H1kjLw05keu8MT0fiFJoGuB0Jj+RwwKXLUal1bzA02A/Mrhn4y
P1ebPJn5+Y534Hvvll66PT7Z1HyJVqkZ0s9go7pCEVAzR/jtFelrY3S2hmk9OkMYqLwWQdjlfQRD
Viynmqu54kZUJyh5RAPg1JqHbKH3CO8G4GkXrEg261WTVQr7QZ9NPiSJ1Awm6JMDiOSlNEbpNz4h
wvl8mD/DtCkiLE0ReOCgY0gxcKvk1wRnpmFTwub759Oguknejn055M3iUG4XxFq15XqRrC4FLtzq
nciP3Ku4Zwf1cY3zjBz17w+Si2hqrtwPvuVxnGPNX/nbZij73PS2XP47swXDf9QzPZNO34MFUT1S
b79PRn7XxZo11G4je3zPgw/QJzaXgiXazWASGKdc/FcV1Y72bI9l7Ny92sj9MGiGC7MhKqnEOTcP
gIGy3qa5EKiJ9yAi2ILRI5pMw8wKvXeZ6phVbXmLmIqw3s7rEmM+7FMVvfK9/tD4tv78Eo3RMJwz
kObIW1hVnnX3Xcn72T8LTlBwI28pktpIN7sNZI25CEiE2TwgqWWx8Y+8cUZ/XjRnRAr6vmkDyUv2
ShDuwXFsAioH79H4cpnDxt/LGugZdQXEWuguQAEQ/8hHCixn9FoJNTtQCo3a0c8/RahYHiWpxIt+
z8hBTAcYzEpg4d7C9TT/X2eEw8Hv2YFLOkt+1KFvlvHsMMnpSH+V6P7pVInJJzbMeSUkh2SP949l
8vZJ21IvV2fJl1yVlXb/BjPYN9eHv9oYHxJpICq17DxZoydbjZFeo10BaK9fRyQyqh989LfOmJZp
N5sK5SsZyhSARxR1h+/oM86j3EPJ52vC2b4dlijaquhAl8UhHlThaqRUM27pMDCA4TNfyH5lQAJv
/80J3N1EuOh5IXAefdly4K8TFmTPbO7t1sQ9/j2n0tdV6whjSUmdPKQvumWh1AQd/7u3I78uz0ym
m+SAT+d7lm/tJf4WQTCve3ouIAIHWJg4y7AxtScDZOYCm41j6ZZqHFZmR7LENIMxAK0EPeTVkK93
r7RwPYJTJoMJdzW338xgMtyrsBGzTQbMJUQopNpkZYcLXKcsEfYYLqF79tKO6tKqJHpyNdgyVPZX
PXyauTlTNFshDMsvfYjAtvtR8ISgjax8YWrhHN3Cc+xfbEHTt7bK47ZJNwJ3TDm1m5QB6/G30hBL
ZvqX3smcYRYgvSnom0M7B9n2pG7Aqet4ZERmf7Wl0QDIh7p0d6CGM4THtSGhYLSMjS394g4vmDjF
EKWkPoMfAYID/iZ3pVsLYlFVYcfnDFhnEPjX5TI0/PbHbHkMbfa94DcJt664sXi3xp0dbv+R08Hg
8q3bbcL1WrkufabqFFa2iyw7dtax2iDA87xoeSaX1uGDxof6n74LAWRM6dWVjAx0AHswVhqfmJuy
YROZo+fHZPpqseGoA15b7xU4E0Lq9szqnywhf5pCVfscdUx+PUDdoR65/uEfbk6PZhwqF+ob+ZUG
L1KZJh6H7SrGaJicjzyQlYqOGL6Cm9a1K7cJemHHxYFTe232LXf4fP1VJULO3rN7l7VTqpbSG49G
eb87wwa4yVw65jjK1DsA0PCT930QOWfJoKgR7nsiza5mQM4+E/Ee7UgMmideHa8hx+Kskj4odnvY
fNYULKTzDcZ8RfOB5rSniDU2kYGfGnBO46jA89BoXxcsi/wm8BnRycgaW5QxpysmZzfMG7E0CPF8
0xdNOiemqfViCJfyvc3dUjjHFKhtHes1okIV+t2cAvLWB49pF0PLillNK5LErwCO1orXLmTIIfY6
wr+kC5qxRVpLAdLELaiMQ35xG19vKNRMZk0F5QVmOJJb5/0mZNE/DHe0gFAmfMMgybOXU7ILrwpH
hVq8ctSxoW+H2fGKBLsFSFhdkrOv3ybR4CzZgq12ruMh4+dDAmvt+lwyZbVEQPVVdhyVcOrG+hEB
36p9AI0+HuSwBGKyioGiaEf0Dj/jVPwt1wio/WNRJWt2dEdkcGXi0bpIhnRKw7DGY0nOP0W0h/fZ
ni+ON4qwj3oXfmqqmk/J+ot1Q7IVPIK4jO9AH3DxMH0fiUvOLsh9wE4wtDVQf4taXlYJOc+On2Uv
X4/Z2OueRIWnLZ6rtgHlSS1Iq0wWcqrcotrhcNasFj5kyOtMYeO3ohWT3+Y0naqN6Iy7npEMLxkJ
DhtkansA7P1B50LSxL2KES18w8ReJTRw82bYR4C/cwHnPDbY9vBYHQiu341ImI3dyACVqRl3C6f7
+2p14+aJrp1SSzEQbzqjN7ESEmiSF1BKPIcad8uXv6ChQqeX/KkDzul1KaNalaHUW1XZmRu7K0gl
M6ePJX6i7vfIpHzaPDx6Ab5w+zzIR+283DNjHlQkYfcaE2webgRfHahfdsi9XzpSf+5GqQBM7i32
Tm0IkirhZet9p9YnBImAeh56tqtdkwLl4cMo25yb1mozx+1fL7xNcIqK5GPgIKmAxm+PGhD5ON6N
xVbp90QLAZw1alYBoMGEKbsLCl/l7N0Uwn+HkTrPJGFA7BMji55ZRtWCCaPUeWH3s+tswENqTMyQ
/nF1mhVgy7+AWXvRYNa9dw6jujzE1R/TBWRPJQO8MHKq6N6wD1zecuf9d6YSsS7zjWAHVSctuwoi
Cd1LA0MBlz2MV+2sXCEZtbQScmQFiR/104FhRlAgQnPNN6yMbgbWrqWw8sgXaJrMqNjVAWnI2M4+
dRJdmJ1Q5XuklV5guVbVHv3VCaUSFnIOvg05tGMFMLyavI45UV1uDF4x1ai+0GHVs8j7vAhssSEj
N7oaNEGnSkYWJIgu2uzQfCkqKMHlhhQFSSGr73Qpw99WwoVc/01PhjlWdXPzim80/RLfvko67eZZ
G/LPuwSeQ0zbar7wU0HGtNfeFy98mxK78OU5GwoMgj8xVNFORFeNVX5u9H7YdY8jEC0CPMAgvYEa
Kf7ZOWgvfksJRnwsiIKPa16bD5nKkS0ZOo3rUm8ycXo9voDvMlC9UKjWOq8V15UPW4uncMmfFDdO
f8cD79AdMDVkdY+b9ZM27fLQN5SiLTx/f789cSl2k7g2kBe87zRmPFEhUMp8XVkdVoumolxUdwz5
oVvedMxuJStSVRo3bAglQtKIBSc9QLQkYZHsI+tXHyaytxhnvW+OMxv+I4zlbBeYE2c8H9rEqc1W
ck1dd5zq1FZRMQCLkrRtbRmHjGzaRIWDzXJUMVPNe/IPdAbmTpJlQFx+g2MenQAjUGHWMxDmv3/M
60CeWQjkx5rs7Xcy8SbW1KNInIgJFVSWGSgO8VE6IEXTkQYA24ydiPkOKJFMrGiNcXl9kDnSiZ64
LCsQtAORE+vqI5U3hYQ36xHVBowSdcRy/5P+UDOHdvmoa8WJFT8WHyHEoBFUExo0JTgzp3hICQjo
k3gM9VaEK1TlbcIKdfS5y3EnT5/pXzX5uUQeQyZAP1EA8f8vr1mDEKpsro+2not86Z4AvST7dKRE
6nnspxld8bHFOX2XtYeZaZj5N2ToeYexo8r1eiTV/ZWC0L0xGgwjgu8hH35tWR/LHTYVPqKFDXXH
BL+o/6qSSwF9bqNWONajeMQbO6OufYTnmKUL6pgNEk8cblwUTPLkTrr21zAbF2AFLyGgVfCzurtY
khFHrZkCdTxRU5bVVWWQexICl/TIllf5fAgDmNaIEjYIGCTmRLOkc6I14FfrKAke6L+CfKXYmhXl
krMAokdeLoMrHNSO/viycIqBa7XLQ46dNtGpxoVklmxZ9kihg86g/rqxFR4O+tOlgC/QQRwL4nEF
P2VlYUTK/kx/cqhzVUUn0IEPcPlxz/J18wNycwlXmBmkvmreSGtGpN3zgTMzCeByfPbP4iN++C3k
bbMe7CG29Aqb4GFrftz7R4cqiizadpzHUKTGaWZswVDmSw0Uq0kHj1Uiz6/TDAg1gpPnmkpkxWmX
Q2YVquK+PxkReAm2Q3+m0gBp8dLJkpqW3RCVRxVlp3c8QFQSsvSqwgvDkkBWzWMSRoEu7wERbMem
KIDmzqJsqqVxv7S0l+Oupzy18N+WJs8knJ3Bw2ug5+92BXLVQKPYsK2bY01Zdl3IISsnOzozyaNM
l3IsjoCGwa0lZVGT7KBrxUZ6IEyz0JWwvwBhsfblhxaoj6kTISaV/eV5Vyy5TKHq7nTAv9LqWORP
GTuPaVUjZ7a4eSI7vNH81RJa8YttbeRK4lx4rKJBOtZoBjWInYAgU9QfM5paj90rVaNy2zs1Q+1b
J6CiTuqSAZIVILIVKZmCw6iZRJcbL2CjQonk7sxfGH4QbCmPlXb4vETsSz+iOOFB2BBet2gFbKKg
9LmjYdHD3FGGrcVoI0V8pJjYCtywlqY10BvVdRyah/ESApN/KvFgsT+ZtL1MCQcn2VDP92FeOYFm
r/RwlAbZNqiO31ScJ5DGojFWrdguF6kOPzsz8kfwoT27+0BV2qZxYcS3nVg5tRQ7KLl6gLO1Mrp3
s8+j+6pUcSr1F8D+vL8Cb7RxrU9DzPel6/SrhpVlLG77yz0jB1ExcjVlkAjeIJtDoUu5zveVFTSM
oqMZIGTOdZVgSsQYL685BG0BkR9TGR1uT6iEb3K3+3zaymKuu1CaXrkMQh4Tx5jHt+1bRoN4EjPo
NKMbE5J9968PQVWVCGrGy9NMoi4ryhLN5tBUxkZzxX6OP21o4x5Is5tb21EED10e7ulayygWJzrE
vYUBk8j4wp0Wi1daO2Y9Ge/jHcLEb/VJ3yTbcM0bn8i7K4NhOFZ+ongpUxZK3ZXhdzl/YNCKs556
MPjnuNh2oWVlcjmjcQQWi2ujZkBQecc/7EZdJk83qAdhdByAqIbZBe7fhs/b7M5hp6Tpv5AewqWe
Jq5RhrCnYcsB9V/8IiD0zj3KKu/zyc+srwqpm+0Fl/jZ1IrLVIVo7Iq1/NCJML3SIXB8beF9sWoB
Xt+Iu0n8BW4/pBT4j3OQe3bPeHNSgVqDv7ezNTvmDU0GANtQsCcN1AIrWLh9Lh7QZVGeSFnRAbkx
dMI9x7u5eTSahHTGraTq8cLAX0OVhtdcGcAdyAT73rPl5W5i17G66tEj8+V1wmSy2sY8oU6mXCP8
SImVuVdJnn5cCoWS9CyG5QYgH3e9IyyNH2MLwClKgDSmODRwgyjYySZ/vMx66OkF1yrpgqqT5phY
FLhJxqnb4cYA/VcqEhdcYsgsRcFNLpwUQfiQ+6eT9YTnKGGag6ZgvrFTh0fpOAeT8pbb0PZRQt8J
K4vc1QyDOpyMq0a9JEEhCGwaNdkgFMl6BoZ6QKHD5AOJgCscm3Z95XvFNTHq/viAn4trgWLX99j9
vzOKJwqi9k1nfajvND+v+SQQliBsc6AkLdy0/sfeFylaiCh+N/lOKT/u5QVEmvha+/5gN/ndlmYF
PnN6Py4PKzkPSHUwiCzu4UjbrXfSgwPPoj0+w6uxlDMwgyMDlBeK5c8VJFcl2SghFtBWY6mhqi7k
DgnoEUgYRmw7Pn/IgeAteseX4PdfLiIWJkVoApFt71PpW/P4vBo1lH9Fhc6h8wyS8j1hYmY66RHT
YHj6iZD683ZgcnfUZttsPfEAkOqNNCI+D8b1UYuhLOfkTAWwtQ7Guqn6kXSV67x9ieoEhoEqmXlx
pZPDkgfyD5UMu1A7IGmiTXFn82GgzhL09ZhnNNAlE1nIsJOl3zBHjVmJheLxhIx9ElMowZvQoMGz
ycuLvWqR++qSCFtHHOmCgRMsqA0MCJD2awleR+pfk/RJ4kjL67aUcu3Bs7tNzdMSxCFqAWV6QT1u
edOWcVyNcup5vqnY2jlfPYPQcSR9Z+HQtPwADjRZUaukXbZjTgnG9yGuVnuGZ5pqPZanZqkwCId0
8wwlaCVogd4W9X4MTtfyDYVeWJe7FVkqBk14no6A/xIV5POBkRmfcfx2pHxIAswOqeXy8ExETY4+
/qdE9WEZ4kWO2ddnEKB4pj3CEs3aKgkKdUgeXrrMkNaMr6AJqHE+GnHMdeziWvNTPIjqoVXpDsDw
aoaQCIrZmGkKjpcvBtFGUegzHyo86WJJ7+p2l29mZfs/qTeF0VA+n3t3th+xboPJuYpKNPuzjqs+
OLW9JWsDERzrO7mqGtJpJfVOppLMWIPMTIRhXfi0Ux8PHzx3True2jR4XXHaV+i4+PSbGDrAXVd7
1U28L6zutab3CtNvXP74BBcMS6cHvfUGBtd1IswJKNIOPyAtndenX4a8gzQDjZvDHjtnOVMmYWmJ
B9GNP6AnXrG8biL61noJ6h+aK5p6JfvQnCvIUjgB+4iyJKkhyPgJIJLJxAfpmLRP1rYkAdySa7wd
2ysfUpFBDp8e9ontO9VqsyT+e6bqXQ4LQfdJCIIpQfbHiSjjSSQwvJNFBA719chcFtzD0BDGebEl
A4N6Cb20GF7mR9Hy44RsNUVxjlPg/VjDafttV0opx4kkXQc6EaSgwDUGD1vfwa9ByPOabhOmk4T+
lydpKabdxaE2W3zbtML0rksz0o2UmvvL83ygR143zAxl/IIuPyvPo319Qkn+YbHe85m9/QBLupTk
5sUYYY6tg5heHgdKUzL6FNfugkkY7qE/5YQ2GYWD9EBYFq6zxMRyRHeVFvXeiYzkojqCSABuFXQt
sNf9cc9WY36SYYKYi2J0wqpdV7g/RM/WaV8JLbVvqxSICb2JIv8/+QhKZhUiBqbrIbiyjSY2hVUU
QYADSITNuahMnU0avCecFvrr1X0dA40SkfJnEdWRmrdSsDo+eEflUPHhd5+qx2yRuON3LxW/oiiv
YNzXN0npUfPtMdL8vz94TW837eSCd9hdo6w4k8nNRu+zwHPfp21oQYVbF72V4cVxsu45nyKMrWBt
SElR1BcQhX9Cu4pCOyTHrC5gNWJ56B/rrNbn8Ni3vrc4g60OJeU5ckjS9acXFdJ1Z9QHhGz+ZfJl
9axx1mHGK6KvgT3b/7RgD9gE4ow/1qOLFvwZYGlQ0K4QCZssQsJOZExOy6WGhuzyKHF7tT3Rs5cQ
jJKmRRNUFewzaByjpeewD4C7LVluVQcX4F2isLzUPAWspfF4cxSLsLUy5Wi0iyikwdBtKLAAFKcz
e9lQoR1t8YrXeKJYOcPMQyE7Qhbb+9gITJpNNx5FGNGOqCXw3h1UWS0wZD547vmYgqjc/3fLBy3Z
SEdqOmCRO5BMKdgeUlTZfTXQDAQ6mZprQmkGwTSPn5fDqAulZrNUtMVLoC6T2+brT/xjl3aNMRoo
DZwJOlKY+e3tiJLpFdh2D2m/8BB17kjATxp3KrLl8pdEsXxDZOYrmqxdlOd30EgwV9AK61TORP9b
MCQLDwj3/5Y7d+rrmDyGQOdwWiPLSYgPoICclL4aP3ivkbDl8EakEYxRe3T3VGT4aiFYDP13FVgz
OL6y1osBXmcAPlYkTz3YY30TWWChskJ0BvXqz1cSvIk7kfgYeTypbl1cdDwNF1BxvC4Y38uooGNm
6BJ8evboCF1bLRzz0xBDRiQ9hIt+JX9vMq4fYAlIr8IfmVZ2y/6Fe0DIL7XGJbie9SWAxlMTQuIz
WbhzAIkFglSEJkE1wYAfVCZW3dZLUotJJZ/tjXJdH3uCCyTHT79rFh/SP/f9wO1xC9jwH4t65PgT
/fEz00zuO4G7is8c22ZWuGQwyR9zb0ypwRPJr+JVSVJ49LLkSKhuV+EsIG2jVO4nTOEzuY0I3rer
Bfu4WakjYL63v6I1jUwrNT3Mfp9LT02DtEoB4uFPe8W7s7vDbBwYO7eBWz2r4U0Czhi25tx8kZnw
Ol2YQdFMdTZFGmWOPqKMskCxw5R31raMoigewQ9Km4PoPKmWWsGJsyQ5aH4nqT8oFnKCgWP9Y3Go
1NfJd/NbpfIWLktxr+sr4rStfuKavUAv82IMHqJ4/YVbco1Dp+BlBSEo7Q2HwZ5QjuY3AJ/sjGl3
pcO3PSGLSS6Uneox1HOpUKVkh/N8KJXv5KpKLx4aeoyeUcYN1yZRAecwB0ttWXeL/9ja24uwRboB
DOfz2gAtE8EITnyB62xibwptSI/ojYn5YqyplMW3A8ERUvUVJdDlOiLgnLeQciwg3wM6TvEkfHco
2jF6esDjYuJzXP57cGzAfFQMBmjUQqmgXccq7uMJHQcbzUpY0bNNOkzQeHQBvmKvD11uNOoLGJPx
fenrSVJjTg3eX3+cgbvdowQmn89Jg7obrfbAV1lR3KZr1cNV8A9xHdExdjQy4b5tbjxDcwxdMTEg
qBzmgwVM/ODTphVbJ0qcn6+k9xH4BFlf1oh+y7VxBsLPuBCJ3ZThwo6WPCRd4YffIFOwL4TL0JT5
LHtfKVvmuEaBBeBHOEdIEql8HP5UAMV5t64McgaSd0UPD3k+gFMnhrBiP3s9OunjZv8kVRFhx+JR
M1PtVhxOfumVcHHK/0ip3WCrsSBzlSTMXArOlXsdOrELiEA8SQ8+SdRvpvburCw9w2YFd1Pk5o9e
lI/lWefP9AnARZZqRWZwlRLqJ4vkGM5rP3OPcNQ0J/fxddObjZ9u7OZg9skZnn7DGNb0wRaYvbKc
p0Xzkk64P7z2L8UdQezoDKsQ9VJs1MylTHhZeYJx+VJhLAkoS5UxmsMEon2PpVrzMsE6iKiAHBmt
srQ+gyys8EvLyBUG+2/wgzte3+oqvYRirTVA7ZJ1Nu0oLEdoOl6LxZcA8KvOjKTscw0uRM9Mg2kR
fUosDjbavDnLEHnn4XFa5q9w202Nd9vxhPibJz/uNXx3eMsNa32eiZmLmxggvXp+3T9xa/X+PJA/
76SpbVFP+bi+oqMqRCpAAB6JZA2yoZQf7OAgC3AujNjHH27A/4IxSAxzpT3RkaP6L8tA/RslUGch
ccLP9Gk4NtoDt1HmSgEFcE1208cWZhmZz0+ssej7gZtiXbHuTU2OBtJZ9ONKbOcK08V221xxNXcd
X1O4MMlRF2iC7y7jYkQPhcxnuN3fzz8lfa4d7uYDFCAU4XwjM0oqpDe7P/r9VWfxkGQ6vDSL/NfF
WLswVmQQv6IrVcb5TSY8UmaSWkUq3b2aP6o8XLJvloVvv94MtFcG3grMIQfU9D6qdJ5Y/cKNOGjV
k7AX5XfDwWSip7G4SRRHlm1Tm5DejJDsP50/AmNYOUW+sUhTr19g9vjvULWD1ns2xZx9mvqhmVi2
Fa+beaGP96zRaAoxd+ZR03nIxg/DBW+BbNaucdcqnJghSKMJm4MlkNV0+DK7aklkBhjN/xFukA0q
hUyheF99NZIg2Prkj9VoELmjGb6a18J/Zm1yu1IS3V3OEnaYGnflDzgGTmla0Di/TSxHiimlGVDo
XIb2+2YQgZq8avxxKkAmbye2kpPuFC25ovN3va14VasGapq3eLszRcJG2SQiBhpehRaNAcPZT+kh
cNOevIgwRogc0dr4OY1nr8RTT5PPTNafonwN8YCpWmqu0TRr9TU1gebSPPbTshl2Z/ypp601YJgr
81KGChXBxfztq7kwCoLKOX0t/TK7nEzOPcjU4WXBnOqKumAKu8SeNt5mRTczWRXjLpxfGM7q0rH9
2LrvZM9uobueFNd4HPYaVEvfcKTv0fAkMaEkcUGmIVkn6h7DUPcbOIEVTZ4kAJJ/WKy8JFrmQKzK
edxWf4ZIr6E8JxDy4ZWhqFs5BIoWjwwWYiUvK+BLG1M5kQV840V2Ju2qgkOG12NWTPP+gghEw2Hb
iTr6Q8Ucj3TnQh0DaSvLNubAAWEqT+bDiRe0eOPq8P07x/uUgS1de9tvHDP8ib4K3Zz2XiZpT8WU
bmOdyC68S69UGrtb3wnIjN1v3ABQUGonr01wz1DiBHjYStEMkm6BsosPKkZ6cW1FOMcgHOocg9qy
19RyYKFj/wSJqW5iRFlbnWmXjxyYh5kskVGXc0hfZLAyVPYDjJYGBr1yGccKxUvYhN5OXEuDpCLa
w6SN2uaF9ws6u8kLk0U34pmAxdeS87+JeLaB6Wfh3pUTgs31gd8yMzRed3C1GgoKvPkf5v1rbPwL
uIF9UkHWD8kP3B6OojaQG1rBP+JM02XHuf16YDwIDwYRvq8zOnKYOYdHLQzzk+YEQl3z96Opv56D
XCM464o7WgFV6PS5PY8mojpVRcMHi0IWYccz8Js7dZ6wlltghaE3eq058HD4OfhTCsa6xtLyI3pS
sIKYk89EXapzoU2IGRlpIIVJsi3j77swqF72V9swc+phAmJL+T5Vp6WSdia6B/6Mtd/IW2bbNqLU
j0zdHxAsoyw4H9JphSx5qrPfTo5t6A51oPYc9mAxkjEikfhGNUQt8eDXziAdYUku7MUGVqMtztsP
4Bk4ZuphYa9DiFqUTTHUrqOfTC/ft4slbTgiOx748XgE8UQQ50cNGeR5t/3Y3RusPmBNHqymrHMn
VO3U0GdxVP8Cvrwa8hpWIjm3q55MKS7hqFEF9kYVdW3vx60VRM+wpi9T1wiFXTuxKANquPy6D8L8
14FNbonDmwthq4dNjNR9eH7LZ+HFRY5Ji9j/4ptYsLzqStFfMvAKsw+kVoxnce83R9VlzUN3bXH+
slxy4sfywcKe1ytinrFEyTTL3vAZ6Zgtq8yrJdYD1BJKPVaG40MVk/GwX0XDdgtQu5YRm0D1VTMc
1LPxv2h0HNQjrbAaTsl0EWJrSG63PWiGTMBJ1pFp5Q2sflbjvWUlXivVVo8fGDGM2BUShkl/Wueq
VNDXC3bmi/pJXm4ETDmEpeE8xhcPL18BbYdj55fb5pYyJkfADG6nl5U6bf8a2Er+kvMh56hp+MKo
Fe4qVsFxD75LoiTZRtv2XnAW70hVFIpaGhLQUo1aQwuQX48JYwdD8kSFX0QAiBf0RT76PcJTPck1
wZ8D5cUOdNaLhA159P1w2Gar0pizv5O6oCg4ux1YZqP58GdbYxxFbuJYXgyMeztWvVIGwV+ypQc9
IfkFoFvSzoH19LmNpix4tU0nm9hu/f1VYqGGfQzk/0tVUqbRs36OL6OLF1+44C32lfGxZp7LIVu8
ZE1kidIaKud11wbgzU8b6uK0CTWClNc8Kd1FtOfBr7EqGvTxsf1giU8gh7HoXRcz/31qrNKTobeo
GbJLi9Cl0BObG54LWfcK5MFCS2uj0LFzenHOfoUks3WD9Y/hHFsNweun19WafoX2Ytl8+xI00k3r
cKL4GcKwIZFtkn6smvDW1HYV+Ypmp2uiAI+/M4gXpSf1o5BrZW2z1TYVE6jOdjpWrd0Hhvv32Ae1
N2Pib52jWEg2Azf/jt2VtfndrhJJQ0XcZ7+1TT4MEVcBgxfGoAd+X33CMeZKhaEJaibwzQ6kSMpK
JjV03dDQGN8oeH3NZ1vRa4svsZG2POOaONUOg8AFwpPrDRi7plXmSjqTcLOILzsa3Xv2exJLtJHw
wvWcoBLaD1nW4Bx2i9thNshtbB1t3Mcb3ZYHPiFQX/EFjL0MJc9utENIgXzzfBOtbPXub+cFy4qF
YsRALail7LZTcTURbv7EF7rXhH5M9Pwd/5FpBQP2kngySjkjck9uZlys/kZ8dpz59FdCZ28a3o9N
lScOGmAAIx0yP2OUfTmiL12z73lqoSkA4OI00MMa8A5j3+fwNuVQr/PaiXbdto6Idq2RAdVkonrK
aCK3t/8RMEMxo1mNlLdPN4RZRqzciyW2N60rwlKBg2nvbQS/UAZ3c2ifY2mDp7KT3bUgBowqI6SA
DNeDmIO93XtKIXqswexjq4/H0tqfFL9dB56jnT8lQDWT0+UdAVpyDqBR7Zweg8aI6iEDw9Oh2moS
V2DcQI+F1c/KOO8mqepMgSweDr6pShqnZQBuKSfJa1LHF04/feCZyYRuel5OS3zxd/3wrzrPeZjw
979KBKUu1CbkwDGuz5zXT+oDJFToKaYH5K+vWEIDXA65CwftCPLnWJeSmHynD8dn7gb+NAmspX4o
3G/bIsldB7HZsvk0FNv9o0DsWJD3fE6TCpjGo8IY3pewKueYQXBCqpmIYKpkChOvRhRdOw1ZNeZ8
4ru/Nf/k8WzVziM+F57BYKrRg4Ua7awupy1N9MkOR/C4f9LpB0hL9q5GBcCtmoPn3N3K3+ESF0ai
qY7oW9/BcwlB4NIYFmrG8zvaVBFdp24Ygw1GbfxkGOdUp/cV+8zyOc3l+PAkijrIXsGp+a/qwiIl
HwMf0LP1ZrezdpQNFxIwoLS2WuMaP5RGx8vhEu7IB8JIcLHw023il7bvyV8OZCsaUwfknlt9qAMb
UhHfOwlgxhVfSohIyLOtf5QmIqtRoHxyPXt+IFT5Xl19I+UuH1MlRJ9db5z3L8v07OHEeTzPBElZ
Xl4cSh4hcbHhoAabNAwmTwQJJSMnj5R8hzZsKNOHUQI7Zk5fiLyLh397op284RMRH77l9X0ybZZL
Y1iypcCI3THwKl8Szj3C8k0qvk4h805xfPg1csyvvBn2+HB9CSUIXftbsuAfZMdyg9mDAuzGrV+W
VYXxWFUMjpFy6M2KrRhsaiWValD91Cccjux06uOYy/Bl5EJVYfA74iHPE2f/DBrEBKbe5sWpEZWt
ZhCPI5uxOADrt9r36O7v2kS7kkJsY8vLlOU5N+o6KtkP++7AZ4gG4koOfwiwNRbgxFR+umJQuk9R
/NFbD7MXmbpWFVOAKNQEtPJCSo8QHO2ip9w5Gp3fEt9fjPx53TDVqmDz2z1k8vCq9pmP+8ZkfBc9
4dEBssEzVpifyYzlHC4Ccj0wobdm8kpV5ACZ6OMX11MFsYS66yOln1bPwt79FmpReRW5Oq1z5ejl
iFCejmylQkJB5tBGdnXdrmuI1XA3QJR8zHn7dKhJBLlLnlPcD4I6+0QWfwq5usv1+rUsle//YS/x
aMOXhJgZYLqHlYt+RBZhZL58IvJGhA43cdFoqFj0HCplAlkRuRhVLFVklY1XoEYuyi1DIuFdynbb
jIIle/hqogYWtonEQsj+SgNjn47igjc6nU34fLDsx+/IjQmA/DJ6eF0Qa+x1nkAEApyy6OjBT419
BMy91tY5l4RW418cfcSjHWIQ49VEA1pGl8mCRSIo81p212zUygZIEA86nbbTS+UxjDDxYdMxar24
oSQaKFMBklc8p5NtGIduSR1vWPjLJAAjIJVm8UnZqvh57x5m5VD6QrhfhukGv1t9uALoL/K4Pqil
AiN0F0vpYAOLn1JvC9mSggdNIcGpWLXqZ74/tX9l1K0FWaHdno4FwNi6IjxteIvHBHwkZwx+prwv
tdOegMBBMCI80oC2LiEgRFCt92bX/LmLvyjrW4MPdqdztRYh8n5tRp1R2bm8f4bZlGFOyB7yhOij
lve7vajkbNZ0od9PjweLbhMKnn7oxif1Q3EgUSg2EzOf3w2bsQzZXQ5NEME34nvHb4J46/cVb3bN
Yf5ph2q8EyTkNhaVZZL+ORy9SdkZlPdUhco0bA+tbl0r7P/7owNXzvalzdjaKUzjzzfv3ntNOuDV
opD4TgVlD7GKs1TwFllRWqDf0Po0/pKsllArurulKOOxd8EfhKaBp6JAx+1fQkw5qUnpY5fMKlCf
PQuGN+ugoS/00FOVMs5MBB2hJ2NkfI9G2ONmR6qra7/PwOwnRe1iEwfgbL/R9p9iMHnUt6is78aE
xmggb4CspS7jvBuFakhT105qAAc6annsE6Q765slmo8OB7bp34AVbY17GMt6HPUA9PuHj+kyqqfd
gB9Tm38bjKVesZdAsAi5JG0g2r4cmaKY6UuMPfov3J+XXCzlEpmneXJO2kIfE1rnogrLFhOxEMCs
N/ql9Z7OXEHybd+u/HVz0FYguromleomdFpxJtLy6WrKq6O1Bn3pFu2sI/NUYB0Yapo7b2Wr6ByH
Ahi6Fxa842VA00zBXv53ro3PHbzt87NnMH2avMVPievwENphJIUMU8TQ39vmQt51Q2G0A5IM3czF
GQ4pCm9fz49cqqJGttw10+dqv1uqq6qG+qqRR4w8B4jeW3c+cIzJ63IGRf/EVwJu+zFPC/o8UKHx
tbiK5mQeN2NdbTP/tlpXfniGLhi4kdl1hIkEz0yDBlkhTQoM5FXphCYccvWpZ+eiGqhb73zFPLKh
7SC0Pkwq0wzv5mj7fkbkzNPC5fwYaOyuGXmSuV/sZm8r4or8U8Tzr3/L6bFEGxJAAWpTDDJDWiZ+
hFKpVgweQDUE89DDAM1Ib+vy0TrKZMZvN4wW2EUcBRrhWDzniJ8ysMVOWEIuvT1kgmOnmR6dyBxB
Qt9tLJmBKuSoAkO3ayEY/n38GhDJ+8BiwFUJ8Xa2PYMUflxOM09zqmuXtP1wyA40DtD95Z5gg2+z
FBhbwPGu8POH9Bb16aJ2vgxaeE+Spc1/nPECvDAbQPn9wyEA3Mf9ubJN0nlSRyEoeT3s0cHYrf4o
xsMmOf0FvSS4iRxS4jWmEuWPJSaaxh9powfNzQUkzjQz2nk0qu9xB8n2mdAjPRuRsWOGcQlN3R/7
3xDLcME3bTgGZHMQ4QJNG4XzeCUpjWPrqr2DERzhGowzdfKGxo8BTKiCeY7Fm2ADKAjD9XzfkW1L
3RSOfuQMnz/pqbFN+U2Fjm63kQCphhhGKrgVzMIwHX6RTAFwKImJeZLdL0bs77su1hBKPhq9nw3x
K8eDOOLDiR/BnLw1b1kb8zSa3B/h8DKrSIM/8Ehxyl9m012an1UOO3uoyMOIIZrsrD5J45PhJASB
CNKlYXd7evzHxewiWPIwDbYfNuVR1KZKoKg/EL6/wWofwztJJYoUCrfN8rbug+/Kph+2/0h4rT4G
ncNwlHBSCcLokvfqeSp8htnv1RCq7Xnl46lUgps0Dpf45PyxWXNUyZHR8Zs/dKN2bk+++A9s5/3B
uDEfKXvcWZhUb52yJ0mt2Cwzru5l28r2+pYdusEoqdWNZYisnRLeXdZvVQpU3Y3NnLQoiDgxEguN
2wXKzEDjq3TASJUtmlIKMeNn+gcbL0r1god9lcJI6PjMsYRDVg8lU4EOnxWFPzhp5RPCVA1pOsow
vMlbdK7ZW6KpnDYD7MlPwgZS4xn0sKQEzCIzHeBx9ItuMKmH7otcWI9XHhw4O6rhvu+wsCsppdOl
VnXS0lGkHmypeXouSqKwbtZPiNDnhFpHog1mMkMChp8Tb5RHC8H/zT1BU8HaqeXUDAFfPVnF08Sg
39Gme7vg1ydZlNQu+OF5f1uHfcosAADTAQPS1GLE+8ZGF7vkJDkRRGeVFAa7ZhgjMPO8CHRAsanE
M+tp1dMt7rpcgiFEPw5mkocPjcOXYV6Bijz47Dk3hpLud6WtWtMWv5+08uWkPxBktXPKhAXZMeuq
Dh6xEZpuDPxLrwBZ0DLAyrYNRBILFtnM2dWWpGYRi0QQ8yfLEDHG6o0O7BNOX7/6Pz5DgMhJVQ5h
Q7+JJt8cuNjVHFhS0h2uBwWMh3MC6afLwANyMlig8PKeMuo+bXrg4W0hmNbEHEVUsIISa/v1vPPw
eH10oJW3nWnfYbiXMm/ep/YsKrdiopEPWCuorZxjJl9ds6nHgSbnI+NTWidOBxZEK0Cfy6NDwRsJ
+ZoHH7fZOrwE/mRt4jwTbrdWz8zQchH4ilZXVDll1Man2HJHDleRIA0jWMW2LQyavoAohewGl0Nl
hy1v8ZqXfZtiErLykM9zk5tbaEfS3luvaCPnMI1mFUju/udbXTj6IARDfT7GgGcsF2j28xAdO0yX
n9EQgBoOXdIakqAoc2/vZdHho1g6MSffePjc2LeN7HfUTNzgfcFUvaCypd4ndm/mkZIrg9tnZTEj
l6AAxDgqtzOAOXr1S/fsWFQtTJNh3noy3jWDXsRnibC5/bZlwTW4mnteExejJVEa3Lk113XXvF3E
YfgH5qVcDvknjSYwSW2ho4MdZ6JzVjWm8JR/ZQrKTzBe0noKTJX1BXeupaD1yihyx71QkCdrGr10
EmRHVAZSVVMyixIZrjVl2c3nPVRkIBqbkTLM5IpWmevS6qZm2p6wqaJPh+fTyWrGdC/b6Mok117z
q3vOGvXB/Bs4Pic2ojgeeO7xYvYfCDubkyO7Mq2a/34ybPGY3MW4FJWLFwoPOXvcU6W0XviWPLBF
mcb1bjmdS8tbDcr3NPjYnJOHBE6dAqfnHQKOlXDKhVbybBTYXTC91tWH9kHwZ1X95qVA8X9Nd9Vi
RB4So0nVTrDYsLrzVpCvUapfKr5ZoFCzSb4rTem/XXv5t8CJfViWh9hl5iQUqTfeVMUXVSJYNflp
O/dR+74WReL9elUChHfRRY36J8RQqEotH+VEsmbJ2CVhyUuqmTlWO33HRr1jU4uBcIFdtCn/NliC
ZUpD/tT7cCljksFKeiUSirV+C68HnsSz037OJAU2ZossfNKOqMR3/z7vNu1Bc0TwOgnpPKpfSvg/
mPh5SLFaXS/CkTV6+apT/0QtCPxvigI3CyAOCAlQReVOmq5nYczMP5eI3WIbdO4gbBE2rNgUd9NC
SfvEBhaqWuGlL3FpFAQad7Gt6gxM4gVr5/xPnVl+NYXGP21+LrvEc/6j9yohGVtySu+Teqvek4bI
+yp9+pq1YJ0XTayxiA1C/ezERxGId9X0URnI7ftw689uf1DVsEGzq/i9lZMDZGdOa5sDXDrwZtPc
2KrAhbzElBA18tybMNtXxzelma4t4H0F2OHXt2aR3HGiqi0sCGEW9XAP4Px284amWTqprP/JfxX1
JueJ6sWmyo7Izuq+T6/bsBShrEMXkvVwREyOljigSaeJoRlgxmDdWSjtjJPtXheBIFCvFvnuS2VT
RiUWMK7g3cHq1BVI4ATJqjyRJU9qup3gfyfQ2YTACSZlJR2QISSBFG5ZHeMTpbWVgToLql7lrZ/V
BtnqZwW008fVZYGJEIm6o/+NHGafy2wNuyvudFOUO4FEWgOkTgvK44dyUfsdObbD4fvKL0KBIEQj
b5BpuvEYoF7cOJL0XZ0H+Rg5PrM0SEX4wBijHe9ScuqavjWQSTRtSBhfEBvG31N+jcEOSJVB/HaU
QjxbNzj8tK52/OS892iuOJjVekr+rqvnrjmYJ7uE8H7UYDiHdh4reFxhutRaDXog7MD912GBbN7C
HbjZaMiTfZVFv7FFrXJScFlarh6DgRNfYoAWTJ19vAxq27lbuumFnOY2DWL5qjd+rm7SFHS6y3uM
mlbPGatPuHv9aCn/iDBgwRjsdIU5KzwupnRwgI6MGS2aqoZ/pLHlIOFLKOy8ldcrBZUdjVYcrJmr
V4CWND8LNrdgVgI9TIm5IQl+mpkFJ9kP/xR192CZHjbxmvDYLWnobnTIgcJAlx1BbHstsRhASO8t
k4FzfLJOsHzLLbcWVHAwgmdUlkeoxnGEmdvokWTV1IaQuV3XjCSo4am0rB8MqULTEkGnMqnCEN85
NUXCWUsJVr1NO0k/gEnckxhm5LTTsLAUu369W8Xe9xz1RKQ6Sp73SNIva2A4+eC1Y3dp3GZfsfEn
ua24zQmrt5OulKgPWNa/1Mt6Qy2dZp/ABlozf3ZMV4ClN3ZZXXChnqgMbnl2OYBTBrNEYr8jsYZg
rSJGdyKk0mhlWcgZmA/iYHZtF6Dkz8e0Uu6GDNXR+ZUXr618BCCkevXefPl7ArIQO0Synq17nVFg
E15B38ocuSR8OqKjb/BNKJdEaZgl7L2D56dRFhFRug1TKZFea510mW+4+3KAvroZ2UcZWHiPo2He
VCxd7zIA7Pi4kN2EpQ7ZCKKpch9xBzUt4z/Y9fyK1qY5C2IWxPhYQVuuxA/Km01RszIaExlO7465
ptzYTEouSx1hQ3Sgtv2UG8IbfBnFnEY+fXSOcdFLEy8nrhiwLIagr1OCTxXWPllKazXQ6Ry9amch
kw6xcpSizsDQuAQM5iEX3EOn9mFRNfTthHSQUizdWEf5gI4qMxscny+FXdWJ5aw5hW2vVtfUdvW2
TyO+ijuG+TZc0KLYdXJLIuG3sZQWpVwJGEWaWPElbsf9isI/Ljyq8o6J8B56ERF1nSY7jJd8xgV3
ZU84efdJDkWvrFz+IYv22vkPxCH4GIwHJEmbChRoeMc5fnrFVQGKZ0GaPvrK2HsBeMqo6KAnOiB6
/0hgF2fMtQlnj//G8QZ9VJrRNbMErP/bhuPdtSdFchYZpRKPryQ/9JcqVPKZpA9343o+XHiFgQkU
s+bhusytBHcazeTHUWCNO5vknLNYazhS8ZWLDEPDkuyNqfx54uslUd7xykfXNPxPRkdPpR1dHAle
Z6dyX/odXainIfO9I4dsvxs6RmMIGeZdYn/FcV6jda58AMS4GOYl1jGIi1ve1Aj7ITqI7iuTWlGu
sOcjQNCylC9Rc5gYmdbR0D5oC+oXDOayQlKtgmzp6tpXZkk2ibgN2zcxBelPy6mY+kQIOZUhbtbS
ZVuo4+RXqDJWd/wE3i0vyku4ORF4EtTU4TLT4OqdpA1VGcCURPR0tI2yrFm65G2WnAesZkz+H1+p
pMA99AkX7k2oomOBgbAidW+iHd55d1EpWCw37JbGYjvKsmwvBstK2lQoeb5KWuS1huJHy4TozdAh
bj6CazXjKPvfQeBegCPxlArJI2Nqeh1yVFxfXFjxrZnhlfKaUuCWnV80BpVrJ83PWhtH9qtZz9Yi
EAqa9rxsk/e5DuRGPeFpZ44W8NL33claGORdpci5MKaptm10dZhVKWa8Tr9irwdlay5utCIJ0n38
aqnkiTtJ7Ko1dexo4BF2umsS6QPzCDt4s7MDMDP0UyGyLnBfEXn5CvBUWS2iOTjK9KPAG0TCg20r
0VBxxqoxFh4co9Dga6aq0NQlT0dFFyDvIU58JovsHchliu3MuFCKObv0S+bEvUjSUKVTdBVs5S/E
oQDmjrrCkq3eFBz9R/2LA2vLLpNj5lRNAiqQSSsNTEYlutXXaZWxyanLXGHPphXQ9qk3MevuZ2MV
AFAf7lngeWScW3pWjfTkuUBUpaAE0tnxfj5/3VtvvhjGwufaibtAfxAPPQWutC8vnFmtAx64lNP5
FrE+QnCGlaKnHCAIxmdfFY6L7RN1RZ7WY6AgxlsukRN9iiuE2ksB+m2ykvJPlSQ4gT7vZ+Vd01WH
RvSe5EXW1ii88455HrDZ40YZpOCQtYFdU/tkXJenV/x3sQ9I80tLa+2eyIQmJ0EBYTQsfSmqjud3
iRHDohw1arNz6qBlh4R0ChrkNBSaGANGExVsDByVel+aVStucON7ylIqDq1kM2VVRlyKKEkGFzHl
s+DUh5gKkiTojLblU6YQ9+qQ314/eZ3Knfny4Km96RXgYet9DryDCT9Dx20rslWbaWm7O/REshEA
ioLvQXP/GdEgR24JR8e48evNtBhAd5S1yfi6YrHCQAuOdt3uDlIFbA+dD2Sm7JsNYC2hsou2Z90k
ZoAnBtajf+9JDKg2wWqROED0MttePf9ybYDwIuFbgqTg9y12bovw4xvT/awLdN/HRdv9i9kOxvwh
ei8h/SaIFdRWzXeKVb6HjOudK7DpUhmgtNzzAGP0boXJatW2RjkhMyw+k1in1W02n0rKutH9S6/d
l9wg/mMbs6YKIja9XrCKyfTrLrC/5B//1b8Sx4tSjErSdrv5aSaHE4KdtymcVG7WWo95uVrd2mAi
77PjHLrHPjA0cEFPQhIXUsiIowx15tL4IxJLsJ97dH0LD9IAc7ibZvhIp4Nfh+1aCkktpWdXLb5O
iPsYqWFg528mLSb3yzWdojGvvlXdsvyzJLECLI4C0ZmvfFztOs6diyv5acYyZFuondVPxWhTqePH
Zbrn6G+Gg033lKkQjelJoZ8bbvyTqmL92KZmSUqpGUe2KSgBbmo20MEbeteEjoqhbHd8Emlxf+hK
wvPOcdVYYPrNC3wu1RRXzLlOz1AlyAqU+vPYaqCrIyYt/+Gl6q3uScL4ll1VAtafXuXsRbYNuZMf
8Qg6eObDBDGVkGKiGd+xVzwRiaSZhT57c+Yq2GYmtpvzzg4KTyBieBaJ4cBBGEEA0C+gltCX1sHy
ekzcSJg03HvLPFYsGzT53CSaE2mZhf53YaeBQNeQsbatsaDqoPwAqyzW4f+6U0qpgtBcd8aX7PgH
jt4BDYkhetecbbEd94zTwjJx2yeXXCrCsHNJFo7YmSYBLmwFG+u/jL9NuthYnN+Dm/KcwcGA6xSa
YCWm8eLGU+TDO4UBe9QoGhieUGL/plc4rlwc/0lgwargfnvVk35RM61038j/ISJRz2HEi77XFxwI
2csorsRRzsPzEnVhaPWyILKLEDvu2TvHTUgWhmd39GPuxiPRmCABPAeoVeKpcnnDM7iJZeV+A3JW
k34PYFUTxqpmcLk98f4NRl9G9iC5we5JQOioaoMhZD9mJ7ZOVZ59o9s4VSoCjjJI0iyGwIuy/QR8
s5FtQm749hE60H+m679pnACfFA7KeR8wjh0dIdO1pNDr0y5w0KT4qvbY2lqb5my2fC80a3rTdNUR
GTcBfHnwFWHv0sAQ06w2LQxESKHZ3MKNwYCtiLh98yqYvnbvEgvfezs1i+FtrIwukKYRl0KQRIS/
eLs/uyY05HySoBgbboS5gCjS1c7xlwD7VdDSoXI38Q9ePaHi210DegnpKKI+kopoIS8t5N2wXaO4
IO8bQkdyqlEgdXuyTQclI61DGAHqZlY5XBilu+GjfkhU5xzrIQBow3eLzKsld9pTnLyJaV6YGi43
k8+ECoPg7Wu6IWiM3wLlXxB5JnCGOnXc4H9SwXd0SwSrroT4ngh8Cuvk4AQFkTCkW7YwNQ/5gbcc
gy0RuEkv8HybR+n7/RVKT9PcLyE54aDfJ7c7tR0E4uWSw5KJUq39Vyj6YCTp6+95bOu8Drjq5HBQ
B7P+ou5nT+p6/YjRiBWNCiyMXkUiDiskSkAwos6nXN9r85TxmxLWs/C2C7sXALtUSiPbGk1GZPJf
739TgOU5KlDCYwrTdRPny9hCRf7Yg55ldqC4CIUUM0gzT18/93r00SGJyiOJTL25YGvNsrAaunHA
uVLlSy0h1WEsVG0c6jKrkWZcAHmSwoUtf2XwrhFFl1L4g/InVML4kLIkP3r90llOzwmPUQZLVoDT
IcGu1SGY5+g6YbhktSq4N+dhqVvuAbHnprSdiKKitLQ69BX3bofB86+hEGOUL9/86ifTKLgBpzIF
JPmhDfsvyT1+fJ1FJtTPlB9mPqSjDkcBcFvdei8vAcvhP7jzp1QQAV8HDElvPq+XLhZdcYdgcZM+
wOUiGppuS7yU6bEP8GGAAZ/CvRBXCUksa6Oms1PEdwiDaDF85uFIiLtjWYo/PdsMIOgzzXiHpSHM
LRd8yPsoRa4o/+6DSeN66LajNsE6FupPD5yT6RbfZF15OM+xpU2c1ES3ABTftTNAe+30xb/1nEQQ
CROeEvwkjZFmXIlKM9eogW7DcsoizEnfJSqdexBdUYDEYTn2Fl2WlHTF4AlMfqsqsgQyrnEWLvfl
L6vLBabcNQo+Si66vWmmc2X1UTSMBoEKLfW5cS8j9vomd0yBlIuAQR+ObMBwcI5EoKBz87D6FTWD
hVbOk6x8VysBtwl/NVLH1zQltSXyOS7HC43V02f1s5WIdur/HQeOobLcQQo7hxeO7yzvjf3R1FIk
5Q8bBwiLMFVK5/1myjBK6zRbl7+SLMTtKsTloItlkhUVjWHLFfXcZ4NXur+y3Mv9r3KgRUZJDKAo
tjEHviFUYBaXJ9yIQfpZhTXE58vQgOltGs9leXWjyf/L29yNwIfvm9+UuAggscnzM+rOAjje4b41
iWZUA1R6IRMhxu8qIJuvjQTzTUnIcc8GSaswY/zV1OPwY458fYh2bf6KrOnRKTiEZ9yeDbYYkc0L
yqoMpYZNUSsqKlzd8dcKdf0F/jpJm0K0nXC1CsaXHhHovBhr6UnX/T8om8ecw2SEyCnI0zKNTgU0
iQ2Po5fi5Zip78DIG1BrYGvJ8A8DnaeZPr8wCkGrOlg3JB3+PQUZ2rVG+nroG/oCIRjI2QV7YE86
GcBvsz/eVvaOIGrNYAQMn8F99d/0Oa9wRaz/EThEYftxMGuB0A2kGxW4IKFCPLYTGzkEQYp+nrko
hvndUZHVlAaxSd8rJ1inJd2mQPgcMfmqHmDyHaIOfVu2rJcbnc5yqZnOEEFeQ82cbWw8JQHl9qFg
pYX40qVqbBDtr+ZulVtMFaTf0dYDScZ5FGXMvQmfv6ABmOkrfCbiHvdi7fvOonfgKRtBewpD3mWW
0xav1Zco2I2QRxtGmg3XIwxj+NRJL60yFV4Gn11c7D5Qmt4skKRaQO3Q8pekPPhNyhYL79ThbpX0
+lHf2Y7gq0qZu1W6DMMI8oylaHr4Af0UDofvY/OFie3xMOvqWGzGB5GNQmGQFmC+w4WukKnofDiv
dFPe6UChwHFqy0Ce/gyvl1bKbp2KGe9UDn66dZf9enbTqFkuXOf+wsY5ezdrTQnNXuLEh7i67y9M
vrcTX3Mipt2jHqtgmtE3mEUTWarArEIhkqEDaYVvEtoY1srARTH3+1Hr/Z9ETeEyy/i4M1l1k1BE
tMpBIxkNm0kEs1FIgdfDxFK+/Gk9gjkq2OWbwWNG5FopchxusdjYJc4GSdTdXaA5pw9tiyhE9aQr
unD9UMxuISLTblFIXQFP+je56JzPXCtr4LfW7q31zP0NbYf/6+owFTRR6IKauo10milqav5tZkRQ
HPRQEArKtmKY1gfizrbEUH+UmsXAnkG4kTFJq4AUR2A9ZoaxeYjDJOyYD6oE/qxgJnDz7tTGCTlo
0Fl/+8cV6FLiClltj1/vFcjVv/FQl1sa8SN4XBYoEF7A1SOZ/gXJ6qufSDWV73kl36LNVHkHLyxr
o1DfunDPMKTaSTVlIfhd8GSJeo650P5hbPHp71P5a3CaOIGW4G27cm4erBqofbwsRyqKxJY2lJJT
3sNR0/DLWlYZLr1oc/cp71Tx9TMkUshl3LiVVwWwm/gYsggdUsBJja75jsDt0oaS6Mt4HZth9OiW
vl0y429I3h71+LwKr0Sr7bQlAWzHMmBDdQVPcB1wuECiVKn7akBU4N+QsQiEEH069Fr40qjlcnSy
SHZfbzoMbgwA2lAen622+TlKqYoOkzx+3fJnL8k43XvXsyExJ+QAhsVd+0ZRzBqpung/wRk+MbwB
EunUrefVxWbT7flrPe+XMe9LOo1MIwpC5bmzQoEFMx18uQBXLezifLZ73p8hi7Iz/e9toeOdxk8k
1Y3b+n0AioxkDyPZ1z5fYQO2vEEadZtsVzBtXMajOC/LvFHBcR8Hx0ksdrJaVRdmkKDrEVshC82C
hzrAFU+XSSnqbu7tEh5WJJW5ZRmTx1eg1CfebzWyDYOUcIAAPPfkFSgSI0SeUY4Wr/leOpad44qo
b6eG33HJvMZ8OZTYmfQ2eYNZmKoiuu+ZOPLdQcVgRSPLtEqDyn3R0UUf9Y9vRkr6cqPRhl7H/eaj
GbTv3bDZuC37pTSgFZ6bkRVm7/nPlBHDM9fj8vciq3ctXBjTIKt5h0lW9Vb0w1WuXb7CTw/Oc539
fkZ8eSm7+lh8SCRHS4FWBX2g10KXMGJXvN0U/GL65agnv443dvjWzcqcswm0Ae/ZDt3yH4ehAHVQ
g53y3Kp0pviOtz8Lrxvk4fkTms/PMRBx/bqbHWTh9FdbhMp343JhzZGcEcLA8sPsEHrWuHN1/H9G
Bm/Ntsyo5RYKc9LsPpeQdVSGlBzVNpqXYt3VeC2NZ3SCj6NeIJI4nlMD+wwDQuDHVOKGKEcUIW3j
z7Gnyje+Ch59S/ixxitBU37JxVyl7GplJSv6fJw6INsqwGg9FX1hFPCNj3Vdpj34wkVXGtgRDPgJ
0eKZJdYkr4QSpdUKa4cd91WvR4HqM8lJV9yyaFnhjb7T1hGmN0PsApbyw2vhct51OVgQq827nRTB
NQXVrTYt+3TkMO+cHd/nDIEeRSRF4soHQLkBXdtBC4rBdmE99q4vhwZE6KHK4pKIgLtPorw37XrW
sHJFssPSYxfsGDPVTsRRJct5Ttk8lj1m25wZVi3a2bZdz+VdMWDqICIYqIQFJRMyqcW6PNJ9k/Pg
Rr6aUj2p9kTnGakypKevn8NNwCzsqziaRNanWle1pe0zE7aWobz2Fg7E2YBU6nLY6vWrxzDZ4g0u
Bf18imgf/Vm6NARWBikVTEWpeC8ggL/uCCyOfag3jlc5SJRV4FzLZW1gjOMQKM4evhpDIGCl5XQN
med6Ut+3nFvn351JTSg1fCDakb276yKqUjajMH3zqacladgfoomHUqnvd6pwW1jQcwwXHmdBblXP
3+SuwnRRSjxMbPZ3qsBmekS3OxfDXAoAsTqynqgPVopFbgd2fqbGBfqRu4mzBSiVFbS0HDHAk3hc
1SCbqfkj5utZaiaW+VR7ZoBQNmJGDvZM2w3FqrbR/Tm7BDTv14OM5As+EFAIkqR1fLMVcmC90xun
g5SjaS7GWwomGK9ht/naeDbK53S4g8gev6Weg9opLZwONmajswB+YavHb+fmKBHZwx1f7qmm/ln/
iukpQ9V7ZwdalKI2mmMKz5EAPHCxHDIwA+SA4Os6StPg20vhbhQOTRCKdVfuVX8oxMzLqe3Y8EwB
p08e3YyI+MomG9cbld/d2DMyLUXDLsojP/HAqvVZij+POtb1Qw9498JMz2O0ZM2d5HB1wS1TNTdc
7kQlQ8a05LSSAXdzM3XEIG51raxK/Em84YkyS4lcaS7kB/WayK8gsRr0kLwAhHQRYNHLDGAHZ0KJ
K1KQ4ec56nTEWcyFzfNE3c0l/qiAb2QBJ65dkFtpVetJzaFX2DpEpbzfVHV/XoUD8xLQs3bdsaSp
osDYgBDU47ucoKUg6ITOhm5IMRNT50oBc32GqA+fn+tsmetEaZRrfOouLVPsesK8wYtEYAuR/ZLY
yY4IlV5lEqbAVRaR/9RRoi7wPoVoeLi74pwwLU+FYg2nodavjrPG8KLdo+N7fsuy/QW+JpE/gQFD
pqNByvsxwdgHCBU60Kclfx/t0KLMuexRNunzBKh9b7m89oi1ihPlEIQoTuQEfNxZszj0uZpGZRD3
Kr9ooACKR+odbmeJi+D4ZJJkE9C3BIEQmNejFvUM/Fg6Fcf3Th/PsHEPyWRqREUmB/Eqb9LvzZgR
sZRlEX0n4Exu8XN1WwbSJycOz1DIOzLa52HiNdLboAWhur0tIHR+wm1JGaFnFLk0TArNqc6vQXf7
HC/K9MeWAVpARyqPAdJLdP4xQIfuYMyNJvYHKaQishUdl+f3ekYm2YMdoZ6ibykMoD+W7ocgOmw0
0BDIezbHhFhSvznf+QjFCRkr/hQOMgw6O51fpxkwoy6rdyUgmec+uI0v/a3dxpi9oBS+dmXlyEzy
GRqhE+6WsNXBUsaGBFvgPQOLdVQrdZvj+LNJS4p3YRfXX7YE2Gp0INZOrxb6r83ZCAwOIcnzmMt3
+DDARBan1AK2gLzvOM7Pz3wxMknuWzfjREbRkhO7bTABW4xu2KhMYgbSSJdL/fI36+ahIVlsxidx
QFDBF9s6BsCVFdADYOjM3JQJFfPHw4bmcIr40are19vJHah3mmdN4rWVMGUjHcdtg6zWXYCuZVMx
BStuY/QKLhAZQOL7oTYKJc6Z0ifJgkJzN0yu+UxlBXs+g3UTBu4bKLgnbyZzv7dJyDJT0HlxI5YI
b4/8wPr7qr2uMWQ5cyRuy7M5yZW+n1peVz4Q/Dboysr7UlxPpknJbTZq63GyE71gRSG4qOhcygg2
SGapHC7grlZuUFhJ7ChKlWm0T2SnvE/xhuy+/+vqilQd3b85WKpXef57h2/LeKpUUg3iWWC3EUFn
llJDImA5562nDpSmSQ1TmsY8nccmxJBzxWB6h/aTench938hkbJS92R1s0oPMsQgXy3CStzoeshA
PHTOzniR+cotqL11jZFIiDAxpyDgoiZ8TVXvGJsQotDIPlSF6QS2G6pzOzE1XGbSc5XHyX9F9Hmo
u8VO45J5YZie3esmakFpP8+NwunNVvIowiIQkryVrzUv6uknKhRyOOaj/8MlNeJyr/SSY+E464o8
87S1tIRa/pWNEcP/Knlfqr/gohhRimHi7jTtMkBfiEDZwQYy2CsZ5mjXSitCCfgJcI1TkU7ERR7D
VnpJKzFWqHcEGpPhU/62Eyoi36c+yNi/qYrnPJlZYBme+/i8Abo+evaJR2ScMsHHhU6ZxhDSCbWy
1yYr1nnVGIyXMUbStxo54pzBNr7I99G8Qef0UOte8YCAnydDXBHduIZvfeUvW+EB1Tz3ZQCkY5F8
B0U14+yfJQEz3PbGIwQfcZDjEetVwWMaHVeJ9DDf4M4Bx+IuDCT7cqZ7bLKuZ1dOI80Zj6+G8HUA
MtjAitGiS/IH5u3PJAKr8tcNrOxkLd2SHF5rhFugVgf54ILgebceJaCcjcLavrzKvkvZ2YfCviQt
1e/RwfSQukydmM5BVMoWaS2jUoXQL5jxE0oaK+HTHxQNHZSk74+7HwyS/ak6F4jdDBuT7fL6bsut
DQr02zAog1cFBnJn7Bb3CezjTVJ4Nbu6UKh5oqGJZu7SGlZ9nhwZngFYkHmuQPWVorJu24F88gxs
N8dsls9kwUOKA07NKCJIiAulv83fHEoafMMdUyBiAdb5at2rzP5WlvkFKvkJmPwpKIU/IlY/nuhG
dgTuvl0LJY0YOXde/Sz31ovTVxfr6L2S/PhDRaXX3wpP9nR8e9OwJ93IyhJ3MHLujjIa7oiA2JLu
90uU8ljf/aztw7zuMm1tDW+sjjTnWSDol8QvVdDTraiPwjlj7r250+4mwPl9m0tKnRne7XUB0qvr
gt8rmfh9+W6E2RW6wRrQiFacl/xCBD62eb4Rcmfyk6kdnpC1KgkO+SDkhKEYXfdhMk5Mlmk4RG42
HtoSVAl5JwYfto77UguYmDZAS+LAaKOH05Ok7SKZuJ3mHV/4wXEF+cAYnTEaZtdYguiA8b0hbi5D
MOFaBD5GEYXxveHurEJU+JxFHeIgMxK/Il8d2pryeX5DAFmCbAeKHpkU/g1+K8nL+7cykzsGKht8
qZLXGKODG/EbxeUGXY/EqT58s5GXY9a+69lageTKa1RPcf+o/HbTWFRfHu8zqYt1V52WK6ZtwH/C
KfFzENGvugAWWiPPCFWNHsZMH4cCxZ8HoXUX+wxe+ynwF3LFbgSA6lmxRW4ljPcQQYsHkp9vg6BI
plbAj2O/LuWszkZ77uRdXeWAxB0ZnCC5pVBFOr6sU7t8t+MyvwEZlC8piVP3YTAVr0pyYEIOjTNT
+cl+sit48MSGvIqC1fd8hAi6eEjbxq+JIT+qb4T9TmSQx73C5yrmGoeMx9cnIhRW4CnBpcCoAmJm
3Y9gbytbNlLB3PqoEksFtDVL1OUAFyTEVYmhlOHUMUNzhXuHto0FIq2havxZM7Q2EfyjRkuqWIMj
XOZ6qC0G41FeGgCIfhLsQ1+UnSuMKSyu2TMgTO9Y8/JzmG8zUALkgqgSb4zH+ae4QQmxOQHKasMe
VFV9slVsMpyuizcc9Vw/o4Cp2mHFUumUSYGP5xN/bcIqoEK6mF2rRRPeX1+7PXEF4v0ozt2SL5YI
e5Cb7xks3PYhdoudKK7Ie13hrW/EeSndtInstRTlpWMwqJ0Mx0N4S9arTY8BqipX7MD0/8rgSt8f
ssYZIgGIJgv33WR7k/kef7YaEYvT381eZz+jizvfbnpp7jNieNMRSjEdFcEY/XUvtiFJXXevjOb8
Lh6YNPLHlMGZHvBBy0Cf3seupqPDNCU9Om84gmmUS80vXQBm7n/wao9lVexlX0kztn1vSAq/nJhB
ig6jhEQ0w4EF8QHHWC+lznzRfxbLjQprYFmBZoAww/xV+pppu+ma9bqxV9JrZvj3ySe1s+5o4Z16
mu3n6kSNTtxOpENZzCCRhSscyejMapPwjHgTF6gKfEr1VSpoa3NLfXKG7YKUISmERuTxpxptaV46
G/8cHQOv+sNK5csjWoCdtbIYKKCwJvrIWd9SdsW33PN4YOR2hWTnPYsJUyxFmE12H5YybVDCMzrw
G4TUabCt9UtClnh9nA4RmOv/0TdxPqRH9Dn+GZGiQ4vn7Aogotgd7VorhHvSLR2pv6vJj7UHyupC
NpF+rJji3UfRYVna7GziSd+mJPOLqWbcEPZRjA1imMYOZ3mNnBGt+8UMcQo1rgdAd08g9cuDgI4H
b/OS4+qHB9EsLNG7GMvpup76so5VD8DJ8NJEOEtY5aF0XyvRdzThls2Kqu4H/JYbcAuQth430Bj+
oC/ufzzc1bGNTCPEsnFt+7GT/iI5LXs/oVU/0kqigWqsQs1mfuwZaWgibGghkbwqmswTdjFtfkj2
vmNOytkpHmE9EFPwQxtzwj9I1Wg+zsSdC876ZU8caxwWpOXTIU2AJEzK1Dzql4Mbvm/nEXYpkc31
rGdp1DPwYEWFEldXt7JSJTIVkxkqRE67Cq7nfwLUFmNgNRwyt5FArCha9/ojTvS2o6hxpONMjA6K
hNCgCuHr+3nOZgTQWyZ3KrzJ7CUHyPrVXpym5B99gRa2RbPldGsAdYKbbKcplV/mDiTKBo+5RO9w
yyKKoGnIx0zsKQQ7bV++dmmbjb8wVdNzqWw7gJhkdm5j6t+/4UKdfsH74egsPMii0orGpurFJUgT
+zqIWGiV9jIZjV6nH+YMiUK5jelMuAUcaIZ0QNNjq0pxahpY5uK1zcj7de7zMo5n3nimjqid0QlZ
/1J1nQ/gGkATJc3G4/0SlNeZ9cfPnbRJ+NDEUvA8aN3ymLuV5XMusFaylq6W0tYnSp3n2sRPjghJ
Ezn0tTedwuW/CeGU/VAHNj8lR1WHa1sH+z9B+padesf4CAsl/1lkRHV3J8WwRsPKinFioqMOIiX6
+K1nFG1jl064H1XUvzS21EdHlwQ00qrU83Pg+Wiu2OwGqZ+qUz0lWB3DpaQs5iq1gGUiz6W+2vsN
a5tg5YIiUqhrtzazuMwYongWA4ALdae9jR1R0hZDrt1V7rEXOrFLn7uftW9qLioI8yOzvqD0xmB9
15KXaWmS24KV2n/zLTpSkc66dHfls/HneNjMpzYLRJj69AsW/eViAyBKw61ryX0LZQAM5iUSf2jo
0k0571Etsqzrc0CMltAJg0aJxgOcE2gdH0F2+v0ZhqA2G6GE/Za+dk3H5edJwixy5jWXm253quLS
meKE3WzZidE+hqsGwWaXMKei2Ge3hxU8jWf3SFC4Z3KdCBIrY/maxF0KYvY+X5Zo2WbZUaSuQ7Mk
MBv+4jnzMGMCcbXzzILMscsHNAWIV1KaMGg8rSRjcxIQ45CcM84crqm1kouDqD4xYwsySgH0dNgD
h/PTwstBanTs64oTv66G6m0FIKyhmeI4wElh1Dk3JNKMbo4g6Lz9UItBdeYz7w7z7p5ayV4bcjoy
sfYhkATKzxK9sfxd7z1KjU8gk21A9kVsRuwk0vcTWmUuDdWwqwF/+e0LRYxlsrrQblW6MznPHo9b
CW927zjKreurc88OzR8vs3IRe0TIV3BsE9KQAezKzUIWv9I41LkM9ActN8iYTwXT3HZjmUn61bAc
Nxke7G36AoNMujVAPLd5f+6sfTRRYJdmPLRfnaSk3D5cAZFnLjKoq7del+BnlpQxzKSBZv5xTniB
LbWt4FHXboteCwtjmoJ/Tbb0D+TQ1876e+EqLwH73XtZwmVKSS8n3iKP0yThXjNZ/jwmFLaTGPnd
T3yKnjU7If9W70AKd2tNJIj1HYY3yQgnnDEWlI/iWYbjPqtI+fqWWrQJ9cx+GQc44xHWdbuF2/QJ
wN73b79GkonicKhEam4I4XfYeNaU2ohD+QXcNdoB4wmQeTaoURd332eoF/LZn4jEcIkRJOLlYU9Z
pFsCU7qzbID5tToKgKAPKPeZndWfs5ZrUT/SescsPLuzGZGegPOC7uXVVZoqyJRo2dfddfGhefMz
0vw2yEa/0EsiRC+zJvMZSlGajvaK8NMLEBFptz3sYf8J28E1darHod9e3Ne+0MweEuNWiI+GH3LN
LZbLcR65jnertA7gFawH6S4qDBqKgam92MoeoPh+xn+JMqXzdYRnxOC/T0aYxc+aK3MtUYsF35QW
npAzXTfFuTNsIsj4HpA1KwTVJ7B2RrtC5I5fwAPsoZDktht8tfHEp9pC/8zwuG+dcqQ8zLmrLpPi
WxoB8od4XDHHYHqOPiIH/doe4JqSMFejtncenS4sFjsbEFqr4CvxtouhMisDOi/c3356/eF2S+er
Pyeju6vgEKLmxAu8TI+SiCoPK/aBI8wwg0BNyQmj50kdGwm04oX0mTfdIrXTk/Ehk6ouIDrC7AsO
fnhjN0p5w7TO/3zejZWtLRtkAT/CqXXeq6PgEdfApqUhG7T9k+lpaeDw6PTvCukzeHc3uMNrv385
Kfqv1aSX2CKi+rUexuPh3jy02xWgB6Y047ARcW9vrOTA2Fx2jy3pA7oi9DHD01y+M5WCGcCkrzmd
WuhcJt8h6hrMMi9kXtpZYJTAUOz9cK0aaNdJ5NDt2JlZsUj/5ajS2R4ZSaYKjAtaMI7poXTL8FD9
xiJKuPaV1exCPNvDCQ+JyEJrW+EueDtqBkXLnjWe5IojV5bCMT3hL/P5dBxc1oNuuK1vofEI/ERJ
93gHJoqUwzcQf9MtGVUSA7pok+2tagMjuNnHD1BBfd38cX/vvMItfJCNvecZCZk3OXIpbEtobFEL
0uWL1m6up4/qdSp7Q7mAaq/9UN/Ap3bwkVmR1/pGl7/qYmPm+jA2qnUbeyhdizqFvRXX287OhwCW
gZldhOxdDLs3c29csCnge46NffigaTTH1icvlq919WcQRoDJMKeLyK/g42rZN1yMXbCW7Qr8OZPN
dL8koR1+CJ4gpVx5ujmkI9RBxAzcHwjDMYwmMjtkRTymhfl2g40zCD5hLJUYn5u66A52J9bvsMBi
crszC6c53tQp6dYpekE4KCyzcaXEEDsAfH7/6KJ7JH3I510zvU66sc5cQzzEpSUBchGc6NT1OydA
Peqlyu4AwX+01BuqISdMDkoMrGAJsr8ab9OAaUjF0gPVYWhe9wu1WAKxDyae/+rHaxD3sWp8D+c1
7fzO9IxHLWu3kmy8MgHkvOQteMOrB/NX+4RYgM/y8YugXJz+TehZfiJReMlteFTWekN3zVP5//ZO
+x5miT97uxUS2enFkZRIDiFxnWZgFQUb42Vz3cskqqs4AwzmKe7iG8D/tfaq2JTtxVwxiSGRgChP
zGcavcytpcssLNJ+1CdwAaB0oi+bo+EokkLIUlIkHJCHxrfsyt+v0G57IS9VO60a8fqN73RzgWxO
CsAF5rFbXPaJ6UcFkmGTXBHEeiF58Z0xR6KJghrpWbRIBIvMAkOLVdFNAN1RfZQ3B27SZh4f0a9N
alxT2TVJYuIbNYwpYeyebdcZfzRV0UD7v/Hk4zOPNHqFmj7P0Rx5dJ9FuAtVEjVgch/ReEmH/YMQ
YUrSE4I5psC/niow0n0sf2sEXmQxZDiWZkKU/c+nCePFCev0YlFKE6Yb5RzepxI+GvoIEFO6Bxwe
RqXqedh5kLzALMOE6nW+wpFGEtteKt6Af/j5sRaSgycbUowiwPlXWm2QJabPPL6L7HtrpGT8sGs1
hbWy84fJEyTQDn8S1zjw7doTunFCGdEESe5r01sME3cPrvu+auh9uEEw0k+GhchxV5Z3+MKUrA3a
/plP2mrVikEmDJ2afVOoygUZv+qLX0r3gl6m4rXEOieftMdnJlht6YAzu4iih3hoejYEEKOr06gv
Jf6yqLwTko+Bplu5Ii51KgI/z/fj0z1SBAbStCehnRDMEfbPR5cUSS4akv7VX3sUgmiOpsqAcoAs
dyqD/gUgNaeadYSmOEBsEPmUi0TfhININJ5dG+aZGDF2DJToxr3MDaLJYfmQ0D2cMtuf975LQGNr
30pooUVxCl2AhSoeLdUMD69rI5HFkd1BiWTykQCt9DITuh0lAGRNGCZLoHjjiaVHDoziw8YnRhy2
ZxgnNlibMqM9kcJGE1C0kHmOes0tDrGwxNBHH+3OLX1LP0eMF+w2ungRc5hTjKEtqTVdKjFNXkYh
yhQMPcRXm70b3Uh2rA9sjy/qJEa/DeZd9pzVYGv3cSe+kYlL1IaQq/dyzIVJU0/wyk5evcBBeZ67
XrKDlFrZHiGAP0WV4DSK7RtrfxL3jqaiboIX569cN14Cv3ACFWo2kCnvdFv1J2rZsAKg1PSJNxTb
vE+Qdf6xSiZ/CVbKoBwPKwMIynPd2XI6nzRNB1BrOuQ+MhzJ0FUyGe0JckmGzlciz6FcFst9zHgX
hnsNJjqPqjK2VuseTPRYu5WGmhA6aSU1XTc/yHnDWELYyB1HmETSwEvHYNsUwWQdB5hOlCQc3zgJ
R3uDQUZysK2IdLUvF6BZwEHt/mF47WxPi4vlaA/uNe9uM0lHbSg8vsxbVA6XeSrR1PgqACrbc0oL
1VmYMteTvLXBnrg1AfbqTZ7ChW2S1DRzh2gLwXabPwAzktQwoqg9G6iOXV2+4kkwgH5ohwYads50
qBRj/At38zCKZfdAOfwpAAUmJLZy2MJ1CrkpMulGc9XbkOXO5yVCdO99xgTpJLwZDmWPpiVE70fT
msAX6g+P7OknP4ARRYTENaJzfHmhyFbbTeCHLu57DssYU84TIwh4/0IQX0M9otQUc7kdmmTe0Pih
efYLmyiSlH/r98GEzzbqBM888KgcbvwHDvGgI+vZyqQX1EFywCE4+IdvJQlFvN9RszDhpo+SWoS+
RRqAmPit/rjwzoF7y/A6TrWEQ6uSqor3zAtC/kaps2TXmpKCHSBcsaR0lIeNVMpXwMIGe7D4lFEj
X3Eo/G4CIoS6HqId3UV28qwkEJIYDip++Dpa432iahIJvq1ucifL9s4EFm+ke5iONNpiOuZI1RsV
kbwDqE4eyYVtL/vpSjsI9g/KkMAY/lZnc+kqK2YK1t8F78ehajzDoLAOSdxcWoFnPcfuXH8sbLC+
tHclgsjn9atE9EmpNjbiuUlBTDAOtA4GzSYxE7GYByTPZNyxZggZ0VxxuPPIOZ0EYRhqnZ3Cj+SJ
mCADBVVANQQcvjxEGYtjQWvTfczFYeyXxuGdgpHzIZJvXgfKXvsnDtnnTJGdRd/Xjr5lXIpNd2oO
3rtAwtb+ZEOqcxaqcmyZFcV3zt36yfV4z0V1xoWwjbVaqFXN+Q23kscX+fhMuw7/buxUBYakBpYe
MtlumXBrvcIKu9Iu8ALlWk7eKHyXTV+lFXGkajysvLHe4B/n760CGEJzThNPHod8Sum/c2anjLhY
PyPausPRX5ukhtmw48B6ox625kT3bO2TQo+Tm29Ip4Kejad/Od93fe9yOhA/QUIiitL0Q8Y2IHMY
1UW/bZYP/0BaTk0KUczIMPYpnKPhUN8B056u4DJs5ZGoDREcpJitnGbwNK9MjZ9y7CkttmGKcodt
B/dJH7zxMVfZhnDNhXwKwoVXWqoD+iXNkSYsggV20CunKGvv1kD0bueXvtareBjKSLJ4vqTYOAFU
SqyjNf5L6coVeHovrmZNAEtYLHhCZeIgiMBH6SHs5Z7bTjGYuQIFj2HLdL68crJ2zobJBY+0VShZ
gw6+8EsX8TYe15/N3Go4q8cn3JlMZEcrhNBbX1zKr/gAgj3xPSQaQUKSSwxuF6tC4nURIazjxuqg
G44ZvvpWpTaz76iw2wA3SJBLLYvfXn/PHFgBX830w1ubn1WgCup9S8L8w7jDEdnv8QANzZ710yNI
0Ekud0qC/PPHPDxPmHd8wHVOo475Ak75loibmzaoZvDly6wipVDPOOvhbiNhc5MdDrHENZPEmptv
5+ltI+C104rRHvD+2CuNgoKSoVSkEIFqx29CFN0OKxCcE3iVM5chmp4XxhVZdoss+z3C6Hq4v9WH
SmiuXlCZmzyuyiCUMSQyrYYYx8rkum/qoXSMY+0zrBo55hdW0MmNczgTvTDA2V9IHLcBJkoKj8lg
P0M9t6DHM/7+ixp05Yd6+2KqLHFQ7gzzEnL2gYS1EMEC/SiMgRwmRh+B64E6BGMYsxmVvx8uqMRD
/eQjP6toyKB8paAAbfPHDtDIWIGXIRZTUE2APR2schmYtc40WeOhgxfo8h1cmQI1+tpD17YMVx9g
lvlTu1yCJEXvxSIjVxNRxgrGoHEauNQw9Yb31Gbj2oRwZxS1cNFqhTNElilTiMw+CaxJr3Q2pXiS
ohY8JH+6+bLxe2+XFU7ildZrwRI9tRI3VtNKHwXE0UcyYKQ3hl82VUB3ZPsWu4c6005jfnCg5uwx
BtiLWu37rxlhvVz/WAUccISxIoXQuoEQlseivi9VHE4aJpfr/iZP539b9sFlGSD21bCggWQvPtGF
i3TQ6k9IG7w/XnEjlf7g9KZ5FL0eE6MrKm5rMoVWIvWTN7ycNQ6PP7kZTskQNe9NuEcvztjCz7av
R8BEsfV19SSFt3dU9hZTKIYx8h1x/POEWojTWOTWWWphssxKkY7QTXF1kN4DjK8ACAEnd1/ki+cM
It+rES10Ptjbo6PnK/86PCw0Dep3dwft0rutVnV59Jl7n/9fAsyEdDBfelHWS1G/DFoFLb64Nhhy
63ilzcx671Tojn6jkKFkRIGDzGnEr+Yg9pkrzmw2HHbxM46632vZ3wVpvShmCXaq7OxRh9mizNEa
vp9Hqa68KryEcvE/+Sh6BhZQ1ydYpRz+GjxXc9Oh55Dldr2xqfvVa5HbimTJi6QAAuI38aggrWqt
YNLZGID4cIAXMfRtVyCvLBHVQ6Rv4bO60WrX/lk3Qe60UXmn2xJrF9Uon5A7TVl2ioGVrce74MYc
t1++7APXv+KC1Pn+9t+u4pg6uXzAb5se0eDRUgouwoKyz8KR2VduhX0t2UsoDZwUaAQKpI0qH+sQ
99dDRQk4WvZf/Dg0L01qZspK41iUWPwxwwwoAjXXTc0+XV3htTSi0oS3J2Qpg7A/TprsJQHJiDnR
L3on/q8+ovyRPnx1ZISthLx+yE2VQVO4AUpuzi6cHNAJlpS0KOW3Ss+BkXy9ZFpJmWOldFaASTQt
sXfFBejZ8sCXBKAAoLEN6RUCIlYSOmDntEneRCDT014tj8F6UFu1yufN+VSvOrur50TEANh/lvTS
kGV8fXLdkKYDiPkD1+f3PY2+xOgm6yhkPWC9ioNmy3qiqTdIOfV54Ybfcfd6rZIwAIv+2N1P2epl
TjURQwNSswD+BHkjBlZkG9O4Ae//+n2pJlQTxkYEJ5pq2fxIqk2F9XNkG0Dd9B3ELIpV+ekrai6g
ULMxHIoiUYyGKaupQrV1aqvCOAPCb6FeJokOM1OZ+zWVm6PQ4RcwDzKzEqIzEDW4QNkAhRPZoW2T
vXtMi/XIaZux5CN6DOCRyYxgLzS7/wsMcYELGQmpET7e1s/N+LD+TVd6qeu3bON6p1qSCd4wyo+K
6hv3K9QBxfBzNTyn3LZaoo1eECPIrRCoORT3DqBbS1FiYCnztxwnyl8TF6KGf414ssAqxDaZe4Mg
4wB57oigevRVY4ThLxPHcnAeMGE/gQ92hsx87wHEEaUEkX7FI8mT5T9cfMbtD2CutWQ+zESnZ7ZR
zwn3kAKBh5Ygpi+SlPt4nekxrHevCpcYlQCfGCY0asq3aDFPDD8t1psm+aCunOruLSXzYM0Ajmka
LrxjlourQRw0WCzoy/eQ8UZx2fvNLwUSDAoh9BGoKdedYxDi7pAQ9PGPX+Lem2YgPXvZfDEp3+GY
WBtKhj4LQLFRUMxW1/djSD7uZdn4QWW2NjnpsPP28NASCjf2b+wsAG5wAvug5Kz9s1OR8cLU9qS8
NFiH0Px9feXynylgRxwALYc4FPAcJVzNVsDBhr7K2eW+S10ViJ4eM0u2BsFLgAP81nnv3FbkXIyi
A58eVduSSn/Oalbg6Zt+zPwjYJIVbPQ8BHZja9hwWnUx5BDV90Ps82vLjqtqGzTN+A497n0xvRHI
/QfIGURq/SPteARw/G48VgtbXIDh+RMm5v2Q3JRAM4O6jbr8XF14VCn+OrnhAMUi25I6krv8eZUk
07UJKH4BY8rLVQBjAFRoO1Aig8zlnJXLqU8gCet9OI5idMjVlC5BheVR+zoMTeokNz4Zs8XZtBxF
OPi2C1I9SSC6MYwPCL/j7LGURRZMrwTRXrL20u42tbs6YZa2UAOYDgV0R+sWxLcw2xCXVl9O/TNp
znDLJHY9O6NWDCcaWv58/dwGiMWdlq3/WpKtk+Tot4d01PoRJ3TJRJ6Wy8kdMtXuJlEz0yiXktpJ
04xWpq2stylLDC1sXJratwHzjz+y3GK47tAoVX1yPcbgxiHYp0RvtU0xiEVhgi+FKacO1u5KbU1Q
/9CSInt5heIQHokj2NuJAS4+vN0bMkgcEITLs7+UZho6N8fSh4n4ThwUCvRMvcmQ17/XskOPcQu8
lsJdtL4eivvOBkN9il9N1AtY0L6AfP/pxawvgOxgBxIpaztRj/yFdmzZNmnl4uQcka7Jv4t659i8
mSdrWGmOt9SoxJisI7zOcjCigyjJKIpaGEDMSo5qVY7cLvBW/ANi98N0HC9kFBKo5snVIjvvcXRL
T682kkTvV3i9cArEdKvJOqOJ6XFLfK2EPA9ilTDbM9eRErNn5nxblnIBqp4ImAbSJQcvsToyvqD6
U4SPdc/kKr89xiDoy+rTiZFZZHFsCK/7LcFcJN9dEr55sUSGx/lG1jAOSJASfAi9V68U7pN3TqL3
0+e8s5HijlEZye+EFpvs4uaX2eJ7jACyr/Ai5FIhGZluKyYi8eDCk3WPSTb0dK0phB2AnRo6Apq4
rUdTox6BMoQlV20SBkJLo1LJkHJQue6ggymohnAu30sparvm1p6AECSZhRXG06WFtt5JNxLVsUqQ
y3K/zBATPNLh6FIDgMf4SvDp8b5l/6A3XEDQDJRJe7G7r4h5U919+YZEU9KmgjGJGP0iaQLEje3t
2HyT5gWvbleWaUu/iTVAThUh7jV9OqKKiHCI74SpLouaKCRBpbXCvkL4dQUeMR4pSjgvVz8KWr2P
79yWUzdcETYRiByHjixQfgyNruP6aHDRoqi+ZtFEUv+iLH9iyO0VpEXw4fFWaik6UO25tDXmRgNQ
aQ1vWNvLObyviw/B3NlInqm+sCFHCb5A72ti/fRTZ14NyhFFmAJaf/TwNwsvM2NnqSqBcZgzOTC6
8NAyksHhfKtc7NPbXKBlp+Vg9myupgjKaMXlhlSfcC8+ao5NbMfDoYn99a7Z29uJo113UtrxLgN+
BoLaZReTW5LS1/LpgQRh0k+mvscCE0xW87XamgfziPzuvQM+2tN51fLT3OpcpjGd/gV/uWv5qssj
kqPNCrk6aIPj28LaeYi0GzfpLjepHROLLXkBJeISIyfgSxQ1p5L1b8JbW1K9HMBwD5VOfdmr3ydE
i1Dre+Ankn5FCs3PRprUeE5K9MneRTPuGqaFqdBdbZcmTn10JFW0lq3lr03y57nCiiFYuNHQZZaz
pjK2/Ul2IVpIuMSLfJLXc4MXGmUhUY6NpszAskgzmd00X+vl010I0p49uE2theYKHFLsUq3wh+Mi
6F/uShgHvpg+33qwZAwRib1adNKRbhIKaz8RGD0t6K4F/28iL3fvhqe2qpIEfAP4kdJcum5gQfC5
ZMtfHS2BgpsFLi0fz0T66nEtlP6catfoIyz6xHb3+wMqltxx9nW+T9TUavmtFCuNNcUbmZEsa7fQ
HqFIa+ERPypEa8GXraocnDf3pOPyC69bi3g5QoAXafItW3/hZqexJwvxfMd5lGcmH5KrIaZ1aEwl
IiDKttfL/AWLtlXdVpfHMecUG+6PkUW8HWQTofxHYKTxaKOGh5BnLogiq6vGlxaWIdJymXlZC/MX
FapW9NQzTLA58rxE54x3ynGS+Tu9D4jK7NQqd0Rvz/NLEtcDY9B57RYzzMeo+lQ2ywoXnS3nJ2J3
Fz/1yMtcnplKR2t9fjh9o41k/gzOlz+CdQwaL/wRCDo444bkKS+PQwcGRamKVlTRyD716OHc+Wrx
YfcDaPhTR5UgPjKPVofCRwPzQ3wrPAMeWgiO1fbmRuROOPGjYpNwnbe3vwbyOorI/HIz8AlKL/pI
9hHhlL62tECStb8SAW9opcrZH7Dg83IEc4wwnIuyq6LFDKlBBVV0b1Dxyh4hNcOGzLYpauUauNjy
OSKDh2sUjQN8nOU6vHpoOA9C/5bQsTQcawRe55Irry1rfrC1dTQtVT6bsi1ir3sq5gxifWYCq8ug
AHTA6Ruo6BR3zMPu2gHx4aLum5qjA6oX4iLbVE14Czg5Z4pjve2g6FDRfPSAWA9skil+dZaEcWlI
9K+nlD40UCcNwxGokoxpV87kQfnJPMpfG6XuRaWYISLPj6GXXqEYUPow9eRIjz14IRPu7r53J5AP
qrtWl/lf6SWBMWGgAH9QNAPA1Ni1AvqTfjJEELkSDGNZP8HBdBQOFVpG3oQ9XOME2Ljhy5ycXYgw
IN7+1sbJsCtcxLARhrKIKVFDJaGUvIgbSUcU0BkcPrMw2Wc0rBFgvURcFSPJqqrtMDh+ZsHd5da3
UhkcdEJqIJqVa3zsvMHZIGF5MqUSYlDS2OSTTxd/XMuLtVn8Mcpx5NrhwewJmuFiHELZwBr/g3Db
6SDjNpAE809D121Ylzb3AizoLmlDh+cbMq03/xkrb586EMiTXvMxJIXztPnPTarmQcN4Cp4NINAO
t9JosEBTUSZp+ni61/0AZ7ShFkVBnhH/asuQDnJ4ZZme+syrDst5rHMVf5omQJky3xDIxzl65wAs
RXQ0FcmPlq8ZDkxk1LLxuyn8TGwDtTG0ltqKLUxVwb7i0sQnEm+P48ds2PNEkNv/5TeQ5hB4pWkl
HTTJuGnqOuHlnm/TKux+M3gENJgXtwKAYF7MIruJ6QZBE3jVpJxmh0jdcoq7v/KvF6jwdCrt7HVf
qJDNl05jiIGUC0EauKhZ+SKkZ5Td24wQPZFnd44KcF3zfKW4GNegd2RNVgyzkw3luFKxHEfpKD0C
v4dQYBigJT5FNYNzfovDdT/jIcuzm1BNM1RxWWADjL27l7Kuap+oyvLUvfZbfbwsZgV7IQET5LUU
7F6S46VBW06Jz+nAdISEYCC9itPXS/6j8ptZfTSuXS4jNFtpFlEohB+A6U2isz6o0If5DEOSc3Cq
g/YWxeirU/VuWolDdHM/2JHZzOjZMd6RB8YqHJm4hhKvcoXjoEHoZX4Ur8CXjeQ/a/rUdEg5oP1R
gE2j+72jVNAk+asEM2+dYOBWkZemJxlH49sCfNpIjag03ShT3QmMj8DYZBMs5QpQ/mAtPWNpq9Of
watuyvqNBdXFj9EPq1Ric0WSYjadituSJ6OiQYA+2NjMMMHiR+E7xD5QDTqUNIiAwrYX3N4j3UnQ
e/m61yt3ltjIdoFyj2t1ogWz83fuUqiPtnFUR2233Yl6usMSRzHsoaIRCSsb1wuUCy6Ms9LhMidl
/noEzbvBo1CEzgqzDAs88XXgznV/WMI4z3cM89LWC7UGnpct5ywTLwC/2xfZpTY+GKx/wr01lITj
9v/Jg2ok1ModN67TgoQxoSvQpW0iExsH6uuBnt1TWUBlo3y5QukraDN/J4v7+o+e1HLYrUFuTQ3D
L6NXRn+NVQtzJkCicyB2eAIOMYpFYD2SgP3H/0BJFRZCEDsd6/B5gE/uzUHP+5NCtQ6oIN7Daw0q
Dq5k9YDxBPwqCwy+v1OpXvvAjccvcQMjtEpUgcYPFTvGbHbeM/MdUCHIAvKuPczjQVzdKc8etY3e
whk9bRZAxy4kk8U3poajKiGPH2r+avlFE+wJ0CzfXqgarkEJHqxxRT375a3wPVDn/JBUQFnxm9mk
eiqAJ5pl5D/xBQlRtpZdH38iyXfD76XP7sZrEWb62Kb1qBBs+rj5m0u1wI+W24uoj5mU/kaAwEHL
qwPAxPOnpM9gRm03SlhAWqAbYvzZ55/8yZruqS9nl7P4IdrCNYtjZyos24vUafta/4J9rZos67JB
3ImuMKndP0JiR1FvNWCdGl/IX4oyUBAlBM95UT19/zypjX0vQKSVJ+eBX6wR/znD1Xp7LBXfPTeI
F7eiXVU2U01Lggu+2F4/kxOZ+0jA5EqNE7sAtl6UXoaJx0cXDMiStQ2iomEmKF33Rq5BtuY/OtdI
REmeQLKLnbQq5x6pBReftCh0i5ytdY0oUCb+VpcAA+N4oc/a2pCnLoMN3PYlA1bygmrxtFfuRE/k
ty7/Tp0hOH4fjhGVNxqt6VuJg74E5p8EtLopbKQb5Ki/ePeDnruSmFJbpBmPcZ8XO255JyYkGd9G
fEaVcHBac21xr01TTUqQEaH7W6o9V5s6/eWcFbB0Mc4zhiqr3cSikklDT47d4Qxd0JxGIQdfcpNl
1HOwT3k//urFGoHhz1DKlT70XEE5npXkrby6aqrWjmmb2XdTxNKXdLfgSir3DBWCG74NhEK3HHy7
driQXGYe0IYdnpW7Hr16t6Iqg4S2EjKlwzgqC1tqNOGgm08/Acp6Y9aQYOU56Cd0aVspmrSYTonl
XjRG5IV3b2B4vLQoXyRP3gERzVdLsur+L23FVpUToUUqXzYawZtPXlGNBJFbfLmqKFfked6GU7KW
LmmorBAyE9ZIyY1auS+EgwdzzpoyDsJOHcPO2YIXeEyNarU27QhmzpA/24+ULkivTvZANykKCDNk
TPL/W2Of0BF0BihZu6D4IF3lWVXa1i/XLsQ8L1mTfgZCyhpSxY+sx/Zo8glrr/lvQ+QduPG91+zB
WKtDp5eThzPCl7W9mX6rh2AsT6xekl2Lazacrsz1BmC2N4ZtB0HNMM/Ja/0E+OtxdB81iLRHg4C0
kp4OZtcL/ZFnrX2c23IYTuiMrrCPG0npYBMYQfXrGMcUxY1U+yjLcXlXj0tXqCGFjSnyBLCF+Edn
VQs4ShokdEBeyMK+V0+LQqbNYX4s6A+iCH0mKedHuHFq5KSz8MJu9GSGvLUCbVGHmmqrzE+1tAU3
l7C5RhLnBe6gsJPL9CLmdLPOUX/olLELM1w0YEBr9HxgmRqXrU6inxKvAJzLFwWc/FTQdizMkCco
QhpG/ScB8VJzvlPBdjKVGpqGMdAoCBA3cD8a3jqpDZwkO98ZuZgXwOuAz7OD1XmA23DY3ZjXwJhA
YlbjjBV7snQkJQdxjdBrZmrakSbaF04HR6t7Dbg9aEdmlmh1n4lvU2/p9DDl2xQczWJbwWvNwsIb
WRLV1bnDojJUEoKGwbTt1Py3azLtv++lV9rmdyZySbn9Xbwy9tr4xPEQ/4Q+/6s69kQRxMQibU/0
QuKcEC0V5/DS4njELcrpTzhLSv2WQnvI68IuC/plZM8B0bC7bNEwgOJcqfhUNEcFmcS1LC5PH+5i
Zm7Y9+qwX0zxJ/643LQzxYt0c0nfmZooiS9wy0qaj0/JvV5NLOP726lPTMcrJpz2uYPQFnyuz7p/
zC+kGQEMTTZU/b8DjdiTi1QniRLHp7CLVa/mz25I/ieNN2/0xoh2z7Zy89aR//52q/3q2i+xK13/
Rq/7vaAfEzmY0CsYqMr04tmrzQea2UVVjMrUv35WkrjRapsoCfi7NwlI318KHeDiAz0JFMZIlCDO
bcLuH5wAwhx7wQcI0y4DJq+R6GFpUOKI7fe5qwWVJDn4SB27P7B/wyW6Qj9Zn7y9x5IdSicGiNBt
OThmOX/v1j2dfULkoBwFmAu4fwCaAcj+6RcrIiPTbmd0u+WutlCT07rhID7xCIR1Ml+WHUb2wMmH
YzhSNySfRici7+Q27wWGssNu9Trqhgys+sp5F4WC6VEsN1lhd7cLbuAZWlP0qpFH/ylzpoVO++6p
wVz6yJuj2vsxjOPuqHkDxlsgVM64R2rdC1t0970bXXZnE+3J9VmxAuncvuLS/pRSxAUJAa1ha52j
ETpbix2K4okgtMCdIMdn99YpGcZZbv4iSxmCMztLkgPdhMnB7jCirEdq+tTOBIlhh/af79m4sMpt
+qBWXBEwLfVOvS7goF2HXb3nHTNKwUFyvWmSmTWkiqoFtG527uuJihm5uSlneXrs7J7y5d4PayQY
bhEpP34Nk+5bVsTrqI5rOTStDean3i7yRgjkb6zceqn2IyRNPQb5h0OzSb0PTQMxgedDel/eU2W8
Wa3j/bMQyZ+EfcXe5dQ3ZrxDjNzkqCKJLfjeqCTRhFEhzLOYZTLVURxPlF8TUUGi00U/i3dJqfRk
pLfptwxL85eYUwNRa9PqhQNcH7bOQg4bPQ8UQ4Q3LzzasBtto23s68qgnHe2ZOe814LCvx0CGoWN
s772z5T8Osx1C7gA99TsPS4VJq527QLhyIBlO/SR/Jpv5Mt2th5yN9KcyQ3KVXLwm0uzPISwVije
evKFLWYqr2LvNCUJC/aCxYIbmxGsTyANjT3UgYAJipTBpPMY6AbFqWgMyKNGGkW5pA+Yd8KMgkNH
CFwLBGRbI/kAM9qIt+aR9EcNvV3yQ+Xg+3RdhjICDGwNdUY70qxkwhgr4nymTQxrit3BKPA72G/2
MXazmNXYtZBp1hGHdGmVgpjs/1Ps5TrNaGv2XYbaq7A07sao2UmvsI8/iUkM2sw9OOafQ9K6Xn/t
ggbUWG4h9mHHnre3bp5pjaeQHXQ37WaAvoU1fnzhOj9O8MxuDfcYnT23L9Sg3ncTdpxN6YZgzk0B
gVhyFuAGMnmvz0QycW7a1+7TkfAQLTBhzvibNs1amW45SYXBc+Lzxg5BdSbhdxMUtHo1xl/z1+Zs
xvPTMkBzIwZdXGG4O1DTEyqBdkljvxrtSSsBGpFbKvs0c2V2PVXKniOk7E74YrenPzhhoSl2gDMl
guS6JcK1sLeExZNPqvKoPr0dTsf1bZlaL9AgDsIN8sW9LIyLEB16C+/D8Wd5K5Cjq486drLNtuoR
MlQ5QvUsPA2j2D55QgVLScLXE5rMsS5/AafTth/GB4JQ+BAint2y9inD8ZQB/qqbSLGzcIUeQCbm
lfPeWb5MT/3yPuUefuf8cN3lZGzboSx1jkDJ/hhuC1duJoTwRX8+ML3RSzwW8qustHWIo4BAC7BT
iYXhkkwAExUTPE0UDB1VMYecT4BFvf58WOuSvorsVA6zHpG9k13ySAnn5lVK8bdzNm6IXPpoAzAA
qDuKYftgfrKEgU/vYC9c1ick6ZLImlu468mYKaN3GpcTbgeRAx/Zjtk7NVRt8pbpQK6saVngJa3j
VpEuiam65Ca6qx9EdULU0QGyCnyyvg4Nuo7NzmgdZbEpZjpY7hhoCGjxaGdClQMi8tMR2yqZvYSa
pKvlZjrr+BsJ5KhO6nyw5r0+ejnWDb9iVnTKPHbOE6NLy6XI9ao0cbk9qNaj04EUydQJVOQQfMbF
z7rk0xYW/BKF5TmqOkCzJm1L98y1o/cKNyE98qt2YyGX43sINc21yaaws7VcbUnmnq/NmwhvkRtZ
X4JHlMmUIWEqukQd1v4ZmWTr6pLJxlTiPjmm9RQDFJ1mAvO0fjk1RJ6bCimTrvegZlDnCByMcENp
DnT3nMFyCOZj7c3gPvQuTM38Qf1kSzSydJT4ean6B/qynmio7IgkbJNbAqWqdfpEd1MeePP9YIab
nvpKQ20rrwGfesGu5aNzURxu4jZk+aChqQFwMR6k8JAXm2W/iD24uurDBCDB9r8WykzJNLaw4Uhh
iOy2mhXwXU23Is6s02cgwWbjqTGYeqNU/qVBuCwNe6fJhxvm4hm5NxemM1PL3bK10xyN/KuG556B
Yu6WqIjnLLos+o81J3QDSnSWvLCAnVOcagQHFdgxrhK8ng+stv28P0edvryfzh9DPSyQv37Dc97p
zMCoQM/0ux+YmgtmCvDREToYr0aqex6l6SpsXLHrERVpzq21uBHQ6SIton+u8QANjLtWZpXdoMF5
dK4z23Ddg5wri2ppilxRpmjZnwmqOfLjhDDe73Ou/miO+J16r4sQlAFp+HVZMGAWhOrUJKp6ggxc
6D3ZjH8VlA7SkPqjXyAoYLgR5d0clG0ko7CE43f+1k0aKUm3wcs7TRb+8b7rJjaXiFrLX3wAgt17
LltbzrwEKsG6vOk1hVvvGyigfloBhXnEINMge6/tpcWwk7oPSvCT/WfcpjiIKX7ce5FKujd7hayb
c1KtiP0bKkbSSbfzSEKEFI2XwvMzYQ4lhwW0xIVZKbk8M4gJ08OYEoQVKdpe98A1Yr07QvEZ6sdZ
Bznj7Cpm6nnYI/kE3TstqiBP6UT1pMaUpfqpAb/z+/TgKAk3axPnVD1xb6SD12jmNLfWRw/4rbLQ
FDH/azEZ/Tuk55qWcZXTbjV7ELYtooxEJv810mmi/LRRt7GZM3zVYzK7XsXe7k6VZg/0yG6qoPb+
Z2n7/Zdmt4jsiMfuQhgnc52car18OUa3y9B50ypre7DQgsAX96c0W/FF0rHztYT8KAWz08ws/7P/
3wE+XKNOqK4IX2FN3NyKcmwoSr47aa6m2Xsdzvy/v2YjqlPUes4ntGKWMhvlm732RIzRynhU+iLH
mQ63fd7jMG0bY1PpleMLX2FEFvo4UDxArWjgVTzHFvzwy5qevbJ8VgaIDoDSyMdIVWenS2iFWH83
ftk58WclxOWt+zKGgXAM09h5N4PhgzJ/1Fp/oSZK4kQJAuNL7ya7a8z4QIkl6b5GE7rdw07On3IQ
7UEi9Qggj8Z5boHpzuOssxiQU61XRXbu0udsb8JO2N60lRN1siIM6NjmvKFhoQCajRQsbd7rNwg6
5UJByCdKK5Hmo/7i7Lo54FEJrUCMnaMX3wnF4QsnuVSeRpKHJTxIr09jq8j8JGIx6U+WXiKCrudH
jFQIkezccQvNh9MjOGtZLFmyf+qWH/g3bZvYFQQyQ5TN9uIDT3vgdACwoXwA6/jo6rMTgaPa0wrD
voRa7kVP3fCsRAxW8kOnR2Y8V0T0UmF75h0LrwO6zezGdxDHbNPos7+IwUd6t4hjTEdwQMwRe6m7
YfBpS0cQDtqkLZKv/y9eonsIma3q1tIYWGeSn3m91Qg1IaQH1BUm16sKl5sw3FFRYlXVqsKEEBvu
xsCA9CcAT72Gguvkzf7dmysrfGkhaGui+4Jq3zXdW0+NvXaMvpRKRBN6Pb5C4X61iiCzSrNKzf1v
+95FwByunoxkKG/NZFC8gCjOmsG1mKRwj7G4CzsWJr7iNJKM4fmelPXxTYrTs5LF6CXuQNBpNDFH
Im+sgTMn+g9ZNAiwcJjalkKykhNnv8URQ7ZsOvk8YWxRdpc3KTLwI+lPA4Mta0VMlsNdAidrTjkY
nMe89WECw+r+7y39SPaXUzE/P+WN+Jj2iT7f/FZCMxezsy8QqweInnr6r3txnJU4t5EdATtgHc7Y
iTupoJubqH0iBJdu4e6Od9VjG5JcC9WkwiYfGp0mMjAxBOfY8R/m5PGr1uEogFR10MTEPQspmyv2
2X2c0mkOUPw687dZ2JYD4m6XkqvY1vWOQOpA/SmsJWc9JZo0H3LB8/pmaZCJKOtoa9H1uTEdZFpP
BGfgYPaMRihTs6mF7Bh8JTk3faBSBCoItaXCxWEeL9wCBLkpRHQk2NKCShbitE0hrhFaDHBgNTgV
a/cobsT8ED/QSWrt3cuXgu03gJ5nWYKX8FhsX//8bc/qM/MfEua92agGeJ+C+z0e4iDiEVgo/CgO
mFrTPOEU/lB7P07lq0dfcu9NJv1fpgr2T9LptGgQtxAiAcwIzodGERtmtXm8FMVtJWnP93USP2eb
aSAjOiFLUDS4XnclKzrEJx2oFt6OnYQbMq0PrtlT0evlJ4KPJaiF8A81gmXcFDfFGpRC1YmLEHAP
L5LHwvhzzdfMdXtQsRmZSaK5W2rRx14fbzBgtaeEBI5kuiXpqGDDacbe6Y8HgO9HtGNTyzQpAfTF
ShUUnZZf8PMQDmIj2ovzm0m9euAMPhJjNGcuG9A+RFkTrvBJRVPggZr4AlvyOki2z9ohTf/P+wpD
HfVrAg7MEge3A/DRM9x325bvVPOWz815WTan5L5Ra5KI5MhKjf8zTvjHOGG4g61BYrRoBzzCDOSw
gmq2JwEATTTJLLUWvEn4oXlrW6qn+b/VsO43D4g1ESoMeDdA97Pqec1gqJxX8rMW+9ZMm3BbyZtr
YDHyyyQIM5XAeEsyfM+61h//7xGUSLPLuubGunm4YBKV4+gj8RIN48xL2LjeVP2nPiWWh6S/XP59
agZujScKMw5RJREnq8dL118fCrCUJh9A86Tr5dtXZMFE+D4b3+eF6IZyuqonGtT9sEetD9Zrnv1r
Yi198X6vIAakNcoQ0NH/jgL5jVxvemleyuiP6kKssx1L+cYSYr4P0i8Im5IjBwcRgEQnX6DTZGnw
Z3qvywdup4d9pk14pAeXa+vPU4zzKoDieAgXucqvy6P7kHDxX53UpXyf7vhfdYVkUizYxf2jtzGC
CvHNVDpaUcoQVUg+AikKhvoX7Jruso0SK/JmS4IP3UsEt0ZWHuGHDWIVsOl/cnN9qxaPiFNrcqq9
zHpLpHv6hgF+8Ti6yp+z2rIz/p7J6qhExyv00hMYJJa6ndofM4I3UJ1woSQ9BUseM4WENEAPDw48
ZYs2tr/AXTpHJVyX03VOss2CO493WQ2HXyakJ9c/OOGdvHR2TRatIlalxibuYopThm5cd30Wn0QU
SsQtjzRJ4LX0BYnMWmC0s9qTMyybYXGGbH/t+7ffZux3WgTtw9ti+e3ES94Rtp7017Mapgtxsyr2
wtrVIeWFkQG/kDKQwdk1oFmX90BGRUM3mh2vcUK/K4Zvu8NIlWgbhyRe7EIiKNsa/6YAtetblWVW
DY6zCoEgfQ4hVHEYhCr9KwijvGq4gtCSJC093Xk31AqudEJcMyJ+IcQdAW/QRcCmVCVHnjW+Q2Xq
84Ms7/a+DH+OJ2Uz72bYOEo5vCJy6Ej6FU3Osop/Yd0q9juXVlfw0PI9GUXBmwyN5fOynaKneHcx
EBQrhRYiIO1PNac0B4c5zzrtLTbZivP86ALBePtVj+9DKYkPOveVqmmbrELRbVQC/2r5QxnClxkF
71eKnMfFwz9Gia7rLUToQz59q4uV5Gtv4OuyKWLFZk5WE2xzeaLgvBw82agaaZf4vTOxxAmR616B
LmALytK7qQv6oEQiB3z6BTIKTLjrHqnzlLETfp1qMhssFkKHNzxQfsErwOwbyrVrcCwowfGOXG3M
92EGCUIeZrJCBws/eq8rW6VzGPu+5rpg/wmCXNTM3t5K0zOcqac6coaYTbQDP1hdZYef4LZjLpxW
lXplPWRz1+m9p7vElNOWPmWLfJJbNUU2nAqDpm2DkYowB4N1JQsPeNk+Uu83Euc+ELQTAU1XTByB
O+cKI7p+gymikggqoAklGel8lWzVcS3qDVIt+CXbj4QBqNEfQj2UG9OJjTMccsXa5qbLL+hX6pBj
hrFyUpK5tKfmrUXuSf7PlqDmrmBAveZEd5mlzOUoVzLssLuPcoX6XKZvh/s85cqIhp8Ya+UIAMb5
RDpDydCssgVK0bvezK5HS75rpkTLX5hw/aVnnY8L1LsnaqTakxzoMwEnz2NhU2S7dnGyCm9w+fSS
Crsq8IUlvaNat8OxM6iZ4Vbw6og+WsRjUc3hbCf4YEccwagtb982kxrym6XJ1KxyZdflfW+hNQh3
p/39YyP8cVgtWJ0V7R91LBSlbjZIgoXbROjcu+42iT+naNW/HksqP/OdLjgBYPMsgosvTcgGIlSV
dZwuFPQiNO2M7a6dthqfAuLUS+F4sMWhWzF33P7z+grJMbrHoGOf0YJJojcmT3XX+V4u8VmBKC+k
2s8PZzZKs1Fxs++wiiPTuOsekCbL0keQAfi/8xaXc6xYrtzibZrhskYXoIjr+fJ0vS7PFUrGky6p
byiV4e0l4cAqyfNBoSKt5wTWcxs5Lc2omsTerWAU6HJgOaFAvt2wTqUqqNJ99Sb6d0Qv0e1FB8Kt
tk5XszEWRitws0xKS0FkBD3WWzhQh5pGEdW5QVpKb8wp9NvwncKgL7yWJuOx8/VZeyEimdBzlWwX
m4WsIUFb4fdpH/pj9dM5cdKH/scDFa5uhWk1AbcVUlM3hnNzdcnvrzrgg4U18nszb4kUrTGlDtTF
pJFidK4r0qiv1ZFjtC1z34AlEcVUHBmT2adquro0m1yz93vzPYb5ow/agtnHP9gj8GaES3ujdiCf
i4B5KuvLoq2CZrTnEdPOJL0pxRRUbqVFkLUVVOxKtHNPrIfBlXSZcDWGP4B5Gz4VhAxJdZIqPkkv
f/MyDrTzH4RKaNrTiLJWN0e1uD9KokYtWIPqMniVCD5q8AgMwz7ONBIGVpw6nyOJeDHnhD7MrlV5
sCMtYWLFkpX9lPl7lgtVA5qJsQxj0GodDFRUtzWFA4sQn5GNx+it9AgJK3jerhsxquc3fV2XU6dN
8+fGLHkxD6svDqNFLnNrTmcYxnwaDBM1BWJNWFcJKAAVhT0uxkzW9cjXDDOXn7AqhHohypMoXnwT
elDhX6AUFZNneqdWxQbJQQ85yNW8XvXC2bbkTbIEGds/kbX5zI8/VbcjeW1qKq+Ip58ZJcWk6sc5
JiQZn7TyQTy5CeLKdC5SJL1nNXo7EN+rFLGkyqS3AKVBHMNdzo14swqLHbngnmQ+wHhm6ao6C15e
Tr2mc3C6UFqEd4lroXbqOUFvHJzk2h3CAiKb/cdp8gzxLFmIS9Pr0jiBBuzjO5CvVO5hNR23EG+R
csyNyw4j5E82Eq1AdAFVo5yosYcV5O/oOdI+CvpYpoM+n2wgbxSjJQgcuWYC6OGxVJ2yx9GT02Rt
zsiujYzQQVP5DeU0VXFmKzrOLgEFu44ykbNII2q32v2m/1Hdc1qdqb2VDMMqM2MlVr9MNLC4rYCb
FcFUoPXlKwxUuVPEAny9eQ60NSuR11p3i/BjgkyPCGU9R8QiDPzl2RKqUPJ9DXS9nUuwppadHqjS
MznHsO149+k+RAMkrU8cfdCXIAyyGY/ZAmfjvSoSbNXfWms07ZlqLXX6gjhC5gxMPxqwGriqmT13
FX1rC+lZU0P+X01xaXT+QjywN2QpF+wwZHksUvfGF87NdmQibcQRuUIRpvuI8ETkAFBpkKZMBvGP
ZJ8S+ocn5wjY8tYe4oqFJ8Tmt8LvE8x6tgsvz6W8YhZXjYPLua0RP/YVr/m93+7Ua5Q3Dqd5tJa6
ai+9+fTfXuH9l+VsWq6EUSyYjW8/skBDcVCamg/S3nnEI86jgDvAYvPbmMeK0NSqYXFvvACjBDhc
Ygod44JJdatQoGU5C5srIjP7cV9y///aXhRlRgTci7QgpCNby3MhzHktpbAQaRpCsH3xH/fYT1uL
E43wydd0VJlS4vPA0GYrNmq1BxKiBbR4jRZGG0k7m1Deb914dQMqofhNAZkmCFOkW8FZljeMvXCY
im85B6PBKNGDrUGs7Dwwb/fBvE0DaDPM/zqDy6C49UPIvGl1ULBtCae6KPl365deaizvtX0FqLRm
M+juEzFJAl4Qj6xgIvljVc91LUQdUUx5Ra7Xvbq08zlLvVZ44dH3q6yRIe/O0XMnjG00RScdVlRy
1vLy2JSNL13V7wZXGvaUMpxdlIVCDjreU44jr91kZTwIp7Cgh0Y3+fQ/TUYuTyWR4M4k241LnWtX
3hnHJ93H21af+MYo9KNuHL5CxZJMKE4vZFBg7RzLl4hQqN7/+qRoaioftMYjGIpxLTYANH+0n3yD
yJvpGp9dSZyKK6mBaaNzs1TffXGo4qDD3BIz79JXhTO4zoTMKh6ZADr+fkX76vxPw1MUvmDmGv2m
6OhU5yNaFdYVrFsyPsh4R4kp6wrUEqcBQ+9cc1JzfhvTvJ23da/GxhzU8OoJse3f4Dlp+Tn+9X/J
PT22ubsiPEJ8D8F8G0MJRBc5LygyEOzw9dtl4kA9zOAc+mCCDp1dju4qxwzpLzB++pivsRnL9idr
vp5BK9oYAaLKhlFJLTbw+j/bxHz/qC3vgXh4IeWAMzxw0lBkhWWT2Bzs2ScrTEuKdzFz+3N6KkUr
RN+zRaqOg7TATohHUE03Jw5f52W0pPazK1CSTFR6bN/2pH+MW+tlekFIIlXl+bypztJu8McfJZNo
AlJBCPx8E4fsSdNtJJwsDtd0g5bZrmjoLealaHFWSWyYHSdUg1u8weyrdP9xWeFqjTr1YO6+/Jjz
Hd7zVFqLzqnZq+Uyr4b+PIlKQYlnRlTszGzgtZKuz8HvN1C9s4E7/Pzcsbvh4S4J69bHgP1Ltlq/
GBTCVaXMDeN53VJTYAmPYao9gBFdPnpWh176j1OuiIdwgHvbwUtt8dBKEIM405tRnrGHplNZjJzV
pgv5WR1w+ah+roLgM1RMdncmU03t/oWWup6Ze8ss9beAhfihLciDgI3IiEAQFOAbEDHtSxaKHjBP
O8NF1zNTeO24KKZpDR+i5mO4bRoWxWhNU2o4pTfpTZ/1fmdWkrCY907ibUuZZoCEIBN8yQeVroqD
39tvCo73N7rH1nB1f9w7nxNdq81XdvPFmhq9o+zA4Oldt8E1nyDXic7w7zT1VyP+Ky7wx2tr1jHK
Ov3ol/G+nUKCEqDsIKP6p8WLBu6nhaisPM87tJwSFwyXfEiYNmU0xfNBsMDDdAyhwESq/2K6W9/I
PT3hpUfy10O16b/zBSLa4YH4uI3oTZb7OWIzLK5u6pb6wlhhzV5YiIHP0EMoqWZdFzyAJO3JE54q
0JbQNz6XZCLccb20/QKF7NnqaN+VuYRfKOuvtdzdOGgyWJDdcDrxkikiPaLvrfOE86sqRFs9zop4
iSYTG4ZOPXP8TamioICR+o16sg0+h31xZEbvIxD4n2BR6LRaCg5ZGzodUfZ8sQF0dM0oQ7fLWxIW
uLrsUe6zdfmDoADhE5pP+ep270lTDpKd3zskbGOpwx59K0M1gwcLE4DdsWlFe3b7juwpQOQ0FQV8
h5X3xvD9liJtsb9OaPKiGE3Jr600IVPG+Zr+GJkFGbfQwaxjFshtRV+lTknER2qG20GfncW2BSfW
CxE6CPaCMNBDTaQuBzt6LKRONvDi5/aun5ftKrhNJYlDQqxWLsMFSZIs+mpia4S3f/ut2IZwYHkx
tJBsb9o1DMfHPcXG5GCa9TpzGLl3biG58Aqs4CLro8ZTd2wfqLi2QUoZ/g0W2/7oSxFL7HM88QZw
8+MR5X0wRN76bN3i5HulcKhLEqzzJJq9orTilqyKL/yPy5YWbPMwtKiEG5V8BFmLgLgmzzDFhOxE
PJ8QmKvrcPpsqp0tqhbwV7qySNIZPyIi//R2xOCcUzAWM6ua8rR1OdA4gjyxtkBG4UrBLjaP/WK5
8bVqpyqRYgYug7u99PJ48plBDd470bHwfxkTB47GdqyCte2ObLX5PEgmkccdvR0J4Hjx5m4ARhXS
QEmJBULoo4BHI8FzUZk4Fu33xgOO/KRqvhExlfzXBpEISPh65PG90fk4USyVOv5uAvi7f8F4WuUu
srBLQJGjUt1iPylHJkIHN63RszvnhvEaPvrExJ+UstlhQbzT6/J1J2e1YbRvrBJB3h4VTfT8TIbG
pq2/WjzYLuHiggEYuTSELHihukxSGJle6zd1HdpvidYMbamO8RcWYiE/zF0ObryyolcG1NtSpHNc
UCuRNLE5ZA/WT7oq4UCn/J7yGN6YaXtVv338Qj0UM6Faxri2tIku8bv2CWBB4hnqbUV6JH4xFha2
OPrnPur7adixE3UfdYWeeGal2gIgWq2APwjpkniB4tu8UgfuQxiRZ4VLjvMLxKEcS/NlWd3QIPTt
nwouXZjI8n5reTC3mzCcTQ/P4mtQ4Xqsj8od/zDoHLPOGlVShaw2EFXUEZrfxz5AMSOF55r+K6qz
jn/7ifyoivMBai1CmWdAnCQfkjLMCDP0itogQuE04l9nu/YrxqTLyC+jWJGunEMOnJkwJiqVVE6I
FGdLQtIxVjIXUI1fGDQa/IFMFasUO6JQqTnqJdtJsrJmoxM/6pf6tuXXKcLD5M1/dsDyFDKSxLMu
4EXQNBNia20/3XIKTo8e0gST55Jja4iVhIF8GWvkoqrWIgicQjX8OK5M2JlV6JPPoY8FZgGAIupk
ha8t1XYkjHYYR3x7Tdm9/+OsaO890AU3PpCgqQaX52xEtGKxCzMNBXHatQ7EX1TbgU4nwuS6VxRs
6ey8ZekDxlyXTCICLGc78IJVV3YyzsL923cjtcKJvsp7RvI4+BRf63pfDtPCMehuYXVBQ7JZ5ZNS
/A6+H5JA3JMlgXCnRQem/b6zUGvVAOA5qtaMKBwj/PIIJ7/5Q9CIAgSq9Szo6CdOA2tlwqSZeK0N
zE5ZCMWBY6JtmMnIs4wh80rLQNItYHUTncnliK5XjcwKg4g8JBOxz+8ym1IAr1ZIC2wgTOKd2XVV
P2HdsBH8SmFwRqAoM+dvHxTt4HFoTmUleu0F9WPxem+7f8GOMxTzWriqO3GK8yYAlLVMK5e0e706
fbVLT0VnUkL336SPvdD+Kt2yJeauFlGhohCy/RZhrX2zOG79QkLMyEYsoVMHxlo+ekpSkAs/6XCi
JP+wG+3zjH3Vkf7MmvBZUKuw5mJijGC8YlaLnkcnBiGqC5DMQZ+z53KnntdW50daw5UQQC4TcC99
u6TvW4XaDmdGfvYxr6iTtEf4hPLd7Xtdmw/+lnpoEbzb4ZXcK6tHZfb22Yg8fyuOVBlV+7lHzxQr
JJZ+ljOgnmdtSEClLiB/pHfx8g0TotKaI3mMO4X0mIANwB6JSeWyUtEUwHoia8ZOwzF1lwlU+Xmm
LDQkhkKwfnA+HTbgYncV7QqfntX0AdNZYcWBynMb61T/kQo1VlC+H5S11633I8bVsAt48sRucwIF
+MiPpW8sERe2zLY/kJhy6bca8ngXJiQYlfIRzZdLpjaQX9Wb2xZrTxuvJPpGlEMxmthA0aIkuDBG
+nhDpOaK587IZnpr5OpPjnwl38JlP/x5/EDLNBxozMj0q6wWg04oMSW59dZ3mOZekJcNI6AWVbp/
fmDrLxKU9f6MYl/iBSfQvXMfercerTVnCLgmvw6kCLrjpU2gyKlln2GXqCRWL2CAfTDmXoxGM/2s
3VLicXVfaSuZnrYaH7D/iVBauQysjHee32VVLuUhI86YHheiN7orEC/GLzOVlB3m2NNL9uOsx+CA
wf2rHazeUwnxgsYBW/FnaBvHwkFEBAnG5+ledZXPmUPl5ndHj2vSD0S14xuA8Zry1dytmb0HPCZz
8lGxLCzs36WXJK4UtuDddEM1Gdozy974KpoOVBVU3GU/DSs0G68MSf8eicAGxKyEs9eFVeKEnZIl
qhMWljAP+pA9MuZ8Ntn0yVYjdPyQDq7Rwpr/Lcm/5nZEKK+lxmMf9Q352bt6ufaNzWQvimfKEyMI
4IKa7Jgl0aP2fzA8JiJgVPtH6uudP3s77QA5WUJ59KYAGhcKIWOypGe2LtpTVQ4h+Lva9XfFatuJ
1DyDO4+4DMjeXCwAkTYdDp8IMFMOJCmPcBD/7pxCJEmNcVau+j1N0zLJE0orGQw4IPOk/A0fs8fG
mwRY5hxMrHUQh2erLBWfeBZm2/hRP69CdI9UTWSHYCp8z5MMvrT2iSNDmMNOUPdBqp9r2m/QE7+8
OIK2Jx1twbYfOQfKvElAJdJHDu0/pdKag1knZ2ZFw/MGJZ1wwPh2vvoYzglvhgqDhCWApVHQl5Zb
T5huU1UnRku0ZXLY+3ErI//cdg1D+Y/9bY4vUSZWPwItcaxsPW0QqSRLEWcYkzU0SFF543v/+6JL
37SRBL4T7BRJLLbn/goX7aNvQ4GtNo+pd0aUMh6rBMaqWW0Pj99gdFml8qFhUITQNxT5vklRZn3b
N0fLGD2qiapIadjEGevfTNCBMSLveWCWy1PpJsRF/BKreNw2xn4aNTbgZIJtSQGBSMhi5/nTVteW
PyRt0lDKndcF+3MvCw4RbXKrT84z9EZNmWIPaJdeElgvdgO74KrBKTYZiP7f50bwxQWe7DfgEDOD
Vk6lEzkb7JA67HCllWzYMjyV0qm0xh1w1bRDR3OyNoD/ag3Vxk/0yhby95FywOSw2nMjA2wQyFZL
b0XKClLCWqcwBfnu8nFYPB9+U0DzPp0Gq4EG8qd8Yn+f/rs1x6TJpJoXaW1Imx9tm1mqtBdmfLKJ
yW43vj0wlgGirEwVemBU0IaLi8jzc9sDtxfw4sfOPcoHJFtC4Uy4hFiH4EEDLtOlQAFKu8bb48wY
FY8PpaN96n1Ii3GzlvhKxz9wShzF7DZe8c+VaHMbGaceVcL1BzfinQc4CfKitd/wPf6bBFvfTVHe
d5LLlutbsqhFHnKUJfHwDqHMOwE5IWYpUOmV8xf7IO1htXSSCnDwwC8vPpVPM3Qr0pdEXTNcGg1T
31eNLEWoBkGJ7wxty37x2dCkLyEy4a+0UnOS0viMJdaxss3ecwXmq9fC77BICBkCRnIdQ6gd+org
YL4ewMAr+uNALZeNgTGLvcmyEQYN5lulxWWx3jER05A1uX9H+4Vra8HP9lpe7Qx66JnnMxxblfGF
s7zJaXrUQ7wEcRqJ8VTG1C6ZZ63/06w1vX+D90EFIz9HXoIcXUpZB16VP2RJdxKE+aGmg21qYd2O
++Wg1shkGEHKmH8f7wUqzVi+sccvrdInZQ4yv9wAVXQ3TZs8NOG3thZM1XISDqWKckToDODyGtfM
5aFb6ThV0DrKDh63MVzXrxI32xGrRS+oHf2ZasFHmKbVccZHFlHAZ/o5Yqfa6nKe18cLqaJhYtq6
Pl9fRp+hj4Lwc9FSgp/poHMtwBWo3x4amqGUvK3IrFYPGgpPSjxbqPB+ty4qL5BXzyEe9t2YRgRg
MkAbMRnpeV4xzPuFqEZUAu5m/a4DCcjJm85g3Cyo2rdD7sZv2X30eWSgL4d0m2aYypjT1D6slc2f
kWIEwT4X5iMRMWrzdZwgYhjn1BXD5m2F6FCOswzjp3n/qn1ozobaBhF/3coyE7lR7P4oLi2TxisG
1qupIc1rAxo9XOXJp4/0m8OGh+JS306YhTY1VD8kp2PXSzFM9zALfhmkiq5YKMGzxZGu3+hYlWLQ
XW6hLyO+YO0hpaHqzxTZjXuXZ+/iGi/AVjjd/bkT4ohCN60mflZcWz3e5jypo+zKBvRGzyouBKPP
gcS3nRVm2iy+LJ1hht+c5ncdIDOi0hLDtBDUNv6Cz1NMBX5MLH3GZ7QD4X/lbWqRRnDBneiALwga
XgN9xzsTin7gWEkxlCHKgXUY8qqmo4uFDL8IXnwDCDampBVRfUUBXZw697SE4Ej/Oz6+L/0C3cK2
ZMQR3woLRCPa1H2no68jSf2ALE+lGoqumZFBMGDpU46L+G7nnI8I7HhM95IrT7Y6YzsZgTVC2Lom
6eIxinxN8cdMoYnxOsn80H3/VSOoFfLEXTJu5x+w5ziNbACippPHBw2l8aWOd6QbXTFCZYA+dEzM
sj95BHC7VBlgm4wwoKDD4YaHAUeULwFA6ww+NZy2/2DCAVtSMv+Oqbm347UvtEsCTjtaude4QGfb
i1XtICxMTH8VPE7sy81WqmZqNuZbvKaYABBBLm2kN1JtTckPGbvuoxcColcGQYRlp5dUJPHjU6cU
jd+uLUAfGyVuKUvsqJqPJmJX/4grxClgfZ9eqCC1lrmWcg3PK6/ovVQsk3BiRvDlDEsE+9iTtI7I
GopaFGPXntBfH5m9veJ4CX/jmSVwDk11c5ap79ErJ4qJxT0pRYCCMh+eMQBGNBYESV1gGqS8amLa
cljnS0amRRITsytD1ZaLl3avMowLr3bqsr7/aDntooTZPQxBZtp0+bTGyf/wK3qK/0EXzMwcehZQ
tacpiHnckqAH8CBrZOAmdiYPx1QvMXwdinvrvdzLzdX/zopBEjKczi/EjFhaQdWSGraoNKe8KQHX
mJ5W/UyQ68UeCpksoD7FPWjiyMQuW3szRdOJxOsHpMogu7HS+TzFNOvJCxleeBGX+2ZsVGiRIbyF
pj8Sii3BSdAMyFlANPMoqbxSGLDv1dZkH3FfDqZHDASJHwsrI3PSDTBkwzOdI+I0/l3BqLd/T+51
BPqhGgDT/9PDvvTTrlBMwRvzo5f4jZsP/x3jimqvZ39JpIoMJDvTGcrNpTlLbZn2o6D31Unlp9z/
l4iz9vG1vI4ns0XXOkuuc00gDqADxFTswjiGz7mF/2IFl0Yj4kEAZgMp8H+3LIJXVj8X9YI1ryQK
mlMzf8Jngj6/BnpfRpGbBGpPbwQK6SX3XOg3FdDZj93ijqFrcq00UCqc8xXRD1+Cu2otGRl/bjPw
eupSZvdb7DxSgD/15qBrkwoxAZCRMH479Sp95Tx/2Mwf084mdkQynTcztO0qG83wfAjN1TjDp+1S
mmSUSIUGGds0vIbc54WZPlT5pxDTvQ0HMWiX4Suh4qrJmNk3+H8XGTaL8AERt2+bdii0sV/6eGIy
3QCiYV+kX0NkMKnT7MeqRqux/nmYIRPuwoIUM4niCQCvdrKQjDMhBDM7XUZtBHIFgvmza74AXYjD
Vyf/N4qz2sZBgQNAPba7PjCJ2xxdDjAi/pK0bY3odM2iahZpPM7TvWS1SDo48/fHKmatodXZd/ta
/jPQMpXf02yL4/q8BahuLWjzb2MQOIv/JfBYEXN6xVlOouy+G2/m5TLdvQRaH3IV9WME1yIic/65
chlHVUPbTsfrIjawVSPbjZdbFHuiXhXf0+AfrMmx6zFLytXlMXJJ14fHxgL85Xy334pxBZ6ETUAL
87kc5KtMzXnEiLnp5NpCtl9eq2gnMB3ce6UEdFmYvcRy0tpZuhUSr6+RcrcGTUIhT/P3wLjH914m
ViglF1WDQloiaBRGwsS14Go061ad9/cXm6H2PfbxUudJ/0Gew1HM9dz1nJtPrg/ffWBK0dXwFsWo
/ahFfCxcDlnWZ3kT6HiVIXp1yYMrktO0u3xEbDxtr/ea1hZ+ELKDsKnN4I48RI0iSIm7c/pZ8EDm
TD+MaRRCGIYi6y0sl6QcREYGASBZtLOOHS+M3f9H3V9Y+7lBPVs5R39YjQeU7Cw/WLGOLMJ/MZet
7txfUpPs9hLbDumMzXvWxTtclnqJ3GQD/1BLeO8KyWC3qmkAJZ9pyY3IssA/3mEnTtDYKFentEMG
jM0devPgpxJSfYkUJ91h5QrK/MqOSt/+VmiqyOnUpl5gSkQ2bv7h91OnlNOOLOtwKqnsAqcnEPE8
dyugdwjx8iOQszZyKS7IjqEnv5a1AiW9xEtEB24reAW138e3fXC5yof3hgXKaZgBUf6QUlmXEQps
VtapA9RC0InVGn78dr4X9Q0ZlNoLmdplEDlMpuhC4IwJ2C216c3IIAJT7XtI+DcLqaagpOLCihJ4
L4cT42daJA6o/hcUpQU7yObxUFuCJ7uc72TMNndQIDzE7nF5IlcjkiK4UwYS/dWoGGMQY8tOmsvv
S3jrKojZJZXrzs0oDav1l/z60jSUQkByA+n6p1O4I2CGYsQAUUfoJYVqGohsSgMQgWZRhqT/+7R/
Rs4U0tkLONMSwdmS/tROh03Ty5qjKEDtqjHLap9tTs4iSLXppblqgRi+iodUVlkeWGIlvkj9l6OS
e9kIp5t7pNabK035eQ7MBN9Caoyj2ad4WVG8cHXb5gmfYRHA9P/JDgS5Z6Zz2TX0w6iSq/nZ+S+t
jbI9TOHfG50NQR5B1t0jpk71IAFCcDq+4h5Zd45XUqBgWshx0Q2xirziB1kBDZAqz51hnw6aPil8
pL+C8dMlg9Dp9x7sgo0wsobyI/gkPcHJUnBcKq36dZvUSIp4qM9qQ8DQxtDI/zu/WmObMFy0/Qt3
8n1l/VxAJATXk/13E891slLLEi+ljQtMhN40FOeZBHgAsphAGP5VvSuUQ8rxxiVdd2HUqNrB29bj
4naiRZqyTPVT6SFRDAqH+OZoAqBlclD8NBGt/Kkzor8I1coJJty1m4glVx6B5wo5o1NFzwROtBXw
g3xbyoQs1cLYqmXYvhfpOTA/+NMLoYSV9u6hDOoLryGYz18UugtFDLtraeduyAzt6k6JDNfqUbO7
ONeusvHZ0m1G20rt34p9d1dTwd4ZGQ/3JwYh+tFxjqI4JLbA5k4j/WzsgkcqsQFraBUGoTpFJRAn
/u3mVfizxFByS9V5tIV+I02RzlY4te98W+R3EAHEbPlSZ83MkuZ10oRvYKe5JNWDvi6ny66W8Dwa
PraCTyH22fw96WoBCcxdnzYmBlBjvIwrE4EtY/Y3u0QFmx8F9eeAtY5Z8lLi/hwssf/IG+3cTnxz
jQ9MmAgrdwx5f8GSvyVesY3WBTStzZgQcMN4LUSCDvMeynpwJGsTEcka9KVmjJQRWIcLjW3utE4i
FBHo2FIMl4F5F/L/7w+qFZKM4orN8Bt8ZOKyRY0P4gePcmQckM7PdGH6h/++I7x4BYqpReNHe7P+
J0DsmPxsj02hII73geEVtiDFDDPvqzYv+fTjwt73arGVJcX/HXxdQ04kDfwGWZxTSqHW0RbYvDUn
FIhTSzGqBo64StimbEGV6OZEl6+sYJmcvcUWl4fvoVYynPqzcUxmtEW2noyqrURwFsC2mA3ffdmf
t0JSpHM652IAvxHzlR2FocIPC+g5GxuvZ1yjevby7/mxb/NAAbQjvQXKPoZramcR2vKmaOosUvJq
uewFP48ilw+lyK7RpJP4VnqfLmtwP/EFuuHR6RdYyHVpl3Dn4EaKke5kmTlwRjn/JxG4BZXr10pN
CAeoM6v/keK5CPRd4SWsmGWJOMEVJbOaZq9nPsbjGoTFrzJON5SBZ2Jf+gyDISFSGPfGZAiGbrzZ
LVcFJJKmQlqT6YhUynSJs+Dj/afBrfmqNITgTlRvnIT25SpnbN5q6FCEYtnCZwTQpLbig57YqRGO
1x1i75wfUZ1/WtmxNOhFIIDD++i8uXCFSTNHg+DKIoBHYBbr2U5tBdH5ZbtepPO/qCWHalABREkV
Yhzf385CLFGz8xgHFxOWLKebJCBHCQsuwZaAwhow4VFdj6rkkB4vztykHlUKXNHABAdWKINFMXFz
DeERvaqm0m+o5Eqfx8387auSGSPXF2xSyD7wAWR+ee0yFdlaE+ozsYRfqaJqBdinIV6Ui6HV7IEN
yBVsePDMi4wuuski5vf7eRUUQWaOD4NphAueUDypxJcLXenhRT/vooC0VKBz8oNipwIdoCL8Mvh3
ZEZAOnH+UW90TI5P3+u1qEpoHEvH5Y2eSAZ2E854tyh8IRF9XOhbJSkJuKbK6EdYLr1744iMRvWp
WR8ojPqXm1/ZXqo6HQsDJtKXQOLgGdzDN/CA0snGg+SFfRkFb/IEMxgjnwe4le+a5Ef+f8f94Cls
CNirIqJB4iOElGJkKkfxZmVh43PWSzQblEbt3U+Be242jkooaIoOi156iBI6HaVLpX7k4G2j3scl
IrCveJTQ8AwS3htHX+SKZ7ssdfwDo+fovxQEKj+BCvKDdfiBm3Pbr5N3ZLAgSb7m82jfOHaCrHSd
PoT4a/bRZvLmydyurF7pXMu7WCeKNn6z3s0TmiWb9bsYTfGY4HRRoLMnJqpBR7J/8NlKomZmBLjH
X+KtEHnop+8ahlZ6jBcpkuJFiD/CXxDoMysnn5orklMYTQP0dd9pxmASwKt61Xx2zlGaY05tKb9K
sHTclI4UvcFMxebo6/wf1RulZHjqHpEI4fsbpBysufsQuCtIMR51/0YdKCB6tDqDrrUaAXJdz7GX
zVq0vB1YvqdQ0fdzayTiUX1HoCL2pHcMquxwfZK6hMd7q5rpNYUlf16WSbjuRjmbgqi3yGJQpaL+
NSxCmE2tsJK1KnyhVc5YTJ8o0+4AejptFzyb2yEs9zA22zzGaXQel27/nbMb9eOsyHBik3kKqAoR
rcMwUtfrrD/AX6WAqUF5bkSUBTsCSnhCjNmmWYK/Tysw3nI4hEy5A1GyiRGOQt2Sl4ynuz0YRmMd
e9M74QukXFlytZolvCJUPto8+1x+heHeaophDkXVo/9Ss/RnsFmkedIoQ6Noij/4/62Z0T5khOBs
CqUXCZoReKR5yxqGdhHMbluxAPR6cEPcNs5Cz+j2LROgxdHmNWCYaEfgiSBcwCjW6Wfx1x/8jqlz
1TsADtRbNarNC2P/F104scGGwi5sjSSXn9C/XRiSJu6jU412wuJ95+NKN5Sa6IfXS9T3ldNuVaPw
5QuqvFux3GiWNciL/zDrlMK2gUmN9CgW8B+FoIlyfi7LEwv7dBAycdJhN2Pg6oLqkGrjlQLlg2wp
FXR7YulYyXd3T/WaoddmxqQJX/0RbhGnB39W+2wYBt3+9knAugpobwZpWhzHJR45yfUvKJPf2dm9
e+YKkj4ilMXZsy/UeLJ5Wnu8IKQCNLs9hLNKy3yjA5g/4GUQHKbOKonOiyGPO1qNVe03jcuHHBgQ
ypeZ2Aie3h1djj/QMFUO/BtMUr/jVQc5F5CFLGGsLlunavHlh+HlqkdRmH8JTWOWPBsDSK16xKQs
w/dDLzntN51+AJTWhjVQsX/zRtw64P6AfnV0wtEmlv1QlHqMCreliCtVsq/2AxeK2WBAm0I2rmfC
7ufDZ7HjINST0YvzSyXewZf639+I6nLEykCjX8Sk83zRASjcS9/JRd1hLoq6aICwmFu0NuEdarKK
EJLY9kBr5MzWxSMxZobzIeszHGx8Aqyymp0+gPc+TFAEA3V+0BVgRFFJwFjGwenp7fDUJkKBtoNQ
2tUXHuSEzC5NTOaTGjnnG59EB2egwgqWmyINVFdRJI+1IY4ZfdWAhv7ykgBrYxKp/eCgcc58zSu2
boG6P32MrOk0wZzH+H5PcZ6Y34u3J7BelQxX7ia5I05Xq50om+f3A/lzLnQWkWU88u8+P1R8D/wW
ydyg7hkGB3qXOZ7FjWzS/R7dvK1bVq21IZUA/nZUDUOegFsJetbrOw9U+xO/CzzN7bDLm4fzPURu
/vDPfSPC9XKzoUdFerQHW7NBTQ1TmhMAj5BQF8gOAr25r4YCzzsd4MsjcPtUDtY8FUW1AdHoVu/P
zp7+BqboRX1ryuUrSgabKsR1UIFG/ThDKzBfSA3xo5M4/z2ilrgiQbgg6J+aUossZK2LreiOokKD
/JarGjfUCkSpuVEqfR84b2ojJAK7Tk4RDZkNnqjYDDiL1T0vFABSpMuRSXp+EIKCrWjtX+N4JN+U
3jBDBXfTLRmcHhs8S7XaWUoPePGhpOtv+zDWY0Z/rQp8qD45hHICQeoDUK+1s5h5uMKEZlXeefKy
98aZ+kvH/9JotS0u5a/pzTr56qPVtrdvGP0Hw8U6vP3/Eiynci4opFYAH+bnnxLxQjZtTneDcFo9
N3aHoGBLf6vtE0ELTRsuyee/Pew/zHnq1OLWTgsWyz9AthSGraQQopoKIG2BdAWciy9zyJ4JEkBB
Z731AAqz+YmTbLeqcJkfeJminEVTN7PnkHLLJszY4RYw9c7zIawstSTIblrZp75cvgIoGUYUmezD
SkJxGIWtIlx1CuhLh/dkJ+hoto8AM0afGgNUITGMSJiijJ77W4BfhAh128B3BrpN/JNOuk1ouvgL
TzmRH0EAhzqGScClFnEWGHx+CLfgAZxKtnoLLLbjCVVESm1fsoPUSxlGz+a/J06svsyEZ+y8wU8Z
zAR6m8A/7Qq1DxuaTloiSOeMXaw8/15S/uV2yTpLCFqzjeh6YmCabsa813qOtdyaA+XjFLtOWF5M
2isSMV8+CP90/pXIOqpUtOfWpbKr4yY3eTnH1scVIVbhKr91MJWNFDq6TzmjWpUQWgOmF4VvZSFE
QszTZEmw6qfdD3BBmqkCsmQH2vGjA9ao2/gT8RDgtDImSh09RcO3HU9P7NNbY3qfC1FKZKFeMrKI
xuuV33P5UqNREgkUHy0lAlFO0VfjGyL5C2FGvvB+CUMw6TDgYG5IzcAzH/CTuhQCe5TWS2/CM+Bf
TM4V+Eacn2YMm7F85fjkFQ==
`protect end_protected
