-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UflGsPdxsCVOfmdtzU5ERan5dP/tAXBlDOsO7J6dlZGYBOjOKW8rdtnVCj9lHEAaOMGxNMnhj0Dz
+ie4mp1+pGeE/LTvVNEvFavjORgcyLASm0wuI6lvbzc3eJUte1/mda750PkL/sjYKghVUaivyHWS
gcZGIwpplFCCkybvYsjkKX84iXmPk/spqgmp3wTbTnZUWkonhNgK10BwMby+bQJSpZErEOqlbdZJ
ewwbWiiixcUov0FF1HawHrgAA54qBepu0y3ozvf786VHihNiuVWQMUTaJUmNvu+fqyjiOm9HAUDL
seySgNEjZUhZeiAwUFCrbGWEdQvSNL6n7PRDvQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5296)
`protect data_block
dCp9+XtBF7pcTcyvPBKoXKvx2nLhh4P0l/g4xsz1PxGaglyDoRGI7GOG/tKaJIoBUhaOC+365l6m
RBU16WG9l0uQ9B7PZ5Mw4xnnyhQfVFT7F98PhFgb+/40qMeaT44UZ8SEyzrw8B2T2vQAcbkyT4Mf
pRe2GwyioW8wJdIoHcL8Gwmm6bm0fXlr8keRbvlcrTA3TUaW5ksrvaC6FsWY/Gkg+9tVtAsm1+pI
xK07Pt7RzZDOKYvFSu31LF3h3DxO7+EV57dGACzbYajTevcLQZTVzIKWWlCFeG4gThDGHNYOCjqq
c+/elF2GOOYWK9N17IzC/GaBxmPFc54LWCL66Ne8ASkKfcjGqLBoNy6zaIu6T2AdD8dYbMtpRT6b
cTxTtxHorh2QgYOxZPitEebch3sUjO+lzN2OQxdIWws8IOgbNZ2Bv2ec6wPoPhdRH0tuXHuPiDrh
O3V0G77AcGQtXR78GbXdQ8xP60lQ77/haVvpbdjvMNlx3j7leWM9pFlrJ9M3r56hycqXlmddXK8r
pJKUne1qrKd/X3FFxON7zCwqfaO5xyxtllpQmQjTxQC7dD61KI7oDcVTQ5qblycFj1yLb4CUr3Il
2YKqyVhzDNXFTqkvq+C8dwrfmo0FPf0xASYm9iEy/0hKrLA6tp6H1voQg7L0YuYKFF86VNIcbTPV
t4kV1kmy6IgQQw2PK6yfWVxpMApjxVSPqDdMyz3ob+fq1hFSftNzOfhw0EBhlLcWm1gIA8cFXAn5
vuEmq5mici19Tm9Gh7nZqX2YyQ21oO/I6c5Zgs6gP6ILUQsYgC0yDxk2rC0D+Q3ay+NC4ffsS7Aq
tnq4FJj+NyhDu9oaDtMXR5u+GLGJTD0Wz49GKVIqLh7mTO0m0esNMMhXYIO76F8jl4yUxctq2s3+
XBQXH5lOkVNL59cz5yWtmenEy5hbqBq12Gccmn+/+1zk01wbB0XY5iqrJrX//RttVJeynVOmwnHs
FIJa5ghhOONJgWuaCPt2kxzd6+vaPk/jonwcV6u35a/0hii3PEzakCj3sMpsCTyGwYtaU4gr0udP
2Gfo6JRGtbRcnaUXa3Hu/FJpOUDzzmIbCApTuXq0PoZ09xu/D36wQk1673/NFdw2qY1W03I0z1lJ
QepJKypDJhBqf25FGMx7Vfxp+IgVYxLJ5I5eVQBrsqeMsRHf/0CZapF9NLxHrmX73Cr8Z9Re2esW
yzBdOAyRhM4WDLlXA/JE0/dQ3GfALuMJZVDSprtbncGg7Bp+cz6HqhOzUO1NxYqZDOKUxOuknfJA
5mqgMKxOuHVCRqQ7gnwkqnRBxTzBZmFOzcZZkhel5XxBd1NvmeOkTgX4r4ynzdLKFNkYaADHnKYt
PfQxihSPyrumHAczrx9ZB9lW2h5byj2w49AO0a4VOogzgkiUNMX4NQWlMA++EHwycsTZAsi7Tzbi
VZ/BsGV534Hjj0TUF5Fy7SbC862US5pGq8HhQFjG7bHdaH1ylSR76wTvvdVc1/RKzH6PigVR2t87
/28Lih+vZjDTqFVLeXhWyi+74+OPqcseEgm9oa59tmDYSVm5eHotAaHoKwPm+N0DjdWLkaCEBN6W
7j6Bd1GA0uZZ1Xavrx4r4SiKs7RC1U85QOZhTtRV4/uRqpeO2Ed09LKH6E14XJXGJMidQqoEcs9E
0KxZ+paSmCRtcFKxEGUgPxemJ5cj1czO1HEtOe6yidpoKPHoJPcZ1IDfzCXIwjkcmgMKzgO7Ndmw
ERf25OsOYZjVXMTEZIeRaZY+TS3XKNe1NFzoGhkAD3VLSwioPIaRjIVs5/PXhtuzUNVlqEYOTUmj
hPyvv3Va5ToSN5mdWclSJRBYXuWxkNlBoofP7VCFCFJB01EmrH/sBwafeV8AlN44ZFBGEvuSnCD1
M4q7Ma1b3sIDCrmJYF4fyg3FAYgvtuLSzcPNRrMZDE0qcRquJVns00K/b49X4oz1Z3HlpMxIQRCW
Hn9V47dB4N23nIRGQFJ8RJ9q8DuTuH/+pAlJTvzT5nf0xKVArzx64dPonNuTpMwllvPyA4fo7WRc
f0VkXwBPt1v60UNjaAI5aIlzaGh5x6nDG5SDB3FMXmG3ztfFECzo1O5I9lpgva0k9PWawLd7EjiE
c/aj8sW6+0ulZkddtL9iwo8IbTU9fke1EQXDvscgzquN1gLL7CtXy03Cw/DFZDMbuBnhWQBoHii8
RFCviK6NK6L5QepLyfHBqYOI6U4fhQmqjcu5fX2srBrTJl0HSqsW4y3MxACwGkujar/VfZ9VxKV7
RfZdz+Nyr+/aQLt9so3UbAvT00US5s+XI4qeKgVqSi5rl6xVtfAWUZ3ssR8pCVjXEqGH4USjjk+Q
X536XC7LI4XE13N/64NivTxGc6vu8IfaMyMDV7NnrUU1MGW8lsIl6xIF3wTWIq2CTh+PGPQpPBBx
3GrfWPKvHP48TQrQCSRR4JPjfUM4T4hMt+dr4zv2tVfI45az6dN+NriqstoLD2vc9Gwp3PgWFt6c
9rgpxdttfeGK+Jr+EWmf3J8qx/sguaCPOsVUoTifYqqQCUS5wMBasZwWiLrlaB3KmlJRsf/B8ck7
wx2iSO86WQ9q9cFGYcujjgg63m/SPyrDulxSk/UXuk2q8OfvjXqxU0ab964riEsqZREM52Hh85Nn
WDL0/jw3p2RVgm+vvekKJR6U7Fdkn9uG5hoBbv9iASHDVw308ohISBCnBsXzGi1R5H3bxqqLVKzU
5sZ53bKeeB2Cv5o2Bgvi7dlXI+zRO6SBixpiBcG4GUO2nonAL0vdBJ8LZhAKsLQ8A7hsXzeBHYdE
1hW1q6DMsA7Pbim722wKLjdpUE0Ct/kmJaSJ9rL5Dc5UveCUlztK/9vCbu7yST1kQ2Yl+u64Gs8n
20LodRXGseqYSj/W/OcNWsEb+7yR/Qji3INl0Pq7Xl1dxebhceb27HgRAD5CBjuzjphiFQ/DMkT7
5GuceJVAICsstb72IyDfJGA4ojX+y2LIdKLv9rJCyf67LPRFmIAqqRSVjOWY29AcRrcoOLqfgqf1
2ug61MOZoFpcJOjET9jG1QYFGJgsXG3v/32MUk5Mn/aqZlZ4OtJO0P8alKpjlY5P8Cem9pCLTrhn
tY0qevLxw8FAlDZqwMwrmQSDKpqX3JPgkKdRZIS2NvfXpYh9iPlrTNLDR6uLoAdVcMpzA6lLdFVS
z2/DG5z4RmqVBTthMJoH8TAVn006GsmKMDY7QtyZmj6rxCyShb4auWe+rW0bf9kS66kPaYDlwMo/
/Frq98HPJq0qTFXNBonnNnSSfz1gXO21G/geQ6g+8T47LJ+C4OZNlNnC6W610sV59CfKu1mIAt15
cw22Vdz6149Dj6aCThF+dvuy0d/mqVE4k82GJSZkxDpbf9FOBrrGFzupRbXjvUgmq50URPlUvbx/
tQWjWWFaEXooiz6G6fGLuA1Ue+MUC9ZZaC+7IlmSrlXP+es9LCANmAIBU9UN/971J3aBJXTQpJ4J
307zJvWOFf3jvOcuZkq6SsiZKOpOcIVxvsYUR9LwcaipJb72OHscv1Q1M6fTkbqmk3IC7GGG+CgJ
O4SaZ54Q3NRZ2c5YG58qZRtnpS6pMKEkPfkdJN4XG+DbRxiuMJ1nKbuNdw18BfGxoPUr4dcY3jLk
KT18/k2gGWW9tE9FOESQjTWPc+MrIEgbG6DrS5OXwd9+6hsZnffLwi3iQR0xPvMQX/yf8KpmJApv
V0MaY9eMypBLpK12MhWaUd5NhAvegg3peZ57VvpK4UC29WCmtUqldH33wycTxaqG0e+i8v0zuTsj
g/YL0WFoBY4SxsQ6f/RRQ5vnokuzV0GrQf5UonATPWY4J1Sgvn1KJUkNputdnKFbNCn3726P1ZPu
KRuw/aT8k+3Z7I16ecXkfit/SM892Vp9XZx/TkWxjQPvhs/6nnk7Q/YODe1bDFRhew92oqhhnsnp
qQuRPdfMSbE67Kz/VIR6K91GCn1jZjvDGCsY7B4YQX4+5RPhQYYfG/zCHFY0G3oqhvGTuJAUa0uF
TqUXmhEvChK89dVYqmnJX9lzzdrARlv1b0gMylbyf4U1DKaiJnk77R5LcABM5S6LR94VuCPFnMjX
NwFyT/VmJZ50cAQ/lumFoZI5eAF3bGX5o0/Bcw5nMYTc+p0NzwyFe0Y++WjyUJ4/C0qS0vtmCeyl
B1UwOstYL0SsPZ8GHC1SsP9Dtkbpnh9fGLBbcssybX6uE2EfM0qlk+MxnHqaCzvn2f0IChPbyh0v
dPnfHpeSIl4qxk9MecDbuRT5oXee9g5TL8o4NxXVjjAI6ZlP0HZjRTFoLDG356GRUkLt/jMyBTMO
B/1ptJ2qanpnKCQUEsnvqgnJDz7AdJ/zbJB3KiQljfUud58iYH//bEbCGtemAn0LHX731zSZwCez
4Jo8CMqG/ntbeCOoDPKZX7nVLpGZirkDuCxGG8TB4B0buv2qQs6vg2u3JwH964cqMt2675gxiSk9
y38yB9yGpipRNfn1P+r9wTQQP8Y1BcZBbKqKaUNgpwj3cG8rLaIJXDylBJWeB7kAeX9/gtwfZS4L
w94bGHaVRqm/Bha4CDrIlAp3LKe2kQ79I9MSO2mZgVN7v30Z+EuWMs7U+AvW76gs//0xXSKjT21f
Hn3oO3EhuVW4EyihnKQb9ywVOTsTCUnqGZt5SYOZL2VN+6+D6tnXdkHsBM5xM23B6gfWybIDPwx6
MrKlyxgfA/nx2QE/5GyoZisr0HBU/4AEHQifk22kTxj/OZTyTCpAGwCXcPAIhnuV/5x7OK8fIU0z
FdxI6PH0RDit6EzaEQ/8buIGbzdPJ+zcqrWpydq3GZFzv6fl8wEVup6CD3okIuD5fLbv3pfWNxFX
Te1Aa11b0O6X0+FXa1605XxV/c/0VFXtx7I5GyjRM5lhcCeuQ8nhFSxFnKatC1kgMIdFfcgc5mtj
8RYbRjpJ0sTBoNymW4yeVZ/XSeVHcNEj0qu6MM5cByY9K8/pisqQTAzreH167d1rF9UYC+nOktEQ
Z02vTmKk//tchi2WxPouFHQFMkhQC4rBi+9lGW4TYCY+QKZihuDhkG/FM7tZZJ4rmSoyjPtj1d+c
a9WTaFG7xS4E4qrofE7VWg5jC2iElcbNDCQfN+6seruOkH4oCZpr9h7T/0HKHAAmmOM8Qcm51mft
NsI7fXKUE+KNukqg6ZNSK8qnwWefdTbbaePi2j7TwyJzHtW5RIOHPhmZBkvQlRdr9T14B3//jASF
id2zptYlC2i5sYZWY3iBndaCdgfrAVPq7RTotUH0y1AHLzzgzSIbIxUU+jZRpUCTTMIbPRkCjTpq
hdle6YZZ7RidcppLeoHLJwnaB3f2NW/+uvAt/MsspWBkJW1w1Em+lIewNCpmCfoFACzv2OOtTkfr
6evjTcSNmZ5/vT8xYUivtI9olD9qv3DY23Bj9PIvj9C7tdEvaJnsYxfgIsGYskivOGNCrTRrARXh
8m3TbN7dtwrPn2ps4q5lA5gPOxQEeUCczh2NyaezvTJ15utI7JHs5HVU3uYu0z2kAFWP6xqY4Chz
NOQqPIOmmiNI3ou1vvcGMo2y4iw1kWIW2fFOAXj1rK4q+4WDTbkZLNqwUeWlUQv9E1xHVbyhiu5v
t9DzsRmThFYRNjMpZk/O+SIkI+kiXtci6BeTGdky7w2F4uk+9HzrZxKhyBNba5pC2NC8OybPHpsE
sMmvHlIoS09vMJAf3t43M/RRYEXbyeG1E267aUysQny5aPDRimN7vEDIWhtPjBgiDdujHZRoM/kq
j97sUvKIqkJU9Le4CmfOlNqQVWgMEiMUSmalk4KTcxREpTq+plj3rPLX0nlA6pwG+5X5N9IZxBxn
8pQxWTWyIJw/Xi1+LJ+EMl+tMK+swUte06VyiXcqQ8NJ6yV9bc+3zlbpljHhYSrK8dezqg/pOgmr
UEwN/7qoSB9hB1ijrRmoKPM5D/lqJEXSa/KTpTtjUt2uzCm3AtGJHX5YQvpJjXp3Ef/S1Vg/NvEY
tIo5Qus7rsmihWdIuzNKqm4FaORwo9fNIG7OG9qXOCYTseJoP4+N1m3YSQhHsL339XL3LfZtdinX
X8hl8etLxNkjN0ZfKZtKKNEwlhZmO/iQ6peqT9nCcxp2PygzlQdf5jFIIFKUq7YzHxICP+AVgjQk
ZmC8MtPzOSDB62ypOUDo+hGGFzM9L03XgCZoV/qQB53vR0cwTcuuUmjjnpyjAZ9YNW4BmoRzCHmA
M2U1a54YjEfzsPionUJTjE90quMjvByPydTGU1NiOxXBbOH8FT1sIO2tVf6xEpq32grGRAYhT2AT
TCd2GDNwX7Htt8blvAS0D5Z2YiQLT5gdqYFJn9vwuhz/LRd45jSvB1kfbCa76waeMNWh4pxI2I+X
WuBwjnkV5/Q4kt2D2zyV30vbc0kcnC6QOFQI4N019gcmscu5RoFMzdjVoYsjtOJpxSI4dVLJDSok
PFL7lb/ocj88lWhVl0adosCjgF5ED4YZvqwamyRiAElZK0JURewyHBKdJw56vsZ4BHagN3nYTylB
egZLXrHT7oGURd+UQsW6bz/0ZawlagkSqa3cag8uhFLRxcxRS7Pe542B1o2abJdFtcUzsbOfZ4nw
czO0Hj5O4IDS1tU+0q6n2liOmXmNW6WKtdb2HxUMATqlGdznOgAEMHE2veorscWBMcSWSHkpMYDf
6eMkUAQdivx0Xi9U03ja6iJUJOMen5wH4ruqYnACcjZoGhHNyhGGHfz/T7CTflS6+ft6UApk1Gdl
Mz5Vl5lHtWnoMFldO1l1RjLaabWQ7FtLeACQxc+4PRTDpj5fgWm5jvaQr1ZhcIEkeqgd8DPMFaku
tnlWB7yoUvbhGTaiQC6MtJmchSpcN8e7TC683L4+vHgh/1/kV1uhvyWZXkD5tmIIPArJP4DOuIBb
ZiTHWQx1jn6j1HB/iN0D7n+b9wicH2gnftb+Y4jQ/Me3oB5RqRyWsb5Jt4CzfmkV/n9kRdWWVEpR
2sqBL0DsMiX1HIGHvh+U6fFDw5zO9hXusMDQp0j+qWeh/eZRbWv21yTyyJQvcYsoV3fajQ==
`protect end_protected
