-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lLYaOv72DHLtKFhpBiasACsxbEwR6o9IquFVEVGju8TeqYokQNDWkZRK8OW6uQroOlecRX6KnQZN
H4Tna4B79pk0qcCtgkZdglYsWo33MFcXA0xMZjQqaXAJktD9JNJHgRzdMQ7e7q03Q2RARHlFJiOF
6CswZQTghLy1QJt/+QJ+SdvS+/oFtomGVWyUedzwiufeOVmE82bl74gyjLPLhve6/2MO7V+FVjZT
HORnnVoygNLMSPT7ZrC9TWswBtifEPO6QbFpkyGWRaNfuF3swUMXgWKQ8FZTPD7rGa43RRrGdkYM
ybFt5LL/ILSXH/Ll9f5cQkKpqewTS5ImfQsheg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
Ft2dlXObabNVQcQETat6feVmVVFXzAh6D4Cy1FkLw6nfIXT6f03g54AsRMwctxU2kPScZHgHUypS
mHsNXmbVQ1apWPecC4pTxGko9OkjVKZHIQ/ZJ6ARFjHcZUSmSlMIjoLxjQBV4aFUs9UAOQIHKNuQ
ncusPfkCg9trXZ8c8h8H3nkONovmuEQvRqVGjlr3WN/uRdsoUM6UHmdlrWStRgILygE1S96yuxf3
Lx+vvbcAHXBJtzwCuftGXvSXBgWFlutGCza/TdhoithHjfk0uX+puBAfBExnEtiyZePuNgXhPLRs
J/Ce82D6Hzi8OvHNpiVHV0fIW0iA3DUGpIoVTzBxSdM6ep4lQYOy5rxM+YsZeTigbJwZo8tUteh7
QjkNVxoKSsvPK6OMNUpmCmwAJt2eG/3b8zCC9wRxgJv1CtvMFdjR/5PfeWZai8zwfaB6qdF6lZ5z
OaB14r5WxkMAHZGQnkUZlkURho76exUxCcfT0Uy/3xl3bmT0gduR24E+Wmlg1iyVn/9lLQw3+eSv
NkZomNn7u1sYdxlWkIi+ObT3mB3x4sCzYqXvFYfFlfYivBAV99sCHYCJ9YfBPpx4VaT14YrfpdOY
eH+1BKT3E+kXFPIokkZlIrCxMu0kj6YP2UEb+TiYDDdv1qTw3Uc4zH5b4ZzKuewvO75HsvxMzjCs
9vwmmxEFxsxAdR4142SDMf3zg5LgqCZgIufuZvsGdzOB3DZIctOgNGRovUaZqXWOpx1mh3/6iYlX
mWKinxbfZGY5TmY2hMbDR4VJqESqn7lax/K6P4x8oHfYvzeV2hZuDo4H7g5Oy780ghkycdP+SEJk
FrImtXzShIEUvnXBowkQfJxD2uyaGWVl83AjqpLAHlyqbaHmzhl8WpVpHAbbVcJt01zCDtxCGCUi
SYUJBxTfO10iyhTYV/2f6RiGBMHs6TKj3IpmEv2hc6GOXFZkTlp2vxqJKz25aG0GZx+N13C7153q
IxeW93em2j2tCEqGnmLL5cHHy6dRN4JYhtItNEXJlShiT+gIq6HxGB363NPmrbwGXqVs/Xl7HmNN
EejIb8F+Y/aCrehC3YZbjsa6eordZDF00cDXiba1rBXyp/+Y2bjkDPozDWYHUyGOdHV1ir+Zcan+
g4iqp4BgibB9wGdrEgs99z2kEYvfcpas867VpsnG+xUutQLv2W2pTpDMe/6cd/yh+9ouCN26tWpm
pfmnSftuU442SFqPTNGJiaLEkd7Oo6tfv8CNBXOncTCbI941VgIXL3gxFvZNOULUS4BL+ZfwRSWg
Qp/5FfRB7p7NvzFOb2hmG3av0LK7/JH3lqsJje81ZRArtQbtUgvaUaxVSd1nRZ0DNiEy1tJYqOfP
YOMK9SWQbu2HMWafaaQjWJdbRIh4AQxWbOD3g/hoAwVZJGvm3EVfPEPTx9MSItRw09swEod43rAy
KuQ2VHc49vy7dJKqeNfs78mBKSScm+cG8ck5qmFQVTk6mokLq7fdHQuCPCFbtTLvF2HLetq6FL21
tlg8BPJa2SMivm4Cm+FsgMAevy2Q64XzXuHYSWvt2AutuWwX3BHP1ap6zqlYDs02SNWSlxhujfsD
g72Y027OfPLf2KdPuzOzlpvBsaD/DWwDJlVOUH5sdU0D9GEfwpBTLbtxHwjf7cJhkrs7ZdP1LsDI
Hl9f+HEj8lqGU7yD4gwEEz4ALoxo4n64sFRQmP6/b4SO82CrcHibrT5PmgdyO777GLfiQo3ED4+O
ABaebVIQA0pefHO78wynz/aEHhTSdjSrczqEo8zt9gwf+zR+erziC/cv0+zZSl7N4iru0VaaRXxZ
Mdy+9YkVs696TWiUyoi5QjxDxk0JNZufHqcVjfY2s5VGxSBGzkBJp2wXxSNAGQ5XyW0lvy4uKoAu
JJi8B5p6AfQTQK0cPH8xXYEeBrr6Ehi5Ex7uOLBacsR3zp0aYsrZdeQJeRqqa3t+DFVb63Jfj5Ws
upXLCjsjQtVb3Nnlm8Sx5pohhQrEdGdykbIPoL+Px0m1d4JySgnvp60mJEMPhHC4lpwBT74rCy6x
vwaLEmalY3hQUPnd8plI1e/EPBwJd5r9yut+mAJFeAohO9sLClGSedCd4+7raZkK22LzGF176ASG
EE2KHWlVpbb/DYsSUgiDFLeJgAWssu8btDwGGDCjtkazeE1D8CESSDIMv57ftDq703/MGnAEVJwY
sDDklq+tpDdWQ72GXNs8dekNsz7ko1pre6mpPVvv9OahC8iDTw4TNYJD5AE8AFMiHtmNAsUOGVjy
eU0x95fBdTEcvkZuA2Y33Ef+nYLA5OKNgOidOxZ1t3Osir6SVoAK9p44XmRgQJPdEFgkqgkmCdvH
xXe/GT2l6Dgrtwi9eddd+TrCf5TPuGQ04F6bexgeG6CUE80dWYBJZ1Y0tJOEVWZ/PFxMSFT0m1gh
59PzLarEhjhqpJb77616jruJE79w9DOx6Tm9S0qmfXivM8xn4rlJk46jnjJlGRDH7oo1qdEJKq4u
hjuu1R5BqNej/k3KjDWdJ62XLIbFo4yAz49Kk6pf+y8D/tPmg2MtPPz86hvHSUfuFEvSeDi+tR7g
y7ZZ+9C9l6SgJZTQc1J2w0lEQzuucpyZHq5nmkCOqLU7ap1WgmKxaKDqbaMaBiqkhFQcZI5+bX/l
naq7Ny1aOcIlzE+NArHwCGb4+60Fpr8eFu2D/MInboiyH9vbsM5VO1mGHIGlxzCjh621Mm924VOn
SCagnGIY8KBj2Mdz9TWK2AvxgutYrtfa62DvJ1uedtZCjn+y0ZDjo3YK6lUg7TbD/U8elHfJqVtR
Kzg+7rOEWiEuz7aFCbDPnqqoSdzxGXaTyhNLnd0MMMOnvoz7sxCjB/QS/ks8uf4G8nbKQOHhjokl
j1jtrdL0acgk9PobYGExrIPXilohYgyEdlZpYs+bYMdnBwGq9Z5Mxphcqlnm693yCmCMc2XXdMFc
Y4eiXNuxg/oSrv90sDaD/nMZ4CFiIswUMn93yXUeoAY9x70l4FFPclR+TKjchXgbj5X6RMHtvR3c
e+xKaXmi29alV/S8TOZQqSkUqzG+VDTxaZxobROB4pTHB5aZIzQ4M2jAT+oOyzXVCWbSy3SDcISb
x5MZS4FFSivdrpMXvLtiyUydXTxo94F68TPu9kZr6OXlsv0aD/U08rXDJqU4q6CWkk/nK1uUF+yx
GCZPmz/qYuwFREHwHrbwV2Es7y+xJuZeAdrnGDMjCvsV4SCDWl9w3LyD8mSAgiSrklt42MO1nwBM
KzIriaOJYOoZqb44JxZNJV4XOMKm06XmWH+CS1RXZlln9Qi3vO6j6uhXjp/SCZXYtKBkA8fqL/1t
J8Ttbw1Xsm27RxpWZfxV4Oj4wUYseEkF9X3Ks2ewUCGlXSczuOZGXtmZgkObypQHd8k/pL0Vt7Yl
ANXGIMFb0jFSF83q+nZTzEbo/Agy6b/RCskQiL6NIpzj8eKTmwxbDP000i+ArecO11L+lnK0nPfX
16x3GOFVO2HlNyCd3IjZy2rBaucAIMCXdXzt5jCu+uWYLztzfI+xQEd3Hsj+36K9rfDQ2y2Q2Eno
o++6sN4/51cCpiZVzLSKa1DKBF16ykQOMXJfRd6MdjzYVV35GiufQMNbmpdGMuzcGWXAa5zrlwPT
2ev5/wtI05Zpx4lUj1Ay15hMIZX5i9INBtXUzAycuyKTYZThJOJ7qrn9pX95zOqkRPF4vLKOlvab
+n6Y2bcipbRHCXi651fygMSXdeeEzOFgoQxu8yGN3di2gXQIJxl05dMv63LjGVE492WbaesABOMP
cNP1WULQOTq20efF8CbVyJ/lSG2AZWJalZ6W7JGNV6bR8fVc2orMCVtWIlVgrkQqvNBm1wFBFmBn
OLeAumcGhAAp8i5amF+dDFROlufNaomo5xtL+gN9RqIh6pUtC9U5meVJw6T0jNwhN8w6pkqPKnEP
rSh9EeSm0G1RDY2h47+S9wLGAtYyKuB2dvlnL6GRjzBXckHqhUf0Qphnol6J5XTGN+da7Kw3EcjB
JjG/1DXiXqf6j8H6nlENDvmo4GJUVumNJWqv1cFyJf/yNSj3alVQ45elg+cWTyPPSI2y7Lh5TSbW
L/1Vraqz2NWHFS7NRhh1BwWYvNHVftr77vIJXpggMwHJtylnZ7Q0+hAI25W7y0ob/igao8sNynTr
B5KR1p4qRYQ2ZE4hoq6o0I0tpVLysp/wMM6atdJTwvt+g9wXALwlObMeJj96WCIJ3e9bKKNktcsQ
hQoo5B00fxYvF2lZIjtlFTfzzWHd/MGlzx48t1JHhhk3XRKxdD/v90ywhknuDAxRnJB1OmKRmA9p
H92GsMCwBa/V/2ZVL4GoheuvM8po3In/U6FLNvmGBmcq3yjGaMMuhJThW13KtYe6FGnWIbasfKwN
yJhJud/u3txxx6d8y/BX0mO8cqBtvoS0nBje2VoivlE3uaG+DC1bZXQjQlikonbJgAmhHTx2nxoQ
ZJ338ZVc6Ny+Vwd8rBcbPm5g7O3jVetKRsztcBOYcN76GF1kLZFafdMAgVjMFDRF7LO+CsuR4Jy8
DRUvTS3xE656w1qNL2X5TbLoeV4JFHpjPzbo8llbPpOyZfRq28SikjMY9IAJGEImu7bj2o+UusPX
aTNo0qgruFJDhgkKDsVH1E+PeyekqyafXWZliDYmt7jC7Q9zOkVyITaeIsNF7h4D9x9/pSDEcnYG
rj+SL3gStafC1CIdrVjiZrWjGsTnmTLCZVJlqm+hzFJsETM1HjoZKs5ZkV/5e/JR79KVJL79R97r
p6+4GXz+EsIzCH0sdJaFLiS3r8UBiAf+1FtTHGqUzIuAtl31Bw0yJ9liZkOWkhkWuqNL7oooDcre
bNw10z2dAs4BT0owTFED3KK/D937HGjMz0pYCne/kJvnNJorlF1Ow6ephZarexaRlqrYQ7z9ZF1E
NjxSyppGadbA0lvfKcvTAVaM1ziZnalYQrKrqdQDln1FbyBQA9Wr0PGRVZyuwNX+9n4ETVqn9ocQ
x7qqJdo+xSku8qJQXGeVEtBptqd5By7g4ev9h9+3n3rkpXWdktyTzeQyuaG50XfEAyNwphDkZFFi
PjutuxlLZLrwXHlCp5tEZslQdD2goOFpe7bbFHklec8rvp4LETZBQZ34Cnivc1E3azBXVKXhwAye
13z49j8SdUBCWDZO2QK3G6+VzR2u0/grndjWkLZ+f9rMW6zYGZ6G/JqxEz8RUmfibvR4Znrup9D+
pAkSn08mzrgwR09NbG5qltiv3cCuhd6QOxOj1sPkHvUSdu/6eNNE1lp9oBb6NgEvUnxehTt1r+Mu
TSnvkOwTkjoRmoWRGmoUMCYnyca5em/tBYSreVVptsE6Bzrh5Ad5fdAGpUTY4w1O9fmfJboqfeVX
ynHOcYk4yFkbhvmye+SgwRzNKliXmVeVcvBW2HwE3n0zeByY3VhCbumydbXO4mWlnSN9bj+s/HhB
LzWrZ8FZMC7aLKpJoqOivtGQKXxRQ54Qk7N1ANLYx/rbsvL2cUGckuAHXRBEyZIdJLTAJz7YnN7Z
HxRn3YwR3rZYpm9dgQdI2LoAViazsOXA52K2bYDW//hfymT1OUq1Qq608c4Z6iMWUHqCaFhXbgjb
bKIlMADmZhpu216gzu9U/2PIs8ccje721Yn8cBSFZQFV1hwcszA/nivgtnjs3oG8UmznBwlytdAC
beMGCrQkXjiDT4HsdGLFuBMZfU21b3g5vGAOYhlRXfClD/+FbCfBtH3jlItv40Tld2pEC6tSDUfQ
HX+yJBYbMrFFmx3ZvgABQd0qQSS540llUmwiSKSkvIMccKv2cGe+TqW6KzZik3TURtXjbsTNee9V
MSkIYSQvRduV0RhT3tV1aDNi/VqruHhodt3r6EcAzfaLUR/IFYpYx0CoarETLZB4Gw1Eb00gbzE+
iy14Na/BXVonNSwLan6tzDYwhWph9/3DTxGAQ0cBxAs8axRxkt2udj2xEjWSVmiLnHk8Eiwu9Yff
B/BLHSf4cu5flk3zOgtoGZyrSxY7h9boLdbzFSpKSMs4NsgEi9ZVhbrLUJfW3Arjn5MX9OKU+sLK
WzHoSwAkyw5BNB02wgg8DsSbOEB08b28gHJzzGi/jxHxp5QX39EVQ+FwXyJX+xovs52oLHdcl2nc
ZfgSyBv3iIMtqQllJcYU83jtXDhmWrdZge6EZ00JQK5kjs9Npm38IWtsWTb8Ln6FnD0AhUnyO0Y8
22YF3xmpCOfES5CeKmfJMcKO84fRmeG4QXPxRWCwYRtQWIe5h456y2t9OJuZ46msjpn0d0JVAK40
ufrpR32WObDcJV8SuQ2hMfOUGp3xoFefm36rwRuKEQlL+jz6BlqWUD8YDmEa+U7AajwpMjbWR8kn
8jsoyPRHrOgjEntBgT7rvCsMLlwad/wg4x3kIcV5h5MwiwPDjt2cqYOxiOsXPQNRQgeRCH2XmSAW
IzMLwiiJ9QJFBB+JLamcoUPxgk7q6ZI/mqZjRRTpUuzu7IxrN4MO3wyH/YeuC17YNu43l6Vekc6F
XbQhyGpIeqSJKDFSrmmPF8wn1oYUqAMjwO5LQgHzpyyj+7EbHOMKC/Vx7LNW//nah5wdf0AvqNUd
+TPsCL9Z5KOMyutV0LwGh6KRalnTKtoDuvT4dt/iTIOKrrj/Q3W85ckI0ALqg3tqqRSr6VlNaBlJ
iVI4yEhYzZaPZpu6n7qU4O5k9nXkrkWszyxtfSrj2PhnAa0QkS0cP2/e5+RHZvR8iDLeDnBdOAM4
RlUPUddy52Z4GoGIBCehNR3p0NPBEzyXUZwMD1J6B45KvesET3T79QlRKo/V8oeWPh6PAXLeJBih
spRiBdsJHxOY6x2koGr/UCNWxtBnp7QBiZD7tm/uz0dYNbR0M1NLiiRSS5Tu/MEXJBk0pJqVZKyr
5DskJQjzn4ZJmz90nRxGDVcpBNrl+FW80htPXgpU0aSCqRePAcUZphGm5DuUvHn5LuVTLKJ2ABcv
oRiACy/q9QXMY3Aj6gWxCXOYsu0lNcT6bZFF/ooO4km//AOj2EfUNlTjJi0fADFs/pOJ7uWJBiSK
Q6QTm7rlWIXxb17V2JUpK0NfqrcB/womq2v3gQ3aCSalw0eE5Zm0HFlJE/vSoeXhkqTioXGNP0yq
o0NyewG4iQGSYyrgXuHLgoD9at4ODoW2Xda0A+GsXNFF78Q/0Btswvm+MNE5qyvuba3f1O/v+CUm
eNcOQuvNvCt8uIg5w09/z+w9xk1e/LNdW0JDNhpDRETzkDQSPeMqPvX6ASJMui7hfJ6ZXhVljT+L
C/oJqMI9NyhwRiWxabMYjlHHahnmzlcyxwZQCONAVfKG9ezxRV0hWhvlV+sgAMwXGQnipEcwjq58
x6Rk0JOKqdZY5BufeiAUSL1zfa+5O5A9lL+sY+PLSMF5QP3wSyXNxrE3Gf3fCMLk/gUXM/rf9Kxg
y77tvIAv3dS1684Mi3vlnEQK42A7E9QQG7HjwsedGqBeGp0c6Mh7zajISos4yjVgJPek33DhWf6n
RJU9myOyzQhvZ7yWAaAnq/nkH2sVvgi96zlb23NZ7HH5QnyDGwYbnBgsV1ZRiVtUCIwLDvchk0g3
6uYLkkpmn/5XkPhdwM4L0mMqNgxDFKntKPcu6ffuQvoj3EwHL230vOgUuUrwRXZuOJsopBE/mFwI
TKi35i85YNXZLjNzITsgM19i2JfFMUWHAk02bxKxslkV88JyOUzJ/tLIAVPXy+fhyx9C5MeKF/0q
uun3HWVuMKRjua5FYFQkPO/G3qq3beTMlyB2PkYeEBSqMZ+iN+34UfW1xvGq8PAbKpZkxPBdNRIM
KW0OIyDFrg0IkpjmJRDKawKF6F2GQyW8g9+uw7IHL8c9rsGPNJqjbR7vyugRRzAXf0THYwpU3uzy
MBYy/Vzxg443/B2kbQtGsLkY6x1a03MRjfi6qBYghKZ96MwpmoKj5TgknfePokjbYQewTtUW6P/N
psd0qZeYjl5EcoK7PB8nHjZEUmN31E3f2AKKoCdIp48EUrDY0VsUyfWGu7cJtavu3O/tr+Sbgp3Y
mKtWGp/6vCUeDEoJ+WK/ecrfOsHCe6LpwCmHLfjDgiHEjQTaIOPakkCpRBP6UYbKqbBeS+M44ZOL
i0uMGZuEz7v71Gl7ckCigNfi0p7PV9VOazA1vg1UHd/VCDvrrSU3JD/SFmOH8sekvT1GcSsL7c2G
cfHwqashKkymmkFC6nAegRzKo1aAEBfZL7WeXrkOfq+dne3AY8nNgXHc+WqVXoAEb/eRsH9Dg89P
BLt5fdrgzp9PwpLbikkWoAVQIg02Fpg4V9tXVMfmS/fXvqqPUfk9HPSJUQhiT/sVZbB4q3Fm41sU
lleyHycDe4P4AZz2pZSRfEzCszSqV+vFKxX3jtdPwNGrBd5FwsmpMSGffR7zm0X5HJkZhjxa8KXY
02LnxQZ9fAW8Sdp1SlXFSs0zX+DxcGkRn2jegom83R/LYXotJTFV5hIcnzZoRDkPNGwlP5Bhd4sH
mWJYAvpwG7v7of9CFyWWUwBOfYbXxnRscDs2lwatBpsJoYHepjgyxqSsmbZkm3py770ibqqEv+hA
joaX4/rmj3bzTRbRc58fQbOyyRZoGRVD/oYlbmU2vSbCI4POWbMmWvlVNvX18YVAUq5uArQWuqbr
9Y+OZCowWcbwnWQCscjE5TR2fCznGnVYRJ8gMkD6v5PUSykYOEOIjbEOf4oOHFac9T+wg7QxbfeG
NvYuBuOHxalEUnb/LhTDhqPvrZELqLVYkHWxdTXVPCj9PvzGQ6MVBcToTA8P/2iQICBAaXapDdVL
tYhkcYEoelYHysVf0iLg5jJAOh9/ypZTodCiE7ZAZzgR+6P6h5HDQnvAUbN1jj7i6ZVXA1iBwjPu
fELKS2pUu6UCMgRr3yDAMRmoVGofxaHILFsF9vcaxPmMhm+qjhI4DIQ9CIH0ru44/dHtsWrCyIxP
MmEO2smO7haxS1K8h/5sm96tSec3etWvxz/2PVYqlpSO2nK0bIuvhO5h4VvJL6AKjV+rmCnJBBNv
IqEdT89zC3nMODSqyBgoit8Yb8FFyhu6iZMnkW3r538TSkBm/FVeNjA5RCmnrkZMqW1auPNJQOqt
/T0BkctqaOP2+jFL971vBKH46v43kWVtoywKUGsUX4izM3TOmdatHYh8tTsMjQJJDiTQnK1OeQ00
4NVO/mrcqZaV6am3LMKXX/6w4K6vQ4nS00tMrxWio5FrIc6ZRCzE7Cgx2BTVfyYqbl0Gk5QuWy0m
8J6kStETiz2t5q3lhkUmInams7s+bw4LKlGTW8VZ8ckVE8ofxAj3tf/B0z98XICJSd0r7aiYfaDq
S8LS7SVU8TD++eucF0GiVtssJaa+tggr8XGI4Od91Fo1xbprfT7SJk8jv112H/lUPwaXXcle9iRU
36llt0DEdP7QJAr0Gf1oLGo0ghRYRh7VxEoh6hj5BbTNWLkcyFf1v84lm/b4azbN2dDrBDe4oo82
RXY51xrD3mrI6lVu316e8+ZVp1UTBj4TBGy0h1WR5qQ3lbH0XreQZY+PN71tU/aidrhXzSRWFZmo
gT2zjQLLrh/g68zvj4GR2Br4A4WQTIh+KvxFCCSopokfY5sEnLix0ipoECdKmU/WTHi4z+aDXXle
vzZDnIVdfy7c9F/JWIxYg+pUt0KF3I/faU/M658qPFwk2/5GMtNcSRGQ5E5x/q2hmkaSij1nY82U
snZgqO/1S5kZRjTE9fTcHB2Syv8h87Fw3U9Bu1kPJ6hoCWDQJCHbxfGV8W6TgqBgei8Z7w28MTcp
P9tjX4Tx9fHoOU0pm/cdIvPPHEVwRhb34s46JRWUZ0U9brZOFfTVQQfmqkUGjgMfVhMWNsG0etpc
GD9l0zUlJScGVWwwVL2ESs5VpxArdsLnon+PZ+gvzVhCDkq5X4SyovRjCKNju0yThnUcZp6uVcef
BF/Y+DpEoBX77lchzrcQW+0mGjNs54NeU00tQiOKcUNImK3lOpZ3eYvyWcnxC0RkuctRTaL0zJws
By+qnBTD1B5SJVPhFt5wAsfvGx5vlG5m2ieBGF5aBNlbIeobUAQWQSkPulw5V6LMHRcAhl5h7vNO
tUlpFkgGdBylYnD1RmbId62nWDOc/pxBROnsy8R5fWtdsgIeZMsm1h82JxubaDXBZm9X1Lp9jprQ
KsdFi6VuaD/LiwtqhTh+fQ9oNcgPaAtvbPjoBDrW4RBgmAPKsxgldhgrywYFPCONmcYuiM8pX5bl
NK/uZ+vwaD1NsCEEow0t8kCvkJ2G+42EmLig6TseEaCf7CZdcL0ztK7RFtDmgz1fbVa8YrSGWJ42
HdUObEAeyEFn+Scpxy0oW8BsjPtxgr/ZMJPXot1nHOptGqgzxOtrBLPJjwOTxGY+3tK7IgCBbEI+
yw47O/dxR/2rcUdV8VCy9kcSMLoTOOGnLZuv++jK7ldOMO1Cbrsf34UWKCgUcYV/QHXXl9MgKX2q
e3g4XATThho+pWf/4K8AFT+XnaTXE23NyRjhp4xl+5qZcRPFDT6kKsrqJeheZ39AkU9YDKJQpXpW
VKLB454Sp6JO6jAv5R/X0DbK3MgGkNP0Yo4hREysjqfRSD5NS2h5UW0HUVg18Eap/t3bOfbo4MX0
NIHpOmkZT8PV/VzAa4HvMcX/lcM6Nad+/ZfSOwAVV69Ac1+dzAK3/ZW3/3Ay/KDFB9n/tYxPtnkf
6vOUkbMDgjrM40P4kUBBc2WvD4ToqKDrIxDWMfWEwlOVLYMxXsqz/E3+PL865Uy39t9CX0gRqB+H
e6sPZ+k4GZKeDOfZftdH0dU/xKzOJN7y3FAqxnX1jwNi5UvdiufHrmos/2fbPV00hZD07nJdNYNO
8868nNaQ0zaa2jPL6r22X6+1OPLQ3qBvYWkNO0XBoMapN4WldLgmW4hoNoxAy6Zwf1Q886LcYLKA
jTqHgU4wg9svP/xPXdYhEDoZp3VpbiHRtrbFh02Z1kd6tRjAjjW8G5hS3lxboYuKgecYpKjsd4cD
WK8hHbDrTb7IqQQ3dwKwUbyR0x/PHbTpmft//Z/kxcpNKqAH6DietatQP+z1O09EqGRsSDeCV0yD
tMWZ3bS78Ll8gK6D39gDAMr3hzKEuxoMUZadwAzvJjTDKunhQxxx6ayJah6YfN9BifWpiQ7MDhKR
0EcV3C9PGqdn9CxPNSJ9MsQisPLPI6w9A20kgnzo+T6jRcG1BhcOdECfZgjM9EXcpciJzd5KOYJH
lMbaP16MFQFkbU2sJi7PeSGgswprCjNzCWHhn8/6TqYrCiW8I7S3uItx9R0dRQyK1h/9Q5vdAhZ+
KwPdrFZHCnjCzp+4cLn8cjsiA/GUsERBx5PtAJzFt+IECqg6fvbHgWhaNkoirsr/93HC2wYEQ9KU
+dvUS/+9EXaIZr+ZsONjNfGlCXtdpCKjKWAEhWyPR3MOk5PIjfP6kqqU1UaIAIcMFPzG56zuBKYb
VbgB7uapoAmeOWHcUdPPqFJKdZX09PpV2Emc5wED3J0aQbC0vco0OJp3dzUdjQFCDwAtmigAb3VM
JvPdZ+DRH1D5NmWO6ELQo7r3Td1NXjpaDSlatU8PmwSa+/aMODpZ41F5DBQBwIiqlGSdPyE3Tgf6
ie64OmcB56C3z0MNJS8DhVQ860O52OomKzHPcCOA3UaB7MMckDuXd2WvyMnlAcH2sJgd7j8ywpHb
3Zs9OjHq8CgpLrEilo1jOFMO9WDtPCWOS4kEFPPcGJNvDhSezmui12TI2jsOi41hv8s3MDBT8Fdp
/W9DSv79C8PKp6RxeM8swGbL2F1pmvjAHu+BTSnC/C4xPnZRv77QelkTIVVqDH7wNjYv2Qev0kwM
cC+VcOshSeniet90WyHIVSzJBEQphBKGg+I8OpqLkv8BWlEBgvmvShR7l/7x83gRgiX7aicYaOoZ
C7qkUDwRaKtVruNem7AxiIdWHuHnIcOZPTuvTnOcv0UTULQgTUC/8B7pP5V6MKCa+B3F5Fm//NkI
QrkF5gN29hd3/dozGP5JLqS8b3IxHm4iXtadXS2ypGHusV1sw12Re+nztihP0eICtQX9nP5bzvwm
SnWYZGErPJu3N5c4MI4nyPAEFcG6a/B8L0wTXsaXrVkgZMGH0kizxDNs+teNuTakC7B4EaNjtmjx
+JNVPV2m/KymZ/N8ED85No4KxuHahwRI8sZJEkVJRZBouQ+HI3U6Hnegr8P67oroo8F/0b3Qn9N4
KgPLUouUFZbmjIKpeOX3Nf8mpNvLgwH0rh1xBAHObPOB97xNdDuUNicJI6Kv7mFcZDy6/Zhw7fQG
WdjgN72WQuKMw/K9OIalbMASOtn84BEcNYkPjlAN0koWOdEMEvUfyxDwRpKZkwguCGkOmr5xm7Hb
JrchaWbzPf1NiKOcKSxCj6ALqRXe9g/zJOzIV5m3iMeOqmLRX3rds2q4xQ4AeNsifrnC/Pz/5GgY
WVuYg3GhKz/16HnyhrIOhjL9Q8yJOONJ7Q1kXtquhngmzd5ON6sD1DDShccXMf6+tombMqRfPzzw
7Mwnu5b0uHWZlRz6EWxoj+76fW8Fis9ARYAklCMv3bnPfpEzVzYpMy0g/nFguegRvLc6n9/yauBe
gtYg0g/fJXJ4ahPADF0YJ/aOjrtpe1n0D8A7HJ763FAzPamq/xwGZ26I0HtMg19EkuZd6vZojfhL
Q5QDWdUe3nCNuwsQZ8TwDR+x8GcxMuVh5EOvbeaovhvRxnJ0qXijioW6bLx+u8lRAiAtN1tRdsRR
RTe4W8njRTVwBImPN8q0IeL02m870PBBx+TTZUEX1ElkSJsDWMYGBprWh6ZJ//AP/36Ci3LZTN1M
oLONGAZ7He5WgAw1nVHS46PvYjZSX55617dpqkXbrqgbwT2nLEEATeZzeAGxaCtIlINY0C/LjKFo
XQqjspbt+BqMccdKui7Jwul4TTN2zFH6D9OHe+iqjK0KdEhBgnU2a3SmV15cetD/qFakn5cMCVQm
9TowgyN9tGj1JTlg1QRYnf7spBucJE6ranpIx9TlQPECMLe4hUxK4mvkQo/X+AVvZ4+jvIUySdf8
EZrqcNyz+Q0RBrsupmgE133F6BQL7K4cCgpOGf4zJI3UEqKeLRytVtK/22arhUgyh1GTzV+Qqc/I
f2HOt8F5rKeW5b9lZzi+pF7mJ+NpqZmUnqREFyukz6mgmkdmwYsthOmS2T683ZFTBREfj4nd9a9S
s2wHuBRSXu1t8onGn6V4+1L6+bRyvPDWPazQGdgZF1mfYyVjhU5Zw4Kmv04BEyBu3iV+0wkcaTDU
7A5+ikP5jnoUWdYQyXcYgxlsQd72jCa/8j2awSNTW8DBDuVHemZeqz8CBOdQcK1QyGLLuPSrshyv
RUW8aPOJuKI2NJqNuLCHRq8gX4QyREQ0hoXR4aXKpJK5CNFhK7kzzvzQQhafehy2IFZAo82w2MFv
J9fGXPFCFLiWhxNJBNL33gw32qZ328RaKX36nHQlwPyTWjEnpuJhgnACYRTbsN1tt38ki3u+L3R+
5tmXEppWgNdpX2s7BTnACjxWptopUDPjHgMsn+hfcHJ4OtILV0hfpv1if3rfCdIWcOuP+4ceHMsO
hgcURKGXkLw9E944qAIJbGSoHohMy19Hi/gxIsYrOQ8/hvW5spY9KsfcnX2kYcvjOFzque6f9wrl
DHWOR3bLUua9Wvu81wZX7faSernB0tpCA9YmjvhsaTArHx3bzWzFcYOTxYR5gCehaqKc3EbxkJuF
ZrfcWXYjOGytqI4UvtZX9xpTnF/iMfY7NY0zZDP65n1khiz/+Wqtrsk0zrO6VNKpx0giHfUeyPWf
KeBCoOe3CuViLorkDNLGWwRk5SJGRXXQYGt7JNnbcPf7Gk8h0JCHt9UgNZaSAmRjJfCcupe086s5
F7mHgH9kodIBdRhEimNgoevPpA/sk9qjmNfuez9ij/lyerbMlYVSMAb3bkwWsM6XO41EnWu8ZRlH
px4bpaVswxsdZMgmuhCfvOupzn/eQ/J80uENoB3MQfE10XQHi3ZOULcMEhCisMVD+//HNTVe1Scn
Iq+PNNmKhJ+M9Xdcnd1sTTWneudFEnKJhuSNP/hXH9A7yvdFZJV+GEbepLZTkQTszevSKj1qEMFf
9soDL6KzlIw84+YhR0ZUgB+RIpGyce29WRfaBCHQdvXWC+kfLzfBNYREXK7gMKibtUwm4Q6rgViY
wFQQaPOnQrAaqp8hTnDkwiXZyttkP1P+RftwTivTEOFrbyLbxZaN1fVisdXwL88Mo4QHMXesp/nQ
ZRXhbu42mMeILADBhfCt1LYMizVhS068qJe6/OfDN9fVBebwHLMGH8qgBGnox9GTejA05rXK4X5e
oFiRsFhLNd/3y5Maif4v/Tryx/MMG0DIKPKSyqfBwYF0O4DHp+x3f2JOnCZrLDgPAYBuJYWvJcF/
nWggrWDz/02fmWHEQP+J6YnuqiHgcE6fqJsu2x816q/dxzL8JFI7rF/KJ0uJ+5veyBbZoHIIzCSi
7oRaEE6dyJyG4cceJtr2Rn5r9H3kdT6Pa3+m8DxN/YHrBZD/ODdiJGGT4s5Bo0+aySabnjEmcvo5
B39lC6EtlG4yJdmvquQhmPFSE0P4Gcfb6ISbjFcavJnnhBqmezD2mAv1NA+Adfea+ESfERiM/MfN
tjwt0if/yiOXwjTlTHA0yEH1ZZkgwTXf34zExHHPeTff0hQCE5iyrdlrZeR6+4x26fxjV/nKc2qL
K/OZ8y8dFJ0lSppjKysJIeeMaYjbuKtbHFtzH5kLN40puZnuaFa7D//MRW6kglr1OZeK8dG/IN8a
aIVzTqbmkE8AzjaasCAhqKjoDtDWBXV0YiN05siAKNISuZ1Sxf6u4N/RZDuROZKPX4cRGnl3GrES
PXrcGTXvWEH+iKUYD2k9GDPivfXz9M8/9IfOQT/qyYgSoxeFpD/y326TKpJrfP5FbVfGslZkDzVF
ZQvOWqP3yIV1k5fRnCkh/+zkofm+sy878m/Npi+jE1YoYIs7Kb5b2Dwsfh0J+OL7XZmVHbdFLS4p
IdsJjWYwePuTe/8pGM9qKwIEw1YX7ZAZ/ur/+Hd3lfesW34CgbpObvv6SputRVPrM0SRMitXER1h
S9DmPGig6uw+8U2ljzipQRuGdaftHygNiNd3eZ4x3LseVzqQabXHbiEtx6BVqqY/svENBk08x7Uh
tiaYS6+HAz45v9FJbQ18unbqgtzrEE3a3HnNsJZ3lt4d6clEKxWeI+Pj00ihYDY4uxkGisGP7JVQ
R0lI+zTjis7cStEuHpqk8xm69DyUUPmY4nRnDtdEwFz5gh0k1Apj4MQEogP+qnMP3ONYHEX/waFB
CyDEFJpq+/j8hLNlw6u6ogyQbdAbw9p4/Rre5sKE+Za6owJgdM6oc0Ldr1wWgr5TpXQoS1kimkvm
rwgdL6ZfDzUPdZQnl8/ZJTDNbzraiJKvh9jVZ5ZLWuXZlvEyJX9xDnMJpupQVGGti2a4g3f4ow38
RfVhEK0VPZAc4R83vMamC/S+H7cthXQS9/9IGJBdyUahLemVh38K7wB6ci/3n39/9EaLW3Jc2yww
FhEAgBZ8v3d80iIiz5zSM501DJCeu0dubY/8RzNevQyAGYkeGVpZdiMTMxTMAxyU/qvoZ6lGvSYO
WIl0d6ZikbFAddQATwuRoPa8C458mctSIXsL16TKzrZbE7FN9ZUsdZkvbXdWk1rNoID1IfdTg3m0
W49T+6MjE5Mukr7aoGt4vxRssw82HCgWnWH26YxNUrXQ/ZQNMZaLe7KAT+Zk/8jtbWYR+ENbygFN
O1Sz8FKeKjkDxs60mf7pX0iuaNZB7CiXOXQ1/kOq6EFZT1nhp7niLfaROG1su/h0JG80JrybKZsl
rNhhcvWJPxhmlkvqWJjk7K1V+CcY8JNooJtwF+wEKgrPiRDPTKU5nmWwTzcDr1spdIBOB8+6+D7p
tQyxlKRw5vKfuCaOW5dOKH8DDeYSrlukg8mNq3fFqzHYND+VbWNKRqhHzg9CWBABYe/QCVAyPYs5
qOmbttRT3zNDjPx6aYO+UZc+H5eg2yoW+Z4qZNZ4JQ05ECPcSat6TyWVIbwaVJIZL/GqoLRL0Z1L
uayTpzfSLltkXv4sQ3WFplhn0qE4dSEBHVQut+oSHeCJDjW7fjg8RmRwYSVIFBzUr0d8Jwj8Ep8V
FPI8uSxlbg/60qFiZA6tHIboCYWeV/NGSlOD6ArLHF6TFOoANCpSTQGVaGuu8+z8qdU25R4/n0dT
1cV68Nwqg4a9dsi1jJahDVqZiB3SyDfu4e9SyZB7YPrkgAe07ynQeGQnXe4gJhrne9yBNgkQ9H8v
0XF4pQ534l1GFuGzRMqfL8oaSw56u4/lu2PIZzp4QQLne4aIHjMVRZFkEalA2pDUu8P7/uTcHPp7
tYmEiXNU1lfUlVsZk9kB4v/OqDemP9XqNStiSz1RjgtKgV7DdSLX9cgwOm5wKMwFP8LJWrJ1JUuo
hQviHGmIfjv+s+R/iIqxQ4dXX7I8fpOZ97E2VPXWqREVhtkPrW/wuDX5/ErCpZthIsmozphkgP4G
LwYh0MwNBZ3Msxa23eFYu/sahVMFrZctYe4Wphh2lPUOr6NeNmRnwoljORhis5KFL5v+PvxZ3C3y
ak0GJmuXoAm1c7hZGm19S97hNUKml8UeKr2UyXHi/stuSCdoHwUTNEr1deOhS6QqXHKq02txrYfv
XKgveLWNsWnpePM3ggkN862/RCxzoQZztcpNiU1LPxcuPNyHLI+oIyCfG8dmR/eXapLPNB95GePy
hA6rih5+pvHFAWv/7Zr6vF38PblHwfvyp/D3zMJYgUi5vgEAv2ICYoyycSj53Mn+UhIr2SBKAUOA
rSNXF6wGdGuAM70Sb9CUJF00ustSPWozZYCCSkf7jeY7tgE4w4taDCNfN2ZnQdFrEpeGi62hQJ0c
hNOXAn7DPPS4GJsCdixvBKoOjo8VEreZ7FU3oi8QUtDTXWFgtyvSJ+N2t8dzqXM1NokmDoUyNATU
aHHn5eh5isfCfohhGYRqDJEaEiWZTapEmahe0tuuRsYh72t4w9nEiFXKznoCxd6h6B/LmA/IePZn
mmICtAGBTDHaX4LjLkkmQO7AsB8omcAz1GjcEiVUjZAO4mWI6wlKtUGxGBKp/pwPvmO6UXQHEIl3
hAjLMKsWhKAxIIsaKJU2MXGVoEAaTgOUkpyAUQps5owKhODyc+1mewZ1hHAIoVUK6pbWQZbT0fF+
JV9cfBzzwsyYfJXGzCS1SM6m3+qtQjAVaLL/Y3Nob3if12T2VmsUvV+ViZBCm26oLwsu8ZGI1Hjh
PMH5L1xSwhsWbTQNWdv36jEM+Iq+m0HCZHuCoZas7UjuDJvL0jPuebPETdzDdkWMVFIjwVFZEtzr
2N8tEumUQZa3tbWqixvWHF3Kog6zgQqde2sG3spZFkuetC86eUs9lBCadyKVz9UFMg+v4T6gd020
jCIIlGXv3nqtapOKfNOBwVILFrWu+7Ie/vxn0E273YqUTzIhicL128J770yzc61dBnxaB+hJJCSd
1Tf8fvYurI0MOlvYe/zMUhwJARHBnP6EPa0NcWx9paAvv6euSZOWW92jVmGc1BCJc+Kw4iY2E9UV
xJbnSJKwx/6A8Rq7Mo6hXkunV/IGLFOIGF9S/FXbZNoVHL4H/cntJ8vS2pSdLphQArZO7PZc3bn0
sdcecDKnnk1LnnCz02182j0VTg8f1wsw3+xxt8veSMWGBesUWavPP4MU5JWWTYioYQk7EAXUBGgo
yzvB2DMo40tpMNz5R3F4x8w7+kYc96DY2S7AjTyhusHRaad0HTItVzSrlF6KtuH1HSc7qSYBgsNz
ChMU/FvkGPEeEjalYgTWxDx4xiaN5MVu+sKTsDvfiKHjJBshgwKwIkEPSJS2fd7LQitrFKbhL12p
3tEWAk9JPxKrFuhpS1S0PBI6K9tEG7bCYfizDKnEDchbJ7WakqfR/PeppUQVVFaAympogef9s+Le
PKZfDbmvkZyy9hMJfpeHExpSZmXkGM1uDIRUcB4nu/RC6mn4omG3kG+rWaPikNnmv7om3uE3w4x2
lVRaKXNYCO22x7bfBewHRF1SQ9UhQE4UTAHJ9G2nxeHOf9PJQLdbGFe2evn82fZHuZxIuBtC4v8i
JxP1VPMI7GQXKbiWISbC3JRzTbMqFtAm6ys0HXUWSwG8aSKuoxbB8wNTNjkKJqAL2t0AbJP52NPf
Z4kgmXf6UPf4ooQxdrKkEkc0GFW004k0eA1A3NnXkcJji9yRWTGRdSPIsg8zWYURtuqtDlVnK2ER
7+fmWcq26NXP+bem4BVn6waQhOc49COBM0HdxtRo6iu0Ifhf8pCCUrMJvdQIQVEOJYQBy5/z10Wz
sAUPbMA3a3mwRVdk+XMxZOItJCrkCEzmLjYBgIT44/7ZMCK5JyAayu/xoRrg9Op9pvLS0sEfxngv
70wwEKHYLRZbnDhKhcjcx7eJPak9Ic++c/u3L4ZcifXavaKgw6MbI2LgXomYEhCh6rha/obgJ3R+
9hDhgGPg7xlCam0tXjp6ntITjSFifPaJ7ep0LFbahuPIWlckZD/cFDpZNlsGOmiIznE+bl8Yxk9g
waK0oy38zeVvdFOrlt0EA7ZpYdE+3RDt5MR30H+e539VgOzmIdw932828lq2q8Q3HYjHVGjAnUoy
MUepS3Zn2KsT+Jh0Q2kCHz7FxYwGhkUfl/QC8EQEwSQWAvFVK5Y0vJuQOaZ3Fs60lyiGXPQ0xEUB
uWwU0SBSe3e3xoOt87MD9kajo+cl4Ot6zsVjoZ/XAGS1KqntbzCjktbmgfQYbD8njUaOrLodHPon
z5HyCCLjTdJ4+/FFHaBCZ13c5flAxMIfiB8BuctDDdmdujSWJdgfMMpK8L9nyHpcyADuzZrEGChf
Dt6Sr1S/4/GWJyqtqQ4G3U3EUTXUeN64ZipYAFu4myQAVTCVB6K+FuzN9BdoXz8RRyh7bY6Owavr
6sbSTOWnPuFzSiVOOINuMcuQ5d++UUfkWlshezIdpvrck16ir2024GS423N04ssIQvxJzia+irW3
D9u7sMFOr18Ro6Ax7pGXLyx/1WU3nQ2m1RVRtpG4Zap7+uu1B4wbeLpUbruSO8W1lpN6Mf9+fWIH
bvtuQw2jtvvzjctb5ryHm28cWo9STSosKeqwBjeks/aATOJ+r7KsVKO5IvliOyiSH0RGyvWzFfeZ
jImYBEJlojARolpOJudXZYBDqGZGxcpT812h3dDmG+WIebPZ2KnG1tXh+6I6tSBCsZQeuMg2s+xn
t/udZDEHjOhyRczW1EPIDc95eGP/2LF6kk2dG7ZnWWkQo2Ic6sYHxAS1k9vafBF5tyqHDfzgtlrD
Si7mXXW7fZs3TG2EeR+PvHmbZHbxw/lOz4W7eh+XJYWtPotjD2OFo4ItULaCBwJTlppPq40h+O4L
Kitg2CZ22bEarlL4EAF6+78/VI3tjBrlAFVEXyT8S77IHsDrft5XLFEEIoDYRhXC5O4/b+ZfV+XD
UhyyQ+MTXVUTSPm9l7mIhgjPpIOnd045LqdV7+aVa9iUjA46+xG+p2r0htUBtA3OpDD1Y3DgyWEa
0nsGdU8p8gn9AP/VVkfwug7ywUrthsDRHwYjhqIRexQuL3gF09wZj8xFROO/saS2eXgw2Nv9kL47
X7U3ydk8xfuPBCzJPefmZThjCxFyR7eOepyjXrqTAmKmLxEMDn09UcHe5R0pCgdDK0kwWeka6qVo
jSc1DKg3Jd3dB9N++67Z8/TdKZRZV6x1qdcMP1KgIUs5CBe/02rA0c65TXm/7xwebIBbgLEQXY0E
QZEMTfxaF8G083X3vyGWFFOY+Ci6qBkDahTvDQIPNLQX/9ZQAnMpSTgx9d4ryOj1GTJFrCMUCgOH
qeA5TsGH8dgHcc4d20rx1gYArJm3l4DctnPVFHTJcEUqT7+tWiXuhhLdSd2j6SU6kShaUPl4uItr
rFlEqBYoMHI6l4zNaX0RTXzU2s2N8Ml3nZ9MzNc9Kq8BP0w8oNbLonAYg20Mbg/YSQ2ItKtWc6Mg
F1AmW3bIHDZEjczcCafjbasqw/qhXivdCr5yj2lCk1/XlFInF7nPdaB4zmKABp7m/9/oMryWisRw
JrwwwXRCQt+axAFysyxvtInfMPFaSeW6prxII8nTfv9WIlKIP23KPjjCXe7ic26cLzUImUaEG4Mi
EBZx14WFlyi8wthQuJefANOh49i9sIdL0aFAODYyRfEcFosvJUtsh4qlIPBm0FgHIg+fslGpQ4zN
Be4NWEJesWnQukCwAsCZWqWP6QD1JGNuX86HBJpZNKjDj5k46Ex5F2rhyPE9+qeIGKLbHz/w7uyc
Na09nmmp6WxAqOwnwg321wFl+EBr+QXMnKAUABlccy8U3bqiUSHOokWiAIodmHqhYFSBK6rklzlm
f5d8xBxGJX4hKESZYJS2GVmgA1HhCTlGHKATVlECu5KyqRZVGnBlPt+7dbELrSjb7+oSBgoWZpgd
e3hssxxGhWaJl6G2dj6HnKTPnhKqIjmGQhJBp7mPesjxkuEoc+CRKvdoXaxGltm4nLxg/KxAR7a1
AlpY3N3QaC2E7Yz+jtBUqfRS106u6uG6Dei/rzxi3GT/uZCpB/rhwNZovCtwB3MiSwVhCfjN6OlU
tFi9NVVleQ+Q2E2BzP9dqEDWad9Whua8/7xuCrXpepoQ4rdeLohqmT87y3bcTKfi7cQRtmRWxO9l
h5pAz9CtxR9nESaXclYfH1b/W4MgsgCEudn1JoCu5UCEQuOWAwSrKQvCmYh0Pod6nMUzc/IGiOC5
m3ibS0nJYXP0pd+3XvvQpPu/dG9V6LTvnb/PCZVNmkt+/O005YSS6OF5VUGOyAjQcemYfO96K3n0
6RZY7yo9ueCvtCc7hOKlRo21kwk/56/JbevLldJvMMKVjRCrV4sAhXswDRKZ+sXUad9AUGldjG3l
Ay8zS2vYC3L8HwXmkUxiS05G07HJXe0XBhf2YOziNaez9wo6S4C6amkf1biCxx5lzpk7mIg/VkTw
PxHeJ+SrGWIFe35BwyYrR0flmPSRPYRFPx0IraJ1ypy5kmCEkOKRlcjMwEMfp5idS7eAey11GqN+
lNE4kfB/diPwpO4A+ylsEZ8bIHyp0vvdvxox3jhuK0fKdxTpeRRY2J4jwShAkP4hFrWutM1eMtG/
gZ1s6wzRR1Ndo7Kz8iDqVM03WQbNBP5w2TQQnYBBX1S3wrhP5rFbLxBlLLK0lh8vhBqNNmnfr7ht
oyIylWPoFB4B/yQpYlquvfqQ0UAIKhoTUUPd8gMP0HR0KX3s+e6LRbVPfAc4M3Nt+1o78Bx7e/8f
Dg9LUOwhB4C53jHkAe3ENRj1XZA1htCPKqUGH28JSpy5ESNg5OxJImscwf+1gHNXokGJmbfXTA+n
FDENvmc0LMiO5+YD90I+hOWX5WGYn9WDlemRgc40p6mvsM/AmranCa8sg4lkev73zQCDyDsiqGoq
4u/3xoFBnstECzjmIijrQIZ8uWh7G0n0lAup79Y/mCXhcw4f0vrDRj+JkvpGkKlYxyvzQPcGwKow
LZBhX91xqgA2hWu2FdEeEKDQ/Eg5L9zK7JOW+3aVOFUjvSkA9q85Jwek5YdqddWbgpx5nOgmQRz3
oHWKgXT58QtaSnp8/iZP0LIZPGasmil0+Wojs8YJzg3qSvNAQ+uLrpDQIl2KVnzbOWIh9QJ5VJNz
4Mt2rT2Ll0TMBajoMEWvCZQfJ0S+UQZWl9iIDFJuLoU7EjkuCBpakL/QzTzf/Og+r2x11qRFyNIV
3+QQberE6Y/G5RSJtPOt0HF1QgKzMqWCweYcExGR/tYil/HMGrAhFQuYEpJ1yMgREiPI+JWH+b/k
/ockJvvExDGUlgkPcJwhoyOWCMu4djsKsBCu/ztLSFD1f5aDtABnNKs0lR6nbWOSc9+iNVka36g/
AgstPOhMkadfhwqiXoXnSB2QVi4RHeQGkP6pGbS4w/C/DNGJbfMefPyhCD95gLY4oCckFMR+8ZCh
lIrzdtKxNnxOMh8uG2v2j1RYJJixx1NUzHsvgvwtY5F6r32mc13vnYeNVDhvgX95zM1/QWatTl0z
7r0h50lktUKrMHLvlgJECVKGY2oXk5ALN950W7rdCtIQooXxaip0I5aPeoy3cByvI2e0i5eHJyVK
1nfYgCEZ96djat4vH4qE6uTFkAkmbpSzsNzJCnuQ881YOda122u5XvQZVhtF7ugQOMpWdSR2bM6I
2v1RqYDua371Yna7yH6i8mj/sJmalA0EYCWxQklgfoJhjfDsfuLp05UZ/rLyGxhKIwW40q2eO7TY
Po/H6Cj+xqA0X/C4D8KY3x2iZgsApsW0Wnkkfc6skesSb7Lj72ofoEdIMVG6sr6tG790IWyxnJ9r
1P+mPL+8nr7E2yVL58+ucSz9AlF36zRRtxWYIg0vHN9D4I0cGz8jvmnSN2ZkGGXTEVYAsDxVNBo1
kG/El/cmRPlrWYm57pyLYD66kt36jslMmycZHLn2jOp2kxIG4oc1v0VhXNeU9v1RzYZrOKJLzULA
+Lxnr/gIP0R9q4AxlQ1D2zUY6pZIhav3XxKcs4hqrNGS/tIaqCstH7fZht6rs8/mVs2fQYxt5Jn6
JGxOBqn8oESeNGK559doiTmo7eMWhAZ94+mlaBeCM3GaxtmeHq6LpzIGZmG47JU+tymyMWR4eltP
1Ee+A5OH6l+z3NIzA49HdliEte+oJHu78kxQGQMKKN5hF2iR1zUGFEVnVFjg9bOMFdhbUf1VrfvH
viyQB651Q7KDhrJaAuVpbCRD8JXiFYYs6yoSWmOtu6hSjZTluHnD+ZzbXxg/k7Ds4KHF/Uiu1590
PJCT3Vis7w2CuNoE5+QOGbR2dTw2LmJGfngYexV2j0afKhhv59JBIYScg6V0SS/18F6yulaNVBy/
b6p09QItryPxwFj7K5I6+vyApyScEH5ih33+bU4np0fhI+c5AE+TrU3HeUrZop0Df2n/IPtaCONH
jknYns62fdLiLsg2EWIL6ILYEjN/l6hi/SoBulbY0OfEjte5mfoXFDUnapvAX9ovXBA2prdeh9HO
s/aIToa3wjbra9laWX/l1koy3uR9l6NlC0TpBLi4cFqwNU/+tG4t6fp35YgyNHZuoUM9YjTTuTb6
gw+w63HSJPq11ayESKeoHW0nOcL2AnuwCPB1H51FhCHixONvgu4R6u3IkbFBPkW894/nyWjWthpU
4tKfUt3sw1jquQOaNSmqzxWMfh8GqMTCKFZJYEUXWowjkcO5w8f8WXKRuj45/ACe2Zl5QoBuee1/
WKyUaphu4DiaZ7pNYP3j/LrRUw6VFPTkaZIlSOYUhRPpD+MkbOWtegZI2dkbSGQcmxHmrVvurWpp
kf3mJXhfagJTceRfYowZ2t9Y9Z/BPQCDFHo0x6a4CEgn0gfGIcQyVlV/dv7/yOT6H5llmUQNPYgI
FKJSEHrSgmWoqRtIz8UFdxg8i15AK4qSOx0rMKOYqk1yLgCjAQA5t17GEK7I4JflC2MaOW/OAbzf
TtIe7V6ExKAycNo+lW08e1EYAaTt3r7ON4rV+gykocbq8Xzvmo+QSJJGNTyJ4mzRrSMBt111O9Q4
QJ5P5cjuDTVvj6wJLTj2kEX5+63gZDKQCxKfu1lGsb8dT9ihWts0kzbUTwUaN79w7V2bBtURD9+p
mY743FbR0x/1dzReVtatMuqF++O7IrEAtILJYnLKZdh68E0Ceudu9RKV9OVBfNvHJTeJnlu0T1RN
VdlqhJC1Tx10Fsqx7EeJked5cUj44UtmENVbQDyH+gTwXCbchKfoRa3H6zV1pKnsU1jWVNsu0pUP
b/baNnIKUBSbJDLFXtXtZ6rrdICiXYq2n55qKaHB0UHE0df+Mfy1olMtkALKsXyfYgGX57VGsYSu
1JaAdHG48N/yDIecOXVv9WWWf8szFci+jA+j2NVn9cmys1oEReI0/3IlC4vZCDJq9A4U2f8+ONwf
K4Ee6VIobgs3pS3PgI0Azyfcau1oslWVTvFftHCGdaiXWFF+K8P95elF+LCtr4d5WwcpO58mmo8Y
JHKk2JpxLzZwWgl+oGGXUvfiU8PE92YVwrw09UyB5PwvNbDr5k1XH0BP+ouFzz5cywMKZTXIoPAu
6hEOahxYLwWjfeQJMBaCa20jtvQvvB6Bxhi5Zdqy4ET5KfkLliSzdFJF8KSKOvzUvGKiSl03Rs6G
1FpvBToWgtmQ8ngLpATaL131T0WeMRxmhLEH/3Oxboriu2JdrXF6PjfuHoT4Iilx6F4A+evpVmnu
CEDUN49NIjPyJ/FKE9ki7W6WMVyS3ghByyI37tzB95esmu80dt6v2apemmQcezFI8kbYVkH9yiy9
u1b8gu4m09PUVg70XPEruJBwUPJwZE16TyO7tFCLSYmSCWVtzZe1MI2Xva/rbREX11gcXrOjRkQG
7RvtRjoCzUkq5NWCLyEwTeNHfof07kP+3FfxZvjdHA4Vpo6gWA4qO8WT3kXQs88Ua/JaVaQfVv0L
8n4UfWqCD9UCrQraC+tUnTDJN1Fs4HdkHVz26agLMeq/7cZQkdDoWYsHDW7Jhrw4UpHJ4pCnA5lA
55Sx8gUibxMmBtVhfB46P2/Du0SgGilY/U3PSxQim1GVq6V33vnR3pdAwYwYm5XAHueEQGLgtr58
wr0d7kmWvyRasW5soJzvGAwiOVRmeL9mTv1IjEVyiS69JwPAw55at8byZ9RV7DsSWQAHXkx6TrZ1
6xooBiIL9IPTFd/XetcS+rbrHL4os/bDMf2QW9VCna+BX1OF5OFZ5cborlNViz4z5kcY5Zw2+qGv
nIJ8sLi0ctX/40wAEn1MMgfT5kq1CRR2hoIRJtm9IBcN+8Ts9W7K2yuOInWptmLh6bowHAW/k6Bo
T9+2EYCbcFkgP0AJuo5PDaiIsGBVdkyq2WV+i6s9tOuPkb+8ODERnZ201GEuNrEO9aJMfFYJkqD5
8Ri5RBCRNTs2rUxLsZBjQ+x5sCJFGU/+CFCeTrCd6+WKHIW6hK7nnSTaRrABi3XzqwvUSd6upaF+
3qSX9siGKdYyCbZ4PXJBDQHqj3wjykJj0K8yXbRZ+GTwdd6N/M3N0ySDX1GPVa47G8CF3GTpFd7g
kKjRSbra6aoqqWfJ7c3Tpk1sKYYyO5pmvOCR2Fz6A1sObk/ehAIguZ9kJzHsETgwKf5+FacjcJgQ
09CaYZBytdiBPqy70E/ljDv2hYRakw2xoLhsRBL7fJSYZn+1XQnJFEBIUJv/In3pPGWExbeWob2D
TV9h+a3Fi+WeZNJs+m1jeCiTDJpCGbmRcwkpC44r1GnsTYI++fQ4TPKf8v1p3REjvlLutKYRSy+H
d9CiqUevJs9xuNvnxPHcf+dW3wRU2iVQsge5vatf37uZrzgZbX709MnoCTzroiXSYCIMRhlSh4u0
BzcqHo4pHn6NAlV0ASZQiqzPCAUwVK2oVKekAS76G+kLHRU+F+eD7ahoPyVto/EgbWph2+/1OzOd
1w868C84dJpaLwuHN//5bfR6+9xZ9CH96DYpEV8o4FHqbzOnIF4qa9/y94AffTtGGL/i3jIEVOpg
SH7bSCxVTioq4E+WgmRzf9hMABCLW30RxxpDmXlORKKJPpeXr2eq7+7KNVz1kv095c5zXXIvqoms
f9RkcpbodDTCBFeVqbFAZu4AEgHKIFm3AKiPVMomHRvqiv3EG+xI1shgLSpG5hUwWvDQgNVAF3bf
ys/nERgDKl8o8dtPgmG1vJKYnyVqFTgtkSm7SQs7Lcn0kDxB5nSkFY9pesHTd8+S7ftURKv9rJC1
n8ghOKQytZCo+8JiqT2BBm7qu8qhhVKzan9HpHVG0xXhzvFr3IivDa+NI0fUYRLQL5IlLCPbuQup
o1+36ztom2fQLrIXhn5qKOoY++7XMXnPZgDsfFvulP06RwG9T5cXSDe6Ez59eUC/TrQGGAnSzW33
2Z6q2/2jrH2aAxwSrndMREk/I2xUUu0WLfFgU1S5BIwx37IUVjCHHJgdMi3b6kG0WIg5J7a6pgvL
nRsqJtHsPVK8pQxyw4N+tscrHrqDiC32awgamNxsclntKIZjI9XvexubRwIayGmEGwQSjoin5zSD
BuO6xwVyvlx2pjakPr4mc24HzaMXA69FAn6PBxWyMGRPxG/4l2Ltx7hCAPf0Utry7P7SsyGwQCIk
CrwCLOQFr4u1rqxJEtxyHrt1rRIbn3+cS6KhfTbq7k9rZL/9kGStvy6hrvuCi7PK11iDIYBcIASK
3TBtaUApJO0QyES7JN8+n5MDkkwruyDyd8X2aeUZh4kRxSrTkRjiWW97OToi56+p23DgKbFM03dC
+J+RmU8hz5I/FcDiZPDhCPdiwMckzjnPIbmzN4P9IS/9QQLtK4GjUCeSfi0VK+27B631g6zHwRgV
VyeD0mZVri1a1bcQkXsUBoyhRydrHE1RVFEXzrW9MbaZUordbkqDW2XWE7k+0nT2Cy0j5UTl9qLk
/KX4C90JLt350oIoyEWnf67XWh7D3YyQtQGAo+Ni1GsWuaJEVLchSbP+l5wA95+wKN/Ymz5DUhtA
2fYbq46Fuo4KmJ2x51a+LIoZBUpJjTEn1ypMXeEFCnUj+g/vrHD5R1zp+t3HCwbufnpI2mfriy+N
QlrXqiQBuZeZtqTiBo6CAwDKo+qWQT9HbFazY1KAD+eDKNjCM+uMelUrRpdhbChlbm8n8LBEO7ta
pbxWZyTKN72hQ0/PcNabjgATwuy4d7y57U8OErCINenQywiZXAaWFkyO9Qdoi9I4i1mUR59yiiV4
EvUGN14AFIPY4EypQAFCAW6KXSYzwWEhWyFjI+oHjsI7TQyCaB3teUeBIi5L3iY7zBwWR6dFe3ar
5ZR32ex3z5qBByVlNO9xGLfUT9n5S7QGID3jFJLn2IklS794e/ssYJZ9CeDk8dUvdnRO3cbcXi1S
xmc7dQiR5bAmcOAMk5aPXE21FVVjcrmN/nb2TBMYSTC2Tb+wNe2L2QN9hIBSc75sQ8NRAJKDtC9E
qvSPd3Hb1ouEYNfrHNv+bHBipptJnPNofveAc7ZhUfhSwo/GiMyXphocySn8th7951U9I/1EeqJ0
ye7fnLvu621XMIAJPh8BnopBl1SwDXxhXCRkegZ6JcCj2DJtojGUJ5Kr0YROc8ojERvxoLc6w37Y
pnOXaXyhV8QLdGUvp4/iyQUaHjJffrJQ8YxP3kGLk3fBKaZcNVnPERLTMtFnSva2RSkZWEVbnVBJ
+p63I+rnoz/3Se1FSI60S53ei4ir91n77CkHdip0fvyuX1D5dE+0I7VhgwI8rJM5lr1ceJYkTi0g
yzYPr2OTiC+aUZRikymegSzJGvIrkmZb1iv00jzxfbYObpbXUElLOB9Iu3fTjyNY62TLm8FX63uW
2A+WMQ0t7un66FNmiToajVUkdzHXxt7AUtc1gbOuaa+EQvr9OT8zDLb70HZ1zrByoqwUNcaK6Uom
lBlp99bUTp2u7Y3tkAhhog6s8gfFXV6Nm8eddp4zbyRJpSTE7qYk9oHvwb3xMRHwbdyp0Bde+qAE
/XIx/BvlZsOpvLKWHMBCLyJCMs697vUQl0VRQrDa5iRymKuoJkL99QE7ivAkv31qruj8wOxaXH7J
JKJMVtanZ2ABraAGK7pVOG8sdNyryHiZw0rr2ANPTyzEjoPwfb9NxqUiPR1GM27d8VWj6ZTHf1Zz
t9ldaIs3VNfg2wFP1szYJTzmiAsB2URRqjVGbYs+3tX4Z7SMeGuLcm/2YxmhizaM5RJXWf0ACSPg
ZzgPbB412n8wkfvdF7mkN2o24+nIR4P/AVIvbWOUE7ObSqGc4ratP+85qMk3cRQOj3MkPhgRQGbx
RpvaWcoN5t4OXEuhXVPk4LMFYpGyHtSBLpuaCNE/kxVJbWe68/qWUraXvWDpwvxDAu+qtzbkfceB
ig2t27nj1W2WRs7mokPOwi0/4j7dOtO2dq41eoljlUzehjKrgKr+goVfnjmi8/wvn/CxlipD1qTH
TrPuzkSlKzf7g5rw/qR593pO7FHsk+epFnewsgqzOrdXMi6k0MyDCoqqpj2lYGEB5JTsm007eaoL
ppzQFbFDDbsPiqMeOalc/CKJN6YTybFGc65vpeU+oJq36s0CYHFXCJRVv1s458iV9Ev/bou+uzYU
itR+unk+Wdv6jonqRcexosuwnNlGcpwQgGM/QLR08bCsGYke9ei/RFsAxfyB+NfV/gNnPVkRHWhS
F+D+Msp0Wf6gZn2vDxBDoxvfNlWkORJ38S5sUxEOeX0AL4fNJr4tafizboLSIlxHOwI9D1rW+HMR
VOvR1CY2laeryxJYb9bQr+BEtlDGAiG4tdh+bjHrC6pSbSRVUK5L/B5bij3GdkQPFpF2hAu5apf3
pHZeGSPwYX5dKMb2r8IhpXlDV6RNI3TzAoQXdn2J9tHZmfeU4MGGh+Rzd9X6fYgrISNNi04AN+Zv
xWAJc2/O5AWxMCxX8Ot7K/cDCA7dcAXDGvyQdZB3e7ar9elYOv7SA9ceQnmdUYxJTacoxSwB+wmI
UtRT6lIU0gXyFRuMFCBwhGkRPUCoSMFfmNAOyHgmLciVsFje+vfGb1xk189DMWxdRS7o+F6T1LYA
I2eYKRyJ6vPD7Ye4DP0xpIyFkbHFW4vIZ0ePlo9EhCLJrGytUbAtoYr25/rkju8h2SsP6wsiVdv8
cG/5YncjKzKR08bkty/bEjkC1tVREg/5AYRsuPvg799tUzvCCrSPfBeSvHsIbnj6aUDbMi8ABTn1
efqBQdMJ7/FyuktPrJ61FTx/eTF2NvxC4XEK87fvkKXk3TxgJ8ZT96TdZiydbr9bU1wwW4SilLa+
bCZPUi1GSKcT336TyKSZnJKOpd0ECDZUaNcw8hSfA8n93FbFlYn7P7uWhZtJ5pbF/no3PRu7WgJA
p/YbvbDk9baNEc9ltsGSL1u3Spq1AWkWqaUIN5GeD8239ZW/S6oUKG5p5L1GTxbAckWM5K2Ld2v5
fYmd4Cp2BYSmyu1oxah06aIb9HentwDscxsip5/NQMva2kkxJ6q/KyOFZ8+5DL0+7qrdCtgSPZlr
0+iSzhQnO5Eg0BybTDGpSGQ+TloCgp+mxJ7beDXFTGHexGvytZq7zmPKk/h60at0GalUFKh4WTwH
JmRVDy7QsFZ/SHo3S+j8neQiLrpFrepsdH5S7+/LvBqJmgj0D3bmUe83zspgjWG/ahgnlJo5/7eV
GKyKV1q9lSv11THgiWQ/nF/tOZ6gjKI3O8ZnNQzZ7DTTPLhbjlJ3xw7z5LecnkpEL4as4P2dbpBn
KbUcsLi9peVTVpudIQixoHzTGMaTGiFRZd1Yv2vSh51GqPc8Vmz1B9Zl4mI9SC+Q7pKO0PFOMbLK
oWcYnNQN30u3eB7d/dV39IMSWduUdNhFoRYOpy9odQy78ERIy+5TgKP8vWlYiJYxoM3P6wA3L+dr
ezIiIJJbQ8TAMiw/sHZ+nUaeoaNxLAlJhljxvwjk+QEVHq9+CN6LxFNaqKLW7Z5u3hwFMF35eLEN
gQfcAYi7INUE6b+ndqNyc39PKZdWlA7HQqHz0tE1/PpBIHbqEZD7dK5mSIqIL2/kEnhVAS2H5J2W
DfQqZZecOO11nOA9Eh/UNKSmStZA06x2Q0sVWHLNX9TY/e2vfd5II2sCP8nCUm4B7pAfF8ByN41h
GUv7gcHqONXebIcaC1r8rMnf0sRMeG70qs+cdGSaMOOsK9vqpGLhho/ySLXnl6lJYwBl53+Z/0Fo
hPc29NfnR4k6a0P9FfWLLOftGrUJ6ASOcFB2UrlzJ3JGlW7p8YXyDJdfUFxhw6XB3I6f7l28t4Uj
gkTB5OCYBQ2KOvC9yo/BaaFo5iRIxMOt7bMghFk5ZtfKbZ+96rChZiNXCu+AUroJY2Qspxc1CZYJ
ilWu8oPmcjKojQNcay1DB79vi4UThMp+yWNgobMXyiE34XqXKtvRTjrS0lj7GzMmYrylr2WomFSg
aw3QzNCljcvIzGuJDr0eDmjTQqTXB2obqhRqci1adJ2QL8/8E/0swRFaNymimzrHRP4pBWDxcxJs
uqMOvcR4SDnMrmJA1plfa9o3xbZT3nXD8yLoIfShOHqZU9d3nAU5RS8Xd+T5Ic76T7jWFGcUHnBJ
fDxkRChGJPRf+l5eI1XJfzC28jsgCMl2pmAoDLWa/A/XpsV3S4PJ6EYFqCEVh02voF7UYQGpg3ZR
6rHfLQLVVP7H9SlMxaPJ55DxEeLG83XrgODDENVVz+0egJGqflXuONxe3kPUyIX+H1gu7VtcSePS
K1fIlHGyfY1lyEEaof10/mxLWX0h/6B/CO+26GLUtngyBzoGYLrQlFq9RjK5DqxqNVKBWpnnxQ76
PehRM/RBgvvwtm9Zg/z2DmijBSbYdbkQDgOH2YOc7GwlecLCdENPQPgsKWLrZF9vX/wORwI/qb45
pu8pWU1uSPdWnYP34mj8sF1Jk6bOPLy8vi0DOEFjyAeqMzQtUDRYHqhFqC5haYtErSDDCUjl0cyQ
fTm8/PyY9Q7t8KTZJLsu5AWe0UvQVGYDD8aNtO3ShdpWjuF/NXPUm8Zdjid9hb4DCJgkv9h/GYW0
WALXFYI+FmpJF5gchylkwC2hsZuiKj7Z/t0XgdHTDOsxw5fNWNAOc2O/zLd8t/z+oRZO/BA7eEfN
tRjBt6mYUHIl9CbJE57T5MOJxqE2LfJfMwyhMKld8xnSdr9q9POxL2scO5XbvmeA/95cd63EH76I
ZIbaIsZAPQVJRJuJxQBLT3NywHRWmeIdwZDgf9EyaOV2iqQokM8ove0QmnTCCkWFLaNZIOY5IClM
EHjKLjNflePMTmyaCRrvMBWhXF1NpaPJPXdIfwN2DvRvvg48XERIuI1W20lZc2s2eodI1o4xNKIz
yvgHwZeYEIZMIONxORZlpLiuK1Xc/9WynUoh5b/v0Er+7tPgb/q9EUSA9sdqd++hEsJAIfIRcvDw
1y0QwihLnFX+N3VH7mMiTTIk2vfg5rzOuaRnlXHPTDcETWcMdE7AN1o359YzS5IhXe9jB3fWRKic
QeCM1vbZu+guTDa+BVH+sOyTTMqnqKgmqpGgZPGwUT2dOgrbb6i0REqLt4N/o80ChSdtEp0vhI57
irk9x7imwT2Agw77UmQXmng/sCfjiwfeBOd67Jo+WPYQWLRKZPaerHwegMwiINo5fKo5vKn5+dql
dUsx4LTsLk+6xXlb3bLEmFnMxet2DaVM48qS5tIKVt697ugYZcU1ITSSuqaamc4bnnYxnyIhkZiV
W3uGKXqEx/dSW7PHepBnQ1PMoRSbq+ZdQZ9cPsFOgKOQ2jmqyH6SRhXj+e6APTDSLtVaanyZ00O+
QGpmsMZePxVqXSzt8G58gNw83xLaMyt8O1WTqhcafai2qT+uo4LIC9RDS1kST4RdholOU8YYMnbh
liXXkVIMwK0b9ycp+Ao0cyyQ2nGYT6TekU0KylKjtjjFoZILFQSLWNUimvjz0l+9pdcIrYN/L/i2
nzpxWoUkmg9RGzglup1N/DpbSfYuxEspgf82fY8fQjgS7J82WS/sh7I8owvSIjeNdhGtBqbH2tsG
D0qNGlWiUmQgwkTbpakUpRssyBaoim7dRfLasUhfx7qd9iWWcjzdgM8iaRFFD/cDaOukQC7KGVBb
FtnMkvS2ffRKba8tfsPGVWBg13mT5mUYQXZSIx6Ih8l0M6zYWPqhyU36nMya4RomaQ7Y7fG6waJJ
mjitRBuTZ5bbPfxMUbpjXhECTE5ybmceNtye0FlaEZBt5bpvlWP9T9yDWyl0Kne+Amft7VK3+e/a
9vkgR3+MtWxBRHrJsY7qBzKLGXQnmOyZ5658WyGhmzYfdVre8qeGxIaglGelm5W35wNRUxl/Mtzd
0B49klpwnK0TXYKCeFXAh/j5lJ8Vsjx3Mkbtn9DK6Awyhc1d4mqw7Y0FPPBHLZsEwYHILLYbC8Rn
XyKT3PEQ9WXilh0bRfsv+3PqrRbXZ0IC3r/bsvCRI75Co3BOF2Q854+xnsr+Gbdolw85FiBNtkT1
4zRnpueN1yX8yPIFhPS20q5Ba/hCaazOQpTixDiejV988HaP9LL8RpsImfm5OjfL7izvO9HCyqaK
fp5wvOJFRqZGvROPNd6Wwczm8O6VmrvAUGDnsKd6AIQNuhnqlLD3agavJlpwnV5BvgGWyzqdF4f2
A/1rUkXJLbVx24Kz815mAGx0uULkAwCt9zhuZ9ENhuoBJyxB1pd4uoglGvI/T8HZk2e+Z9vEyOnl
gItQTsUQN4yidS8AIRAHErYPqkXQjhQwS92QydNmnaaVubFRwJDkBR+5iNeHEgdrL0UIRfA7uDny
laQNjeCqyZXqJxzpl0bLns8aBVNsFmpvuMdhSqPqWnDzSUJSqH7GOTtVPYRQk0AjQKI85/rcUsFc
n4Q1Le8Vji58GqZjkiQhqPp1zun79bYd/LyRF2jLw6QYFL87jGP3lLDqWTjZtLdqZzUY3wUO/npz
hZxx/LWVgn/F8zmJAC3Qvut0Eq1LCABz4BmjXJAmJ6FnBrzVyYGmFR+B2nj2kcE6nHUgJeleNRjj
Eczll9+RXR+6TbYHhhu38k58+9QNpMnZq9kBvrlzJByUNAdMMv+t66LqCEIVUKlAoUxCcE6+Ikpd
VoN6Pg/0n1swnTTsRYWAe408S8wWSL/7+PzVZ2HSBU2ALJ8d7ia8Im3dTpYn2hllPomsh9eqCEvn
mmTF+ptaII39qoZD0+Do4dc3COB0aOwVxKH65vQAu34j7iAyY2Xayb8q5KVJ6sIEJduEAOCPmiki
tegBg7PpSTLGpqDiIldCOotMVt27NCmhA3esxKMwLxiqPkiC1QkAwmOx23qTBlFIkdtkrWK7nxLV
g6KL+CivsEQ6vHVbJuipKBhteClNLHSb5ITSEp+wa13H0AOi0Zr+iwHTuUWJjG7KimLAWdCpvYNo
y2WwCyZfmf6xx93MRlfeWmMJCIjemd6PMNilkC9iG/bcFAUDd0cjd8pbVC/ywS/jY7EVT8NuBFlW
Al+aYiEd/BvnL9p3zDteDXxoe1CjJPE/J7C1fCNIA3CUd4AM9EPvtvk6tTI93Tj0Y6j9F6+HFZVj
vOk4PfsHUtrvy+spHxlRdfP6y51orVHEnSchfTpH9nt7O6boxx+0kY9ZqvGVWvGaxIinaw7D793Y
qvue1bq2x5Tdc32oSeXPla2b7w1p6jqnojGFBiLYKkDD8zCWL1s8FMbCLUoQmQqL1+JSM75ppkSZ
kixkKKbIfCEa5b6Gf7bwL/9pJzLBIRGck8pxKfS2/+SMGOUKX/t8vKtqcvIlDlyPViIIPTUocPFq
IdZkYmBPpLWs1HHkcFgvvTvMsZEjiMroP0K+2h9jW8OOp+a+kXmTWXMgV3lJdqALXcF44QhAQFvd
apU5OMqBLLi7mJOgHesEPD2YE0DcmDxIxbHhDCh6QzDzNbo62HMkEniNrrBA4fbSXy0vfGjwxW2d
87yT70jSzJIZMdz4blWul6QWTcE6ZH7qmKNaBzUhyuTIEFstE8E0ZWYHwWc3E5+FNf3cEQQDbX+f
j69KcrN2L648dwYcjxWzN0V6AOJwd6UY214aLIRpVFpTBeMwBwjYDXwDof1PsNvks+gQRc4aaoxK
74YzpP+C5gIvCdLxuNrUXh7oX9I8qZBdEvRzNDF3H+WyfMhdLA00CM66P3MGk/EIgLk2cbcLZKan
yCLxN2zeacU1VowuICsfZX5baNjomJTXtGoj6GQy9bI9l1ZqosvxwDCEP/Q8hUIEDNA+/uSuIWbK
cubo7oC1OFz+1x/Z+80L10bXv000DRiiO27mnH+6OAVDBjX1022lLIoGV+xp8H6MR6CapoUaqyAv
mMbxhtRXIViSlKD9hjPJ27OpPJQdgRy0jthZD9Hz8N77f+pq6pRHfqVQKXxML5QA1aVLzpF0+Cg5
n5iow+4oi4xXcLJ1wQqVLVyPnajQXXrSoJs0ZvtC1sUSKv6tX9QDvtKwrcV0yji6EJQ7VZPY9Ip/
Zvy7SDPgezM7uZPi/aNYFLRxorFCvZ8+nmivCsfJnheIxNLwueDfU5uMbCVZTqi7QJVUDobTcTJv
Zavc69838SCWgeRp+n8laWumkY4K/V++G1vrjSDyFs761wogMGfs3dWVZVfqzFEmj0+/35XWU0IM
4t/jmHUI3/lPFHwdykAgWqwOg/GJVORcMt/2OmDHfP8ZknAbWAgIGzLENBa7vcMpfOOVPvjMHWH+
vbL3G+sMWPZa0kROroRngfGhayaSYTQV65WMAdB1PEKr/4xmmMF27S1EYdDLH1XTCtlj94WofL8k
W/ravbvaZsxvsIN4Lcjq7lHLT6R0ZKddOwnoK3v6lU4JiTAXXOO3QLPGtMUQ6BAUL0186GW45jhP
MfIQcF6OLx6S93jQW4UvmN/goInpF1kHBsNjojG6yKtiByhbQBB8JQ8HLFrpjrCA5vh8C8OJfNo4
r7m9uYCw15l4gUyVDn/Ny4/ueNOIU+mak9tLVrPU0v0wvRBYfLz+w1oTjfrwhEEjXPXm9XZxSXd+
VBb4jkvISkQPv6U+fwzNJnAQILFXT7othmpPmDKVgOHGlU6/I8G94BQBFfkSru9gJm+3QFg0uJct
GjPlIC9m21z9fZUdr8ivW8taG06bUCTTOHGVqBoqNoi6AefTrJRTH5bkH2nciJu+tu16MONWa2sh
UNQkk1xgiciwCrblMXkCov8T+NdBQaRF+clnfIknZpSXJN4Xo1HDzzVuQq7zVc/h8gtZnmZ2U0O1
Full8sgm3c/DaLmEzgJ/aNF4vbfresw/niQrioU8SQdoE3wL/m3RTddTp15rc8UX6wBjx3yERVE5
zmIxNEmUfCoJ3YN3wA8HMKBLoN6cEiSzGkMDd9TJS7OHOSt5w0x3H6n7eDTd+Wo8HP3BA24jcoXW
A6iRti77UaPKMhqLJj4ROJBD7CvqKgAl2mKkdsLwAQ+gV7Ny0ZKALZn7BZlDgfqBrVKNAaT2OvOm
+6brxsme281QR9ZY29N8Qe/Umj4IeF3liR2FYFKJcFXXiUfRmIoLGP6zbO60YLP2DRxcjrCR8Ehp
SjVN2fVluovTn3C3oMhUKTGIH4LfwwVWddjxPNA7hyVSBvyqg2Vt8uCaEef+asTk9uSOMMr9260z
kmpniLrrlbEYSiJlIVYM4OGFFRd4sKeBV6Dy5j3bL+wM1IN3SB2ma72viMuh67sHDTGdrMfBUoDy
CrsMmlaq4GOHMEWHyIw3XAy1fEqhKlNgd29v96vd244FdIXzq3C3z0Qoe4pP0vSS1m3V+gJd9ChK
tjqJAZ82GEv/nf0Vp/11ly90GBvzsXgUFid4d1cX2dq2CP+hCAGe8u+RBnesyNYO7TwFFAtbSl4f
WZHrgI57Q8op37SNj9UwS30J58H49ilv55/BYh1wHW23t+HM2ASO55NBte+Eg8/2iHP2warpnuYi
fRLMrlmeJzovCGJkGF2n5cSF/PUYzMkKplWZVJ7g6gzweN1wVg6jBgVhtJ4cPo5VckROur4ROzCy
yLCbKwAqKYU5UoG4ko2NCMdpRDir9EtzJURjXbCwZu2YYagRnstNTr71hj61/aLuLV9qZG+eZsWE
G0GC56nRbxGuzRmDDANrIQ9USnVZlTX5m21PYXaR+Bt4r/s9QIllhv58xUwxsDHGd7/jSI75SF4B
ON6Tu06wtzdUv7yob4QLakgN/w7RwCngVez3PCm2f+p6yf8LjJuXRe/oASHpTOjQ+lcZkzj4IrTI
fOj875BGVcG7s48XXjqDKsMlUJV6bB/JLHLdZCc2WbWSqNKWEpTA6eLt5ysqlNAwS4KkZAWhmS1Z
BymRYDxgOcm17g2kkxECX3OwPiuvRLk3uX8TSHO7zx34pBois20kY2n9X3PkQ0xvUT08xmqjLGW8
pXhcqfRwYL/z97uvZnQuFnYzQtHL/l1/EhhLLLUDM2apNC4Wxjx+8tE5iZo+J0UvjqABxjEESPBt
e077cYG2vG9rOgtITKq7TukbAMn8AUpd4Xv+yUIndJy/wpKFzzpns8fWEBZKBzN0J/iKsk/mDV99
uXgy/f24bTldcVuLGn9iWBCxLu12XnkPsi+HVrJOQktH5rZ428X6X7JqYL2WvYIfnBdY1BzarYeH
ClKSTk6flNKVn4qmVWTlrYOIMl69irHWUmH/TD49KJnCOugnTByNUceJy+KMvurF0BsOzFY3NDwo
g9dxGZhzJRO1OHDJwr7TajJxFO7w41yXojgG6BpgNRm36ChOQrChszlo+IVptW6Se0YHS+dI10wJ
odgbB4ZuebckrDGABmBEPHLEKGT7pLERamP9BhzXVqrPTwPTcDUyWSiV4wtLhDOboiGcfqebPWkM
W0MRDPjumTJqHQbT2YnHd/0hiatmgHTYeYxvIci5im0qzRZtRoO/vDLndK2sCKxYNa7BO9j31e0d
6snc2vPkTqze7RXGmU3mTiLXgrJBRLL2+gFAL/MazwRWkK98qX8bbN+mDzyTWAITgLJowN3PJxTB
AwyTU6MAn3MMIRH6u7xVHQq4+NnMI51YIL9vDEGySKc5MVzNPhZFnuq6uL8eHskGwU0KYIS6i7zr
/8UlWPhoA3wkblxOY8mAunT58KHhR/dT1jywsR0mA4bCGE5ItIGGAmTdACyxtZok6xG5uvt9r+iH
Q9KJz94sD4zeQ+o+J7T0LOtDAc5ZpG0+3EFq7399mb4mNewpA7iRjQw4EbVyHQLHbLlvQvGDPwco
RmDNLFPfCfykX7BT+kpFmuRCXIyQK3FFIlSt95odj6V5i2lSKqMwZdcFfMZZ9oB0okSpp7VeLmoG
CE8+75AzM48i9aY+3aiOrKZVSCYfXI8uhXehkfNk88nB2L6vDf4a/kaJx7YjFlCHA67WEyZIDdMv
tgL49+2dTy6PxjENYenL2D597jEhMt7zETlD0yJ8E8QDayS9lFSbhhglv9cWj+AuFMtQKXZN1ty9
X3gdhLmH1y6V0A20et0HjCYIy1+Rvhkv+D/kn31qFV8YBO3BwudhuND9KbzIiSH1NfPtD4cY3wgK
joFntsJXEiMmkB2ylk5xnpUypx1M/S6Jhxdb7ui65HkH803YQVch6ZI+wTOsYRI2AnMos/pLWOLZ
c/m9mSuC5uVGvIJ+aF+SujHtpuBInPIsWDWAsJvXdr0H9+xquLHojh7GAlUpGKMn+TkkWLgIv35q
9NQgVQDsbV8L68hHW1jC4eKYc3/obe97iEiYIb+R97Pjl5s0uP44H7kdPIqdA5+RwjZBqNoNFwgx
r3YIsqDccUM3W3QUk9NQQQeCRLhnmCGbQ8/MS7JiUYboB9uKGnv1KOJv/CQncUU2cgMXZCgAZdjt
2+qrx/ytWBwIZ9pSCwBR3ykH3Sviq1q2EVblQCdxnH3LPBF7rvI27o3UocLGgpS50JPUpgt1m0K4
Gfu3eeKVuLSiiu4/VZTg5g/ymNbv7Efm6aTnGW8VJ5eVJfICYihxEf4jZUW+XAlVPVrMoYp8EQCD
Kf9LqEyR9sZDzbvLvLtTKUpkE92E1NEdL1Ifp4uh3HHig2P4vR1iDpSPlADo+bEKC0eGvMYDbWVK
AkqrJdDS+htg295hENqNe+FEzxwL3hu5UhkwkAoyxpeCvXIcJiyEo+IKcrtPNYq1Vynzb82oS6yR
UzPYt1naeOzA/A2iuHI0qxPpjjFCovXzkALS+kScuJCLW5DdP30oH6d9OEdIDkbcl9rcU8Qjmt5v
wwIIk92p15fbYeSJYZjFs0dZ+pecnpDU+LZ9tLewhScqsh485jlNpdEdXogwo25QaBYbaHNi6sbm
uol6TddOFDS4vyiE2ez+k8YDqvbayd2s6YKGTDsBe5absClEvqvmzg2s2OdQ7EpU7uDHVZhhvBxc
euBW1GqNWffCEYZ/rB1EGY8q9DLEav4M6nrZsHs6CGfb3wRrKqPai6Sb5tAvocU0I1C4JFEwCbjZ
m65U5efGNwAwn48TKGyv8a7xZoj1UsuJT3y22jLM3JomezpU428LuHyEsFrjZX/FDG/EcGMODTOy
U75WF3IL8/6nyiR86iw47otBjNjaZiu6xXmw0wVGaGmJ90eWsRU8JVRZLgNgo+jirb0dyZGn1+UI
7dScenhrfpQtp9Zi81gGxqiPJn62hyaRhmLu5H4r8pq3vT/1uio8uSmDfwItwR5O7jHmMzu4gVh7
ceFZCE/Z1rWSKOXvxn6Xg3RlrEN4vBXt9SVeIXw22ioAHvW28HZ7qXqZkAW5R0Hc6b25pORkNplQ
nGRshzyVYPPS10cwWKSe/61/0t+wYIOCWAURuVdupAgp2Ndldmc8vb31pPZ7FYJPoI4LoWMDWzw+
lK4toOM8ejPXiTK5CpYXrlpCT42zf0dH5vgr325k36yORfdq0J30wio9lfe6RUzdKpiy+O9QTD9h
tpIwTxRzHQaGfVXHDCQYa/xMYa9bqAnTfQ9lCM3wpsAawfIl5+0LGYv8rO++XXAafAvbCX0v0eUK
1TOvYW1ZXKp15Anb9JyBp7d4tRjAI406bUPP/oID5DoQHOowEr+6d3e+aVx17Zvy1wER5WeOmRhc
P2TWgencQcYAj28X+P6E7/BAjrnR6cGpRDSkv5bXuVXfkj4iAWyoyJi5CcF3V5fvwlfeu7JGYw7s
1X+sZ3yoLbhmGce639s3gsVvatJEm3oTRRZ8D15Q8USJ7kjCuQA+C6LXE/Gcb/EcTTpo8LnpvVRa
glgbrPE2vGVwGKrQREiaG17u+Cmgg6l3k5zyKpBmLVdQZNgxgcmfmQ2XP1uZsl0TTd3F+N6/BPLD
haQUIZ7DK2MP+wGxJlVn0BSCOCwBxT5aLqni9/OZZMNmUqmSklTAT3Mo5BvkLqQPwM1kg5icMQhB
z861bB4FDro6qi7c0TWYTl9f19R4it9qD5SrHXVbsQ3n+wAUQzO4g1sTnpqnSgnCzi1udGgC6LzO
4UzrkPgCyqpNz6lsSV1fgRdgV+cuun/Wlh/zzz0t+HqZAuxrjpN5cs4oDqpSi5VGUM4fjDDpmtDD
ZTnxQdD4mwSQd8w5DMKsBRN+b8fXkJ4mvIcdmvW0td0OStqKUDtGYGdVSQlVK8sPRm2/8FSNwyut
Y9TdpU2ZFajlHlKtBeSQXUA1thSAVcHdb25FSXnMuRKgDAEOheGUkKFzwF6H1h93PymroqDZct64
emUKv+yKkLQ5NYqYuloJ+7qIwogRK4B3Dcaf7tBCtU7k51IXAf706AnamGUG3+6qIWpAW0i2weRv
4S9+RdT2wntGANVrLaYcopJVygXE23GxIu5PwrwEKsu0GFdDTXK4EI6TlJTtE/cECOwDWvjIld3g
FpVoOAyXwyoeDMLgGybtK6xjpV/bxfwxJeQ/KOSh++4OCe4tAtnzRNmmhV9aW2OFBw6owDs9MyrY
QubtsXqZbiARnS7PSGyz/Rg5nSlAzBfjDgUxEC3feAxADGu84j8arsPqE3deWFS+EEe6df/3VZB0
5DFbS7R8w68fdB/yXHtRFWGhPgI43XaO1XnXeZQoThU7ikvAqDpQJ+qUBBp2aR/eaJgBlZQeTy77
UMePaCAdPdrYiPJcRri4Fs7VyqkoSDtid4hTjFFoy2Kpac+I+HQ0C+YdcEEzcMS7yRN4a7zs/YAm
HCnL5ER1n7fT3u7FrLfh2Sy2U7B9R+yKvQ+48dFL0RgwEeSsaBYRs3NmY5AawUUxHx6HGHl/das0
BJPH//rLcpzXl9ZkQHBAy2iSsQdNF+C9S2qPhIOohUoUXvxP9czm5ANtQq0PLGj8CK65814lMGGS
p2dLf6AsnAoQCybWCPNam3pP4jepptz8++FWMf24J7wV6sqElp/vPSmu8UDv4JbBQF0zIk9dsmjf
kIANC0Llgh2YvITo8Yydgd2rcbgxIAhsxAU0UwcK7H5B06Xd+BKT2tpmJwOti41tg8tc/9+lv9Gu
AE1B707jrNmFs4lq5MioSFV+lToUpBfQdJ1KRV9iP4I2XqYX2E5TAeexQBbsGNToVDhXjqI3BkzW
M/V1Mrex8YptLQVp4W2ye3SPLKHMbSODnsI9xxxLUPGW13eBmA1pghCJKCQjy7nme8TO0pYATqnO
UFTtAucXQUW3Tvlu0HJbmxv8rXuO1B9ZqD+2LwPMWZgjm0YMJYWRe3sCivSnh2YE0lbz18SefYke
lConTSrnRCyFJrnLgk21amJg/flLi0dIUx4DSLcVUpvhZPtZQLtnb/QfoOvTmUVh2PcEOg1LRMNY
KWJNVYD2wb17x5JubiuKegeVwzGXR2tBlJ2VUUO0zCEjJ2FUEjYQ/nBFuObiZGLydx7PzOSh/G2v
87AdiPFXkqXz7WXLmk3bJIV+4SSN9KlODpHtt4MK2wnuGbyfrk1yTDZEkO2vuzZ5/oHb1svVlCSv
utvdD65JSjbCDYUrEouSkwOLCm8/CJN2BXWK3qAz0VbckyjwB5rpYkwqakE40637HNhGSwrUMgm4
d09eeG4488bc4ckY5wwWi4yEQ+cE/q0UjQj43BrnI5mdKXqDeqKmAjd3FD7/exeG98/klC46LN4x
26rSnjeO00tbL+gAvq7QHOltgwYVOv91aTV7Tv8go5vRZkGmmlaDHXHsXTnieIjzdMzqqz4TEoJm
ERgxHdO8dybkvXjeWQchedMdx7HXNZaIJa2JUPG1EwfsitXfH9DsnQxcE4taIPq+FPu3QTrVh9ih
iMdTy3mhQKqb/MGy9pchJhzkE7rJY9SWczKxg1ioQSGbjxlkVYlQwBAOEoroUvdwmqI76yE6pLnA
MNe8TEbKLeBw2XB8dNaE9kbGenSnB8SmMGmi96yYysmVP7lK1mGHClp4Res+KjmdfkAHWdhgLKMI
gOEuQGeL+leUTAJ38zf4Xhsx+fnuxzVK+xqs1lrPweD672niJh5JXpWHbkjpPROVMC15TuHi+Mw7
usZ1H+uj5krzndIbXNrvFuUOOv2Dvr/qm188wDgenWIgEpPQqEzzEb/Dsj6LIO5ivravqy0EB+Bb
4OwSNlFTUQ+3RorhCeUwgBJ5O18rhzsYAC/xfWYvA8GpSII/r9Caz+DPikeavYkuY2jcgKv8QnB0
Iom0rs+ta8jfHDu55+TAIrixaSkXCkflJGliXfJdK3KRt1dxL8CkY8VD/LBINerC9bD1l5d5GjP0
u/fZqTM9RamyZ6HD2f8iReqVuYvAKA84j/CMl2HN95/WgSXdRDYp19DY68Nxox/yyNCPh3cWsZlh
aakp6rWpZU8F1uRWsjgYsDYCxIOtOGpBxora88TQMkPT5J01BFeHu7MnRBkwQGle1FW1dB9BDaoA
OypTtD7/ge93rqKBO5BLyOnBFW+KmKWmuIsQtWYEmaj9Yt6NbZVq8FLgbw1GUNhM0Ns3t2viMV/S
GvQIw24b3SkVHI8UfdsrrIbV1EVwPdo+8ka/JMwvUXM/mGw/tFX1Q1fvPTeAm1nxT233SWGXOjks
jUoMpnnYxnJnigFcvWd/2PKRFm0UBdt91fGc7ubJokY6q3U70JaCQD2yudpj8dt8TsURV53TD589
BnZrt3h4WSv5bnaZz+5PMOue+COkQAhuQUA1THF60fGJC9WglZeVmvKEhqSR14gsB5rxtIGRODx7
mJvg2P1luQftt6lv6DRSCMDRdMRkyva5sdPWLuysxzEh4hakVD4N3o0Z7aJ/8lIumSZ+dyMZOi8G
bGOYltfWUxYMV09CrZNJmtQpjeQOgxJsvzVjJXhLHxWbulR35a6dPy1IangmiLgiD1/q4Vdth3+T
8RxuUZQSrGQy75wYunY+HYW30Ht70vY8swtDW6x7cLYzd5MOCKodacjCw/F1iEOjbaop3Lj9txHz
zM23/ENrkGe2ASGo9dyAnAHHzeYIhwaX9emAZYXRw08C5vKDR2m8sNDe6D7jtj4CAeUauYyGj5SU
WKJgi3V0+Zsj0U2KZ5PbNfKx8iYiPgd3NsX6MplnoAINJY+XwuYWxLh3/gk4L/Il6uwtMNrHOV+s
UFNkaZ13ItL+/HZazPbCiZk5ksTwfmX5Wuy2BWIn1hlhrypyE478V1eHPEAXeSS5lT++aNDymAP1
vDBdiSC/ZuOZl3YqcP1oQxOL0P7XyGIJTvMIJOsrtho/5z1Q7DnlcpAY5BbSPe64nbR87Nh/Fuxo
48o+qsjdRMEupqEM2ZBiW7Y7sK83AMa0UyAjUqD28eV17HBz28mxbRA5QVhdAfGnJ/8OJLzOrXu8
GIyVvXIW62lF4W/RPI9fXxnMSbX1P39xZYL45Q1c+WZIstrcNXfwDeMS7pQIpEgmTKqwzwTJCkZj
XAOD1e+rGkVlsxNpIH3/2MpUhRZYPsbMkBCwOwW1glQphwA0fAeGZ2AJlVVKB9khsC/gNdlOHExn
2/fzCh10l4QzXs2w/o1hNHAPyqCl6n99ZXe7SSma9ciH77WBhP+wH3Q3zy7qQGeE+ux3KGPz6lPY
URcuvDTnqaqVPAJR8qq6JwBwKU2PIPc3K9KpMP0R3pYX6+Hl0o8u0bW+S4c2r2gPKRgqslkGHJAd
LZPZYn8ek7JMRvEwbU3MNN/XVY1Z4rOGCqLGjnU+iD9gAMkF8JziU/2Xdm4E/LQ0LCSwrjCyUt7r
XU2cUdmNG11KxJ4WQ6WyIhvuh6GTiRPzZH2S19tQvfCjPcrwk7Yyh8HaHxrclxBQs79lxhZQ+/3p
9xkBbe+t6bSAZdYVYtEr2p2JLsaGuatjma8qoEq7dRlRhvEJL7LnYzPrXcdnNTxNKBra7GSzGiBZ
OrpLvwlrlFyPpCgJ4zuh/0xLvGIi/QTzwlu2884+Pv2ZPs5kCdfIJ38Fryy2PZcuIKhksAnG9ATy
4sXytZU/v7awSi9Lfgty/3CyJ2RVD8Cxc21js3VfgCxh4MzVUvLzpxid9w5/tarPxXLsTlBvqxEv
51drl4HMrew0W/SADX9jGoa1jeObQj78AWOg77ZGfTFRZXt/+rxANGh67W4+HNKWQb+UEXYQvM3G
68n7/k8IKwqMYQ1c/a7q1SLEGfo4nnLy5JmwcCh36BV88Kv0thuHs8/GBeMgaNWgcJEQxxkltWaP
If3d8nkOL0h9jRTuu/EY7vKxDtTs1B0vj/eQBb29vn8yyk/oOs92W5rSCiJGnp6MSqnJWT0ZLD6H
/5YvhxgGXuwCOBlx+PZ+qXQXzMsu+0mPVGOWjycVcN84MlYNHVDPl0LH0pE6cszA9JESzGWyF2+N
6WYwuoRxnm9AHWZtmTKrnfodf1LqGPOtjlAbFiNCMqz0Ra3EkPxFCQ8GpVnKl6/78QnDfqpdKGn9
S36GfmSvtq8kTWlmKx6gGMpFGZzjf8b8mXh0uuF79n02wG2UmCPFmrsSyyybwwEoBbk3LOaUMxqR
0XxixHskMgjezUMFk7+2y5mNDvvZvTUh1fv/NyY3M8MbY4TFUnR+nNF/LwYXj3QTcZ15hR3ljah1
BcVXNOIisdUOWUMsmit2PTCB9KH1mXj6poXevTo5X/zbjCGg418P+XM1E/Wj0FSanzV6nGukJB+u
J5xL0MDEtUESzJvXXqvSFvYSEDVGbsGSsVVWqXnrHUUNA3KgxAbXvxicoOvMFT+qN1GWGuhJNw2o
Zj5ibhzzvtRHs3Qq+wPnF/j2rlVM+so0tqwWFKrjEx0g6WRHQPI1DonwzpIo1r1DAU+JU8eGAxK+
2DqHbsTUQE3Z2jZcnL/QxG88CuooSp4spDLv+BjK1cLzcKUP2MUXJI/n1KtuJQB4DCRNw+iC14Ai
NJ9VUWiOAphvu3qKwADb4+ZIgphLUya2Og/2CNBevLTqXsr4ctYVAbh82u7/wR6oyFu7037gR4e1
zoROBiprOV+AikR2qRFvqxk/uolMM+1qSM4OA4jmKnc/lyoXxky8xd/apHY5RDMe8QNubCoTJ5pZ
KBJmLFZgLF+WEpnlNH4fDMFLHkKI9paMJun+rflphRtX6eEKtjSLTrHi+g0MBqO7j4F4ijJqoiJX
hSGF9ahmoKHwVvDUrTTYI8RLYLv2SIHYm21Zg/MEmuAiHewApC1GqtZhSmu82YGhRTZhgcfddMrQ
G3Keg84Nwlg2aCOqolcH6HoMR1CjkwO8egP53PGCXI+wTPS37nTUf6183k72bcyoaDPmsL6NJddb
yqHHrpDH/fssI3iN/lJa90rRS/usN0KX9Hmk+ZG0ErOdWyQW3vUQxECF+//nv1JXi5CrV64rgJuY
5CPpPWUjn2ViDK/DdYBYxX+ZORFVJs5rYiUli5y7A9LuKOStgg7W3gwY4mWwPNYG3fWlD9nTr+FV
HfoV5YBUblMRReZqOTvIFUnQW9IRdsMGwHAox5cfVHtR3hjVsJGCMQuUSyacqLJh2kij/Uxilx09
pvEJSxTdoQH/bwIaxSiJg8UDOY5Igy9SY2ma6mzdiDzIB6hNipN2BLwe3rcZCnLQGO3EDIJ7JKb0
aa12J4plj+ahQllPNbeS/9NXgt4jy8nMtwqkWCx7ncCvTCUa4Nn6qvxiq6nRQ47zVp1tZHJbymto
tnku+enDWghLyoNocC1MT2EYwhz/NSKmxnciGjg+rwzOrpt7cz8QTJ4ojh0C6oez8o99f4xoma1u
kOBVc5QIFHus6i4zjMLr1yjrvi2uAQJMgvqWIAG3DJIqecVLSf3Vi5ilXxL8ysF7sbNBdA9/LQWE
t2nVBARHbFSfs58hBntYI+yfB3dUvKLfxlAgnLKtU7x1fcZ3CUmeagmkIQgkEh2XWQkZSkcHW5uF
GGTb7Cr16/s1kHzIG66cdGuHugUUaOCk5Y9RBwHjmHKcL/pMnSoxpUWy1wH+kkUhajApAbmX8+gQ
4WOn2pLJCRT0l3drOPJDighGYPUxYx9RxwULfM8JHj1mB0xgx76hXEy39rWpA/PjIeEploINnRzb
yJs/ZhUmNM0wG9nr/ccyFQYIf1wV0wpTJ5kMXwXVwsxFBFO3dOf8sKFymvcohhSMGiF4idOGg6xB
3QWxdMWphTm12jb8MZnbS9Fmoy5gAP7KlGavDZxQQrB8/2ttQxfAO7iEfbz8KGA4ENoongP90bAM
8Y6VMA0te9eWZbwbp27W0mXepR0TDkDqEPKYAhNrGXCBjpChzQ0ScCReAiUvqh5w5xqR4G8jX+Jn
aD1vBdxtYLtYn8mGouQLFjUL7l0poAidjWRD4OE7zAdyiyndFlmFdiSqr6HQXtdcKp8tQHoYkZLG
5SBtrPw8IaavEQT2v9z140Unsr421e5GGeMIy7AegdAeBpVK7QHZT8+TkLpnLKs+feJlvBaT21e6
axdN/GocHndpTP27CBRo2GWC/JCjrkz1mmikCOn3rGESpVHx2bo38JA0CV1obcL0UTw5WT6bgnAe
rCdiWZJu8UgJB4Wo7v6mR8f+BqrxSxmpRxkB+0IDttUvCE0Wr7HMu3Ci2PUo+qskoiUqdfxmF7VH
LVjgZ91HSzdhkHJ0aoeRa+Nh9TLIE4YUQ8DBAnDI+WH3IesOUMQQNaNKN6Or1Tu2Lu3znqox8HV0
lamFKnRyx2rZvod+QnhPiTlBAgmtPymGEW7kOZTCsFdTuZiF4luZsXe9RhVB14U0b8KGJmrVnsMu
GBW0D1NElL9dmQP9IISBFFDHUiqvCKx4Ul3q1xZNwLCjXl23MtquWlCr12cCxvdDYUBWfYTD57SX
BFJirXZMGZzyMToyZQn0V9w1AvGN5UhXDrX5Ec2lgaNYuxULutX44/d1Rf4E30dzceUg0aQj2Z6D
UQMIY+U1opK/aFMLn1VCR7hKfgf/JItbQimQqUE88ws5Iu/ff2sXVJRS5FL+GXXsE5MZUusGEi1R
Y/oQ7gBWewozZGerUFA+oQvVICIuIEBlzGylZ7elmNEliVpWW134XAypFe4x0bOaTC6vIPFlVLoZ
yQhLTJiS/CiuhzxKN0UbFWNfJgx99gT4v/tgoAOrLXcFPMF23Rwc40GZY9vHAHV5/2dArupA/LeL
bfl0plkgwuIxQ3PzfMx7uD6hltel+77XBNUJE80AtwHGAhukpP6IPH4aP6/38Ff2943JyalSwKvV
Fy89ncvXH7EKIpr07meOwgTuvfVr/xabkbll+0r8qZ4sa1eqoFRJ5lE4f7r8MJHU3fBj/GXx4s+V
j/uc0FpHiNeqNjw44lw1tMwEAbjYz+oC0AvQvVr7zt1Ecn6VegwzvufRnqKw127YKCXW1zAQtM6D
8C96JwDt+KHGw4SE7P6mBg1+rSJ5bDrUK3Ihy6I+gZjJudKt4Bp6iYQ+M7+xo8cIcE3TyR91hbo9
eSpEPgEPdpOSiteInm/8yddrnFADeszaoAs2BEbhvOzPO4IS2CR5Lj04tlhC3R+vRCrjIv6y2G8t
i9aw4ZzYhLqwO5FcbeZs0J6TDGPxFxZc27T191l/xswlh849F9NwpeG0Ps+UJpl3KrGcbCDkB3lg
8lyFWgEELveQZjRebm8KK9zypXyJaKZC1cAwnYLsgQ7ox6hNh4TSNUef5qkeqru0TrS0xt0Wzi6T
m2t+taY3sefoSrG5iI91qIjvLEtXgVUMO4KCJrmOqIIFNzWE88wfxWm61sjSD5dbPq8Xq8+7bmxK
s2GsEPJ6rhorIgrfGO9w9y4QW+jgtBuNl+e+W01RNkrbw2EJ+uB+NtLO2MT90vqT8NIHKENJpv3B
K5948t/e4eZ5NlRieH0J1uErOz8toWkQVS8c1vcRhZHgFK1iuN97UAT6K6LdPgi03tKt/YXdOSbe
EfUAbE+SijRxReMNRKpDoCuoFoZ9nIxBAatc8XVRlgSol0SWnfSXMzjvjZ6Kebq/Zn+IUaC5Wyzx
ATKSbQ+/lUP3vvl8dRYg0/Odvj0ukKYLqEPqRsE1BE0972QIyClndmoHTp5VO4t7Wxa7aYn837FO
5mtgKBPg0rexN5uYqFWCBy9CC6tIhcGISdc0oWsSr03KE+SyuClLgEWIVbzZ9yjvnswVRi4WdXtE
DPOo5JxcCtj3Fy7kXApJtfY2mgTf/QSSjGu7mJcEzyNwSXh3iKlfUq22XHmEzFu6WDQTamMUcJuc
fditNwqr5/D6j9blsqgEfWmg4PMUZgpuOsJIciF13N0E5G1G6Wlht5ty/N8wwWy6gyeu7S6PXeZ1
uqVknOwyScbp1OHnqPML/m2++54IXLxVaKgIidIC6j6Rx4Uw9O67jHnAi1PFtvU4HCSljJTIfUvq
TPFYdtwGpccJM2k39j/DcTWNqVtvG2NZ5eD8iZChmbF3q+drtI8T1KThgJ/k7iLAV+5sX6X+xP2X
o8mSQN4r0aGOXshNFZ1GmScQsgFz1ONsAuuADHZEU6zu0swpK84BOxMBayflVbm7QeMpGVan5CC9
UAvky173lSW6gIkVZwJfubGTK8vRC1NroCe+U8CEaP+4yfh3s7CsfeS8tzS6UDkfndoqGmhA9g+2
gQDBUk2hHagmX+ExGsjeKFKIsAWTiE4klnyc+RPX/e/gWayuewI1d3KOyYTyuIff+3rfF+jIx5bl
mRTxqyKLypT3cgVdul3s9+ySc557HGmhWEmHBzeVHXeGvoEpOMRWMee7LFWCilfFUmZnsV1hfJmZ
96nYLyvNlvHC06txlP2kIo991tW1R+e5E4U3+Nz2bHDx/Qv0vIfkk06vEQx3rngdt52lkV+LDo8R
ZSVikRe1kpCmwPcfnAiGkHgDfyzq+1Osr4dJk+QKbwsYXADNeYPWwpGEQrVOpT/m3XixUNNgnCZZ
KeciXSH8wFoNkk5WsZzdUtm5L9ZmNnwJWXL12wDcTRK5TE9KiZl0vZVayFwUwT+DqjCj3noag9OZ
d42c/DV/9+BkQZk6UcnzSQeTuzcUQ+dM0YPeH7GyudxFcywASm86pvhEqoEVimVoEV/owGbt2CSy
tUgaUEdjJWUaLfoM7mnfkRze/lh4YcodJ8HAZKixNGncQery8th3L2THjtGIo7+//9s+qLAzoJu/
XLFd7EGH10ZbRCtdYHnqklxX0CFUudx9Wm6HiUrelK0jpqs4eI+NkCFzD0hxT+6aPYkxYybiitlt
2twnEipZ8mlHBrXgicrdvAK7Z/womt8zi0gJKi4qOsMZdoH9YKhrPKrZeo4g5fMfRhxqWCAbPrBO
9emrf1ytQ93VA+ZR/51e9bdUk7ryNDsn/VmoZ8siQ2ObeOu8Ys6pfEfY6xfia3sx4qx9Wev10EXl
cWGxw4EQOOgOjeEEYIHzQEljw3qWvzyihuAKrPcI9AOhVRvXtgJVBuIkNz10cshbcyUM/tP1uxtm
jB0XUocGnCywyXmOibZ+MdABArYKDEr2T06GKgjUwG33n5508N3SweOwbf4ghJJ9/mcULe7elwuq
8UVpq36qq89o+MK+HiUskZrMcg9/3c1T+Vh2viCzW8wmBAGCQOEBRk25LGjvV+FzpkjAxwOQj9eR
y5Mr6ilu/i3qxOojC8VQG1W7qs4MmATw0FAgg3SNv30H9B1D1EeyUGCB+B3BjHP+nVZVPPImLNxL
diIQ0KoMtobXHjF5NsSPYPi+F9nCrwat8spd4xLgwLXgmvHN2SynOIMTcTTVzY2dDIBlpOPaIUn2
HalnfUjjaQr9fi2FHDckackgWGWIZZLc9V0vDSPmE4SumgvoJZY7liDuHtUgRRO7zvX+zn5ns14E
csPvT5o06bYi1L3j0HOB3jFpWKvHHfs+A81yhpPfYCKU8lktHuplkBfw9rzURmQzRQSNiO1/uZVK
5F9Rl0LZpexJe5cWWzfLgmSbsW9ZaPYGQLt8fgmU1qvnanVgNorueX7ihAWev/Eq6IAIerfQbOSF
NMgDQeHqd0BI2mWX3pE13sB92fcgrlj4ZiB1IWBFc5L56JcE9d1li/vqXGhKnfQoL/yGjFW2SyoY
Bvia44bd1KAmAmmykp1Wb+jo4qT+yb42XwtiP2HQ1sH+943ULBaDxZekwwqtTM9GKMO48ipNFJpC
xfwzDhzr3sMcyIDToF9gtC1KI/XKy87w5qdtjDUQtsp7TFmOjNICKV0FmDQL+S7JOAcJbH/sG7v6
2tx9hVNSZ6bzU/lcKH8E9INAw2XHpA0hgrvh8s0pQ60ztKcFWId19ro1ktFiyc9WDidS1k1TnC2Q
e5ARWFbMGkB9wTLkz057Jvd07i0IwuDzkp/TCCdNwYmyMn8fM0TP1Vri/NBJ7pid7LPeCzWPT5QW
Gqe9cLW2vyc62tp0IxVD/kQix8+I+sQpHP/YcU5xmBZsF7NB0zoWm8fxQgW2Hh2Jip/JF5wFEwvm
R9Pv5RLSC6Opjd9wquBZuPN3dz0CXVSV0yhc29HhDFphwbnJdEA/ckCG9FMmvNUzgVTmc4KskiPs
PgzbaJN4gSXDMsEKvW7Vu0ddCuiGZCIaM0hgAYEYR1Yl3IcJhcAFvZRYWbQjHaSrza55d91cmgXZ
99I/2TOD1wWHnadzCkdTDEIK+3MtEEoRbZ0hVpHinqq3hCirFoH670syAYcsCdTFGHc2MSbNJ+FZ
t6qnRK3zXKewCp9Z818pjpRD1Wi4/gkUkBTw1RDtIEj+kG3lJGmiFfC8L9tnlV1a/KfrK8eFQUk3
gmDu1QYD7LtAU75gldo47+3zkZ3fQiCuPrDnsrxg99Bxyk8hzBvOQeyaqaa5yWW/6y+bd08CdWd9
JGB+6tmhZNqU2MT4HKTZASti0lfIMlxEwB1gkGD0MCBb+lPhDcne5iyvj3wGrOrrRAXQP/LIEOwQ
erIGdNIA6fhCVelzJk527xIJonJPQWQC9MlwwQkfz46v6Rfl+Ssx1DGMVyc2Kf61B4s7hZNfJ/tg
fcTZIXAYv/IVkKmBBH5Vm8k17ofzY3G+znY4ICzZXzV5clyfQX1ydGE5jbUL9IbJd8ZH8epcLaWX
1fRAPngms4ZbItj4mCBsnqWB8bgjUNzllhz6KMomlLVyc2t6bF7s1N7MXnLmiVCR0NBA1B0qHIlT
W2jb9BdpHPyHNAXMkkMotznsWw1tIOrCrPCzBDY8gxhXkUYOpmeI4gChjJh6ciBGSXSpeQQ/rbLV
ofdS3HLvpjpLB0JLdIb44s8xhiuEHwJNhm+GP2aMoBiXNnxL7DrMxVKIwkwSXzqz/EydjPoEVGir
ltUOZnHkUHsIYfZU0d/CZlvGiLl1
`protect end_protected
