-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Q6YChPMn1Ahx62ZGtx0yfPQYcezbexDhbUZy+I+16nKHxwdwW+14DakxW1TMMlF1OqsKwzL929Z8
5MIisaXhzsl6yYFoawVIXn2fI+KO/RSUC8KXmW1B2PKwAE4h1FtnbNzhElu0CMvP4QBBKByGaio1
wJZCNU1HENZqAV37okzwJFmR/8DULG0GXhHVRCSgZqs8lbmyZ1J+K+BDB7nyMvF3bJD4NyiXp6Hc
BONHrv0LLnVtxsUfIbOI9Bn9sOK6zQI+XRSN5HUvQJplcVlp69P4LjpL8whTSmepYepbrrGmZ+DG
oe1xpvxpRu2G3luZ54W/ZCAzVIqH8T913UBNBw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4816)
`protect data_block
TgwRAYN6ZFupU3Z7eXDGQNVAcWdpEbIlLRu4OMtGSYTPyr5XgG6CuSumydUDyROlXTeo+UTGO0mJ
vNmcog+ElD5qZkqT+8pKO9DSUApgeQppvaawsjbJJvbF+eV+0CsNGFYuyBpAQYPuP2HDCb9rHyU9
plAcf1DMIpFO5qGMDjkLR5idcfCWY5w2GuHPYus99YawrDn9p5QH5QsAK0evRXrwiosALr4OzbjP
7DTQbK7RW0yfBF/IhpIH3J8T87PJoRBaqpjnHG3XAzNUiJFfXqL6UAZKws7wXoUwwHg9Iuegc9t8
Fccioj9UvL6c0M7BkfxAjy/dgPoFIRea4jVXXUx8/pcj294ydLnABvGS+plRuveOEOd5g6EeKQOu
TqPBavlUa4IpVuCWW7Ztqn0sXsrPHIaNfx34hQAJOSG++iq7xoF3/OdnkL3gEZFWi25+HI0MopTl
n34T49wv70e85sonnoyzD6Qxkh8L/I00k9Bau1JD8fte4z/SbUzUlg5c7wuiaYtt72h1TKVqZBE1
8hhKdE+9MqzB+lu8CpdKaNQSYpPrMtGb+8hn8HepsnR3wp+eIShcRrGyJG3dy3Kx0df3pUzy2LH8
a8uacr60Z/8IZTrGyRmQIUObj7+DtF8lGbz4NpBZk7MrJK2og/0+yHBRUurMlQlpinuiVBy+wIEU
IJaNzxeC1V14BkYB29zLrB2eeId5p3JXcXfOGd/xTiuZA6UfC13VSadWsDm43sejwsaF6v82nPFR
ZsQ307DQpDvL+KCE2XUYgzBHnUXlYCn8x3fLvf1eldIIe3TlVR1yaSUFzCMPcWu5pcLwV/mEFPtf
GyymHv7d1hF8zzDrx1dGd9diRWPF9G+GXvpsNwIzFj38YFhQ4V2rTrOj+O4OJlzL+iJqeLcD5w3E
7kZ3fWsm2pUMoXGN7eCzAzw+GDiHCz5CS8SPn3KOP50xqCGkPdRYVAwMIjckR4oivuhnhmOMlDFU
gt5pgIZxgakb3GFK9fGFIFHlAiRPI7rJ4Mx2l+IbdkRarFWtEFHeNtxB31bvpW/L056JOoOTvqAe
drMwKUBLK2Qbq6PFqb+0keSyCuqrE3Zf5brlnpOWW/xWgzK/zTTJlGZFPO9cBAQNgcRs/bN0YuTh
vRcbH4YnFdfPlR7EOf1G5YaCfpyOdS9b3GifuqWimSleniiFjzJrqH/twYS3w6mFdPwffJTRnQUm
VtQi81aHunC3hKVS+jMIW3eaRV2bFOoB1s2lhoSNxXnUM6DDsGt1sBtfR1cPVVa91gP1a06443AI
UoGfyW5zr2AZj8CziIg4PrJ8J6ugoXWe5YGMkcr3hzwml2tGFs5Ol8GmX789IGYu5yDGe8U6/7e6
Hz3RRWxaCUZWwEhWgF0IqN9UlufKqYFkhCl0lBMa7jLx+7xIGVUKhsGfRQ0GOjUqkbD+9ZqrYTAU
0c2nl8gWF+Nji+xLV7mn7FgCK1HxfPta0ZMQ2YQLM2O3QksYNyec3BD4kxuaiJfhVseIr7cyFWZ8
9kaMRHnDa3yZVs6GBaogTLfkrdVUXtAYuvJpYfWZ3uZ/FeMXz2kWbONt9wTu73eKDxNnX2poWYqu
drk/gFOpHpKjhjTQ8f3WdttSn4mS2S+gS0cWW8F7aX/nSnqH0ry7xclpDUTK473EAsvJ8APlVOKl
yoA3OwUaSRlqScEFZofvPDjMrHNTfyhU9mB9/bYW46mULjx8YCxiW9W8F90ALC8D/uouAU/LLMN1
fVL+oDeFMAXp+C56xCgXt8xd3ZUnDh103QEWG5vRLn143Z/RGtc+g6aXTnaMhkkUvtR7vHyY+qMy
pnjn1KQVKsI1ND/TJVuqr5Qnrby4jHnDjpNiwn2F7YwjGdnFR8naVYmrK7cn0tZHAGa4VhOPe9Yk
P1Oa0jM88AlnDE30CVjo2vyvOuKUqdWqdkSOsOi38FW0MqZ8keoIURLD4udJUo36B8gYytjQHmLZ
QrjknKNmEsx6ho8PppbwihiYfrQCduBMVlP4v/0n7viKOLL7Ed5Ie4T96/upX6tDdajCGnlY4YSj
98JbdQ5yvPMb0fAeZYWDD2I55eg7qIxoPUlU+Fm/IPhNSGkHFDXTftzmDhzfehn6/1BZW6I4869h
SV85KIt9NCEQUl/ukbwH9wj2ELXOvDKEZRuEpOMF/abFw6AHMZjACCxEPbw9jfvIvNYXEq4XSA+L
C8paV4NhScRCYyi3ld3kwI8qOnKi9nLvsCrhUfK63EfddupKOXPaRAtyHWaWWiz2owMIO7gfZxjF
/lIWu7X7kUGnmQYXkXz8GdixYKpyVywdGIJPm8jOWLa7jVJdMlUHdUbDs/pYqU/P8FlfxOFya+e/
lLFj5x/AYt0m69nlJHco5UOzbnccFwehEt/NmULq+xrX2tZRLXTuRBhCBWs+zKUXKwoUZdjYPKgV
4lG9gHB5VADxjq1KnmIOZA9Zcvzzg18j4USl+GyfoRngg71wrh5UwZMZz4VgXkTTCCwJHR0ZqA8P
qg1fVXXsm8s+tLBMB2/Wp5Gq8kxb/7mjQx4GRr4dh1/iErimukoQvarwuS0smp80zlzxaWe5RSf9
c8nRp4mT8h9HQRHPkYR+ZX381THdwIsVpfvtYgOzC/A08aODz6Umqy0KwEkmGfLRWN++G0Qr7ut8
fVbSV/qn1Twtj9iJKp6owCzntk66OyHXcrw/UzOk1byg91wwBjom6cGXNHerUtpGX4PvJUQdmMQh
qzVwgJM5WRHM1oE+qwZNG5WIJhbN7mshIH8hY767x5ubsWoAnsSzQ/4dBMGmKO4DhwJ+Kg+9Vyou
RJhV3ytkWJtxezvP6hYkGhPQuTtAjJrj3vXUoq6QmyzKmv2YMlnjBE5FyQgAisjusWoUUWneQWy9
tD1jf6fxKuZxM/VqMa+s97S3R6hCjkJ5J2mtF6F+IOq19TP5ySnKVUp13LfXTLlFeAfJBmvXm+b3
ufiQ9WaR1wYtFx7lS/fuobG0CN0xq1VX/iX2tpS8Z1eb/x9wD1fQflQ7p1h/W3LtDln89h7OBIp5
F3vIVIgKK4N156G8kVCQ//AA/FvDSamhar6rhaf75oldR+7Mz53CmLsiTstPUeJ7LpNZfM1mGkyr
zJ3IJ3LEzeiDCIe/H04YPhj1DbNi1KBvSDUY2jx3SYfYiBL6QRdrdo37bEuOk3wlqxx+r/n/shv9
T5rdObv/JFK7Ax3/zk0LbihJpSxVES8d43lHyanclqqWtVM3gGnuCYdJDylzczQAKzSGdxcqYxBJ
IJ2TrlfNq/OR54i1gB72pO60jc0m0Hzl0Bjj8Bnc3LVR2W+bWdJs1g4GaQzr9dUIX3loB3F9L4pg
/RFUbBrCAJUgfP/T3gq6RJjFBhFfbM4td7yn845vWASHTXayUGvh6Pg6/73ze21plQHZL7asa3JV
HfABF631dLsPZEUjjtlKvsJfRVHEsPG8zz65g0GctNRhTPez/oSlE3EQ2Yi3vrR92nJmJXv+23+n
Yy18yxiPEqAyvtM+DPQJ3aARJ7TOfPsyloq3/7e/05hjOOsWHMTPLuxg05OR+hlb9xJM8hJLPsH1
RwD9LpjR5rbVetfJctSXvDjuERsRBAezhFLxzvCZNSKo3VNv6Gct3feBfj4mi+4XXNyfMO66qFe6
Pr6akCHMmFZPwl+8+t3bXgf/WsQRxJ/q5TfBbXEUZxEDXOpPyB2Q2NdAsLNs5EHkLAEqfi4ftQne
bI8o1oQfawW6vCG/M+Yqv3vUjNaZ0vDFGIj+mATj/eHo7Uj1IxPKy1pwOCViojbgbo8PZe58rrH5
mXUQbOSjllOwoYx6OQ04FXVGWfSxb/qzgU0UvlEYYFGphvcbCneYNa0kbctPT1GaUZd0JeZ7xrIX
VujUmX/yofyo6sPQnPfo3ECwEAgl8Or/8SMri+EPnP+p0pApn6GCUep3SAwZBrtwdxxuxIwM14gU
zGjJJoyEXbgGXAPtk0U9ZVe5VzSfbjD3uJgEoS2MpJrzHXLygEBDUKuItNdL0lHrp4vFIvHLRFqK
9lQcSp9w1LKXWBNS636KXFMOtPnEMT2oQmexzuFiGGHAKIw/H3riSqHQsbm6WERpxdWPPVSu8DXX
xWdQhYTNwP95KiOnB+6ccd/MlohBf+qwOWpC1SmgJi3AY9zJy3eE7Yripo0gQqzvvcJ8O31oB6Ct
wfO7vKtgfh2dcx8BNOAlCCJ5y1XR4kdd1BZgpuQv6pCko02D28jrZFT68vpj1YfpBJdATvC8KdDw
KaLClkXt1uowRYTsq0xICMSpmH9x4WP7vJwU/3HrrM5g7INwC1ZEOg1L7BjsuQimrcCh1eeuVf/j
hDXWTJ///IusfW/yZzfPasRZISvpXtqKxnQQ3mTdcW1ETTYwGSLdmQY8KjAdOxQuKsqTjMbO2Vxa
8AqQIeVJEEWXV19nUpXZh361/jfbvTLP9dWXsUoiXESouUV3HoOuEequ7vrDp8Rn65oZdMVoEaTS
caeK0RMMK6yYomGFaF/P4YvJczFhER7md+odCm48gxYnMQ8ymSldF0uAlJTWimtZdAZTCVZFjpNw
Hs5q6iD4QZMGLvO67w5b+rMnWXB5gi9gOwjolAUn+ApiRnGuhlg20vxoojjMv4gGBO2QDovwiCWA
o8LwhV5MUnW2BnDtgiOUY2DkLPWzPZ4RjQDMZYtma61Es1KxrBjdxJtRfy8ZCr3KqQT24H6RTkG7
/k2KR98NEwgPIsrWwQMiW9KdIcOZ+1tyOMbLETZ02kGW5DYe5WTQG0cBa7m6Tz/gpbiPB6o/QMw3
r5Pa21sNJpygcLQw1DMJAxxwIYms/31OP9nPAHp7OOwejlR4Vnqz7HKQHn8gUTDNZz2d9KDIahhm
fb1asJv4L2Na6b/8I1RkM+AwooYZXeoSThrkYDNCjmevdrMnJmkcK3pyPXUlzPR0L1KDh5PKi55V
mXC6hYaAzWbP1qqBusUndckVDH+v2oB5X1e8TP5lp9PaMB4tOXEjTI9rU7v4r2u6fU9U4MzYiaYB
U6pBHyBvEKTwFwMhmCCBvrYBapwjvBncrFIgN5uC/7wu2RoR8JYeVW2bRD+tJ2Vt0yNmDdiW+Wyp
2BaAWUwGncCmVZ/T2OmfJGGSfOQNulWWUTBVueTmD+jyCqXmj9vVCB2suduasM7aDjPqQxlJNHva
KYo21Jn5/Kf/0iyjxx70YF0SXm6JuOo+RVXDW7upj3sPY/Ih2cBYdXhPvf7TDP/Hm/bJK97utB3f
M+buqTlb6osSkNOffgbrTOmEznP4wcCPw1RoNseSA5VVEu/zC48wLD1tSCZOCnkzzB0oLoX26Cyy
AecYOhdCd2G2VfgPz02d3PQ8KE+7Ig+3E2RJ/rY08h5YTKD0npD13TZQq7kAFq780f7WX2aM22gr
9NJD+TnJIIs7yTQwe4xF3WniqyV9xEOff0U9OjzC86FbF5MNIF+hzfSeBkw3/qg1uZ0cO4HKoakf
b3AMkm/gm2l77ESFA6sDRCJmj0IAAuHJyjreH3T5L6XKvs9SH2XuDQl2dd9OGK6ZaG4R3thhfI4O
o1SnIv9bDMcHukiHWubRESwtAr0JzYfK0ZHAC27DkhB024nTn1YQY64vlJZj8tzwmTPshOUKc2Uk
3DD3JfzUmhbTm1xxSOoeAzea4SYsQ0pViWKtleXfCyHtiVtmeqUyDzcQPrSNp7rf8BIViro/OsGg
FGiLPnQLJQKi0pAZ2LRnCU2zdGsXfu67sYvw6UbFSwivc3OrmqdcVuyJetJ8Xkk2loz1nlpspwaa
QRnm45tSUZY8Wgiloh8AMLdFSrUPtp47N1hu2zKYtxzZfJoSyXyRV50KYc/IDoP7Mb58laqcX5Cx
/rwzWzMbX7EfimV2MXH+Cn1L7RGNaingbxvPpO8FrvyyEOhmGJf/w5uGEjm8KrrZ4Ovloh6Wk/Tc
kcaSax1qcVIfTUTxMpzyPRT8jHiITActdOw7tkmAq4omCwbR8WP1uDbYP+yQH8bb8WL2gLeEAGgu
uTzky1GLGPX9uVlLtT+GMmbXXelUAznPTCe6J3NMH6SkZJnZkRTaCcWYlai3gKiOLle6rE5XFOjj
H/IypV6VQmJayvxluANqBoijcldgCF++LsPL046FczYD4kXOYJqFdrXAdzpaqvL1N+VaXZQ7bkJ5
FEQTG8Ze/e60nSW7HaV0KqKJ9mF9WWhhdCYP/2yw+pBGZQ26d5hpK68FYogMGeM5azUNq5xf/8e+
69wpl+2jxe5DfCzcx7vE/FFR53ccOTDuP5kNkPt/+DGPNeazFB6ki+Q7b5qolHMPEQezhV0zlF+U
UT0nn10yWrNyQn+WbqZibQBvMMCVKPyR3vxr0REjbeW9E2mWJX+nJY7FO32Qc+Jfh2MkSpwPzYrH
xfqyz9/1jwW9cjx6T854DnQJfcXCx7kcE9VMsA==
`protect end_protected
