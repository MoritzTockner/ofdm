-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VqJfjUZ5DG63PFpcnFACjka75QbvAP0uLC7uQ10wLCqBnRdhIqpMgC4rRHSoFdFfZBCuqScVRazZ
jgsCq3iRVM7DALG3FsqK3TZFqAhhXRcRbvE075Iw2fQqBOXVOcdvdwtoYfwdueBHIT7Jyl4dIR7J
03Ohw7KWeSzANpIBHTDtMVB/0bl/ZBejZZ6RUR4a1hrAL0N5AXlWjLPIXBCmutthSEP0mtYicoVP
fx4sYgjYlDF3Ja6kA7Isx4W5Z5tjD74uWisv7CX+hHeqR8gTFX9F01P1ApypRwXqhqPKu9JpbDdi
IGIQ7+B/ax9pHBHJBw/O5K1Gs0H8mXU6QRvdeA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
lXdrA53vozcO8+rWax/QEFUJKzhMDtSM71Pr7FejqKJEh84FOx1bsk1JBAJ/rnibuxXbQMOmeD4O
cvMWAEOgd8ytFFeI6/iRBiUqI7SMqFs3FFn8UHbLJi2aS6CaDA9DrUJ2LULCsbbq5XArv15Dr7ro
zm6Sbsvk/mGyCmSUgBdEki/xBLRHe5hzUEQHa6AtUEVtJ6fLNU5wEGnwqNty0UylqlxvNFoL3dzl
eEJJGX8mdSBJzvrzI8LlEp/boTKcxbaarPtLrYZvawT4a/Cqrpn9pH79E2D+fX1aL9PuZT64QheC
pvYyfpTnHGDbzbf1g+kLA77uLDZl7OrDZoJuPn4Mg+LWtiJ2GU2Yfp4wQmv3QmMS8Rz4IHOEMVPl
HWMqMOLXZ77gM6WrQT87Cx2eplJp5iuIax2vtVhOj4fgB8M2NUE3bDnfwZklPfmRdCjVSVCLz7Qu
OiCeBJKoudDqqadvPJk4oxan4IN5ivaAVVO+KAruVCuUQdpjAX/nJQCwUEfGPNifovyc05X4l1oB
dsaDPoYqWRcaKOt6CMsDdE0G4U6nrXrk/AWRxxFCiok38UFzdqWxJVw4XwPSh/pK6+w4uydyUp4B
EUWvzxewaLKSBOMKrj+AKZYXVN6HT4IkYthlmW+s35ZpzpsAIOcHCdPnChSmzKOSZBJeBRYd7a2n
HHoBATAYWD1PqytOkiqKyvYVaDEXeDiv5Yl4XgYgrW+yjJV7kGS9XSvHQJsei6PwQojT8q3cDzEy
pcKFYmSKH0AECS2WCfivetwDU8KswRX4arM+doOLF71XmYjWogXLlkockcl6mJcfQ5fFzaWnGMCx
pCrfjHhB6qo+4KgIJRbVhl5sUBUoymZmm8LomQxYWarSwDvptD39xriS6+OhQSbPRbNEAocOFSYL
7eSL6EpWaYkpL9c1npom2ysHPFNAsnErYxIwg7WW/V8jX2DgZ3eJRN5Ire93gh6/dlSfVmIsoM00
J4ckNCNmd2QmKbOPEAfPoiRi45u8sjVf/k8LQfSivxown9ZCnXs12CzL2MnWW3mefEMBPpVVuS5c
wKfhYRQb4caKhaS8ir+dw/yi2scK0mZ6zG2SpgkUfItE9SoYD9qbNDmQ/o5p6rmuiNmtpIywNivb
6B5E9DRnBeUR66SZ/BDO0SM/W3BSJlcZdvfI2/Q3ClxVCT+Ov5TMoDQm3LaM0MlR4WviSHQ1Ss7s
MIIaUJ91ZlbBgSskyJaErQXbLWPeLyhL7ODz1lpqUj5SWMBcTdTn78aJBOQ5i/7UrE6f4GTnp0O6
EcXJ7sP/4HNmsQq2MzT2xA7NOOPN4n4Eshcx6/54ts3MPUkrgf065i3QcXOjN2Ia/D3cwr9oZY9I
PUWZ0KoynjFZisgaMH6Kg/r4T3BVm7wraMb6VSxfODIfZp5zCQcn9xk9wTQn+JFkLnNB5Z2fQnAi
WaQ0LCzd0w5MfIhseAy0WowOuo9fIBQAx6W6sMoJfcrl/H+9Jb1AN5WquPh1COUz12TdumFHycpM
MCPVG9fmqHb4Arg3ceU4ex3k0McqEa/xTFzNvyMogiV178i302aatY7QVHY68axMPtKWLQpH1OsK
+zD+aXSb+VYJD1P7wZdB5WdhvQR0E5jHKpv7gN2cVI1zrTWYX+SO7HgYK5j9aOUTkQK0BCVC4sVZ
XGh/H3RwBRz1fbaerW36NM0BCmgRl9+7V05DvT5zK6cX9Evp2wYXlSNnUpvdm2pyYh+XXSUhBi7b
RH91qHk3k8at+8hejyKEFvicVIk2oXbUPjsP5zImk4BFloAsA9L1rFha0KJt233HXoVIcFOGrvK8
iLLyMc0lqXtwXUhHVM2eEzt6GjvRllWMkhIeJ+q79qfkYkDuiz510Isnoe6DfkItay31LZKweJhs
CBmdIpIKHFRqatDsZpOpPo8SZEhESiYaUtrFtWl+X8KzhfN29149HJdTZPXL27v1TPoun2F6BoCi
ldpeyANXZGRgslccu9k7Xw9Y+JQVgTlH6n27GPYm9uCqSvgfPLyK1hpBTcRxR0aVsN5mY0+XNE9n
OoH+hcGGzPrDYVnzDcYQJ63JINAoGHfC8YLofyR6KHSY2h3YuRq2aYZtxzDPAsrLTeMoobrEN9QA
NPKxGdElvqLUuSasJJMG8X4CyOmVikNQe8sSdHYrYCndHYGQQqWak35qfR9WG+vLjYmvhJY1Oby2
ku3lQAbDL9eFRI1DepurhmYs7jAh7R1bXQW+BHKnwAHsv0XXi7kP8dUDxPtJH28pVahEhAqfKyrQ
JJTlAcncK/q0QGXe6nqekdjQn1RAaUn+nPfGkITIU6sS2SnQaSrXHFXGvt9uMy0Lc185S0tBDQXE
c8H0oM8XZhEROkaVZmiFQUfHS/2ZKg5r96K6HYQRX8hAWULKib3krcsHdDm4geiimr05qaXeXrDQ
hMYjLkVSoVBPdZ3AEtljM42gvV8fH6a287um96vIlR/DI4zNPuM0CCTWbW8xMQViOfnhNfRWU3bv
hLbcuYVY+gmJM9J+Dyvseraf8JPAnWiUbYFzWrzRi2W9C6/fVqsfxDjaT/w/ECuyu9eKFXbkfYy5
BekpZ3D2wf6iLHzr0oXast7dw7yg7q2XEfCYX4Ycxcwxm0EiHNix892S3vSiPHDIg3IgzTVO/DIf
07fVDienJvdBRQyzYA4JIFDo8kSl6BYe0wr2hKiGXXwrKsUVg4lREIySJvrYtLsnd8GaYmD7FfpX
pxsuWdOsSEQFMMgQnEb4+gkVNSi1PKhbUo5GklUUby751WwEUYH/P9T7JTSsPkJc3iMWMmzB5w7Z
tKVyUAqOuFL1BkfsxMvteCmJhD+xOFPnK9cBMlDgG8bef9e5895CcY4XKaEH+GO3cEsaH9k5yZHt
9kdQPwDmRUSOPFTpVxTQ8iCWTw1rS2VFMhn5c4zLbv0LgWvsbNm8+BO3zxisxnJm1YjJTLhPeIMv
l9hhS6qG7jx6RhKUw/YgYtZtHaC+0EGJqmLIz9P5IIHHWqoLcYzAahZeSAMiU82jtUNi7wchkVsO
qMP8UnQjVzpPCyLY77bKUKy0IaS8N9zJTPUSZStXNlP7gxy3J06YSshn8d8iEXalLaUESiFLEfxh
yKyFIEUae++1rYqw24vP+GNOO53t+cQLJSfn+2H/vPVLHBOdX6GX2UTpkXP+vfpin+Vwcj8K0OWd
o4GWR8BczGtfgEMrEM7PIn4DqlZv5fabueXNioDzS6U/Dgrd9yTRTX1ND2Yg8XGWOwg4MAvAzJaP
+jnQglUrR7dMuHf6aA8NZKbaIT6bdFOCvVbkjMoUKCC48zKTXfyxYZjFVLdnbR21KpAkpEdGWpjK
VMtPhkaj78TN3V9nBSVVLZi4FcJt0scXdhipR60D3ZS+SE5VYYIjG1/XttfWDHObOqPXfoNBvmSF
rK5QcP7K0w7X9IXs9onDPRxQW4dHhfBiDZVcLPX/J6qawSFeN2bEakRic/Zq6MtqCxEU8KzYnpQy
/yxCeHJvjk2sN6Ruwa+TMKqdXfNtU1E5RBpPnvWH4mZvw+cSJq1hDMtWulAv8an9XQLwnC9Ij8mU
OUhy4li4wlSsemnBbl3idJd1p7wdG57tdroPjmNX0GTsbSA+W+Y0hkXDf/oksYoE2J7idup7Dkjj
FQlpeOttqT5+etO1pVYQkFiK2VO3VeDMkEZ+o8TyhOWM1dWCd9qA0mHhS94cS1qeaN67aVZhSTTd
ybzUVop+twAB6UNyDYe36P2pFlhrC2kflkwW/F3kLZ4AC9H85CNp4b23pwv4/EZBsBQCTHquDbiE
p9gbF1hRCXewxHXZKDSzJIG5fAS9Oi2SL2NqAvGPo56ZXvHyR8j1h6MWjeuBqPQPKZ/SBMcY/2H5
10a4zMhHNty6pwVTai74V5OARD3vWk0lpZXOG/SOe4McwfYqhlaQI9J/YIw8uvPQAIj7qIz/xJAC
rA/9auPVr0UklM0a3p7ZVCQULilztMJqHRrE0NExaOZ/U53t5j/l8KmbmjiK41bsovZhdq9oY+bi
EKhvM4crRI5bKOQ7lmGFM1eGgGdYzp8MiWijxw0TzPzWkVvzZWSkF+goypGAMJmwMHTujhdKiQsN
bf4KNTRsfgloIGwH8p/lelHParZYJexKGm6gMIv8DS6bjLGkvuzdLxyZIQV2PfJlmYyxR2rvjyF2
7JszltnZBsXlxZ9/nMDgPzN0gfHnmQwIuq1p9A1pD3gf1LzzGntLq/GD3EVE0gky7+CsvLd4bqMz
wLadFYFtNcU1liMrUYKphEo70JX/f67Xh1WJZKOBu/ETGVZhlfajhKeJDQH8nWhV5/GMRRmt/t+P
x6TyYk2yi1x3q2lT8AZl68UtHv5G8nx9ERHv4iGjgPpnaSpMn3hfGwOwDlBNB2RaJWeXryZukBny
uZ22s3ACtLi4VDXVrtfuWuantcFMFkn8WbbXkDZMJwFyTbtKmJ4XlCO4dfRx5gXZo8cKE6kOSjdh
nbaKggxVoq5ex9S1woSW5L9/1NFbhj7F+KOuUlN6uDnnzmeB0JWCodQX1bqaV74FlGqGfTR5VuZ0
Y5Mk8Xo/4OZ1xrqx9MsVWSgrggclY1noW+60wV/WtY4omw+f5YDM3SeCOOZF8dv4f3YWWX/LpqFS
JzLgPBZAbJ974U7cSpj720Wy/UTICFsZ1XmiiBZslxFNUO3fUNPTakSvZOI25fXu4I4DA918XDQT
Pwuy8cY30sz4VUqXipDGj+LwDvsbVDGBxview2U7DzeWpjb+EKzXlsppvfuuzK1J4xJd2BzehAoi
zutd72HSTZXTPTGFZCXEbwMDo7Liq0c5jSfgyEmLCy+pcYjmFnnPiw4czYAOR+JayLDYMEX5lJKK
KmoIF23nRPhQyQk6XABZ4oIV9SeCP0sscgpC+g5ED9r81j0pUua2tYZH0SzOZ1//MRYPNceOMlk0
qO6XudmR+YyP5kGNFpsTOZEK505nUFfgzcNM8ov7rbGeftYBO/b6sHNvpRdakhz9vy45cRvVMVRr
VXGsUHj53pLglKhAn1puGx7nhuAqVDNng+5QmZT3Wxp+prFjgNilyHweiUhAjvDr29cb7QWIC1Pf
5OH/t/elGYDLzCFqdSzOLHzF/n7piGqXWs4oFgeJJIO2U6IeTtg9YN5ZUkHik0wf+rO5ZFTr+4hR
0FWaNsBNWmv/ftzb79mmoQQYaZ4Rvm0QYTMBE2bNcBeqQfgcWhVSXjFqLgWnlfjES9qs6WRN64eW
AOsGtG7bhCr6KAcYd8h3WCZud2yn2eldcv/qdLg82Jxml4V8uZ52uJHz7Jvl6uNlLQvKivFR5ujU
8x4IQE0/AGq6SloeX4jDB0TbVD0m3GsreGOW9ATkdTxXXJPhWNDkz/G2FuOIHiFdKfhtZO9ILBdO
RhNgGCJKQ5rpyGOIsIVuY0SDDdSHwi9S/FxrUpsNrUonXRDxFwGLpVvULYWO/Zsq2TOBWbQxKChF
TPsZVhZQvHKmX/ecE5+ujea1kaftOswlcW8Gcgvqi2FabHSoZkdmvHGeBVEY49m6gHfAn2MBebI6
Ow0noevEUTdNUQZbRprxLmrIVUgafX8oahMC5bH2XOPW5WhotvnF7xJrSumRlX75hsCiQwgWKCOF
30IPJke82gaphu4M/YLgJbgaYUT6LtQYE/rw/RPi1yv4tRfI0H5oqTAbXAwSquGDVxE/6LCtxl7S
yuEyMYooJrTwNlFzBdsoAAYjMktD0FZs2BRvbGGoiKdxmu+jiHxyEb+h4fXC3ldeJ81Gl5RpWdMx
K5v0/vkBRtU6ps4A+MV584o1AP4mU0bfJPziaXnp73zDiYSAgwdbNlXZLgdRz1540Tl7//Hb9XeG
vhb/wu8dWSpr65GZX0gCSD35ngrru/gkb6DsMFzA8gO+5X2LSpsVGV8z30DY3ZnPyWyqhpVfFGEg
j70kfw4NtTAqcOJdRIKZ/9LEod4QpofReM7ktZ1iuTSqesOCaogzjDu7g7ym5ljOfo9yNt0t8DqB
w4yQcJO9WqLLlJCWKrXgT4QisJivtVIpgwnb0pVoE5pZBQ1R5aGfXjFWcRiSoVvpTQ/ZnpuqDdMx
jJdO1rxAhe2W9Kptz48KaxQZNigivgrFhZ6Ewyow5bmXMpkAzdOGaLQysr+JDj/y65veYz/zllK6
OkNnNQvmow7AfK8MYrP4KZYnSRB/IZaQP8g2Rf1P1B9Zw9RF8RmoYpelSHy4iqVfR1R3ddKh6NSZ
YL6TPowEqYTpz1f8X/rLiwcIutZSC2G1tPK+KK81y9veLjKnhlnMVTicQX3ycuPPlJuQklhagHe4
N/gDD9Z6lLmuwoy2Shxebl8xrUgAWTvWIm/JAWVMaM+wf+QeKQ9mXsX/a8VXwYwXBzpigZAzEypy
fbI6eVA5QmgmdJ67IPmLwBZ4cQYB7qkIdy7LoTa1l9KwqTGYHD/PaNivdX3iUntWiVmS4guI213H
Np40S3Wk56sj9cWiFhBtumYg+0v1JPwWS7035JjnVRgTr7ONnbzrN5/HXRZ4sCqTzpz9E28yr9oY
zVGGR2O7P3gADqMiNrD//kzW8p+WELi9u1tEh/yPeubN1gFw1yeOA5klOxTtJx7sOQB5TVOCtQLK
DOyrsoLSnBs5nSDDJTiTlwEEX+VsyyPSG7gcU1Nj3ZVGmNfS9iI4z5GyrbJ6RLN/W/CPgTjarRdS
V9YIsbRaVlKdMc15NwZ+6+yZfDgSB10k3O0wEcKQv+5wiLhkRn9Rhaxr7qUJ7fnOj4v75gueetQf
SjTlCP0jLGNCXBQ0PMPPzNhwftJAyVoaYYYDiVjDpigHObLFqoTUY7N1d/ZE4m732sZRuTfsc6+d
Z/IPPLpVeYPmthoGLN/Sf5NJL5+FLWlTDGm8BzY/DUu+uJ7tdB9oUld/wUUmGuYMz5j/5UmfVeCN
+eFWvP2QAJUo4ZEQkVOhrsqffCnjKeNTcw7JDw15Nx2p7q9n86UDNou40fBgzdr6kI1FcsKMhtuK
oE+pXmAhkdkFbVOUqzjdhK2PSWS9Jy73rtLy336ti/1LAQFTEec4PPx0F1teSTATlRd2vwRFcjfD
9qD/G+o8C2JhUFC5Vx2gk9sGmhROWo/dYyGem71ClEeQAsiZAxTQ099WM9uQUEsYAki/BwLlLLO6
BQTcKAYdgRpHfgOQLmO351zpgycwjpdBGJXydixLNyG613NbBQppIxRBOeir2sxMAUfMOaCwDSk4
YGnEsEGqTmjKiNHCl+knqU/KlfoOs1Yj4nS+DZGD9nPeATGTUUvW8AtgQg3hbFqRDTKcW9q3HTtK
FYVkL48hK2rpjTw4WBhKiaWO4hYPa6ux4bG9oPE6Rk7QOzBX8l7gVCcpjV79shxmTY6bKm/nFwrW
JIhVUMFX9hY9gFMOwdF48xYMJ8BAvN+7ehwpT4jCtBV1EvJ0sQYCd8ErXxOxBkneNfjMDjTXo6RN
l01uN08j9RD8JWHoHf7emIGZE9wTLtIeklg+X8WAU/o38vx3uBTJs1I7GzblkEGgryfQGvi6VyP3
THMsterhNwu5CFqNK8NMy/pR+IMF5IxAtdJyftqs8ZGfFO55c97gC8tqpV20YH2YsbkyB0Oauasf
0g126Z+rQHUPpM0hL3oe5Iwd4hQU7+C85Ztj7XmuLsD7lyFFhGLfyfGx3IXBLOOqVH/s8JaEOpp0
y4XQK2Z7dqkwIlxr5rnUIr2Fw4QfEOmVI30Mw7F/QkWw6NsqQhVQ3G/gH4HZAkY5VRot+kZ0V++y
lIzCgLg4hZAZ7HuzZko4Jau2H0Qo9nhC0IJ8vN28CakWNoAD8QNrGSYyOb2ORtc/1v6vIsE6lbNq
NE2qCJomtDjngpX++5Jj3agkpYLlhzDCLHXkgAHHZuJWf1t7+v/Y7VaT6YikivNX82WrgYMaE0gx
dHWgN4B/uECQRncaMtYa+XbBbN1QjQJyWJPiKLQQejXRglKuNqmH2HZWjENMipfbkpwCaHKFTmqx
jyYFmDNUE+s6h9C6K2W52oCL9dAexS1/h11nJoTLhg1rE9e8u9EH3olpT+QUJhwBx774BbibEcvi
AUAiEpEpJmrAfO+eYYhyCh3QGtiTgKdSglS0U/BEum2Yx0oUhBxMA3StENVwjr0U2l9I8SfGqVbJ
c3Fx5PzIuFMOXtGPE3ekH5xh+1n/h0XXEUKwEwO8bvmVuluBHnAp/IB9j9HGAB4GlhtE2vPlju0s
MhRWH34AqKi07HPmCw8crPV0jn5h+mOGBNaBpyuswwLifU3Il3kChCnhH3eXVBaE5h2yslQvRV7C
MdhDdO2Bg4j79TMQ91QyaFESAOcXpgI2ilps9Ml3jEeKy/c//ZMysrCIjvkTVgQSDE7cAaUz03QG
D7iXlpq6f2wKQHjtLYzvkRqkzRosf/7+5Ki5+1T+HqDCFrSjYY2ZjD00GFXlgHLxpXl6jXa7ZJ6n
azc5+jXPx5VBPj/2Byq0n5L2PwWobh7A9Q2F1svrhlc2xXqak6SRBz0YAvXxKb5QhSKcGdAL9OsG
qD94djefawU7KK7NAOK2WVyeFtZqjdg1CIDPeoDrGUOngHeJAWX4wmoM8JzJdSKXNCQVxjYSxc07
zBJ38yoxQ39L6ypzfLgRZMqdsIXsHaHJHFOCEpouMavsn1bn5wxQKvKbdU9EQM+BiVvS/l2/pkv0
+bqkO294tSqQoj5djEN7RQg+RNgwt5uaOHgvQkctFWw9wRbDuvlr4dNyDnkZ0+8H2TEnqvx4RsD/
55I2FiYMNBsDxsy5fMvco5QCIIBqi9cOEd5TC44FFCenlnraS7bdSMhoZ901gaQTvpvMxjZdmfQ9
NEP28Ejxyzup138jvSp/D9+D+JgjH1fil6M7XdDJ19cPrafwLRwTTVRiyCxHRjGtAZf5ZF/hHxxY
t39S32rm9vO7qiXJ4BhYIQXx4A+d7VeQkoB8bwK39EC/OsWDJEMBc1xdGPJ3K3SOfQeD03Ma5IuC
WGqlYxIrrZ5moe+AIDhVmOJyLk/etk3U1bnlOg16gR+w1tLybzzQ/a13/+zHyt+yb8NojelLVRmt
MZRri9RZO68WMyPLWqPYbpcff2t8K8PSC7jvb1mt/z+o72pLpP9WZcV9dCDjlYuOv3Kg/EgYZoxQ
PzfoTsAL5NligwJCrucChtT9Sk2CrF+T2cGRmNKIZiHQ2tS3OZgQxFE748mDeMLzZxvkK4+32gxr
Mv1fP7lwwUTlIlf7L0ZsxKl0z1rVZ7AVSMEPp6ZooUsl2d4OVa48m4zbZjL+te6B5kYVIVLpk/L4
xyWqCnKGy+HUTa3rYJ1qf6Xj9SXllwiV2qlk9kvp9MY9692WExr3NRCXYx/eZc2DKb0tm6FWFSnM
njIy6ONMqBzchRruZqlN4hsVMP4zfnMFZZDqwUxrg5BuzePkNIZH7bNEK0BuoDYRXrEaHQ8wXfUN
wF8S7XkyMkRybg76dXCSMBppDhl7GO8/wcn/EvxRqCDwEzz++Clq/sSz7CROjafMMOSrMOAP6sFm
/2zGAP7R5+1l7O+ZXX72EOG+4t734YQR1G7vbA0Uc9KqZYrqX4uD8lICt6zmn5RcbAWHoMbmHilr
deg9nNpjji/KRq25vJQIId8wV+tQUiwj2Ag1vKsKzoTdCRy2bIR4zJDrBw7DNoTLJxfnr/lR3I66
bHZzq3fKaYSHvtT+h6GkIYzHGOt0VfzoZxo43TdHmTpXEEgyVJRAJX+jYdF42NhnAat04ay6L2Nv
N0UFUTsRAiJwJKiPkILBxOEOsQFoqdW7Y87gEEMoU7ldq1etPTiyO+TFhLGd68tGUU+YfTKPBiuM
lsKzWncmxVvSrL15227lHVfosExBKt3iVrm+SFjkDzQFYSiNVXatB4kDEBC+c2f9xeN1SNPSa8DP
JGMQcixf6g+kHua9vRYlyrEg6S3va9IzmgKPF4GhCBoYD5hYkMqEO5wRzPpICYtpEmL6EPeiA2dZ
MtrcuXWGmglxF0HhZhYclBKfHQ7v2nOFdyQu/k/IjZNquWBSn1XoK0y1iex0RV+Z4Ych2Nlq1/AG
Fa/aaXEcWGUgbqVBZCzm5aB68htCREQ2jChR+ZBK4SpU5VUBQ2mjpC3o7EqOswf6aK2Xjfr6UPA4
wLXgyFW8QK8IzX8RMxFoXmZuHGIY01vlUr3VPyjIVEXzkxjiqjBVIqOsJxEmbaiADConLQLItc1B
87xWbYMYswVCNBC5kFbAKGKdAQCe8vXAr2QhbuJGtiWFcwZsed8CAfvjU7VmwUumS2krdfPHKPZG
TVmUMpPr+rqe5HtkfWC9CDcalnqDocqeV/refmI2T7aGspun2sq6ZAAhG7QAwynYEMmJj8z3xKCC
uMThnZAKz6sLnRXn2Vz/DCvgmFPRFg37AoYJ8/Bk0woVPVFhHG32QEV5kSNrO7ES0FPoB1EB8L7r
igROvXbvp3ZQ8ZOhDzbVFKIOjzn8zn+01Iq2kDHGZ6HScfHGLkHZYsfp9QT2oWZoULGTaG9o7moe
uWL3GbIHm2OUXcxAw+s8jJRJFg+JJDR7P8nDAAzyJxte2t2iPdIKThv13JQs/IWwzqwp5XBCxqE8
Cp0Vg/7HHEBnnTyIxEGy9HIT4MSAqyc0CgRqtkpnCq84S+g4H+WRq+SHXoeHAVXV2h/45emkpH5s
n3qwS/TizDCbJxHeU0ddr4O+uLN1dCKlzUGMt93Hi7ys3VhojxMkxzFaIWxEZQTm9i+BrmG4mBN/
cAbPo/Bd3cPXSZsBQlQ7pTBvv22OMB11/IN9UtQ2IgZzsq4seV70MEPlKhGCALErtBlhRnLGdODY
LoiX/nZdClr5gGtajQyRlRcnR79vSBb+84CYv+uTq9Fj0QcovRbNZfX5mbwYXysMSiTE/X4U5BoX
WWvdN4PnZoJqfcIxUoliw+yeO2cPxm8vSmJ50wEMrc038M5Vk0+AsLoXmcyNtXtGRImS+yZVBviM
0mgbBj6Kcqt7csaE5MUkroWB6x3u4IO9HyRmNKiz4rugwhWWrlx3uF8RlQ0vCOVyzNUlsYZbslJq
B0Quvm53QJdKeHNUfjRpp/yxA5wILklvpQsPkrNY+uhgxR8Voi7j0Orvd2Swvgt+WJNMuSHXnSpT
CZvcSFQpiS0Ibzhp8gMUjCz5fsfrFFm3nmQH2rN16mHdqn8MTGlLOYkPN/h/utb/G3KV7l/hn7/8
ZGHBVstEB8P+25YnbBi9CeTgkKVDIGNY88FxNNNrRqR8ByEgCrHWM9rzj0JykZMO1I1NmhbE6soA
kMltOZltMmQlby1cji3kj+zFjYoGlfGdOz8JqATa2Wuj7xmKtnG+5aQ6iMPyhQQkZs/KvulBczzc
9KWN/zJw3gW4Pm7Y2eorb8CRO3y2DMoPeERGbsM/jAcWq4C7u8iBzL1yDdouviUtEOwBNLGFiwIS
0HgavizPyONpQQwTKfJRNMnrpCFs42X9LtXabejiUgAF01UdeaWU9If23RGVatAc/QTbow8Rq5ai
5nQPpeJk89YYWkWsUloeIcozxF6dEJk1fgHNYPNmQxKW9zBCaw10RE+tDqD4bBlMm4rvDXl6QZig
L1Avy1tenjMqvBv4LZFd26qLlL9VzLHHCBoz3EYbyUn0+4Ec/sb/u4jtxFnJGC4VrqPAokA8BTBy
UDrghPxNzdOgM9VpWdKU+qJLZ7JZXnWZh7qGW05N2y0K/fZ6majMmNnv8XndTnAOoQry1TZQTJZU
4QokAO+wtyaNiP/IHDp3/p6l+tXVwgQl6X7SzTaOj5sVM6PRuCTpTj3VmFVMe85ZciodvjC6goRQ
N1bgq0+szBJWwif3mguu2hj4nKgwGt/+i/UgeksCKbeQurdcfN4+T3qZcLrBAre84qTALa81P3oM
m58WWedo2wB6X43KpmcQ3H+KRog/8uGzXhChl/kq07PC8gpyke9np1tkDOxkZSx2X9dmE9tElVja
9AWhKw5LgzOJgNYI67e10q7lgzn580XGuKcUdjqapCSJ8rf/AyN8ax2vtkSjAT7pD22OZ6V9l/LW
mgZ1bgXJaYDyEs4UfZzoymbhLt4wXEcrfncD54oR77b/8D6FK2w7jSD4ujhKKPoWjFPuOuE86TIA
/riB0npLmyu7Ln8Pa2mJ6SFUEaX1z4wBlOYYj/TUcFH8GBsBWQGxzzwBMBYOrHvsOnDyQkj10kK6
IYi8WezVTDhfL3nLVJTMrYn3yKAZ+KEsXqYwrjJLKhifOm94cSYyU+BRa7R8bvMDQ+HdknoTYzWE
Tq+dBFfx9tyaCSyYzeALzYlqXhyrFPVHs2J/CdhX0nb2RXmdAboe6Bdh15LAjOQLLRbSFnPO8n8H
TvKX4/JXufWJCaTI4oPSaLXKIu6ir1JSnKkAgi+xT4eJXun3h4TBdv9P8K5j3pVMmm9TdLxOwIR+
LLk8wYuA9uQeHPLHJeWa2IRgjBAXdhNOMBsCo+hqSeGdBByoij4pIqHC2sRhZqA/tfBVr3vMpf3F
o3sNQv4DQaEHJ02unRw/5oakBG3N7Za/CTk0Erl64JkaulHpVtnFEhRJn9gwAPL/pLqi2ZNR1FFt
t2nnIYk7wQBu7AjqJuarvsPm6EJi8ekysU5k3Dy4kjsu51VQvi/FegvHrVLpWMoi3NPssID8bZ9W
zVYpZXVf+2xUKbYuU6t2eKb1mTRFJtnV5UdyA8e/M1odC8GfbiIsM9MSeYiEfUNEgT2bLFGu/3o2
7t2aQGTaaglTHreELjbEc5P+YJyJJUobwv4dMX0uGOzvge/9gvj394s/CC46NfQtcl5QmYQs6GmL
oI4EPOQw2n9+N5kei/B6ENo6HPd4q56hPnLW5DpAygI8KVUDNTuc/1xFkgWCzxYVHX0i/PFtgoOT
uL1rABlxn4TzA+vP+jC6sGJ4l/73dsqON5hO5d6H2wjtXmw6CRrKL1UDc8b66UYydrD6QUSX34oV
zQcGmu7HmbBl2x31C4C8KLiz6QKqGvKitKq6ZqAJ1Hw0dDyHDJcPLehXYYde3o9yklw1kJTP8jyk
KWXucvplushH3AuXS/bUpuIz0JmPAEDA7dt7nI8HJFnIG/RF2IDbS89atZU/tbFRJvZ1oQdSv5Bk
KkQDFg0Dd2ztHbHltmJjbN0Lr7p9jr9wby6SF6ygusvA6PcTfh5UZRpN+m0MDiSlMaEyfzaJ6bU6
lGuuruJitaOVK+gI9wf5pmdG34AfB6Qga5PCtZhb3nm4eDApcCMG1wAP2wf8Ihcx6tx4z4tEh8Pb
WUoqicQfxrCUFHxEXVdS5IE2lTo3IneembO3lyyWkDNKBLU+mIdRqmXolxXVJDGJipC00wcawsi+
kq144aQigmG36L5LpEaVWWKXq59/C4fYJxkbsFpNSb7gr0ootqpWId9bR3H6kTxRsUNMJtMRYknF
+FTxceqanRa3mzRqZAfYxqzaG6Y/uQv5MPrFg0Vg5OA2FM4eJPiCpToPyym39bSJuDO8ZKyhsnrT
HgDf4Qd0YHkJQnrszrhp06811m4G4+JqkGt7bCOQ/6KjT+DrBY+9o1+VAVW+AJ/1CQuN2LUFaqWF
qjgOOkv/vduzJf+7EmYU3LHDiRId34l1DpdP8BRRpfMWGtc4TkgG9Ff0v47jZ6W6LMFa7cb2a9vc
o73GC5VCbd7d0heaSIW/hm8au6hEVD0c/oqKdlK4+QRvRnL3fzxsIKtg+E4BBZWKfJoYDsPFFF3L
Xw2EfcUTligCEtRW8MGi96N5j3F86JDYZrfWFIRxDBFjlVkbenRXM/TS0UttWYCU+jpCg8EMP6Vf
0nYeHtOZpuPg78ZcyFUZC6FtbiC5NMGjhEaJDY/J8wjT9mwl2iKa3nI65/20h+9CUSZQrVGihxG6
THJL0C/D20kwZ6o/XPixsOxAZNO2E+1b0Y/gfhKKU8wVyMVY0PH8hQ/DrTnchs2DLtr1slgN2Np4
y1ftIUSQzXDj7aFr773PnBkf8cPSRnCXKOTETid8DtFhAZUhPjU/sIxWlBn+7RPjJf0Su3w94ZH2
jC2fslTiZ2qdZRFKVIMq9HeuPrvpeuS/hpcE7KisRSGXDri5QZNFZ4nTOoejWgiuH8xNRUoULvuZ
YfORYa/bbzAc7xdIeGee8ipl1HCcVBXRi2Hznd0Sj5WQx6Su0YJ6FUD3H1IGKcF91mnujPGPSOrW
pinpjBFks0LCownDN5YuKbMbZgYVWHbRx7OdVs4zmny7Mix44/l2guC4u/EKb283Fj063pqsm9nZ
0yYt0hXmKmFuqlyk+JG/Ad9cuehimEjIvO2Gh6cwbXg3oTbSiZIZurse2vzFNDrUoUL7CV2ntGHM
2WTybnsVB8Kl2byydFDKajQBfdejw77zTb7tM7ddPGEuhOhbFJoiViNmIbs3tXYiG9W6vEq5djEz
2SwfwSwf27h2dAS7neLA/qtZCaz6jHu+xoKBX/6cnZniUwHCGQ+XZuUgan2fvzH4NsQ6ssANnm+p
SGpXTBgr9NhYxFmx5cVtZAU80Swz5gqAV3Wd4RD2SC75xaImHG0KX+nxiDr9iysXdwqbAJ8yDssR
JUJOBX7G9FFs9Pinku3Luw1Y4IzvVby7YUWM2GyHi3f8+FLZdGhwXQmqeKqnKyUpno6IFZEKSkb6
r9Qah5szlJXbTtVFhUB/R7tIlBWlL2VDQeOvvtpdJL/IJBzw7lj/jm8q+rp3+akVJJNmFak+oZc9
3tjKsOnuSuEA4nLAXYuij1c2AnyL0iGOLcKa8g36MdDh0/eBAWH7nAOebsVTJqQGBwCMTk+9QH4o
e2Zla9qRi6TgCkBmHypHmd903QZkQl1BqZdHeIxrOuADV/wDqDtLxpd2cvIHalxObh4TT3KXPmpg
0v9hO04kgXl0uvrJwqmU+lhKRL4HOGD8IsSZkjQx1p0xAL/4mAHh9YKj9zUl+HTKhuo50J6ebhEk
n9b8zOwY6+3Y1vZ+i0LxAyvkpSsU0Yhbqs3hV/b5ma8Hql9R8Fh/6/rdwZ+I/d6KL9A4BzkTOfp4
inZT4mjyDiHaryeUZHUQS/zf9W/1QqlNNFg9hGtOdd+AMjg3rnUL8zGn8Ey6XtgWbaSknQTAvSip
NwwsPPMSHGQa65RPW/v4ALN+RrnmcObHMVx/npCo0q9bjHeGHRgPjYlew+PJF6fn9kIe96Kqng8+
BydUNlmGivmVQbEKWASz/EbejjWrLYWMvAZ1sRG7hgVpgYrbMeK+tNbwMe5u5ebEd016O8qCAuOa
7EttMk8dfys7j9vak88/geibJb62Usxy+6IfWTY3FAiQO539blGiBul6lVilyywTWmTIppHs5ig2
VCPEctUgkZMGJJigk2vugvWrXhB28EPFzwyvfyDKddMIw6tboaGe7v6x3Z6oXyYsQB1gyG20NWjU
Lw3kH+LHruifWdG6pWZsTje+1UoRsXvL2IwdhvafIEYCJxnnvnBU/pA32s5N+9kHjL2qMajM8ml4
2m9c3qK1qmg7vC3ODZzdFC2i2QViESE8otic+Svo7vcbXM+i5RpMGIKLR02NAKsnHOHaKEFwXm9+
Hly7zd+mXDjlcaetCjTLsE3YEz6NbMjLmPytZc2ZP27uzCFBXth6jrz7bQlQGtABhd4NfPWCXSRl
gT+auLz4uX1Qjkd73ZvLbrCSajE0FLmB88+Y5Ks/upb586NdTE2tf0cWcly2R644FMd2RdDO0EKX
LMPKCZrzniOQnX5e60mK9mLol48gtcEmlI+3BIe68VmUHSskeeUFqxKe0UdiMv+i1grUXltaoVtu
6UNu8RAh9IsATo61cFLbtktvKH3AFhCbhQr4SkSgyY0FXlgfIWGyCm7pbmC7WkJ2/s7IM1tYuOTt
md1DTTtTFWli9d4jSbzDA7Hhe9Cl+1bMQhlcP3LQAPKy5E6sj/wYyFfrKXNt5yMAWUx/vu/7zINa
t525E9f32oSl1sJvajG/NHJvPbX3sQU+Y7Zn0a0zeEr83H5IXAvT6GusqYwYhkwJI/s1KlObwhOm
bEkw1CxcTeePNHTSf5OUywMEZoOGLJeUtGYok3D9f9ZZuEyE3WSuTGon1kopmXIUtv/34oFWVEt9
A7Ja/J3EXt6rYYV9sKNqWKuQrG/EaSK9U/D2tGaXy+lnWLdyWDLc5ZHIrAkOsUu7R0NdMCYxbHX4
XvcumSm8/RsIfR/ITi6+kr71VahYhvsQhfGviuDkuudhC2KbYRcBSqGtkRSAfPlTpL4jvzWynocd
OWt3idqhnATZtnDdgRnXr0SHNhMcAFNXGTK+/njPNXY8jhvroG5Ly/DtGEZY38SmO39i+jlSeRmA
14Sf7Y5DMkvOSqpAK5ocjPhWUVk0UuWqzZ+E3DJ9J4P/ozeDxUmdRy/BFeLB54ASY3MgtyAs4L+s
RcTcxq+aW7D0g2u8cYDnNjcDabjrrVOrZA1SEvdUaxrnWBl7xrohSnNq35LuBFoLd1mGKqkAA8T6
/pVfgib0/bFTS3wqc47YseTDbaGSZ0W3uEwPidBEnUqcemZ0sbrtboq1FyGnaeboBsuvGtWpJauR
WCDW4QNHUb9w838vu1d5woupQfQWqzFfz8HfpiNZT1zOZvRJ2lnqq/4rPqwT2A7DBahvgvqtPh5B
n6ffvpBfcP+i1SXjbdY8ZqlTOSIkM6eXlY9EIqs7TshW0qJA6q01fqUMps8Erb2rIks8f649i4bF
FELbT+/NxN7krM1+bUFxXLPigz2/5kj3oftJ9ph/8CGXxKfA6W+texag+OV0KwTeKDIymQZ4LghF
a7XPgDbD4qAEfF16i74q1M+DUWQFTU5Hk2hbkkARZjCiJ+aODCzwEa2iUQvjlrf3i0x7q4Bg0awE
bC5vf5Gck7vqsU+5oj8Z6vl+x3X6wCKpbkO+lup1jUwe/AObSwGPHbHhRjf6MKefZrWib+t6BzTG
Z5R/RnmYPQRSdseXaWC07y3CgbcvVuILjubKUltCZnc6MNlIOSxdJmZpGKeMUyLGWDwcp/kRGTsg
a1W6W2Nek5BoXy1g5W3IvRwc9NhgnQlZivWzgO6q/bphwAHX2X2H5/sfmM/ATuKTfZQv7BHuybia
z093IT1fIjtH50bk6DSM7NusLodKwzoJglezKQzRWUmaO30ifzoQFvMGc/MCs2n85fe+sGmn4Zum
Ja62jrz6lqBbmsXxGenZsLtB+9YusVmxxOMadnWjYKF2jGcsI6L4ocBsooR+tygjs4wf8+bS1PJ7
u2zxrmZ0gR3hOlDblA1G8Xcy/COOi17fVPPip8oqijz8Zbk4yYUq5eQqG7ZH7yyJ4kky8798NhkC
kzQBzphNTBU62cMyp961+dP5F+tlNPhg198LoZJ3B2mFYB4ujU+K3e+1pm+D3iEm2ldviRW2XX4v
mifoVsTwltpmURpoJdV5ye3LxCNA0tEGfxcHRvO4DF4ckELnxc79EAZVLWsnVeLSEYSOViprWWYa
a6EBv1lDvxOl03q71Z6V65F+/IioRGRF0EqWdie2cnwl8qBs5RMHz3sO3WPb7/AWnSViI2igKN89
xVB7w5+nkD9AJSCNZ1R58+tsfkbwrqoON8P4482cXkmlIjLgOIkhbcAoeLtZ2euO6EcT0bUT+B1Q
ePEWbeMooLrjrxWOKM204m11TVsdWFfOyk2gPTkqZ855j0c6Q0xE1A7ClOpWD8+JYBMNF1KCMpl2
MU9WD9fj0wwzfXRaJnuP3iJSUqAm9dyOzP2Edh96IOtbpZXAff7MwVdO44MtTYxlXHFhe+qy/pJe
oOWgtRPQbxSBRwRi7Su04rl/S5l5rVy6ZL6mP0kn7xJSc9E1kWc8gcmEcU+bOenE0qizMfxNDyZX
U5GncPnzrkYTd4K7/LZKyoUA0d1GZOxQnL7R8YIA3Yt6Ux8UqJ0m15MAco9p7THcicW96PvyHTZr
ebguwm96yBLu2MsWEW6hvXENIZ8kje+Dz/61Z/KDAFgIo4QCHe99j65bson9HU6y7dytUeZCeAn4
Pts6GjoRh846Dqs1ctXAaEc7B1Q8bjnjRIYmKJvvLQlUOrmn0vjP0PJVd2PeUqVb6CSVw3bYARzW
6GsWq6HRd/k3p3PblVxIorXBTywex5FEOLKXTr9WJF2KC11xayk+9MAFkjGVbIH7xbE6uK1aQhF1
DWFq30J1gmcZ2lRQP14A9eDE5l9gEo3gGWACAQ/4s8bkjN7C+UvKhaOCAy/Z5r0fmwYT5PsNldNF
Hg6UhT06FKKsLutWMLYLaKYxHRivhxZ/Vck/fPCkB+kG9cjBDvdzdWucdo6V9Ej+MPHHW3auvyQl
rLZV+EKeF5NcxCgS5SXq+EMGjn6UWuFNK5aYU/2KwIqLWTVHQEwdrp2lAPasH+g7YZneznQcODdp
afLPRRIx8ovnLt8/ugcXeFNTJgCx7l4UvD9oXwQr440jO8420plXYFRND/7D+65I3rTv+SU87W9o
WndpityDXGvRaaEmYNXSjnVNYhVTZS2X4sS3eMzJHoh+bHiQfRc6UFWO8dXuNNRiFtXW2UXF/6tK
CwHXtjFlneb3BDyMBRcY0ZnqR8Yhpx4Sw7+xxFllF93HgFkKxBzi+vFyvWbVMROCsrnZRs1ZzsoT
UuHIhdsjynG7Lp2gezJBl5xEjP9HMiw34RcFnmBIXKxSIJ7ve7VWJz2UIaiU4kJCNv7G2Fhl04n2
l9V4/n9nkODK0Y4RK7KIUQL7p4GhtKiJHfUnBU50fvLucK3Fb6eBSSoNOjh/i3yGZdQDZ2EYmDMv
mLBLAc2jaDAx3FTm/+uypKsCO66U4OA+Is8BPq09+UPSNIQueIx8kDonyBs8xibFKi8GYFQP24xM
2NBbJ4oY+AmvEFoB1M0sN5ed8Ze1LVaRkdxJZXrEw1toEsoNxpr9DXY0q1UqVE0eOALaVCFdDDX0
JMDHV5fTup2dZ6/GoVWzzNTajZcRkkOM+lVmPu45K20Ic2hvsr6EI7Cx2GauXwr6SnfVsScxez9H
xCrW03mqxScHunbL95w5JaQPR+SrH9sZ5z9bSx3gBGYEeTbZrS0JbaP6sZO2jtMW4FrGNzrDS4WM
nufBlxVkYQt0x4Ix4MPhQ7JurS1AMrX3aqLEqZN7UbcFBmxwMaZ5di9pHLDO+CLjs/5LSWZtYd0m
e7tnNJON0NBS3tCI2jzB1a1cOtRZOMZOPMEfCTEvUn6CQmXqWsdL49TNaP1z7E02MBLd32BlZlkG
kAf4VwLnYBlP8V+qzkKGtE0sQqt/2ErGJTlPoJJC+F0ech+8i5YmBMN/gom8P8CSaoiWbkOXAqFg
VMXk0AR15g3sTvb17qGPZS8UwrGbQvKL6B7rI7Y+kpcgEcFciphG2zTo1NbQOqTQsKCR1E4SzlM5
FVwJp5qVL8NxRgEweW20h7pT1wyKUiAzwJkktl/1Oe8FvPcEOa7s1ORrTxh3XCNcgeKAevxXlfN9
BOizfh9WC3/1Fxj3/nGDGR12S8bOcKFp84+/b0RWT0jjit6geMCHsFT+qoT9xnMjtuH7p/a81FlM
NKThMGPS+JGK7CKS9+ZYf7fPmijtpkCY3bLPO5AWlVE4RYYozSNgQyfiJFgZwEhXR2Hwd60Mufcu
SPqF1ZwsigVIl46TaruzhmkZSxQ2aEgs/8ucvpl6xTNWr3WqBh1zfjYObQzjIY7RP9QZ5J3V7rVG
URD6ASDjpl5jmDwJHXiAvdxdgfJYnemYAUZKksWjCF/1YGkvLeMkHtQwvCB9wNTTFz6BL3ohDpPH
o4DCDY7MvHtL8AGThSk3BNUyliT4j3PsWyFdihePnDpAXWQHxtgeIW86q6RO3ZV9DDrE6Jd1qQe3
j2XNy1pcrfXi6nk8JRSv64uss4V7bKklQkXy1r5n4uaaHNWwsPUsg8+ZiN7KpSgBow9bI2cWGCIF
YinW4OpMTngYDrQPJeKcVBWL7npOej8uU13OgfbblOA5OpteV0Ua+sAfC11FdYY2+x/Q2ICyHtXg
34AKLz4mUqHQJfUvK/9fjYG3NXKpr5sIGOC5H24W2DTdNvjDrbS7HBD1pyDUB8+9BT4GYdgPja4R
sVquLRZ8vZAAX1HGvk1MsO3jdgNECt/VBoTb1xC0NBwCoP4TgflXHHMtsfQR6EYzjgdqprnT45xK
6q77lziu2Hey9Mb8OdTjKUQgBw9K7GaZm2BIcGGRsVVSpm1rsNXDQvZ63ApQyECu2zHqJ8qKbcuF
RTHiNerAmt1QQL4gX0NcgZql//GyEHOdquBpf83HKNetjZUFG5DYSJHc07DlqktHe4xHAXptk2aJ
JVVxDa/c0se5vghkNTk+eSpZwfV55UO9AD5sHtGxQ49PfJoujvYhbvuxGWTS7c6EzSppM3zXSx3e
1qe41rRQHNtCzBCUrJn0d3sUkHvQXzX2GEuQ7P2sZ2x4E1pR/rkiNNg4Ze+HVzWDKBz8XRdeW5lo
mMMKLHLeaxLXABNBPvOrnNn2nfuy6AnqWcxBQmjpSAxlHfVQbIUxpor21gA8gOvgbCPQiZ6WVuyN
QwsNPktCNQ/iDFGjrjmiknDY4gCsHb8m6lllw0ZIiSHKbSR6AdOxNOmDtjgeXfRyx0lx/XeTf2R1
uJQztr1vUma9vTOVrIQneJIiLNz23khb8MsO9sprPDIO0jBd9wNifCt9bxpdx9T5jmeMnfuTvfWb
n8kh9ej21uPzfLnem8hnLF5HnDz3rNRTyi7yQHETMHjJSXqI5x2byUiIZgyiWsv9/W+E95IueKdP
mAeV6vpcUOkOgsU7B67FZMZHds31oJERETEOCNSyy7iFw7SHjMj+JcYZeo00gIsPEP0pHaY441DD
qYw7XxLOG2yKO+5S/slVKP7YPDjiM1fmU+Co3sqojxEPqQP+TgcGFnX27DqGOJOqpuLnzw7Rs8Uy
szdyZUDch41qJIRduoee/fpbc8R0b1djFEarWP4No6Zz0Mj71mxuRVbyPYWMyJGtVMSif0jvSNbh
fFRhm5Imf6H/ltZZJgLVgPSlyLb66yfQ1TPdIctgBJ4dyrHF0kpyYyqfhyXDKONsPoq9cuKvJyWJ
H3pEm7j1nwDYUrWi5o+mdrrnBtEA8rTT9HGK1nsfjpKZRKXRd1Nl+1KMZdPfrZnSZWOXMhyVWFeO
Fls/i/tmsqcR+Ar7uKG0tYCGNKqMOM/Bmsa3wk53GMdnOrfAV3BJeF8nufnTblr8Ww3lfl2gxzNx
RxlA+raArcp2SvuJesbBRWXeUsHEwV4No2ETB2SqURulP2krg5xxTywj+m5G9rbkGcFMk+X3qTzu
m+7EATvhfYSkouQ9ad941IqmctEsGI58PZndXPBBa+Pfzt75SDplRx30mYLGbMD5tNNnBl1zSpZL
D2pkVpX48oEWib6SAdpUoIJPCUbA9JqTLyHnBTx87XOx2YM60z+vkTAuNvASGaXiLQ5gz47R4M3h
MuT7tFVoyhM2BM5M2coeP8cXQvNQofHUEluOgmctYUrg7Re6Aicwvo0bsgPVNGBF+Guo/QrVd6uK
Mwi2RPo6lGqmi2VgSHHah4W2dAqirihol4xxXXmqo/SkrOXFhVvY5ykDjTe4tgkxm4+8z7QPC+dO
lOhAsxuJvFHTqco5yW6vUlPMBk81jloY7nF5JOwfkAmROq7JdB0FTadl1PeNz3wnZKHGWK41NYt2
OSx5D4kdH9ZWAviSoVTF+/M235rw+Tf8kFRdHHaf1MAdya8U0HrnJlTMO4t0+3D1OvdrFvhVMppp
0qYbxTUkG4OIhXxs9/Sv0Lh+qzyXDLwRg+EKJWTHg+d9HJwaC6YRWomy4m98kPQ1prbQefVObM+D
LVJzkhCNLRR8Ehyd5PtwPVlMU3J9govIBielabgFiB2bXakxt+kz6qZOUi9H9V1dOfv5Xg5cMAm0
dt3zkG76kbV6/8mqsLVgFyqH03qXQ0XVpOUdr7gt1mujPuX74qlxBzp2O6VpDJAx6jpvr0K6pCQZ
zaCA7Iken2il83/h4Rt9JcAWG+dPrcMBN2oZoqyIZezHEJ1jZjBx4ugBvhc9wEK5RxJRI5soaVAe
qbYoQbfVvPQfUkup6TTfqciAdX1LGTwCnh2nf6ogNnxuPMP8ymCXWs0wYJlWqlRxHvz0R+AaJ2jm
Idukbr4aqJAv5pPadW3D2vMMEx79u3Iy7tz8aH/PQmeCdgC/XAe3irYwADl/T164bm7xEyDCSU/u
y+YSESyeKlzjWMShxMIJTJGHIt6DLzA+QvIHpNUxegnfHtoXFFLil4Dia8VxNAGGEhrA1z6DDuzD
gUlUKDdXncvhAdtF3ZzGiN68c1OKtSrS/yWB7JaKdSrpfOLvCNLdI/6+Ei6UKO88VI//Vk2vPwT6
VU4CeLGniYPxvvmT6vS2gQ39bHz+7/ahW+c38XybCQ6l10TfpZL3QmH4y1C6vvZxFXUDXgc2nS8Y
NQKkJ20Y28OGoOATRconKWcdexx8+Dja6hYHbzU85isJeC1Mi2cft95AQmV1vxFymiK/55kzv46f
3z2OF+HQy6U4j0cPcWJbHTyMVsGoKppxv2n7LPFdzYWVFTCyEQA3Gp/F1hcGgCMjM322TOEzIg8C
xO/kGYAv6dsgRxIyf2GvCeF7Xm0037v1i8yOmBvgu1N+jv5kRSnkHjTfJjbi/Q0KheW9gU0jay0k
1my8xurQb130kZ2Zh8Ge7PM3Mba30/wWYoCGZPchKcd+sokDm/yDtbOXDsbIP7+gPdaTg7sVU8wq
9RyZjbNdBJX2TNPrFW++ckVuEQrlyr0YB/Ms1iHO5L5cF8IWSbtipVjqj5uScFbRySinF1HQCdFo
CksDg2MruowSESob78dH2O2ZR7+hl2q4cGjzj/HYzS4ZxJPEKFr+fni78Ff8QHYPIicleU0dgpkx
YEiG2JwHgzY5XB8exBG5dAW5e0mxIiHXHbcHDiTJBmh0yLvXUxojnG/LOu3hIhPXgIWozOjR1erO
GF/dEG0hyGl0ZlYsQLCIGpLeG1RS/GLRuj2pLLLWKtd5kZvz71HseYfpVOyVzNfsA9PzGjYinReM
hs0MmLQ6wf6dQACV5EsuTzWHr6zAtpshfaArL+XkLxpOW7I6bXLUeGJ43E6pDswHlLYFPh9LLaH5
5mI3BWhJL9Lz6FztRR6lZIpVrhv108j+stpBgmsOGi5sNTNk63U/APsenVQZO8fhzDHdMCwAGUW9
eS0uf5vP2N9Q3298ZRv4OYAYROhELJIj7vpnFdEegU+4ulKf+0L00MLjz71Bb+WfAiv11LpS3erI
xEhOmUvsIXlb9Tr6ukTfq3YVGABhVQYk7cYwUc7wdA0WWRBdIrBrO6ORRu58dZzKMYg+o8HLRDpO
rbNunbxYg8qjT6R6Z3h+/cZrgdShWrA5IhXQ7ZTjZi1wfUp5NZ3o5kRAy6Swx8yVI6Tl6vurHAKz
27nd1jeLAza7P5aEdyqfERUoJrrOvkB88YRsG2LBmBbQ0HyN03GRTPyPjQzWGr1TvlF3qeetZi30
8cYQQFxCEOdPMJwf7gTkP3KLiTKOrCHuSGA8rjTxubfnDtLAY35X4+/OBkzGojBI5ag1vA4Z4o52
qWwg1KDCsOYSncGDhBgDPaMldvZLMOyNsBIQ7R3MmWPDKEO7GO9N0qGKjxj0dNPGe5aJmPf1+52E
Lgh0q5+HKGkLaqdhi4AODbDf+CsW/iv4hwzjFvsWXquCL4iaTtzEN2l+4DNMWsAdOU34ypSruQK8
tOb3zJE8oIv/B1pttzktpTFK+rz6NiSUcDYVCfL5BrHzbqS2+6qTzKzbYTM02pAlMM4I2MigdeaG
ealifOkA41OH6uTUzclTn1Vu7wpm3zGt+6vy/8sU0ClEJJEjids8ouo8WOwEbki074YG5jyom9FL
Vke/rOy/1wrh8N8/NjyKPmZfslu9lxJmIU3p3H6nBRn68WMePNYnMXO2LuItZIfgzKnsmC8OoG70
kTgOC/P1d4mZskF1rD0/vWzEnLV89BraCGvfepiLIjSC8DiEdlm0xkvFRMghLoRR1IIq83baLmNw
yvWI6rvXlsx5Og/8DoxIJJGZFrx7UBfjsR2SB/ksaPVqGiDmq4qzgVq+uKLUY7d8KPG7O3SMSDDF
4o4V4xqZRXk4bY6fNdkHDeYPYf07lNV9a3TKYV/3PD+S0FqfpdVy8TVSZ4UmVMaIwFxxm2mm5n4y
OiFtT0ncJYrPKikhUJniYST4gk9S2qU6v9QF4e15LAVHz86hcGauLjoc6pF2S8Vi2C8KRF5DSMTs
uVSPXV4Lo6tvrvaM/D6LHaZtFdlDJgZ/G/4uehzvQs8ZA69+u4YMpYVe2eUfK6cWVAYpvmTJSwi7
vgVpxaoaEdlD9QtjNg8EEAhCydirbblSIpv2TkgzYdOoItMzgzzMAkfYpEQHtZhgOM/LJwOtZWpb
k/WDp3QkpRqZVYgcopnZ5iSjhTOB/ALlxFZCb0rfQ/HyAvqQiM+rJrD3vtLJ8WE4LdMeGJXQLt4H
++6+ndb8IPoAxP7vR3PGNtWq5za/WIRpMG3OkAqM0kbXHwzgyClh+aIRw+w60kY2iFTJhWAMyCJ5
ZhxjSL0/T3OgdQLX6629Y2he0zZbtoPRz7+Gr8TW+yDZtVkqcPcNUb81maeMDkbjyUMLv7zHPBoG
Tp7zHbF0FWMR1pMtXtlKi1f02ieeML4hbcP84krQc0hOyYsy9G1yGCjsia2aHJMZIL2vGfJtuXxy
DgG0tPgI4nQx811T2l99PIh2rQaL0puoFp6kFDAxxHNqQlZqoAroAdAOjtRAdvP6Q9mGRqXqEdAR
eV/JWEC4DoW3zsjUSv8aJRpkzf6yD+MIYn3vuOKKBJBRb1PrPb++E37x2zsVyoUMp27tJVgCvMLF
fxV6YBM17yK66Qng5bYiLvtnQ/OF8FK+z6wOETVF5ubWgmw84EMJaazphnPvOBuezVYlBlWVELv2
/gfskCJE18J2BGHu/C5+TGu0z/pvPKLHD2lYR/0uJORIo27+Q4R7nFQ7gWbT7env67bhFot+Zeof
pHbzVIa6ZfB1U9kdVo/tcB2SDLP4xwyjgF/unq2jzM5A2rowJm10JCmbMNibr5Po1BubYGZibwJQ
flLSOq5wKLxzLhwh/1yxGHBSfwgizFYIg8SEsO0n5Z/YNsW1VjQHlNNALpyeNjIl3HFhuuoyNWkZ
GmkQfmkTtbyCpiDwLFl993gLRSY+2sFOTPe8208jj+WXOIGNoPOZHu+jxPT9g8HzGfXqe4Eny0FD
VqfHoG/veTo5UvgR77bjqCRB+LbzzNH0PDBINp034gYKOkMF7FzCulSYOJjE9KYnlNGk1ncmbTW+
HRCIj79+ACgpNgS9sJ0W95DQgc4gth+uIneB+iomTCPHlZJ7lfVj7tQ4XmyRhwByj0OuUSPr4hDE
7eMVkH6jTZW1vGz9FyhwTXYsHBu+jYLTnBq/4qKPz6YBuAW6Z9CZP5KU9P+Gzd8/21bPJ25RZn8s
LhplCzc9+9ski/QCtmYY/SreKsN2pcww3vzx0H23SZXCLPiKE712PiLkl9HEH/EyJEN6eBWZ5Qik
2MomlIP7f4J2nv2xidGur2CmD/hfw9dwJtGaSJ0q3kvKqPcZxTBXQQHTw1wGEFB2i35VkMPQxunr
G0cI+pRFyGHqvJk6bYiS2k5BymyixR6MOQVl7CnzDZZyiwEqem3igJFgC6YHSJKSkh+J+yqG+u9r
BUlhGWkNAfe+jNb+H/k3qaslXwWV3bTsR920GqJQJ3UzDW1M1EzcEEwAvNZRD522ElSi3jfYcZxZ
TCKieIRlqP4FVEHyamfUJF6dV7reZkuAX18yzR2Jd+gXsfyp82DDbGugQY9hp/nyy46Gp0PPaElb
Xlv+gLTjDytHiNQ+V7wCqryxm8z6l+agv7BfHhBWWJx1xEit8UpL1vQs1Mvlk8DK6gY3SmC9IrDy
mRJl06YUmH7wSR1ZR2hwtodzSAh4mDilBmadhTroEqPNk068B+yI35hevwH+qZkFPwH8UekrhnUD
26/9E2p0QREDJcdJk3s/6FrTNMpxV97kQ1WC/ZYheZZu4Drxl4E062vhMnQEQ68hADGXJJ7pPU7i
WQbUcVMDiXMqyb6qC0FYkw8QkuzB3TCQpljPhbhgVLtQX2ICPMqR/JoIzRmQMYdqubaVS934scXO
30217OSWf9ee5clbFBnHZ80Kcozo0xEGOFIzjNYbu6MXn0R0ubJnt9sNfMvHc4F+OdLiJBPAouiR
0N3bu6Ek29TEIEXJMUPpoauMCXdCHjYtxAZyNcvcrs+Gto6xjN+v4j/TpyyJ0uXWn6IFYDsEXT4+
P4ktzoQibO58RgpkeobiVPJKj2NVquCjx/oWBwuOJf6iiGb69gFXiZ/vfTRkL23uWT5vQE3sOtYd
ty/RPFFksOt5eWJSU6fTtjixMUmAhQiMz+O16N7s+tIHCJzMAC/Wq2NU8VngjYfnYofwmzM4yTue
J8nyJL+P01njrXse2tj0w2eyjBvHSSriKixkX/8qpIaSSQqWn0QCVT+GAq1IABsSv6hf0dSLlqXQ
2n8/cD1DsRq91Gvkg0H+CZ6tplaAJXC9qfOUH+haZur5/PwZzG1tGRPHrXUfLRfTDM1zYbAqK8pw
36e/6ZlzWbMqhxzh/D2y0q62B21Q0FxJAh6Qgz4kLbzOypfh8rIxfnT9tpvU5bFVs0jbmdrKrXKf
rFek3Hf0Bz0365vA0Nxwsqhesg1Ny0r4l6i/QBX9rEG7gUmlQFgOcMu+cUCQXJfunXFYWGjGFlHc
rvUv07nbYNf+PJTTsd/wYcDjnjYRFAM+XcghRHFeHQF2FxDvblADS1GXQj2a1JRlmaUhBBozmfDt
WJTRBxdqo9tpSXiBUogXOAB2OZcnmXVU4SWbnFCvdVeyzyVPaFdp58gD7dzaaihdSeE8aKoJbe+z
IqOMeBVLJ27feY98pS++lmrTKluaPICZuOThLHFI6W+fNzyIaENVSd22Vm/mxlgKugtI9V22b8z2
IcvAWEQO1QBBbyEBwc0q3zwL/GDjfEnDThp+YxqwE1IfajTQL8OG6hQFkfjZIOFsdWBPSpCzCnrl
eucxt1eME+AzEUcknRSs3MuvU65oEDmyYWt+9Q38jDjijTfG4zfFKzPxnUTaR9TG4jo1IY9qGH49
wkyv9pCqyH8NC1YBPyGvciY34xqkOFA2ALJwvlzImFaW9QZHZbiAIOMLkSBNNCzxjtDl6LdJ75Y0
zyqgcq9x964CwheKc2GxXeQ1v42enjRd3ZLSEv/ROn6pdZXWHjvPlrL62J4I2HtYiCuCQAediiTR
vhp4VKVApBpB8w3h9/zhf4uxS0wJqwjFKBN48M0dN0RMNJh8d1WP7lvWbkXiVwHCkTu01NhcZOb9
bkO/5tjokIwAghfIlwLuHDOFgzkKriI4IUwHwzg/9VhihHek9tezSYrmVPgDlkPdMm/21t98Mtdy
5l+hyK671w0Xr1rPFeT9JjGL6hq8Z4pAz/HAfKlTTj0uWlDA0W0EMntXSXdSmIc25074oneDe4XE
NKYhO4NL4Ag0s5R1n1VyOBHcu8CqD9hyAGHTZiBpC6puE7saqpSanq/5zVUxVvBGbTFAoyjqn0HG
Ty2IAf2NM95uSeLO/G0NbIVdiT+2KoqJkYyAcJLIJ3PLEEFWBNkgmBN3jARHrCyR7ADq6zEfIWba
aKL6Bo0PAdyRv67Z4RjdKbCtUGV1Euyll5DLo62S8nuZJ+3vJe6vVNsGPHxs7F59Omntp0c2UlWq
1iJonw6LsqPb2+NZhln44mAJ0+3NWWL9dr3W/5klJvkxWfC8FqGWrYs06mfsM3xTBvTKot3bEsnI
AdIp3miRKu5Jp362/GluE5Chs550olwUX2aKDm+aIJJEU48ZRMnznqmYrBkpQANnw2ZER7kV0fNh
VghUVlLyoDym0/b6fhz0F0bAS7Vws0WtUpfvzNuioF6HzLDnzVyj/Rl/rnuZMVdaRIbTbNVKfOrW
cwC/LX/1fhadnadEVZbVm4LUkJnOmXzbDHLfmUF1HtiNs0tH7ItDYA3uywJH+FIcLGjhy+eNkhVs
Stx2txGKA1WJ6xX4NHxSU4Y0k4+3EuskQsk+c8drxXMb7k8wt9qPx8d53542m5bYmivlz/BgRjuU
3umZABg5GLOdRSaU0vmmUImW8teE5M2cViPMyUoWKtGtDVm9V7K8hhoAWMIIYbeltvUrYDCgD7XR
Yzeb0zuRQcuhxtpXvFVHDH2QuIPgn1ey+1b8Sl20h7W6ejyAzn4W28rAqreVDBexToHHEpwfzwYZ
f6+b9hqJRUjpo0KRwTqofrgXUrvxb7E85EzwdSzSqB1r7hJYrgC+LnfGP3YMqOLpq6etB4xKWAPw
kPezPBhvWQsxK8o7syloeMaLGoCCH6SMFiRtS9+iXstGJlme9Bo1c2MILToH5C0QNwYKZjtpllwK
ds1QhBOkbFQogMuzoEzNAc73H18oM83/NKnvCgTO2FO20r1A1MjdWLuCs9Vexcu10BPtIY4JN22r
uHjdn9I91M/GAxAb5MXtCNnyWjkQ9JsxggF3baUwyEGVbIB9e8DzO1MfKiPCtttWJBuu4WhY3fUP
/uu6fR2SOngd4P7ZP96I4DxL66TWBpDVkwef6bCF+t9lA/27r3TOHaeC7K/UAgkXiQX2+N/Ixjvm
87Bcgim6YBhdCReD0pv475Nfam5vTCqIyZTiUu29z36qdQImQdZJcpiBtw1QW2IPfLyEk4dBjBvB
GZH9S0LzhcrDVCsZYVTc4Gl9RBPZqpffCTA2kvDoQD3ZRUvQKzakEIGLHZ/9uqkAfMjjEFZLaWk2
AGKNKGe7mLzMV2hMtW5r3PJvgwEEdlpGAY8asbYs9zK+cjewMaEcMOkyC1Y59QNS83cMs8elM4lN
TFed8EQ/isWtPY9nxsxnF9e39h/e1IuocgAWD4Y4JyycXeXEAcHQg0lPcdluiSEW5r4Zjt54Cwre
qqY80hI1irDQmxRf4OUjvXNz/9Ygs4QgsHVPyzB9oD34HdWWhiKd3TOkQkt5OoQXUy9x4m671Yrl
l9lYFBa2IDsOluOFXvlh2VkCfw4TRNaruu5pdEmKd/awH+jqeWzC8YoE+j420f9klmSGLXeh++QR
yLoRBIrmQ6+L7uu+3wXOiW/CZX8xmnO1QDrU7FE5JxjCOc6sK7FjMKGCxjJRYr1YFDPjLmkQm2mR
eH739zwrag/f/HVqpgMs9y5bI3ar75iVoSrJSxGS5usI3E0OEH7sGqnGU4CzttW4FkZsnLtkpGT5
71a0O06d4R1nhj2Gbsbo964iK4qazTKbmYyLp2Xhu42cZK3V3V31BqB0035G4cB0rbJbda8HySMm
4ZmZ8oKmDa9BzlaKbDlrr5jVD1vLk8nVDq+/1HFYeuBXf2POz8hDkkji5Z8nDi2pMsBDZ3bHvUCO
yRKuCqe97D1VH/xG0LX93AjOPQkl/2SAf+YeQiHF4l6OuJLJMJ1aedvHAG4WqBFF+nOfFJyuNIhp
NKe65Ng3hMsZZ5mHXvUwTAuUhvqI8HnTnSj/Bo+WfTfe38TGdcfNqBvcCxxYqfngqMHkpQLK5Jn1
ZhtaldlPJ7GhMd4nsYFrDemoU9ji8C5U2lAOIwE+r8eLlnI0Z+3QJBV4I68AtVkdmN7ZujEROINy
jXPbw8WPvY7a0qV2k/4O2xFJARKnEbfxCl9X9Tir/f4Wf0oB7r50Ur0xXjeNrZgndoHb/BbD5GdD
Ez2RGxF8eNlXhRpC9fe5csosmmF4JdWTywS3RBpUntnnRIkE8KFSE5LLLnOgEqdjMYwPmHREOizC
1Hiz8XWjKCy8QHqFXs2eRxxYCWiAgj2yHSZXsObs3udZydpzw0BjoLmbHdWNLXDLkiV2vAwd0UwU
Hew9coD45CxfI+VzMIEmU/i2GDfssXv3euaj5OrjtOz4RcPGy6lMmNgCM14Ff4Z7Qybb/5318iV6
YxN9guWsvfdDtrj5/AXQuHQM70BUzNF6PrwFWr22EbPo96XE0yOj6J0CRqjiH1eUvBkuQsGTatsQ
9EPp9J5ZfQ33Qu/gdKiiCLNGpXFgHNNlCd6pg4eOvci2BqhZYeEUd3k+YPQUr7FzqBHCe+amYNng
3khVwGmaPTsY94DQrTQqB73sgCyIDczyuPT++ywA4HqJDCQZv7ML5wAnxEogVpYEl+xi2tJQVd/O
NIJ/oWdpmKVP+SERnkS8/BdK3+R/4DZiqfV8UNocOT/VwpXqpO+u+vbELAgnXrXtXlVI9dYRctdR
HblP5JRxuWjS+VGWyX82E9V3eVD5+ZT5zjEpUsUUxXDkRMeucGbIwwmi8IH4NV2P4g4bkAx7vGWf
5krIzdEebMuisFs6DWzY8WxWAmPKZ6cUVR1LQdvtsYbbcg1p3nIGmL9sgHVZJeJnxwVSliHAr1fW
mfZByv5sCSfXovKuaI1UnSMwcVza8CJtekw/e2y0eeKr57yuzgKj/ab3p4yYQnTk3zh3YyMldK0t
dKDXxMhII4RPujm2JyBzd7qtU/tTQnGJ6Fpi3cXSgJJ5fP8xtRET6seiv+USoCk00R2CJiB3OpTN
R/Z8qJovHFWZN32Qw7QGcVqscAoYQm+43t02w3boiwgKMqtGO5ApK8kXK09j4e1q5v5vCuUZGdPC
gySzz2aIf4cQ6gQkxGC9XBbGaGqLaatKX4aUFZcP7J+ad8y4TZCoOPqloITED+GlGKLvKWiBQZGt
aWElO4ToJ5Ltc8VW9ol0ZS3bIQaCQji3OS2mMv7eMWZZQBPD+bNIZIO3g1QsXq7qyvvCCCGMG84V
6TAMnRRP3IIHfc1bx6PXtFW1eHI2ZuA7SiH5Is09TcFRtKDtRG0D3O4Qtuw+Hk2Rg3XrTN+Hzv5V
NaXVmBqVDaMxCuyShu2HKBTxoBnZ7gOpmiXDihDiP4xV0Cu3U9LZQJ1G9CEqHw27bHaajOy/PHlv
WVahsPsqO0KeI+MyCj3FABAeVd6BsU/7OIXU848+7MXoNSfHIMXINdG6jDum43P1fI7cDjwkPffi
GhJO9Yr44jxT0Z250w7vcd18iijEsZg7WVhEIdubqWWTsyUS3qnOPEm5+8Upa9PEnGK7tSF4x6bg
ta/eZUvu14xvSiO8grldrBE6puPATbGDRBrxavfFJBOW/v1Rz1hhkXtDsO/UrTfV414Aw3xo8CC8
NdoJolGFVQ4jCm8/AnIO4+Wjvk+mALaigkZRKYJaVI9eHFjCA3rm1NJLlqcyDi2Xr2rsjRRdOjJ/
xTitGWdHCCHra16/epH3lvdQN8CFGFf36pApN3hat5kPoHj1pIiXLK/bzEjWcfq3BQObhCHehDtU
hD4+w6Ehbi1mYdyBtu4B78wDrr2tq6aqwXd1e6Em6eMK7FbbSQbgw6nC0s3bdDZloYPccN/bpPb6
2x80kG4TvCWWPpyNFRnlIhTI54jj5K1pFr9Qc8zyvPBAvld0lmB1xp62Z6iByFpYL9ZXruwNprDQ
FSwkUrAAZiwDnUNytP4Rc9A3G8krIqXD2jEdNiVqS+gbHcXnEIQPWq9VF+jPGeqIW6HY1nvhqZnt
lqcTLVm4pWudsshjUDfFPvIB6b9ofpVKdZAu5PLX9N3s8F/4NHjwfIhp26GkEg3buqxNFdfhnlz5
Agy5friRsZEqt3JqTmIJJq/80pb9MTYUgKEEQqzaSwQf2hWTc6aeg/PrkPIuELTkiN7FOyZRK7WR
S6UJdU1y7HTSoSk1kTYC4K8CGEMue1UekPbuleUzI0fIoGcivGyZ+5lP2x3+nEATU8YQK7kLlysa
yq9tJv3JNWSb8zbxvf+O7jzj9egDwnzRvktD129F3G3pUQQPs8bNZihIFCvxv/8Y1yJfAntXHWbK
o+WJdh9J5JbhpRBJOlZ5ToX576tRewR/A38hku2nOon9JCUFewaCm4f55PG7arBaHRXqaxjTUtZw
wpdGnIDjY+YSRcHdZ589xZS66UZfWL5qLyUzDYn/LgN8HzGT0DsstYKn7MzWHnVvGWyZxhTws/oC
iz4b3uJ645xo9+ZVsfBA12npfQEyAq8o9YJHv8PnBvOlH40UvsyMCevCcCedneQVSlCNNuCkPRPy
sq/jgbZKu42yPbZXC28unWpjB/Orf+6D/Hhe5p2O48vcAKPdm+5qc7pPCOYjtRRRd2Oy+JP9W4Wn
0N9bWqpaKo3zm/8t/mSB4dN7jUPGhXRnUlPbR6oKdaaXHcMmi++YWZ70599FnF7QSOd9N6n6Ri0E
jn6M2pZ2A3cG8JQlQCDZSWC41aFFbVvGhOTX0k93prJFKU89iQ+nDP5l0rZTAmv6y1pZ+aUKHu3D
zpLOjCmMowEESFKu2UghvnBO//a4avUKdy82YZQHSnwYoaECqj1GCGnphgE4WobIQxLB8LtFSSVk
8b/ewhEQfJvF9i2kVngVRHgPKygmjMA71f5kfm9BnNe3sREis1jvVAcSYEwIH2HxsHExHtOtR6NX
GL0hzA7m4ghr/LLsYfWSYiu30c58SEunlFOnp6MFmuwTjv/YffZZ3lTO/P62wsaGxPGe36WG67lc
thXdoBVjlzRdDvp47g2a/rKb9FMrI3uw5X8o8HQXDJySiH7QTw7UoAdqEz8iO0a3pte48E21O0DJ
L9eivndYD4m7RF7+C/K0l1j5awaahZDe1DO3fQo+MataEQD6wRJTMAx0GdMh6ykqKquoH+QNM72t
4RHESWctjViOQVvRgXkGuMD1iKgOc4Kc50V+xebVJ1Ou8uJ3ern9ZphKJgVR6irdYg1Rp7S8PGs+
les7IGSO577ToyBpLR0I56QjpEIEbyiQKCORzEh/t7LaTFQx5bXUGw3qCIHbZrpKI5bh9DvQKA4P
6r7SScO4vG6G9/UlPuZxmdTpjWglFMxBVtXUfmwcCCK6NsvgEsAx8Jz/fdPGUlIu72Fem/LmC7mi
WnuX9spkGFAfTqESeD3XUCboGh9UPpFTxfq9idqkpM22VG0zFgYPhznAZIAQhfzYioslQY3+9SYr
Qj7GfdUz1SlHdVbDit3dWnpx2eOuwMdQgx8iY8voT9WAIolAR1gosZRSYbZn8tRmNNYG6IvAVkA2
hgQZWErUT/J+H2upoc6kEbEMcJOLjy7mYShvws38DKacAWWg/sJbIvSyv8FuNy8POa/CorwnxK2G
ecStJOGDXa+E9nxpQr0SfWgD/qJt+FdkjpklxsyV0FNVOknh0/Umi5ffZkmsXU0V21it0NOZzLHl
gUOOnaPzk2YMnB+sDSfTNkTUt8ggxBMNJj/RlJ5S7Wf3jgTAaGOXqfb4bUy0MDf3s7kT/i4VsFtG
TW+YUQsN71nN+qfK2GzFnuUwLtf9aJzi47SDa4dvyEFw7iu/Z4QD5XxE5qx2fmg16ULczUJY3BXg
LnM+iL2lrmUR9mj4z8iHCXdUQN28xTGATnFXRxYYE01QKzA8G41xFyyN6oFOqUVr1q4HzTJam6mJ
jHwKQlP8fNcmdUZ6Dh202oVU1N+l31o+kF227EcGU08kTaTuKj2q/OS45Z8Hr1Ykyq7kH6XeCzMG
w82K7JUZ2rR35bpowsSur7oA3AM8dgHrlNbAz9kHC5PedwbDypETpTS8ivtPa7YI9EaoTTnCFq0s
8yoR0QIAp7S/VjEIGdANczY+5nHg5PlGqnVqzh9CHUV7HkTe6ZHqUsq//4nuhTBCqk9L/1CjwdCJ
+VjngtAssVamb+2qLjgvdzHi5baoGi1q2MIv3Q/alZHh3CqpQ8y/EULz3UDc4eDGwvm2NgUbmSsL
Ljx7aPWbUXf/10RAYDEpEZHDwnMNZBMo9UOR7IE412U6HGyhNXNRCD3vr8d49k2o1PbeVltVLG6Z
97d+8HwkDiZGFI6NGzHPykxV5WfU9U9CuMp+e1AukU82xFTOk8H0O5HbO0kgjce/AbAyLYgMmPnD
l6utbMs2Sqnmf6Ti3E+9BS5edtq8HdTmZ+8+MpEEXIWsdhGDojvQdUHSDm6tabHXmnY0wbkoaljX
jVPUWf4SnMsi/XUpktKgi86qI4vyY7xwGy/GmIqvlPdUABFbOHGytqA52PIPq+57vocujG+xM7zY
j/lPY93FOI12fnR7Dzaq8FM0cr8yrXZjJdSlbqIYh3b2c/GMDvo/+KR1niznoGBKH3sneWAqy4JI
5m4Pb3IvjieyGkQOJ/K2WAGBNUtzywqtYWus6EYMvT5kx0NLtRLqOqmlRHC6Qca9maj1g6GbJRg4
zv6/+1Fdd1y8v1WOp9yY+1ixCJ75zLwSfvK2Y8MVUGqNfvE92ZBNhaU87bx4/y1HjXZowKS9naV0
h3FQ7eU00FiP/Gkj+c8As65UE1VzHInMu34B9U8QC0dNFWrxseRwRH68o/9FXFjy0iHiWp1LHmSH
UF8MTMw+tsPoUj/I2X3k7aniAHvqk/FS1gNkS939+fW/fparrrFRbU9PfGmGcT2W8SbkEdxQzuWx
OA9jCRgJy3War0bG+wriIHX+Lhx5kX2S1VVJ4BvppiD8nOgqBX7JXugopBbizSCoJE7oS7ZhIYTU
5omZUuqCCk0Nkp//sKIQ9dsCthIoSJ/becZ5lCY1Pj9O9eJKVFpNdIcxTC9ipVEB7LLDXhqtHUGK
Ebk9oDGc3ZCjHiD4/8EGZo3AEWWUKTxnE9Qlf0SZU4UYkIPbKcnkieIy/KhZPIhDg1miKhCiOQZv
2lD30C7QkZeg1yD10IIubfy3s1HLG1o1YNSbUEcNkAc4UrJKjXvZUcdI5nhvzvhrxlxu4yAmJSg8
kQKhWu2c3YQbu/ErEA0Ma7NkL6FJc0kEmEA9+vh0+hDBl5rXdiDdFvR6g1OPbmPLpbesbhw/7TBP
ve+RnTUPyv98TGoEMfgD2KgfGWkOhzbvDNN3d+hyp2wV1cRMtODmZjsBTKKnbsLqaQL+5W6EH4RO
Sj4D/ZteAyslI0KUTSj1YPdHptoJw5RVRJyxXpyTzuOWJa07W2s+5Z4VQk6DPR6rtSnmIcb/tMAV
eoCthYbPdn82WOHlVMuFN1mOBauHXAk9+0aMZC4c22n5e8QX5Vgde4iR/EQrZFRptv/pvPKBi+wt
ApMUhp1BnEY0WGURuXFbcmdx7hX2V0Qfx1le/kCYNipnHFY9ldKKUNq++yf+uEKyjhM3yrfDaOjR
M5rmDhbJskcavDoJ5qpNdUB3vUGWoaZuZyyaVwx7jcwOgUwWNubyR3BafekU7qp/1YitGZHPyUim
s1OgVUhB4wi3/IvZR13Ay7I2YA1blJpDEXa4k/Z8DUcp9ZscjjZ1YRataFMsNQaO2a1XtsMjDfAC
kZY0wF6qHoButqK/u0o7XvOBb4veydd5UVTTvExp44cAE32BEaKP2wBFl29f+V7EZ63YXfk1lA03
n1lyOx3ce4BX3/Wl2tMHEgXGE5eaaBAhfMcXR6aXrEobJWq6hSfUfvYDTZUS6v7yVDsLoPOMiktR
wxFPGMvEP1Hyl1OelAqWzfA0yRooAvu8L6c3mRbxceScchdB8GrWKmdlZiXUpmYgrXeOVESk1bya
0ZnsOE+C8A9aGaloezDl2omXcfb0v+9asRjISRH97Hci0rO3Km4C0oJ5AYggg6exhTID4OltmodI
QrQzDFwUWxj8oK1Nw4HADHJScfuRsA3Sof7ukwaZ3VwwzPci0A7ZkzAS/2o1OC+xOz0HIUUPwJR9
cLU5DAuhS1G1EO4PaUyKQfyaCNsvJPu0br/ODkKc8ZrYea1v7sDnYnKdAWcteTB4vFKrrI/2Kb/m
5iq/cqmkjBevME1NaDa2ZrJG2mbSY4ClPm0tvxoZjWQG3O5etVcplFB9TxP43dEwDx0xgjtwyjoj
WaadXJrLQ36fl0tB5L4xXgFCrpSha8/6jMYVWq6lDl0hC0vpYtSA17h89e51Fc0NWjXwLRwF2SjK
fR0l+X/OsKV/5UyOpHOgzmMUZlmFLJn5xRWV9IzH1F3+0o8i4FZkgQAn7JwujrjkdFlKTCPNObF6
EAP1ms2GlUxcOEef2IB7tEouVXWbU29ZswYxZrU55GApD+sW84tS4iAfqwqLL7NJDkVceWzUUd2r
ZFiL3XNqoTV0IzvJDle1XWG9KubYWUSj/CEhvAskF8ZV97HaF46/5DQXHTkPH8YWPNDKaUXN8Zc2
VJDsWcDqLACzmrVGUpUDr0lHzjAF9hdeNzhn73ivHtr/SHoz/+rH8h8MJob7GIU86DQaMXAu2xB+
Jh1zvxoegM9gtm2T0OADZPqXcUWDcDuNb9daw4U7b3YUX3ACmO2Ofnz0X8eTJ3mnqoO91cRHXN35
3V5HrTMXvDFssos+DTDBc3jMiOhHkgGtrBlmbeJKmzqv0JpOennYH5sO8AJpvL8UgNctnxi8BtK6
Cam0xESswsXQ1h3qXpgwpv4/ZaU2gjJfrCfAHZdUekeymxGb+J7DoRLYJ7ouaLanbCvQKv6rijWn
O3fn/2MbkMUro3bG+QnRxwqdyprVYlqDr7aD+GzYwP/121OFFdSOL/BlKZluy+bpYH7p51nOk8hQ
FFqK4iRe9sf8qqSEOnUJ1XkmbSMSpLb8PXjgEeg+YYdzZ2T+F+U8IrPBSi/4XZJaRNo6IZeaS2m7
ZAxExvBOdCk8Ig+byIi9x3RcJp3jRglCIEpV4J32EZnEcHLsd6PqEl5wVbgc6gy0T8Xw6LRMkMWI
zgPQ60FKgSSZwsAJAW5f/wiesf+nglItj3BWPt+RMQC+s+/nO9GD5ShNonEHWdYLB3kapgNtgbrI
OuHs7eMYiSZUS/Q67FeAV6HQUo89WtVTD0uSDRItHP6of68opOmF4xC1LJMGUmWeVOvbPIGG8lml
6sPHCRXt62W8wOGqXfjuq1w2uUZsMoBYceZyo9XBUOC5D+x30s1F9VucBTbfsV4+qPpQdZeqJqrD
94BrK8FASGc16g6P42SMFWbC3SDwTtyms4k1kUYxd9SxV0He4Qyed8fqJGXNzlCclAf8tfjSdc+6
wFSUWRGNgNdAJ05Q9URgdjtLkwdpoXs0HhNtqmQ7gwuNE6V14b0aQahisnPY6IrwKAoJtlcANiMg
HrZEFNnsW8nx0ycj2+1cYMIEOr718EL5wXmLr666HTzLNvuj6W0deeNMD69KHN4/nL1C5IqMBXb+
EgMV96ku0MHZDcWaakUHF5jOp5JQo8uSJe8Ue2rwGgsaXGof7+HrjU8qUjdskZwBnv3ZbneBLS42
QrlcHvVKBoK8kmqC1SZVvc2ehSrYG6Qv9BHLt39K2bEkOv9KVHKB+4VCFxWpJVoK5ZWxNWVLwUj5
UvoPRf55FqxkUiHBbpljpw2Whyr4wyjoLNavklxQAOfPk7KUDWQCSdJu6pHnJKEYhTMZKobSxCxn
T1KqHDGXty99l7wQPJNiG6gEe5K2mSQhyJl9hAb0JmFLcnXRtEh2wQ5eEfMkN2oVufy3fzjhCiQY
oilLsKrLjD8oevFGRxqIZiubGfttMnmaShiVXoo+xDHDR6uSDjy+iWkZsQjSHUy783mQhUOVmW65
ktskefwK3CjIXw+UkDOXNRenP5A4/lFwgANLqpf3eV00YnNzYV6p6SpPCJzG2Sf1EFkHLYjz6nxn
XZnhIKKrfuVY8AP6DUoya33vrmAnGS5bVsEsXG39o4DkmBO2MeD8l1iIIhdME5mVvWLYtSzm96E5
8ee3b0lyM9ntDpsC/Q4BBUkSk8sapj3sF6PLgCqycAtdSUeR5hqaEUADacqFu7kH6pWJricVbhvs
AC/VE9jWTTpviJBImOdb9DdbGPmNSvtqTUPrVJUmdI4un0IJrMQ0ZjWas4cOlCM5PHJqH/pI05pD
DJChTsSksMRFaf4XBEiek2rbDvx9Gmf6qGFaerwkIDMdjDhElS7hShI8oZyFmpSCK5ALrRxMI2+O
lVWqiHb90EacqWDX0MAyN4T/oDQap2rG+O0xo+5/MEOp53leMRihHZL5mJLfGAmxEo8oulVZZbec
1RtS7XV/XKYKIXll1TZdfvXdbNplEU5AAVOlAoNYaaKpPlvsoeYyV4yYXJJo8VLQnu5yX8m5OqCt
3g/NrflbnW9dFFNU8OteWPz7BcVe2BpZ7pY6szPpLf6HJaT0RUX6p3vif9qsgjy867BJdBA3Pxrn
G6L/2u3rFcJrewSj3zoULFiSfDaK3PN/eDIgYUZHHoYGdPAWJZsIrlyEo5uXHRncGIbkZtl0X7zZ
FgxFLaO3I2ZKZ5EGK5BbGBM+MV5150FCYxHSsGFK99SdcDjcaPbDCqyG0v9mxDwyLTirZdDCjbGA
6yu0lHllmiYwsGxPucMPUkq25S7A5drG5JBpDmQf+Hhkr4e8rj4cOUwBcLV8QJ6tYNL3v1CIequP
g1+yjU4J34mH6rLg9wYLXW1yzqaf0aVBvuvC95g1miJD3V4qlO1KVDOltgyOJK9H2e79jpLttP68
+tRz5MUU5ta6h2lCdJbH6sQLBRxF69gcInXZFMy7AwX1QDYOUWuBvVNVvr4al/IsSGfVgRqq0WU6
iJyQuRKmm/a6KrLiRTob01WMmzbVakyIlJcFZ7I6BpyS5R+Oty0BCDARylgAduy2RAFAvro4/nk0
Pnif2CWjCzRynIdqtflmT/+pZRifuTw78ar9L5DueKUKw1TZAnkBZH2OXqNqjrUmkayEJtDaHz/q
xzQpyD4NSTbb2Ve8IFgzCLlWtFD3z70AdR6zWIHpnopq8Zj+RTxhgsoplfZF5I+aJW7iQIYi7lsa
uzb8wjAWfNrEcos/mgKvFAudTa2n/eeWCQoBstWWXxREt2E0aNC40uRRwytE2Mv147T9n6oNakYh
fexlEiSvpTy0jXxqQD4TGrIDQVGNVgOKKk6KfjJKVaK3yJ6RkJ9RAEixlWF4o/vK73rOp9sGHU41
rQMpc/7DusDap9YcCrgUGAl0aGp0CgzSGSvl0L/T8YzOEUqSlN9AW6aPcPX5VpIjSjGpUwJE8O7z
y8XOMQ5h5VZ1NJmYbmLe80cWw1ZMwcYaXAV68ANnraBxAKrhz3W8Vz2xMODENp2rnWofc1j5pR/d
ZH5kXQfVXyJDvcfAjaJGgDIWYZspzEuIDPGBBLpdSZGCg717nNsFqvPUjbPCNwyAE0mn2HY+FP7Y
P77A9L0h/1Vw/xIKLqCNgs/SytGlnwoCNnkR/U6h/bkfggtBRAA4V7TT9HgoYleaowdRbiE63Aj4
Y1h+ShVJVL7oQimKCrzEhhionW0/2+m1XF2G6zMM1TTjioiiXnAW55/zf3yZeshBDV8ZmFbM9q2I
+pK0zxFxd/Zuo9/VDjiUeqKU7d3yml32n5KuLWnZFaxF1xXNQvsHhrUt8Yxwow21oS9dWxf2b7rE
aP8lKldvaYzbcJjZF/+gxHDdwOSNTOuzPuF0Y/WFfKv5bOj5W1f154QfREyMJbt5E7QRLpC0GQN3
Iknh1dftl2pZbZmfdVGsb4eBjgWfELRcuSE69wmTYyiEuUPEg3MWVcLkayH7qt2QgEhSUwoGxXJv
BdIfhMShv8dBvY4qMKXCPgNRQZehOC73/8/SICtjYG3IUNe0IRVvU1sxCw97gLZpGBElIvJ/AuW0
WKukz3VlkZsDnoT3UehyV2hqRddagZtv9zseXDS+fVYTfQPBYn5cMX0PDTTfBV7w9AAGFRbOQ/dw
0VFMaMFTK9PXMUqTJDiCjvKwxMJa03sxSy01ZkMoqGryiiXApWo7OLTmm9MVTp3135Tqu3EbFOla
4kRMFVoFDM34ldQzSThu0LMON5KBo1C+i8xtllJZIP1IdxSMxaT8xt99KUp39kU/dvMX1twkmu5D
nfXKDY/HmhkDUoCA0Yl0TpHuKQzYGoXvkO7DGZ8syzjIF1+O9lf7o/TWCpiDUX3kHJZH5Ha8AX2L
K38s7k7qDGMp2nsOQlGHNwJM4bIY8gnlpU8C50EX7VkkaevufMxmgKgd/Db7uUNFCzVXdMuTcl43
Mk1A0vhZkgxFMdUFW6MHkM4F6eBzlNTK4VcXcKyMi0zczZ4KrBdnmX/kArZ2xdTtDIKv/zb5JyyJ
qi6QlDiYVcigYtiz7exwXUgRQhfny/kzrcT69gJV39SsUCb67aNI/1eMi+cKp1KcbMP9F0sC+SsJ
ojoWdyRCuVUUB1Xk+LEhtr7eqxy9fIgkpqpSVBWlCRuscNbcW6kUZGQ5QdsxgHjcShBwBevHlFtJ
61AojJSCCk71zuH3EuHg0h3E7GIO173tiITEGye+vWQJLK45KjP9iQU/TRtjiHLG26IYJhwXKi2B
xX2JnF4hlev43JmVuhy7mAuo3ZUQJD5hTkAZZeHJ0/wMi3c1MHOwezSUCFnhV1Rl8KwwTlf46Owp
vJywaOxlq06qlnI5RtXvE1ZdlPfC9fY+Ogzm/Yxg6YPZZVoJkhGxl1E0TEY31BNJhSHYUhMCeWPt
guPgo8NudvbijkXFRntIspOS7TvhSaGtVNX67fEnZtgiP+pjBETW3sieunscT+znCx6lBUX0WhrH
f8PcWynXC97hHhSWIjah9xdI2/kXdhtCfOo1DSEnoRHCv9NE1PAgzb5ejMWBvQWem+BCHXN3Nwix
RSo635vpzub1n2iqI0hFfj0B2yxQX3q7Ogmzeuvt4nDogO+/lY7LgDRVWJO/6DIRV5t0n+gvYYoc
yf4tLNoNdvTzPVShU6Os2G5W4FPEDof1ro0BsDy27NvnoC8+azzeVrDViisb9qSpnwZZulc5fubO
cyWFjt95cm52+TSY4JAQvmch7gnBE8tZo4qlGaZLNy5Cure9haPxL6tScxgcfZRmomyNT9/B91K3
8qmJRY1TR5/ndi11lbM8rBprRa6c3FQcQPMGn4TNYxU36yVYtfhzMdKRPTyNua8yAo6GLH5u3GSG
syBlB+zdpMWwso4GJ7idbZ1NJ4PBvjdHacbidcftiaLlMT1m0iGlvH+P8mR+2Y35nZYFMXCyVr/l
zvgccrXHiIQvPktI2z1+1TycIhlRyElncg5+ke71Or12s6MoVTUe3zOW2NKxgIXA/oECiSPn4Nuf
kBRQO/NJRivpH0Lcqd7tr4EQCYy6czMoRl/hiAg8NyXw8QnA5gnONl6eo5xLoHqsG5jcCQ2xEzGa
ge5/8oAVUXgEJ0lp1OLCvnWozHTS7wncPaZzZFbohT/xWTp8Sf1CxLbI+O6oZ7ZjGL9AcLA9rj1g
uPv8JkrXLBhaAShMycfvduqkPLWMwLvpxxAyYw37lNYZLTm6gA7+ZzGSUxo0ckSxibvp4wOQHIMA
U3YT3X13J/nkEusefhmJks93ELtXSRyBRytwUtoNLbSI51xhsMeF6Cl8TNNAcSPtIYAL96IajnSI
iC7Vkb63gJ+kBcKQpiPz+rtCUPgyZYkkCeRujLdSj86vVrPE9p9VnCVpfmbS4vkRW84+ihziQZnY
Y/xWMToyv1EvneYNCrOoAGX1SDKx6FLF8wDImIoKV5EogtDdODj7xgunnpUTFTL2IqFnqGzbm0c/
UeObteLJ4AwJwiLszdmo9nbfkmP0p2cCo6yAoIrUbtq+MAunROJE5sZEITeN7gTCpX/WF2+7naVY
twb2YWEeYuOSAA5+ZoWI4bxNoHEvJLsGbnLBwEy61JPBRJdn6UUZQZcyCSfHCA06EH7uvcTSdOVt
rfIPu2/xtY61O9IYzRr7lt1UOHTVVGfYlE5f+cA1LRCHbxaNe4ZCTamltmudri7LXcLRBr+R1/k9
ulDxMYgf4ebWLF721IglSIXJnZx/fzFsm7/4LZgxKa8WrH90SSGqeJhYFQxTVlyrvuMmt25Uo3wN
7LLGRuf/cTQxLG8Ur7bgTLbQNFUGCIVDnbumJpxCmnK3wtyGO1eahbMgyXYN8QDaeoCMw9YjSaAg
l0018FtvQr31BLel7SgL1lvfxURhXuPO37bSTmxYO3YVtXHmAaw5z+DUu4fOyiL2NGZP/SE3ANom
Vk/lXFJ4GnUOyYvfY6XTmZNFcHlnxo5PDKlMrDKTYylDFQ/5scdsYZXyrNKbrwIHRt/KLzjhEUNe
tZ6DJ5cEInAYmJWWSwb824OLan7B8wkm3nANuKJHHpmf1g62nyyBKA4mYnX6kzijFEnbWMg0NFPX
7aGHw61WR3mMcuIm1MLDt+JHn/Y0eDVUOfwj0c3b77044H0YmVHMXa+cs3aNnHkQristw1uBBv31
5aa1NQ+DrUEHLF5xglsclzPKPB4H1i+O3Pdl98uHIhMDaA3v+hzuNAD0VNElZxqigJNvRxJKN8/I
DF8Z//SFM1zZWi8dgqlbWqeOiwpxZE1yB3CdtIuoitj+eX9sHUUfyR4TLwynlkMCSiE3RdamFiK+
HWuj1/9P7EPTZIKcb47hGxakTSArV8xAJkokNcB1fuyIP5IFJ8fRg/40yPbjo1hhIy1/ZlTwXITy
jX2J29Pbzx9tsS/KNr+6O6daDcr6y9VY7nOZOw3MKVsej6dqE/VFhvcOpjSdtcOkv6Ou1xKDdW2P
+Sp4GZ7RZDz6Qh/LUAy3KIF0f6QCz3U6f7nN9NeB3DPnYJoUcj8VLLznbqBmqRpjUSFf34WQtycW
Xc/aOPjSLdYQAm3kimc3vc2xX2K/jghwhMxng+MOpVWyh2EIAsOCHEEajT3LbM10utqv44pXAzOj
UVpGRFTXnoxCCuZW5uB04F7wbjqf/d9eD9lnFgIXCEgkTvqagqKMqBSyVdzpau8AVEpzKQ+Yi2yI
tZ3ZTRnnc/0UtK+BEoiI06hLu9me9FMJQhm6mbUlpmYJyrna0/cE//6KmvYt5KGU0TeVAWB5t1CI
0Y7O9MpR2e3tlb2MMYEOzALdVlQ5UmGEueXKoptuKoTldVAE3zFZSWSbZZ0z0QK18AgwCnYOoWc1
z7ie/l0CaCUUQUI5PsBOQwWX6Ids/4yqpBoB0qR/AWqguYVcf/GmQm93kHN09SjqZT295e55ZuhX
+EkBi1xlUdZ5+C91QUYt3Ld+ugxLnS61Z1ov99xMFFRe1TM4/X+FjgVo6yjJ3RCUARX1bOJ6gu8b
95sMK8GFiWPWE+FgBDjg92967dvlXmPuBK5IaXNikuUNe93wGRWjmpjZSdxrh+kxUyRjWwRepqAy
mVWlBx2jg7lm1185izHR6BF9apMlSNL8g8k0gqAHURnLAOOzCWBodPyFUqoHZCGEI/u2Bp4eyDyQ
i9e0YiUNra89XCD2dMDudkJ6CRqyQAc11wJWQdXXMnzC1pmYBdpISyCaa83YXQXGqmdeg1VDt0eV
TuOXxXcn7xihMAcyBJSNjXMtXbMjrYrfLN+tdwZ40JNST0enYf51/AzPaeJijIyZ6FcKlw/zymdq
X8MbFj94wytsmoxaYR5yy73icIr57mB9CDmPP7p08QYOK20vJT7nKvAD7j4jzQMrmDthMikpp/ki
eYSp0lcL9VnUilNH1w4G2SEfQsSw1K2OEv4jCQZU7b4r93HKwl4ghktHC02nKwVFh/JPCF/mUp8V
E/1ZHvEAa/WUELScz/Ddd5v+TMrjFE6LVM165GtjbEUIeF4Yrm2fsQAm0CM4r144cgxQjjWSPJg7
+stoKZMHOcamWa9hoADzURmy4Gmqd7rJvZwRvdZztjXyRYiyzfthsI2ZqB5iAJ0rZGNVuUIyWuMw
4fMOUCYmqH63VdwuWr5LURqhcXm/YlCN3JQnhu3lafD7/75cBx/KKQE3IVPzFNsk9Nv6MZoaejA6
9vMln5WAz6rWwQtKnsLVZAEa7jG7zi/ZRNWRMGs5uP1/GxZVxPETJ/87il88b3dP01GgYrxPu2Wc
kx0ku6PdNDrfBG1c062xWFu7kChPlJPMWAELn4B+CiAtlogLijGLFDIz7sNRGKytWEbsnlhWhuKE
cR43aC7BTUhYomC7tlsrwR/GYqLZTsRWSQB8v9Pv7a6OYnVsXqm1A25f5DZIMdrbJMs6clZ76CSQ
gwUDN2fQaWkWKM3+yjik1XyrnatVNSDDksW7hPP9EHU/MlOwCZEdbemeTI+dLsrLbSyHaPwx1Yyw
261w1/MFzP4UlLQ7FKBGnCLWr4hslTv3QLJqZaR5LIgSe3rgffrsLHpWOyZkiHrnGps4ruQomia9
0L3dXLwS619pANjdkofedqm5NX6dZ1lUMzpw9ey+qXi83yUpYQbu7z1DuAtMFGZ/sVEit9qSIkQl
OgRqFOqMEa199PgH3nSL+VEEmjTI/Sz2Hv+tF98X8M8tIZuiIRihPXdCxEQhBHg1YdWcDlbM+Rwx
V3oXj0XyQDJ9MvbQug80t1Tak2HfHPJ424RSLmQIzieS2/ZYBpYQnRn6PntMI5KGXSUCehOARpsO
QWJP6jUsaeuCqbQbggeLO/cR28SZru6rsacP+M+fVoff/mWo3xvxpnbTgN+N6hp5IuAeSOrjQezm
66O74C2dftg2L1Q6x4Hd+bUKYsBEzWiavY+NubkURxjIEPaAScHNX8a3PbX7eYZSrivo43mUltNn
vtYCjq7Zk3X1EUWbRB5m3E9Vd6Q2T5Gz6daT4Y5ieP/MjPPO2nf+cwVq498cDW+WgkvO03KZvy45
lTumvQ9trImHMiEjln90XPKUtLj9YDDkxybg7mCuf6Uj4/ObOhoqC3VUhTzUjcubqkddi549sC4n
1jnHMcNL7LEH0rqP4Rur3Rg2/XhKgkpn12TF51xMzZCh3brZnblgfokHGHVnYe3fYoOAmq05acYn
cqWfMptu31LqCPvzQvRRZIcworfDq6FjdEDAZ4udWW/Nz8DK2tXpsUZLq+RhnDiNTJz79wrxM8gw
T8H4+wSJ7Mq5TZnrhifVEp36ADem6Yq44F450b8b1zfgYHKMZVgt+36M20eP6G8pPIlZp2KypzCn
GDpCYOKLquEaMDtcKhp/STA1uqg2nzMJklrUJSSChOEuFRfJLtvgOQNj3dtiYlTnoFh73JsCuAmp
cYTdPBiHoD7pJ/tPU3AoJ9qWIiG5kMxDBDJLT92n6vtcuq9GdXbOqS6wp2aSMpmb/t92nVhDAbEh
Z+severvZO44G7g2TgflfPKVeH2zVuT7YRsR/+ibL83a6e92ktaKLP6lrAW4Hm/ItWcQxQH1QhJY
j/p4ZRNb9MhdfitJzD7jNqJR1Hy58IEJpX75HA5z3menSQnwzqEx4c8cp1o3k8ltQsibunAWfFbp
N0cQpiVAk0XvuLQUrAp7qr6Ca9jiokeiP7eOfBwAHiTgAT0t7p2AHrM7rfyiFQJ5bMkfVH44XCo/
QB+59UPX78SXQ8e/eOPq4IzmFlT9TZcwQYoOAAX2vn1CEm3+cHzARyyS+u2iYRbnpY54sa4c8kki
LnGLbw9pYkkhTWY9zSiiMwtroSJT278l6GxcMC+IH5Z/Y/8Epf9qQhJYAdipKSfMRkC51w2NpuQu
ScFt+lHy/a7lHnXi0DGg3G9QOCQkDVek/I74Kg9iKwFYzEIQam12TutJQQyKfB7Rp4mYVZ1UJObZ
zrhFyCSj/db4L0p08pul6Wm3Cs9gbQmE2WshOB3QgkFr42cTYFOt3cRzS3+7yk1Gq1HXWDWY08hF
f4LKkfrSQP/OBSEH2H+TFNqFHf3r+0IOYfglTPy3oS/rtegeA/E3/VQfbnZwuUeZoPqgdZALMu7l
NsJREhkxQKY6kw6Vx+iVH1WyvzmcZ2gxY4dm2cXbz6NQ3uqjwh7VEW7Ie/neEfyvvR/RiLEjf3MY
F6uE8PN2TqwM8p0BqB1jV/9wiVpik3rmW1FcG2qfJiJbKNIP6JkUo0EDOgMe4w8OnTNMYe52so9s
wlKZQOaE4OON4aabgrUZ9u2sVLNduM62ltH1+RhzgFqOBUe0Ao1aQ/j6LdKyk7qTCg9KQCGVLHhz
aNli/disUK87Jjpr1GgVRZ2RIG/JSBs3O2H7C16nQ5Y3YXCn7tEUSZSo/BCOzOOkxoQmjduBB/Kt
+pAVPx+yoWvgx7hs9VA7lowpSBWxlaSUKpa9TidhbTAvnb024zdQqGY0tWd+XXuIi9/hnMtolwPz
GRyUqbT2qMBcUkifWeRNXd31noG9LWOrlk4St1Cni6F5FT76qb05bxdEDHPzV1SrgrlbB2yZvHQx
xv+OxP5JVIOL87J79hRTiFFFxkc3mQh2hTMAFECRnzf8P781WuOiUt0P0lrxp4+brMPQdmZMy1b+
KKMy+erHNhVHrFOumwI7LGDngLtXjY21RagFXIb5AbrAiyNQ8HYGYfBF33jeceNEJ0GzAPRvHmHt
857jSWTBJ2BPDdYdbnbKngfHpNRWYu+tyaOGhJ3LJMpTO1JG7hmXx7oG4a3bY1tAaMTPt4HxjRu9
+mGklQOA/yyZff2H8zZul/NnQS3gRKsGHIpNmnipjB/NKyVro6O6yFb+6s3y+vTiwGFLisrBL90I
JxoZBzlu3f/eSFgJviGmHFf4VVh3zIXMW2RfSKaAoCFcA/SV7TKMdE3gtijxZ2KT763gpC1GwW5+
rEWU239ejrfyIYqRJqVv6fvsDXOc7OAfLNRiY71R37LH+ijXUAvSeR9TF3NhWA77W0roBsflMuyE
JYFzR2E9cCHxtfr4N6dfRJsOcioZgNMFMLjErAqs2OZJ71mkb05Vp0YgcmW+5RY3M4q4RgBuVPS0
rrxOt3KmLc1Xv2JEyJNCM7K5C6KVhGpZHurG2HF93N52KeC1PBP2JGsWc8Kxi9guAwDcgmmhi7sZ
P4DTer9ZjVtjFvsiFG/zdQa+yDmBC3CKGe/BsnAQC3r7RxKHVt4QNXvIwrsSBA0jz56tP2diTYDx
/hhFIXm8FOb4ix/cgFEJ3r5/N/b0Rd5ZCVntVjvZZNRGUBDLTMzs/KgpVHfRsJAccnJWdscSFTn7
5QZrGvTijJrBTRIK2Eqfu1jl6bdk7n7N+A5wBXbPwRze3OjiGhQFuLQLUoYfCqshG+xQeFW+vkT/
JXXpolbnpC+l2V28pA5lH/h/0UXOABHSyjJHvit5F6u3cRt2c4qwyLjTxFFgUFmFVz1n/z4t6n3Y
zvpURCKMnSCprfi1cvsG/ZUyUgJSz/+VDRz+gxlDpDUCAixO+Fnc59czUaljObVfJSDx41vFnIoc
tW9C0bEeM3I71nao1GReLStgu9IUgFaokiHe/enNTIbAsL9jk7cLOMF1YurhRIbyFr64ExZYQfEh
c8FEwKQ+5gBpAGA54GcuDGodPFWKszvHJKONVBogBORdHIHvBGT46P8+ZSjVVuCnHmnaAdirXvtA
FLB7E4xmF3TYmX5or2SSLiG8vqdwMH6hZEh1v0zyNM9wJ3UPgEdpW4acrW8qforQuFp7ruaZf11b
8QcNbQMcXBUlULqj+z5FPDpBp/0XSXMM+49NjJtWUMgkCnoBjpodvo/KodX238yrpum4SCgNyFl5
FdQUjX355hLt9JlRu4whS6c42p6w/Wyujnt8yF6syVrYfUK37FyLDm0BYjGgrpPIvrZ1Dtff3UXR
tspYo+P1UDBEnRV+uiUNPTnKmg8HFq7y072tJLTdhXOqcV9FfZhXLDSua2qgtPwygeqUliBVCGhI
2RXybuQ4t2/GsP7DJqB5199meZ8+a3USaGhnAU0DGBtlcEWo3rNx/Rh5Ec5zJOWJvoXcAv6sqCLL
PPlj1tg25wGXCCZVPn/k7s46eTj7qdaDn0tTqSLjb5YYBGrxNXLexjrSQIo0A+rqY5uSd6ABJpo9
MieItTmNP1du1cu07ojPjs4NvQAsHcGSyePjXPs570BWnAoKADFYYn9tR14x3odZhYCwTmlLaoUP
XpdU3RR3UeZDgB4q7j34Bh4MxZ+8n4kOktRdGKaYlJM+XC2vE5yklYHvC60ku8cBUSdlNUgSMYz/
n7u+iD91F5M+NDyUrxBF+M6OTfF1w+nhTIUGQGM7YP8Lt7MTmp1pR3OUI/W2WybeI/7M7AQRbKMO
g6KhNND0amgkCHJhevKoXm9YoLLuW+FH9xO3CSRVBgwiahn5u5JMsIw07NKmjQz8guFsjRtdgjNN
eERoHd1ev4cPaqmSV/LTkBOCVyos/8vlrw3rEi6MwqD+wo2l5k7TvGJEfijRvMOmMVpsS429+qAn
+2n3V65Fx/4m4V5T5a8SIMp+9osUm2xsHKNWv3XQ9bfRVU+soaQ6iHQ+ktBKRPLtvSCkY15aZM/9
QkOBBxPLOHfLSc7LzAbnS4Warb8xWw+bASUdfPbY4cxpqDFcCW1D72EgbRRrQoBVPqdqMlOmqoK9
yQuvfSqbkPD5o/NKFeMb1IraWlK+pDFrbjZeYOWrEqzcwRm0TJbjoZ+tVEyt/Q3Y79zfh15Z1Gtk
sgvAGL3xm9sKL7O1n2zRlZDIJv6SCETuRrof7P6lF7a9BmokjHqOsYtZuGHsMx/qKfPjD9ce055h
TTPMaLKWnwO0A0198FS+i13O528A4IYtjbYE/0TgPsC8MDd/Najux9NAklbXkfRPUK9T4e7lOLSP
UGtdYsv0EM7SwOTETH8dnYPd6OWcs+yiaokCynZH8PShtnhdzDRpdSKzDhtiTCxugoZ0Gg+mVTQP
ab70RYoZcuqCYk1oa7p/roGpfChDygXicAFaRVvwPHZUbjR4EmGlqrO5cbXnI+3t8cqOLC+E7hQO
739b0RmMGtVwaQ1zliPKqY3qJJxyJ/j6E1lQGErjFFpZwelBqu7onzyRFMR8AmcnAOYh8Gfe2A7d
eGAqaOZ5F3td71Pr6VFpODTFB/DrsEFt6uYACddaDz5VbVe4IPYSxqk6ga/pLiItbGkeVYvaJyef
IHpQunakB833DUxDFD3UeJOeAUtiwvmPVOEdA4Ei0D7glTUC9ljl2zwy29Makcb3d6EDyJOzQu1l
KVI1bjAmtmUPh4aewt+UeLlZ0R7LN81HmrbnMXfQeNPhkpwUoJuKr5/m9nxVEfgf3YZuQY3MjiPB
4jqwmQ/FUly9kcSDN5MMfYFTb/aX6JqbSgQ9jLIrk6Ozdqdp/Lr+Z+SwIvyM/w2qSuVasYifJ6DZ
nVRaMrvhCczEnAPNjLfgYKiEid6gHcyPq7cyv3Cgo9LPAP7910bRzfTVBWsbcmBMzxLGESHphj7l
+8RyGcnNA40f+Ajsftwqk7qvFMKCHXTN0z1umRcCTElRk5Zp7YfYUc2cKhcrau2KRlyeWLLzQ40i
7GJt0sw0bRNVtLfGgcppLG85GyKG0nK0xabc9dPG+WTleggzNAG3brV3Acq75kUbnR94iVLo4S3V
0WMSEfSW3w208NO++8MEEya7r4rr/VAifYBkRJQN7KQBazVMP0IIq1F0sbZogIDdAw6KCEF4OR8l
Cx9sjKlnWOR9IZrJ6Gs3c6gJiDELBnkVeV8gGb4MNW0DFBBBRzaLyHukm1pjMQ6MGPbVU0/IyLt6
rPUO/IhxhezqJ6uvlUvvRSQXZcwp8J5LsZhsGkG++IGuuDHC02vxkYkGC49ZWfeUQpcd2AtAKmm9
LAuHVOmxorqwhpL/fY7qQxzJf8UmzyFtu+loeVZB84ge8eO2Id9u1LGqvATaxGZC8oVw0+ASiq+/
rmdrc4emTGwaDp39BgcZB1oif+iGX0g1KhLITXI6K36He61Fr6H07O3ssatCVp9r3JR6duVIqk4c
7lkJJgxUVgZZmsRJGKIHJ60n+r1v0l08upT1T+u20VqamO5pYVl6YSr1i5Bo/JHN1xZOPiENof19
CFQVRJguGnc8Mpj3eIxiEeHKzrhQaPX+r+AfAcMTReuXFz4Nq+VdHiW15UyAgQkGWN+5K61zp3oo
fuMuvHbNAAYlksInR8aFaiqxoFua2x9m4x4EBk7xK+MQ68TZbLu/Rvx2DF1GZajB6yqDjBwKEEHq
CgvYnYhddGLF9++xkjccu8Qx9TTzSneEWnxo+opHd807/Nf8zr582zqoJo94No24k+n92IifzOk/
zlGcApTTTTG/ocFpOzrReCcC8Ch3Nh0ahB5GiXLgqJ00uDI0Tqb1QFy9aPrF6ojrl8Eg+XTewz3T
auRahE+pY/QEQRjAyp4WPF2+IsBhuG1UAV8T/4NbuQsmf2AxP4wwGnKIt0t91YRdwBgZB8b0gi8e
mv8Ni2CLmL3zFC2f+Fc9hpJKWdJ/CIs3PanouDTnpwsySszvoejfvC2RaMKAKg27ZX2sl8vJL+nQ
897NUWMbhWV7q4hdg/BuqSpzhIsZBOv4KCq6jrNYzxgigjCapHxulpXooZhgie8WrHTAWTMgFvUB
bdKAsxZlN3mN9pi7uWBdDRHhiigSJpeXK0GsA6kJsH52O0iENRylpMy5S4pk+gSw698el8jZIp3M
FEPCDfXDNQkotM+o5dH723hmQsHZwlvu8xT0QD4d7nMjRZb5+1STFlkWXjSJ0DnbTdGGLEQ+D1G6
0SB8jXXO+OSve6cMggO4Rqx3GqOfltKwJh5c1FcSjJx4dVnVzhxhaiMSRlwu2X9hCDyNqaBQwyNI
HeVGsYuylKZpZnEFh3QxkGbMicObv3xQHVaurMWJuqyVqUIxrPUOJOZN6hi8g2osbPqrq7jf+NnC
U2jgiu/iymTIKm4ajt+EcAtT+rqqomlclJDC8vxY/2FLW9chLspMphuhxvoHP0Koqz7n3FWMPXU4
VSEW2lFU3sZt3BbMYLqggKgRk6v11HFRohp64+r6JWT7yqdC3HarCrQlZcF2kk+NSbtomcWGvOhc
C7gyEh3WiWGLy45bQizT2xDjumd/AOElOoMu0O1XXpq70Vs89Z3J78/Z1KJcvdROh7j6auKf+2RK
Fv9GCLMc3ZXPZTt2uyX0eIFEaR5/ozriz4WM9dmSYZpuGuW2U0Kx6p9fEfNHQEIxRioWstQ3WSew
iYaHmCQG3OQXarZEfV6DomcuHPjzBE4uFH6p730irJs9GGPbUugRoKzPWIbEjWUObWlPzVKfuI/x
xRlBYorfNKCo3+pbaqvbuwn8FQhP6PRofq9Qf/fYvI3GSu+Ka8Mc8NN4SCD0scXJbfnQ2n140xv9
57O0nXf4XdzbjcPh9akdF2w9doazuDjZFZdkh2DN30bWRzWYa4W6z8BHu1BDtoFb0igWgbw1myhL
q1tGM1+Jo5rB9/91GyYhG9xuRfIbiOA66JY9ZIig4mpkEk9Sx3FPIjfaOP3Rz5AB4205w+affZ4I
dp3ChpyRup6d+DiPSROci+jWdqVX7SRkkimEw8kRhQ92GMA8W7kKdzyZmxusbgb5KUcnrjUMjA2p
DkKXdEUYqXGYWbvlRtdVPmwsolK9ujymoNABkQKVRjawGQT1Ls+sfOdFTkaNg9sJCm6j+zqSGMlA
MX8GgcwhrZsYvVSVhWziQ24R9bXybg+rB7ODeWrKFvk08Iud1seajCmgTmcixDjYErxYrPPmkumS
PZMqWMPBdUQwWiCf9RupsYp9bZU8Xt/GUp+5/v4HACp8QySb6DmK+wCiXwaYThznKWMqVcN6zM2O
II32LzqdPDfh5Ey0aLDLoPC1cO9Qy0CkGD0ttwjbNxNZkf/iMGH/HXbAkkabIAVKMgdnyc0iAQxW
v0lJx5bpvtRINt8yd3t51/q5/pvV4wu+b6NAFQyxVxnLL0T9mhIJr2nu60AH4RA/aEnacoATJC4d
h2UCXHwvMdDsDbu323RuEQuxqYiPuzrWkKFB2UNnPGcCToBuZE3ei7fMbKtdmHAt6+OATEd2iN31
DdRdsSsdedbGm6i/m1+pnqieRQ0ke9mdlS5nFchKjQNYMCCgotOdOgfm0TeJEfRPPf1BY0peVJB2
p+MdVO72WJ92PmqFDQ7XPf/GtzBRGEvcCnRgs17Skq4QKCn4Gdbg8aSTR1sbVShuzEKD0bt8opGK
3W59e++BVXoCX7W+fF8+qLl6OFt+nFnosXt20PqMAOXkjG0vqL4sn0JKKPC3vQxmEQ5QUuwtqPId
M0aspaNt/5WERcebdFeEsQVfZeEWFfo9ZYLXM36PbXEUPhiP0NaZu5nvvcUCjP1wjTt0CKNRs5Mm
sEa/m/ildVrXnZIOazIg6LMUMihvyQ65PO3mxBG1mo4ba3dpzd6fgEAs1LaQHynM2KfO2JbDQ5aV
TRnFEq+c0up5fZ4xqWnezgFjfHWHjOgy1Qi4NdsvhQETopKuCGWbCGbMvEru7wBKwRCZ7AeSnsGQ
APAD6UwX5q5yyUbW4nEeFLxOCVneL/dcanHxLtGhR0e93iAxap+95MKoteAv1zv4zNDfAlfslUy0
4201544gXmICsyiGGN+833YlklSQ0SZE4meNyzU7AN/rFNYe612XI2FzH7whdj/UHcc8DaNIlxI0
5wWYY/dhVnvD7hbWDv1JGkpf6fU1lmh2xRI7CZjK3OhYMhD5eo78BTigZ8/TYe8zo9ebnTFCt8dX
tgFEdmWlQlX5pvyLDavWD50VaLcq+mzlFf/I9fy2tBIS2+mjEiQoZDNv5HnfmgOHLX5t1kOVrTj+
jSg86MZjwKxvd+p/S0Yup1Ak+QIteKhsuP/+MlyzZEtNyulCtVG94x9p+OgXtU0PdELjIF2UeNTD
eAio/Ye0+wybvy45+8WppKPkk84fy+2MS3R+S5n2oiLZTgij7cDOICuoeGtpYle6FoP48XKvz/qr
wfG88VFUox1wzhqKWhFkndW0f+KsKkZGCEfKfIGGI8WoBR5JCvtSMugI3C81SYpSzmMWIU/6oQj5
DIqjvc+oLxuVjJvJq3bfSd3elKFpOEKyO0tnJee2Dyt5Yqzg4mgjhDSY1sYo5HlrF2WT4yEurbmn
FTNFhdTTh5UgfAsdaNoTBY0/2gBuZnW6qmAkDC5X6gqzPhhJZbaAPPd81fNcu4hW8wQJIsaJIPBA
P6bfrUfQ37DMzd6SQAOAdmCofOQy5i2pM4v4sHiggSZcZcolOWCFcyIkesj1qFhGHIk48sJtF5qS
aP58DBBdjOG5EO32kS6aRx/Ayz9Zu7AGWLGzyP7yQg8RKtPoLtYI0Vc+AERZmzaIRLaTuDIZvDS5
h7Ok0NGj2E+a1E8uZ7eCK4K6y8M5Rj++lpeL4q1XbpSZTfJB3MEuoPBGpkNHoDs82L/iYVz9Dxyz
AXbW4UJiR1ZJ7UrXMin7M80I4FUT5dI+CHtxfSNdUmKD9I68oZLIpXTWtVJatwhzJNUwDNHoqJlz
lcB7XnS7Fm2siBm3a/KbKCLdHEJQE05PU1a78VvSQk9sidWNRxMN8KtO4or+rFUjTybUsbPIEzGs
EpARWiPmG4ICzBz4F6NCBp/F9qauC8Eqdzyymmf2SAMl3iMNmCIGDM2vZORtiV1Psw6MfoI8RPca
cxmMASinzEJdqaUOOuD+OvHUgwk3ufLb7wqYlUJy/o4RNMNcOq35RRDeh2xHiR85JyD/CyMoahEM
3DJ+8b8QZ/EUKGx3dcqfmg2Nnc1Ok///mbM6o8gy6RfznaAYTEKT1xkuxBgZErGf9bjRRo7la6px
n8dsfURNiKRz/BAw0oXef8gl6yYD9uD2ondD55Dj8okRSp2VFuD6AOoLlYZ13X6c7/KAfkGzTY4Y
kQCdvFVjOghtbJXD68K3AmMGtaYrELHWaJpee3m6qKGXJrKU4WlLl4mObZpFqEtVp1JeabrFzfmO
B9NVWaiNUN/RyeuP+yHTaCWCYtEYZ1Zg5dKHdmNs7K44kR7NGSzR+qI7PH31K8BCy+5XRAfT6Y3N
9Ot17/iGWjThZiDcciZ14H9LTk8cX9/H0JGdPdGlhmJ2sWJGRkALsjV7YFRprTis0+Hw2j+cFxCD
0lxZKO2y5Nk4WghwDijsEHHScj6NTq9OdoigdEMq2zf5HHZWMX+Sik1RJVTxJ1/kutCYEqLyxQXM
AoxrKjrusfdN1P+OXBwIlzjKbrNhgrDV0V9hyRSYhsASNfwhPz/UTlTUHI010aYCPJq9DPzyKu00
g7n89bg4Fl328CNKHIf5i1Ik2IZCng+3kg1e9edDFHFd+FHm/enAikeNYkIIBupt4agi1ZyQBPwz
PXZqoTJMJlvsNuiWda3uDhJCJyhsPonMANKLdRgMHOgxSvYUBEqF89m/uPZYgURi68GNQ61DwVrn
ilB6PieFSK3Q+99KVH2qixb9+HFN6KhUaPdngA/8U+1N0hTE278EwLsyewSb5eCd1Erfo7tbKcjb
4ObOKRQ6pLiWy7iil4eba3iZ+TGFM6T7Ufp/xfN+amlldVK6eOpl4PAhJ6cfNDCp2aC3aogNOdl3
B8kuc3zDvNQkE6onokL7+FJ5nwSiZ3+CupdPeqctufMpo6AohxVGWjcGUKIWistuUbIHImom2E9C
tLAMfpz5+TmAeiexI8NSczqfx6hDR+T5IkutCQVEIsPVGpNbQxGZFW8vnxIBxOiMLnUOYR4tyu5B
j6kRYV8O1vuUjzMRusD5rcObcpPWNOgm653dgPVvzx9sUfWkyb1YrZBu+kpIfVFs2gZfC3b4u5FO
5a/lS7ppBhDtFYJ/y8svCIy6/LzB/iTB+iG9VuwXNSNXoA9Boo1V/x7XgtOtLNrHsAYOMi9PnZ1u
2ScalXaG8pXICS4akF4/UnxzCEp9za3WyGWjgBEgBjB+wmZa/cwHFtjZ3vLkIsKp4Q54wLg01cDz
WsjePSdDJwNKkuHis5ZASthxc/YOXR8pxsMCTVNldTjCrZpHbpcmaGJSgez4mf0riPPn82oJQmZn
MHZp8KlOedsBjUoiIkQGYn8XcpA9+CB1VIetfK5spELWb72eQ0gw/UfKp+C63f4tgprBn1lvLu9B
qzxOlbKoaM/dQXmRJ7SInlpoiHRLJFcKvXvXQYL17Q49b37bAwDHd8OSYRBE28+nTS643YoEj3ux
90ixVsvakXTb5xe2ppOVJ4oU0F4KU1ScMeOUhNE4um1VZJ6vSONITFnXFrhWb6M2AC3tZttqJ6tc
XmmMoWphfo2PvipUMwcmB3jNvNhQO1bKkXjUXY4LygQp0so2FO4IUYcE90mQC+aC6mfNQ49qbTkv
utkJW82Vy/0qmDRtiVFwU8rw5NX9lXugJR9+X0DH7jlodFo9DblUQzwJ+/eUgfMdAvrulEAkq4VO
pryVYvlWjT5q4kOTxablmcTtY88X1p4dfc1XQbUzzwzqorWRLb+2rC9MiNwWVIsxVj0PjQ88DpYB
0rdeE5zhm1HG6EGIfb5bCeBGSFgCbWM8jG6t0hrtJn8FY+JZmfNi97wT/xdDHi8ANqcE8Q3/zEfH
+AZLYyd4SDIhL/lPrPTsX+RqrHWei7VBverUP5FyUQk4P/kpIla+ridiHKzcu4i90BGxcrL/8aa+
94XJ0hDDYu/KYJUsSdivOiZZw2aUhrrA54Us8TNG9ohPuuxwmFg106ou7ZUMFOFC+cJJ0LRdWF/p
2Ehn9E946amKqIhqGj7+zum/TkCsyzaogdv5PcU8g42YSjVvLETD+LxqtXq3duJatzDUCLJFPIlE
HKegpsEfTo5nnfA3m+0c9q9ofkpxR1yBXGuib38lcpt30jRkt8obQakeC4xQ6WKiPp8Fl7ergE/b
wKtuDR7YX/Xxe7iW1NVctrgprTnE6Gz9KDt3mPkIMh6FT23rNZVPpL6S5UZJB7RI50RuIjl4S5HP
TnRcL+6lY8Git5Ig7qmuEVJP6Yzhmmmnymrx0iUoY7vafihmzKdGviCpox6e2caaD906hVPCXTmn
uW+1+hFsd/Wn+KE/7cAjODkqhJaagxHp1We/dIVV4qEyHXFfBOiMN8U6LsunZO8Uyc8i3QiwHBx+
a3v9zMdB3ccFDEP9/Hizky/wNRL+OU+qaspzDLuxmsB3MgVgsNoypaMjHM+L1ItYIWyUp2FSJN+W
r1nyUIeut7E5G0a3TvAISAMiJlKeXDCNnuaCpzSZJSVkYZ7QFEME0qwpaA+50AudPLPFdScZW1Jg
OY2NnmPFbrRC3HjfauCBAv6BtNFZhpnwN9DKyan8ALhoqKCKjYJht5tW08WvXcdS0UoJtOqnOn2Y
TlRdllh+86XDeb8xmCX6IEB8QctWm463qILYS8dMROOyMNolfKjnJBP25411yepcN2+UEBFSYwdG
knmOnT9cWlcKO4x0kkqncbDVjTdIcfGNdX1KD/BG+8S0aXzriCgjgnK1BBvh/98a56mGnZR5EZnf
XqVa+5bR1U6LDwBWLd23uNeZ5zbzRqDByLz0Owj7kd6hP8xao7pitJBpbC6rY7vAj8bWLPmNhU8y
ArmItFhMyNLCIlwn3DP4P6yjPXFJeLdTPb7AcrMwkQwIxGPaz6EDLPT1Io52DDiR1a52cxA0p6HY
+gwCbMT9m1MPJKMCs0vBABblM9MIveGoCFMIWr1kUqKQh/EgSSOA+6uOyEfI0XCqyGe0DtsJLDEC
9sw2a6bNDk5alZZBNeSpc6I79Lcv1eojLQ8pUa4er6r/MGSHTNWIJUNT2iWD34dn+FB6/E8c0dbm
ncs52UcTNgsCXZ9vSB5KLBrWJ7j18PloYTLrir53YepboOtVptDBE5X+bJT/fm0QIfJz4I/kGIl+
3/LaRZ13tBz6pKD+8BEEFr3Kc0Jm/Zx8CfaE1AONze+4I5Ed+mikONqbH/ckvINap4IQ4X6xbMph
is1bXFiKEcVc2fg5zbzI7Ir8J6xl+yi4ZRc6JLPTswIdql48IRM6FzxLspF7QDITI6V5a36uNNPW
h3X/f5kDapHg6W92jjXPQBBDFvQJb6fQaskKX5sk67gyHr/6ll0PYF4pYr/HFI8SDNn4xtOFQK7B
ppfEdUPY4lceZPhoBRphooPYfXgiVs1a9FxR+PtZNG+Q4Wt4GOa/wriQOaLQkNT7TXb5V1/vkIWH
YG8waHPSYrzJo9n7/E+kPqoIbEBFqX+P5lwhaLCDMYRxgwpTcPLA59Z0KgLsEaIDtTnBwwBXj3u0
9IZFH4TwN4jidFLu6iCowGDnvjQNmO/WM3SqYyatLdzT0Hu7okNwbO2n0Ohw8fKCAxcYmmq4DkVM
WIQ0iHE/w9FAehXzyeIkxzn+iIhJAg443v1x9v0FWP/aj0bbKaygeEqyvnJSiXlP+6V4l1162JKG
J/wFYy8FINzzEoL4c60+uQquA9PKAVKICWATQxfAte/AI6sc6i3eor+YFchK2qsYbwV0mqHCDfWG
MCWT9ibw6onWqIzxuYD2ppjXEsJciOrEdVixt4YC8/e0StmBmagKkqtVEecJ8fr7hJjpXq2OCb8M
7uvHKHU8K5pCBXLd15eVhP9Pxww/QW58+uG5m/kYjaMXGtJ88KMFope9wz892p9e3xHOsX+8Qk13
Xlu1aIFzgw9Xzxwty/B4yDJHB8/zo3ZdOK+UWRAT05+O8+XI8k0faF8+7KeGdODFKljD6+m5mJIP
rj+J+5exLnQWSy3OmvOt4JWl39wfFE2mRM+sW8gCTRmgAAf5/hqui/VGJ96lEsq9FXLsQSW0fo1R
lxueVk2i5c2ipTYi1U2DxzKSqwB6B0pL/dAkyclVcqRUSXiQTf3hVPGlcqPYUnBG8zbKP07yiNbS
afThNU8Ln25G2u/g0eN7d7A77idOCwqFLZGWDIpcPMMailzu4GYbG5N0S4/fDud8SP7+mvIMwRTL
nMe7esnfhRbfsOV3KC22OKx9qK+BxstKbPy6ne2so0GX9J06yxc9B6gUgdHr8B1hHEWonLBJ5h/Q
LlzDcmrbJ9gzGp+HkGwnyNd3wlb4ACHYCZ7NLz8jmKiKlzds0ocRffd+mWQu+KbtxDHUgoZqUmGN
5bYW7cbvWtKedYSmOj6GV9KZ9YG2PYpyLGqcbID7JzvSPIAQOhV7xqGiDV31f7TSTZNlh0JaDrVQ
+g/KD0X2IXviCP3ZN5/EITiOYKI1mA7fhbFtrYLZOUwqGo6tQ2i2qkaMLQ8xThOr3Hu07VElG1gv
uSgX4pqQzpndJlbrxXw9RFm3wK9RaiwL4Pfukkgx70z6DCIEXVy7egXsPCGwSncslmE0StQHb3u5
dsi97cttiAZLMebaKMlR3t1d8ldViLuuTd0mMzkzXkOOdQIJzh34JXDMRveZA35CfiUhUX+7lx9e
A68m+vY079uWm7iTq/gLhSGyxyLbAq5Ba43pdZIs/wKDmiOXOqu8dmg8EGakbg0L2hAV2L9oNioG
o1o3eeQu+CwTlFJ16WwdMuPsj2fctnRxAhQ4Ff8khpABx0uyww6WHucDVAApvle9q+TuWhrfQt75
vwsmdPDSobPTPzdElbfiywRaD9rtyvJ6K6t7xdHx9B05YwliOlWfnXXKMLM/JjHfCiOZqmhsZvLW
scsVB+8RyxWce1furuGxVh5FS6EK/a94u1xHLXt96hREYp/7o4JBVpLSWtQI1REtjR5oV2QI+50e
3dYfXPpTYu7vE+uOiwOic1m/zVikqvhqrR6slZ6bHdlSrCeIGcYuHhgSw5PMehBRfcqUiHbW/u9r
n7W/Kc7qMf/1ZoRYrr//QHI/oywzVPHFFhNOwTGTy92E/3Xj/1OSCAhZOl5cGTss6+/CJ3Inv/pk
l5HswdfA/rFXhVN9ea5/jDShSEGgzIYjRGCwqau1vBtCFKhH6ZeTzO0CuNXRk2I1oPtyt5ff2iFA
vhHkWQwnWQUI0XUsAdC2Gk/fWZ+yx5DteBSPgFHOrq7F2O3YBnfLrkqM1RqN3TWBN3BfeHB+CBg6
7to7JCFlLusLi35IzU2YPiGfasmoUV5ocO5B4WPSdW24zmtHNNnNrYwO8Vh8ARRIcov+cduWKCSq
1FfC6WhM41m3oH9KbXXjYrGcyxfF/AmqbgiDCjA9/URa0WSDOEktU2jhZ05ml3wXYObffkbBy5aJ
ScgVVocdi9KG3FljHFku20Y0ACjbA9N7wSWTJeOY0O3uil7moX/DsBGIQhRzA8aDuYx1m8yAUfb0
IAU/PXqahEa8V9wmHUJXXMZekD3uth89ud2F77P1eNeRTFCMxB71V4LL0f41VUNPgOQQ5tHsaDXp
X0ue/hIAaheVRRHhIO0mXJJtuZkF3LPFa/IaDGLbQskArrKaGeeo+90sINUYz5AwRGzJAe20MtD3
mhFrHLTWgnLlqRIQEnFDAlaemnXlWMWFkNOomFpstVEc4kZGbofErujvgUAEGC4Nu4lavOPRe4w7
0LSk3wqoe9wLd0aelyQdaH224YLqv0LVQnxoKxZm7bZ1rs5vguAPW7GuYUMWCkdBZK0X2hL4WS9u
obYEqAE5/3tiktLyV21LDK9Tnhns3hsZPG+csMk1k6SznkmOYBoeaiFK7UZyDoEODKHGKwcP1eJr
UDk5fMfc8J68C0rznZZNKdYaRbcI1OKfOZfLYnZQcGfvNQtl8YyroV+cC2OzjUI9xIHjO/S2f3YM
kO02ifR8dm4adpvf4fjwvM1VPU486yKFpOD8qSHdcDCiqTI0R/QOGguaByPtH0uGzJj+VRq8sMDj
eZneWMhWHxnmGZC5J3QbfQ4Eb93993K33j8FwzBU17cBUuPhrKaPbfpaXR0giMJ4Y+w0jmX07QVn
zocN4V17MKOO7NAJ6u5jyHIhGZR9xaDCNdiUT6B4S5LplFEqYDSc5O7OiF4PZy5xh0wMxEYrnsCg
NpWCQHOBgJfVqu9cWrNPrqxitDBcCPIFBjZbGossqfPoZQW0oepL3ZItCBB435p/Vbi9P34CgkdL
glFacyiBjvhd4bqt/yHd2069yfX0tR5nf4Gc1VRSWb5vtYZ5ozhzh7q/1tMsPTgY6Ng31ptGuNMr
C/e5h0C/SoaRo8bKa6bI8rtJaUXfXy8ZCPqoX9F9f7ISxzuOlbzH6ja9ZfZ3hiq2IuR6v76RWbCs
/OyKPyJ422s0DOTYWmIMK1yB8gshZH0WQAwWKdLIV2PJk7eCeQW5fC+hxexG6uiLRTkD4TvqGFYV
s8jIdjoebCNx8FWyaP/HzosAiGCbaT74jvfbxLbyrYYRGwpxd19WqfA3NHFeQt3Aad9wmwRDJRBe
hx72qvNMP1tdSKqyX3fbEAe07vzg2IJhjCeTD6RXSf9wSD0xDdpWpVMTdBzrf4RFKKCq8LgIPz10
2Ihkl4iry4YngG+m6flulqPvIyWzxsYKHSQUaYfY4OttJkcBvQlysuRP8trtlOmwhTOazpjreUKt
bzyKVumZEoti5aN5g+SGSU4uUzuFlrPlUZc7ML/IZIqhsBPTJGFQg7mbYt9LQslcpunUY3oDMupQ
ZcPQljR9opSrDBMCqPdyaJ9B+nNGFsdgqaD9f7eGgyifQy3gy+eJzw2mLH6ix5wgaOdq4jovjYvL
sngGrmcd8G0Qnvq1o/efHqEL8ylH74pZHMXtVnrT30zP8VYWQTq38AbX/rJ27cP2hx4uNgv+vQow
rqPdlnBxaAeH8msEJWelMr3rFz0DE9DHfWycLSuh7LAUG2BTjMvagKtYwMjzc0P8xGfKpTFJga8R
jhV8vgPLXpTVIAA8RzkKdaUnBZaLPN6HaTG0XwGxcOkDFvqq0BfJEa+zC/OBtK0J9sH5Htfop0MZ
ySkIqmXPF66vlU5DRDYRaH985TVaPEAzjCx+jWr3ri+pPcXzTBPD2YUL3SZNTn9P+l/ztq5orV+M
eF6MdTenoFtRQwkdGcuwzSho5ox3kRe07waABeyBxbE7ZhqHjrAhJjV/15iSnj2J1Khxpkqn0hJB
cWvHin/bSE2kM5XLgSYbam+qCYfslNja036fE45lORi0VgOxLtdyI3bUad9teM1/Ncfo1MAg3I6G
0W57c8a03nHlV0ItAbbQeCYBQ5oHS323ecRgcyTNkZp30m3sbzjKc1UiMiSrm3tCIH5oc9e+6w0Z
W3bHKL83UVOAZHBFvXP9NUzZjJiWQLlv4I3t2amSPFGXcFNugI0hfd5mB8wBXe2ZnTm4EYdXxUT1
XFaqpgsvISQ28Hk5ajW95cIKDAHJue6fSJ3KOzGEJosAl6KskNswvqjZrCSL3p9peAAm1Q7zDSrm
d+Ew/iGscJO+doglcy1SP/M8/2Ixle5m/jc6tR7Uf3VKY8tVNWIQrxGa90P+SFXxKWdsEjll07UB
sUkC7UAbk2k4rwXZKi0TCr/4Ey1OMGhzEXILsIE9FgAAVCexoNxK3cIwd4+I4hcg0n8IyHxwLrnX
12hLK6t6jDrE+fjsE9eRqmmjSEUTfrnf+zUN8OjE/x/OvCVml6OAbT7KNuZ3nMPxrWZVV/hU9qDw
uR53nf37a0tjQAPAAJADYbmn4+PHaaazfccqTqJtYdZrLC3ZXU7Pa9u98XWH3pDk8EsEvva42c/G
vbCzqkKtIfNE3fE2QFPpq3BZ/Y7+iuhAsdP4nByMKhtFl2AFTJWFELVZDpm+8Jxpjny4rMWuOZIr
WdKlB9amYvSKIH+WZ+qOPWU65uEdMbonySGX8gKGRuf5WZvi2lhbopiydDKqbtBAyLquBhO75u9R
Iu6QLTbPkSgIq+XTu8s3Gplvxp793RdCUYhF0rEK8H/sWZ2z+/w1ODHCLMHl3oVSr0aJy9oOJ8tr
TScvlaYClZPV07risjJYLN4vHVcv9+M6RtLFoliUZlJHiB4RGhdRnkPEEbAMBHrOTlhL7R7Emmha
d6wlp+/2ERtUOAfqs/MfVANCNjw2Vnw4gla1bdzakGrlqSm65r956kVS6tYkt6YXvW70NfZqm/RM
oNzfMoc2Oj+YATBXt+ecv7lww6q9ExUR+7ridP5YGoKL9R3SWIu0BY2ChT8ONOcMwdzgBxJRsvyR
ixVwqJFMcldY3J+7uSYVZQptOuwKwULnw9Okm8Hg+quIpfsMqV6TDEQiFRtpiKk5Vy/mKPsSXFoe
Xj6G6zyG3VIemrNVUC7SpDFyhrShX9/nORzHsqaYqa30KmvD1m1gfUVPfTRtRHgrfVRklwUrRsPX
OgJ+2slEw1DLtArBxlkGHCnHdBMAi7wAjjzRCNPAlcVFbv2OT2bO41bPlfql5/qEZQU6shTkObVn
n1kj6iGj2qgCCvSIoK4Ph8d7wk9N8KnUxERbhtPYLgf6usQeh5Dfkzz9SjdKZxLV5kCdXcKZMtN2
LPac1TqgRPPCs2zCfz04xWkd9eSd6Vg5zOq+PSsazYsg3unxkIkL7OZfSqtY4ODmzYuVIHKbDky2
EqJNX7AMjFmqiqXB0XUznigfDf5aBMRzkHnxf7LdgboT/2F1UHchtNo76weN6ZUCs6f+sTS0isZY
kzA4HGlIEvHGyC0FpCcu363W1MjuFicx3HEuQ+EoqEuEJTwFvqCXxTo6i8ZKo0DGpRMorsJ1vNvB
shCUuNmk/cnIFEOdxNFLwJmekiKoaPyF1OrigKELcATZFflOYYprchWiWFGOxLqooM16LeCfVVam
P+9APQrNYiyO8XO4lRtv3OBCvqHiuITIVvKx3SsEqgT9ZdniPf+rrlNAKN240mpGcbJECUiOT7/F
KaMUjfq6P0UMwdk9TADJPzwgtoiY/udG+MezNZ/wk8glKdV43MgBes7zUIActDeLUvSZDN/Snm2u
AwszwGht6ksLdtCI2Mpayae172PuU5ktoASw1qLnCTVRxEUYSWmBUuYZIIjKs5JDuNN3hC9Aiq20
yBPK+jJDCkJdMsPSnBDaYCyydr/sg8mXPDFseeLAqGRQ0/aSRoJdWurf6o80dCPlICqMZg1Cr+VS
dPi3DeOhRk6HHbRgD1nAmDQ2RU1wxx4GF/AXnNR5c7xUJ2N9jd2EbUoI9zSokfb7MSHcgsdzJ9pN
4ar8SwVfDvMXo+hqk97rbIkImdJb/4UDDG6M/IZwWS4Qo30eJ5JMKvoZISWqnNDFd5DU1TE3KujL
/3JcuTht6PZloI85fFhS3yNd/qSR/F2D5r+xtl4g1Lb/28oplUe0TqURtZ9tk0V8TU0+qbu7LXKq
aL3xDQs/UZVDMmUA5Q1WlNEgsVFJfTvPA5sJxTTLstXWpxJAh8Rg/15GR0Fy0u6NJIvpuiXVedEB
CkF4ndmvk70u/d/x3fvwhDV7RXQpa7cOcqy+uWygSoJN2aqP/gVUwCp3h5zrvapovdcrmPXYM0Ai
UUpYVxs0LPTxZWUSdeyOvK7JEy0GMyN1PoXHGb6xApZNN6TTB3UHrpiynfmOPhh7os5tfuhz8+6k
wNqmF48eY5KWjXTpewszNTHPuMm8UrXGqMg8z1aChd7Wwe5nLhBqMHIMZmJzD/Pthna2YdAGQVRb
dFlPDFwqeA4WteH6nUA87ojZDKKhoG47EtHW1Iq89TJkh4SX9u7mqOTEzLYlUkLUIevj+3VQjz18
ClX6GpbW31lTEItIPu6+UWe1hU6L6zVxe2qxHrKrtbC6oZfPv9dQ6LdKNNe+SDhD5sazkbqe1Be7
WEuP5L6YlrlogicQUIAwWCiiWtQSsMLoaRxGFZ/HGJHMEoBUHk3BUEqBRq8XCXQnpQvo2bFXVr0y
3SjnXYjrAXR50AGq1SaVN/dwomuQ+OzX7Q5pENrb9rnwdJimnueoIUIsGKnxMv7nktZePYhrQb2w
K+Hv5Si9oBGRBh1H/3ZVpbcItAfq3o0Ir4gH+sNoO/zdaOV3Gnert6yFTTY+ei+xLfYlx5dY5y4X
uxyTjmaF5N6S7VlfK3IHIdXpv+HEsL1DVkGQB7ZAyiXZLWhVKYqGcBNoYqG9eWpfrPgMBsNoLyGd
4Jz0Bw4CkC+Q7Ol1Y88lnM4/fBdJRaIXGZ8XsAB1CopJ1GKDBejUSNO0XUkklu+PpgWDY4FLT2RF
4X7z8Z3JfJ5oouSnKRLqsrin7lSVQJbrtyQ4dc/heLD7D2u6c5peOL18n/bw3GxGXywTGcHKqsna
HzzmcqsweTfMGDeFsaEcdN+EB8kl2nBvyFTX7AVc+GxprYYeN5/GId39UqpgBjuXgnj2t0DrugMB
ctTUB+UiqWkEydGx+bi6Pju5hevshpc9u1RtneGCDx60e+KdliCZSE/+QD5v1AYSUmni+k7C6kap
7up4YX3pk81SJU+9LS14W9BKljEYdR9POZ+X5uhcqgSQ4VSeONnpJb3mnZ2geXJ6izPLnwfCEViu
FMD/luUhdZQaHQN2lQssqTq1Wd4F07Y6a9HA5jUYU1MwBmujWsvgrM9FiAzW5bx4sXcl/4X6TB6m
F8kjWXarA+54QXCY7PJNBNqd65qrnXYAB2+djyMjWzw3FkIpCVPQp4QfehDZ1ku+2KgGwMWcAre0
l/ArFH6gC4B2fbhmPgQXiuvABLkwTypqPHidbjQ0U/VcoJM7iWir+1Dt53wBqI1Jf0MZ4imYUnZs
bFBEw0jPD9gIGpjWIB1uTAzWM1LEurQJL2A/ObiYVLpYlzHTsjyBcoyDu77+j9nznEkx9uJ8Ew8M
SFWP16qEea41GwLNI4yramqpdTpfLO4RDgOVEL+ftNEIkz/WcLC6czWcmrfvMHskBK1RAcshsGav
S+9tUwquWNbmJZxCT4OlPqIvDWvDQ0WaXzycq/tsKIig8vqQ6oBLu6+j5QzpsLvrKFZZh4uXpVab
F9ZBv3rwtTzuvvELwqHebtgM9SAnNVyTswb9mj+6/XBTIqNXAmf68SPW6JV+BENuukBtA86bU5YL
v1Up2aP9iBhgwpOBos5rTCqpgIy1h+7vgmmrRr1LGkru9V4TneNSM+iG9PEHpzqRoL9RdoLF01lF
gUaOAypsEFRhKZ9Obx0z4nGrKsXWKt70QewZ5t7TNcwEzt/+g75CbOYYA/x0SuikqPapsr0CQT96
n9fAgPpptcNxwhjU9WrCMC5oDRi7gpFT+PUec6lTE1JaDgdJuJa3YWHt9uGVMV6tDZbRtfl8E09t
dgAJkPUkUX1dksAwPs4bblSAUIjROfYFsxzT/MFV0MTPpq92PVCpCZM7Lj571l4Lo7q7QwSitlv0
aZkgfnmWOtoJirFQpC267y82jTwQkcfjsfl3KZtTj6H0awaaxnXIAqbsmTS7fH93B/baTwlKwU4e
RG1NzOwJT4iD7FNpJ0EiD1Aj2TT0xPNvo2Kifch3iQ1x3LegRXMX8MOAvFL6oVUn9hDX7Veg1FLO
VDpLLQEqpae6qb/S9S7MSbLZIC7WPftviKFv0ldGlsceZGWE6VKzo/5wcZWgXMyyc42ieDd53PSQ
2HOCAdSJhCAN+VOFJezpp3GIbFsz0YWSWeN07Jo5asHMNK3QNcdl0Ssml6nYVI1IGG7Z9Fz7JOo7
j0pcADn3E3w5JfLSZM0MnoavmE4UUFmrMgCqVBMEDTv1NF6jyWFu2fqWKqt9hS0BzAcIieNAhJzr
NhK8iI1r4IFoWVX2c6qKa5iIZ4Ref5hP6Dua/8Dzxg5BZqTAUnZVhXAtaOnTVrYv6lOq/VMqQTtn
IwXqM9MTwntkWoiT7ahOpRz64q8yr6bMwmfuYt+46FdjuX8kp7aysEg7iehNcn9BahlPlWYAXRd9
1hW8pXK2Ha6+HpVRPKTb30yh7SUZxrtgKRnPK9sbt25OA2bF8JHZX0wsdaJkM5RwU3q0EISlDZaV
jBjFsW3t+6gUWat43nDHge61OuYUwzMkm+VR27e2a/EHC7orGSE2ifMO991FYV8bIPuregRAMJre
nzwl2H6e8uXBGQWbEp5Zma9O7oet50kfL9ftS2a2JvhfwV2uAZcF2WLcQSoEygjehVlK8RNSz8Wp
5jM7S8mcONAUgRT688bjBsBBWloLDZg/4RiYE72o9TdKYfYJ9C9VfS22bG55Eobk4secBupYuhOj
rNIS1gjl3S3IPiMBMjgKu70vQ321t2s2X9tLPQO7PEl0miFyrcwn6rrMby3EJfakHyJDzbmKEO0U
mZiMQ9IIHogsAW4OH4fSsCEvOAxTxh2DdYOyh1Wzz+jM/44LgF5dbnxrx1P/MvIyhJthXGSQGdLQ
+RgMN5jCcJs8UtpGKdT0oNtRQIqNQmEdGWVQLmTHnjP/JiErH6xs+1XJpM0lmDU7IYN4bG2Hyu0n
vngFxtmYxDdGKH0afhw1mHwYBiU/hEykmghKLiGRDHE4oXt6vfYNlSlv65Yzci6Vy4RCWrMrXcG4
8uFMt5PGbAptScWhQv2UMo59IjqheCE+eJHqK5sZ+CEIymiU4i6fV55PuqUo30eLme2rcaDTscYT
Mkwwz2NuYU/g7wFYyjOAHEXmxGeJcoHJv8G+qevnn/lalszN/WQm+oaLbiRVdy3z5C/COIBq+hUt
gtXFM2PSKDzFEQfqV6DArCIqVdyd4HCqupe1BVD+3D3wlv1GuUiwVXWwnQI8t1/EtT4L2pfsQmwR
IvyBhK9fnBM4k47JrllAZ9cBmfMJkPOLLKWy2nhBa08PZzhW7g49Bz/GpxoF3GWkyDypkwYHdHq1
4D/qP6pPY/+gB0MgqtbB4PJMpZAjPMLd6PmwcXYl8wyDAdg1/aEISqDW8ftcy0Mf++QKulHDFsAM
Kf1i1Le2Z3VlvFfQLwdhNTMhgZuaUaduW2V9AfWBj1N1rdE5AmDk26py1BW3yBKuDJfjGaWJ1Gv/
MAEk/Qf+RSww9XRFbvaLtPOPGCnhPuhO+OLYLB7jYYyOyGsJhAr9zyTdTMXeVcK70PanrPe5dg7c
242lHsU/cqQSyBy8j4NCQ+N5/0GaiHbigvmhHX4LaPLYgFZbcXtltza/tUEuM7t/psYoslobsy3i
IT9uzUMLB9sV4v/k3J/Kka0mxR/fAFwu1ohVuhsDVkTq641c0j+HOa5xy3RJROjhkITpt6UMZAEO
rBrADepbz6lzNoVjpnMsBufHddzPBKk45YA+FLZUSDijro/09UjQeN3VBq/OJ8/A8+OQbn2UY07Y
3NlMGxBu01y8Ek21IB2pxXcYuC78gFkRQsciUVzyH3NSpwV4wU+VzHHLFaMdl3gTrVS2fw68ZUX8
M41JGteia+sJNBjbdq2N85QwABBz4Vw0jiBwlpEBr5DyNNGWR208lFmjzigw2OGgVlobO3hN0mzX
d5cdVZ+nvUskehPWnLF17IdgJZaK7Y9eyAkUGCp+R0SfzgnZ6jzQB/8U6Xq598CxoLKk/61YNKSi
c73f6TYVCalwqb/j3yEkBxPITtV3nJL+6HRU47ma1reVTw6xvURoDHSCurtbtiuNKijIwtf8YdaC
i4sj65NjG6YHkCzjk3fe8jY+w+A9oGnJBFkPgQ10s67csiSVRCQ5SsS+4iheHcoQ78WBcMaj57/9
lRAy3utilOwlYZv8A1mFtZicpZkhQLRAFlmWq4Z+BQCRWBu+D5iH6J75QDR9HqHwhlrou3WUxsQG
k8ktVy5b0XCbycqeo/y4GOjQ9ElPf+L25WjNWrs660LFWpfYszZMF8R4Me9ORVOje5j0w34Z4tEY
Ga1uCsgOs7v6OG8kLARB/J7XhW/dTWsF8rOzn+EYtQL2Q5zLEoEQfPkNhSu2aJcLDCsFoMunkcdK
nZAXCNGIpr6lVqDGHD1dGyi83o+tKDxsvDs1utg65w/MtU25ZS1kzKUUpHxxTUhFS3P9yY3w/O/R
OaVmFlB9fYcf0pqBmmsNazufjSwumcRwQBlOMZFCretNH0mg3zMLV0P1/T4sPyyXqGNVw5E3Sa1H
WnmM4UpNjIBT+k/5pQhJj2pXKov693nn3N7g9Zv/zVJFLqPLjFoFyve31uj+a4gjazEiGbqfe606
KNIRvvoOz3wobDBaKbDkzleEzz6nUqWFbSSqrYhbgcu/19eIDN+jiiwmZxlpKUTzLrdsGXwVWgse
5yju3I6d378lK972UPLjQGeMPfxSOk9zOChvKn2Y6/Bt0aJ/94ZUMBwrZf/LjYAIDoTjCjyslE/l
39xas0X7mtrTVUOPddWgGpBwWwavNng2GCEAGIdFNH2mC3/inUzQchXXSHo2kGdx3a9Q2ZhR4BtH
oAwrjNXfdE/mrkjIp9nEdtrVbQfFO0PQ/Yv4B7MOPjwSna2ottOJH8hKN0UhYEhlQjy7Ot4vmn87
ofcVdxPhy5OoBdI8LKMYdz2HpXjvSGvyOFHuaNxhfY5HttmWim1woH9PlqkjvKvkXpO2DSTTES9+
gzPKDiS5bFo2Sow5VqYeu/mvIPJyCrXb5u+D4GFYwU/qo/y/CE5tAN12Z0dqN8dHVGxwmWO7XgXO
8ufd6RsurBPigBXo536fHn35bIZ4oE8qitKDtEhcyoK2Fz1g444DsDW8zxWa+jGElz27GkEQF6Xa
5DFdhhMpG8tYBpfPNDgQBHWCw7LS46vtfzl7X/mjEpOI8JCdAeWPWqgZ3/3p/F6FzCC2k45ybwku
6Ypvum15sIELPBxZzWjd3m1bl0U0D6aiCuquAzPhOg8Hir7CMudkjfiLFWogxGyHsRcrIWiBlDVS
jndOJmI+XYIx41omVFUIYeaNGIqQydLgOxzz6M1l+rwS0ISTg01o03/etMoPphmmddA1g/gIBqRi
cvHCJoH98bPf3PCB8ukN54LiveP3ZVRNhqwifg9vD+Lrb0mFKGL2tuTHigEoYJBmbNfDtIJYb53c
1eRaa5MhaHWYzY2FI7dn85AtdbumAPqL6SB64DoerSnkzoEuRRPKnmTHuyhXOr6/w0B7CH6E5K6h
CvHMX9/vjuGk+vqcvJVoAIJusAtv3BkdBKvwwVX2iBGqHB2yCDhC8+PSu2P31EioNE3TbzvaO91f
RP6GWVHoDHdh3EIScpg77lxrEQnnsC+/wwvbE78mUmEL/Qu7QsHWrLCKLnyOv73H7PIEeuC40J1F
jap9ySsB8qU5rhW/z8ow1NTmpvmKwycSlgzijzBkWVhU0/FNk2cqjvP+JnR2PXj+4U09IaUaoEMA
T5c87ZwBMtmNdAfMCZqc6yjZM4GHP3V64e9XZLpbixLo60nDtDCjNOtQxrF0n9GcyjY5Ojua2DsM
5gkeUogzHT3+Csloc+EN8iLVKqduHTPYY+6XZ2xo7I2Q0+xm20pcXjKy9McbYlNuIQdde9YrSRYa
S4cfErkm7j83sZFCGGhwUaf0MXFprEXwRoXuARx/MyTxi2LgS/1U1vlirt/WxtC0k1LRN09ut5vQ
PIrO0dsTv0jrLlLZCNc/MaLBG+VoJyB09JIo13vgtigey6EoH/sxvE3dCs8Z4ZrJMCn4pFr40aa3
FSMgEaDjihr7ZH3Ch9tHpnEA4jdeVsoFW1iCzL0pTMZpgZpWzAqMpJH9QC94cV0TtjiYP0LnpPEf
OvX2srR9lZpmWJJ5wFJwn/BKsGv4JvMpT+Q9HUmsxkt2KwJRExoStCi8Vltdp3+58HIQOaA5zYfL
1R6OpOfzFs+aa/F8LxaaS35w8pYOgLh+B3GJfdPaEdeydebaC/THo1XVgjR4SDF8/Sh/OUrZXyR3
CP3skYTlxgv/zKUh/rth6gUCJXdWwj9XWTEAuXsBsveoEmqdC9PRXtIL/xQhAan5+nRw0TFjyUX+
FuCNBwijdXg41+j2iRWGfOIlumyjM+m23uZSmWpXYrxqtP+SeyTTjKqe9tsb/+2903l/zjwCOqF8
1zzk6kwXsD/7vPavT6cZe/Amhj6LB3nBZ0x9rFvVUtiUc/oavhuCuBlMcEte8ODCjYX3nBB2eLX4
HcjElSqcvzA3Dhmd/f7HYFWCQKqKun3pbm8JjLJZmB4f+j6XN4irUUC1kDXGGTMIodtpZYx1ngRZ
kHw8C4zc4bvKZFEZh6JZ5AMvYJHRbVKn67KGk1uqpTjVkrKYPQvag/tVWE5NcLzA29fubdGlP+/o
qCrsIHWKpt+LKPgcrLfB8Cr14uEcJ7Yz1txABN3j+nSjywW3/zdJ2evy8JlFX/fHF8FMc0h6OpxV
n7/3nMorSVHgaIwOOZ9mcyvYUxqAZbSc1SO9kysN0L86qDcBtDMIeDy56vUS1HYiM2ftZ6FzcDTa
deDuHIU7fzlAFhun/MPgXY8MZGQ0/5LiZy2Nfqcxw6HTC/78qgklAac5fCys6KOz9CgP8yxH9SEt
QyxbXSrXZ+Fy8Ew3VuRZPDlGbYaahF+gm3Wjnw/qlxvJLGNE/5VunfFNR1l2fwG+/6qAArOfTS2Q
SwjDnsq0oDN8gPQXKzaXRaVTUs7GHYRCtfkpVJvK8+ZqFWjconBC0SRHWyYG/hT8HNSg1tt8KEvK
l3RAFt3oylJzARAZBALIiCbfPN543arvLE523fJuRXc2lYkOez/iWOQjaEFbZCIQNx7vSSPKoSmu
JCeO9Kx51xFuBZtssTilQl94HAto5Y+Io096XYeisAG29A9TX3AKbU2rbhSqLoFvT3uDsWPN+8vn
sr7nsUkPsBtRDV2sfoSr3+Bk5So54gwa9uHeRzzjg6lCSncHzvXX75rzHMN+e2f3n3tU+f93B5i6
GKGviDvcjlyKyMWgc61PfRvsZaMVVJgNj2hwz9QecjhF4o97l9z1SEa29HYnjbUiQ1otGQdKM8bU
K5GbNRuKntUOwNRTAz94ADO+Z15a67RHrUiQddCe8ry7b1gQ1umaq7+RgWo/t9ZSE96C7zi8Vm/j
IsA4ol1s9KWQ1FWJTtV0yv3cj/gzJ5rySjACytTAuy8FyiBfdAtBmLA7Fab8IoDp/fqwu9uubpEg
sCSlmtS3lUbV3WbgZ2dwxMNLTxIoHjFiO5rqPegm/TeTuqs6OGu+ZOQrXFwtCMhhaS/vbUWnQga+
Gc8TEIPLpWi8W0duVa+30sRO4f7PuASW27Bkou4u1W34RqktDjuULX78doZPCtqwgkZyHdmWMqSr
W1RBbLrYZc2axPIyE03cYEEDEkenq7ad9sOjKq3H3SOEQ78KVzvbIzTZ02a7sFKm1qj0Mqymh+Nb
8soAJsKAra3GEdUum5AMxjFLAKG2J3EBAwXbQg3/t9KY2x5mWo/mKJglAH+0J9ekqz+6/mNXj06z
dQ58V6coW6Jd8aldT8bbWTcftNBqB8IXaAl83XvPWF1ZbkJeE9dr39xzIzGGHhjSJfPKUdwboz6e
W+yDlbdUcmHpsuXCz2LGrvnzx0YSZmutvC66e5zLSVrTvXAGVfsEbNEY1oOYGUHP1bLYGJc3GtDO
XF6PFfABHnC0VqrgrBzIydSg0+VojEZqB3nTu8QUNvHELm+51pyEDRhle2HJpL5TiadtB1uJgoFP
u1N2uaERZxI2cHFF/LrdKOvJQhThA9BuAAcIU+uurtyKWht4z8aCSweSot13yHm3fUDiDFJcm7KJ
2G2ggRLjZ/eAqpz9i8GnsnsuDovBB0Ohp9C6hpvvnMdLc/6TIiCVMCkqyRpSNVmA/uXcDcUmP1p1
OHsMZr5a4vcrtUu2jcPXeD1mmBlPICErj8oQXZiMQFIDVwFgnnH6+Ap+/x+wocTF6b9MUVeduB1L
98x5ERFJAs2BXtBnd0x++jq2AVM7L9t602il0qifc3HB/qafvc3dKPtm940hYzT13RuF5pabrXYm
JmfrSj3fhl4kYy3tqeWkz53yX73KccbyfuHJNcRCFCMwBE+sOK6F8Y4TQErLGFn1hFIE7lyfGsE8
Fr8EQb5QhNSJ63Wj5HbJzZ+YPd6T+BgXxOd5P0cYJ3xivwnhzjCR1LmqnaFr8wNn2VXjhGXTqwO7
sdtk9lCRv5avIbgj94hloCBPTzUOqOCv
`protect end_protected
