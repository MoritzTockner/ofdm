P42407@HAGNB260.3976:1639982020