-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fn0Yl3Po+5kVrT0hFbE78DTKcmOEaSl+Mu+rUQqYnufHFSbDPkuSVzll64nMidXtM0k/wd6B1oGq
0cIe2n0aPXhS7OvYjwY1fRcngn7nJcnlQ/Jxv0q8LwCde4L2WyHuAMoFwVxJFW/QQ2W/pj44fOYw
NPgJbekW31hqV+gAk2EfMXEveiSiFG2D5jxJmD2l5QYhM8i7NOtgLeUlmgou26ucY0sXcbNtpXMH
ixwoTOXnB36jmwChN7XB5nJG6nsDhxoJhtYjPgSqf99TIMF1dcbJDcNOMzyfgu6m5X9FBeDTrKVf
i9kSjwmO3+mQhNuYFCMG4acGnvICfnFQV5ussw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
YG9/ob/e+QJutWaloO6QmYjlkzRGZglElAYOZ8B32XPkV5/o5RU6MjG7mTAsC01fhp7df/Xq3R/w
gr4J3QyhytD+MJzTDwzi+FnT8/v0dsT7/7OTzX5OEoOyFjs5Ox7WIKLNM9f7NWPrAI/6qOVVXThN
fyjMlp0gmznnAzgZyyQHC1vXQr61W1k/QURbyADmbjruHORl65q7sRAua93mBnqUqtcf0AAlVGnc
HbEwbT4BhrmpcsbW3IVOvqjNos07cIq6JkntiSQqi7Pb8HXTnQMCnc0ZVyx5O/UuIJ3piXnkvfqU
5KEqVw3A8b14q4CcsnQheAL1k1ShbpbOzDeicIb1XF/PgleVQuPGH87bXopQXZcGBsrIfwbaVnzH
p0sS1yO91Tct6boJAdVmRF8ptAtqzwH2judGSPyNuK8FPqf7nlGQihy2T8cLXLRZ80hn3L4G1Zol
T7SeziQFHSqiR0Q/i2mNhD8t2sKQfHca1fcB8G7tOyzGskObL0x4t3QIK4gHDEYisKKlW0X7wr1m
t3fSHN5zr1NB+I2anYFzEL5zhhJ2qqLoyIHMeqXwpNyRaE5X5JGjIgq8en/Isa0gFjFTJJkxBMEf
ZmkQfCINUSZboTp+aB3jWMfmsn5YGcLm4HMOHFrjjbrA5EBgyZgtbg4G/KlaoyQcVugL+NBHFHFu
5DAdteqGTghzSOKPMoPAJqj2FWNm4/0NbFDpdLjAYol5MpUtYjAVhB4y4hLnKH9O1E5vwPDS/NUc
sWSphIPb5MjzjGcUjt/H/IvD2TSLWDiYdffZnNS8df9IhR/37glP5YBB5x79islmhOIkYolcCuMb
Rc7NTgg2uLqX3Ie+zPLfiG5EpiCfKK5skwkm8os1X8kpo5T/CtS5iNR/5ArPrK7n5yNBocDshX5k
AUh2xJH7/uYQS1/t/t/afNa7famRueNVhg3E9dwyLBGBVMGqnrsSlczz0BBuNBIa9I8nmISDfWTX
Oza9MAQ78HtyF87RECgJJrtk/pS00WAXhvuoYrwXxBih6x7pSDMj5wpboPcjFBIY8O2uLKu5ZVT6
+6wBxLpEbB4RK6T5mTB7VZRsx85+ncoptcJG/IeZNa5YeXY8Tq8Dz/HgrfKLS/F0j/28VU3whNwC
OM/LSF6zWHV0fWrKfraE8RcTJlZCkxgG/bJSpZluHhG65XElBhhYpmoHS/J7HbW1vCIKlg8Wzzr4
Z9pT6hQjMn8Ee4dEVXmgDbgoMdKuXliJWxja2nXTh05R22yg5kFqE/rEh4YiN7P54H7RoGLWU6KI
JwQv5n0aMb1DJxSb6b6n/38FnM3BG332P3bbhmLyyNCh/rGSKxy/GUR0unT2mER46g0MlIpmU1gH
i0RGy4vEdKIa2q958+Qy1leO7+wEhI/SGx79onEV283iCJivgh10j6B9ZW2H1vlJDDiQxOCHdQkR
zXsiJmrKdOFNixzpf5g4tBE1moqRefG3Q103Be334eEoFdJ27AYfCP/D21nFWzxgUYw3YNaLdLAF
0YT1BeBOo7xaSmsJmfGggYNzHU5QmsZGXQ7BYMfxWaENTf2sfYAypUbENZBtdHBYCPYTlbW2Wb6p
nfzklEtR9iDnkfcwuPUblsGUxToTq40IkR64RlTHmGGbunlCIAJILVSerZT/h44DGbyRMdRYCNs9
CGVWNQU5OJwcwCxWZHJBNqBJDQd7gKhGOWfB9Ia1vAoFa9SWRqSTuBrtB7GSqcEp2TmGeyanuVdb
TA5TGmzzZclYY+Q641xfvK0Qa16mSaLEsRZlZfS0bcYf74tHWNzhfORCs8ihxgrm7/jC7ZHT6p7c
M2btvx+yMUfviey9HBIj/vwsLCXGBFhVvcjzoS0wm+ZupnInqIUC47WjdKm3uUSGgPlJLv5S8jkZ
ef1W4itsw1hNTwPa4VAYkqan80w2w/vlTMOBAMxNFyrLQEfansseQ+3eYcDaVEb33iHLELccoT3w
4LwoAufFufKo16uJaTs/7TPVvXwdQYa0ShHP9PBt+4X/ENXTKJlx+8NyMAWBPs1czzG3Bm4TzHe9
u1A2SQiYopqX1InL8IzsLKObpyJOjzEfew0RPaDwZAfhgJvcIasHeCHa9VnlG0fG3OplDJY5si39
5PMnNBhAOytDMgQn3/Afc0O0bc3iBru+/V5QCY3vxSb/yNmyelOiCpLrBY4QirouGLgMYLNy9CFW
3gkkaRIUeYyd8bPXXoD5MUBsgGxQek4C7oiUrYk93CJVa8L0R4+Mn5LjqvMvKfWTLnX9n4y8X3kW
DhYhmW+4D+hGq6HRD0NfOTD693p9oWF5x+Po+z/XeHyZjdcyq9pv7NLRrw3bujbyAhwc2sTEgsST
8sPsw9bI6jDcLoUtuSc80+96aqpiOiGBugrjIWGO72pMSjm1A+oYoDbaQFYalhjffBeLtVHdT/+G
+hWDB+yQpnM9cyeQi9eX+UyO7XFo5tsB/yp+CUnAtXHD+JTisdy9Y2ZJ8NHLdm8f67i0IpFGd+d9
3wli/Vy0OfAivDW6RH1JdAaUIvEoMwZIjHh3OZW6VL3JASxKtiruXX6wXALumnifY8e//tVT34u0
uz1Xj8EB+u3AqfICena6SWrH03306WQVHHODEXsxAFZjuT+aCV2fvWSh87UByPonMHE/M0zOweU1
f7pmwG+mfxDxQ6FA+OnbBW4yu7SJoYUVk09kupFZYmgqUJnZVPxPkgPr4cSWVLoYyh8I692EHbcy
5zCHbjnRmes7BEYgCOLRLlwPHRoHgnzE4Gib3nwFagIArgW+iqH3HmiX+g1gcdiBDE4w3CrvEFnj
mjHSMRlzfGM3p/Rz1L7YhPMBa2MVL9hsWYmkEHbNjKm/WFDon3Y4mFtCbfY9xoOMJ2SasvgeSomj
mhcDt78oefjNOclclSH3keeDa/kI1ru+6K1OJsywZ7yxvLPsOJxLJPxK+7XoTAN/6s0uWLmkbpuN
Nl9J1e1iSlNfWcByXWfxeUdZB3UPvI/y21v/FyrVqH0VLD38/PCWXmDrZWu7TvTJV8eed7w4kFq/
k/ubmUSYnRv054kUb7A7aWLv3xtXEZfU/LyY0KuJSSpmZSfnc9PNVVPU6wl53gfDKjzN7J8MpEZ5
gdE/hQFW9XZUKIX47ddsvkWoW/0gYs0WWWs9WMvA0A7eI/H1pRlgfxpkGyZOoA61HM+SmKILyJjZ
7EGrFx5t8f911oT/9qHYYPhNROvBOvy7jAtZ2DowoQkkRkJ+oR4UVCIhfy7Nu2BjdGMIgGfY1Fzt
E9EQ7leabaA+iPI4owx19472Yj7RZU2CDRnWsXNKfQeYyHdJbAx+AkCDi/SlC/UaOYU15u4DNGOG
w/nByUQ6ClY+XifUHM6zzbj3Xev6eqKkwP1gNu0sBnDTkd2O/XcPSSVDdwBqbXM2ttoYkZ53zow+
PzKN2CEOJUfeX2EyDMg20BbVYyWPchw7QJmUPxZWNf0G5+jsN0iW6TRCCqCDG8F0cMFGGsP74/1o
k0eUlNmaRHPcNKs5r1TffUfEB2dthJj8YnOFGha98ABpgtVhT3UDoA0vFeqr6ZtVPuhFGfKxM0lB
m5oA0ffKznM/iyjzJsO2ALunXLt8NX6MBnyzTR5/PcsfpKiGde4JjTtmTwpegcToIVf24Rdsmmqw
4WSIXfW6lsNRUc+2REHDqU57KD+OvYGJ9MGX590YRp8+4rlthQ5zcXNYBIMbqtL2XIliY2d6oAmX
NaT5dilV7iVqJBqjleBBH3AaJyecOCD4eVQ5smXntBdzcsPIMAYQpNOP+TtzisjY69BPYSev76R3
GhNqkXMtO1EkE7oeJG7OKaa+hwGgaXaqnkTIvD3g7EJZPbO0pbISTNcMe1WUXmpT/MErzst71++o
6vQ1Tfpl4fVokC0q7lSb233UPqO4I6/yNzWcy/1YnZtQiEM+v15CKIzQzx5FHnYR4OFTcl5CDHgj
7oo2FglQInWYBeY8pQ2owzg/URrcnsJMevXvsyg/7kr/bd5L8qjfaG/C518ibdxQ0dQaewJUtS6Y
rY0JDff3uISyaU7h6SEtK4P3iJp+9Sg01b7CPDbajQCqAAGosBr2C+/XGahaVGD4vg+dnE7eXZkT
PjF404B5Za1eawuaD3bphahVUDEQUwYjO1qC7xhtgXm93xT/oCQUkG0qb3JuNwIO7ikp1AdD4xov
ZzugUWhvDmdLtGtMUHATW8CJ7oWnNel/yu/Fk50XyfL5rkakntPzUU9P51+GJ1j7fYQ34b+MjWIF
0zJD/wt6M19qVau3QBiCXNoxTEEbwyjWIPT+aiTyakKMFSrhVt234rymBQiQ652C3U/rC0AehBWn
KCOvrXgriu4/8wEzt2cZfptTxiS40h9mbUA9X4MdHUDWRsjBeoekq/hYuP8r+KjME/5DUKcD5IWt
FhDDBuFETiYBX6pjy69ljBDuRprcKdIuc7oON5oMSX9DPMyDUCLhSwYVxKs0RxQcave8LAb77tDD
MRM06YZcdveYEk2hjBPiMCqufVpJUE6FU+TSy9q3IDet0OxfCpRckVCuKQsAUn343mR/4HuEqxRD
CflpdPtAeG5Klf+bqNpvDv0Yfhgk6kb7H5WTazbg9otk7OcrPNHT2QdTDcPigEDhgpkyO+4YXV/c
vGPFtprcTYqukfHsYF2t2v3jrCZIoNxVsEYLjK9mCFAq3xlaLH3UlbZn6Txt//6K2qMEI0i2w9aO
bK647ZrCXPx2R3AAsd2MJF/TywfIbCcuMbjTs1XKoX7eReMTKI2tw4fZb0scEk34ODQxDCeEh8eB
AXkOQI/qNM0l+FP2fp1T5L/q9o9n+bpQGZh+izxJ6yCk91gqgkxqA/m0/6AIFEmGmD4gfcIA8xM8
637FI6R/CjZyTp7+IFiTmBvzKpyO6E81Vi6xcD2t7ZI+wDBYU6amUkv+WGrCJxjOxNkzPi8UMB5K
f3XCvqAEv0vUhtOMHKhvFW4tue/2l/Xci4Y/WnD1Me3TnqodvC0yG4LGMcB3KHu56KXDgFFZRlBD
C1yINw5Nd9yaFyavOgdo8maZabvZOCajb/ZncvrjjwAwgjd7QpiUpqGzIloi7dlpxKf1XAOnRm/O
MmqV03+scKrchQ+kM4i8m71liWQ1V1tiuk5prp2AUig4YOjIjlcqIrGHg6hHYCpBqPFn6E4myssG
hNmHCjnC7fBmf7EhSqTIIQf9Cb+2aOuvtzP0B3qMEN36/+mHXgFMNt7sUMpb12vRwW4zjy8ZfGs3
wdUGnNHjS0Pwb24lB30L8t6PK8I5QpvMyWyNASi4tCIQgUOjQdVU4ISABLwmngn0Uz7oHTU9pcrH
YaTEw7FukvkXCpSZRxqy1bXTXJ/LPX79w7Oy9ZLZHBegPY8a3xnSs6OfkhgxZul4haTJURwabvmI
zjHdQBoFQ9wVopyre9+2sVIWX+VtXLT+YjI/sPxr7ayO00U6aZEAuv6SeQdRMg+15qaIscRGX/0R
VqckQqnArsg+prefCUQWYg2PZ3z51qrvWE/MqZnlk0ifQuzguTw1hyJdtojuwwec/jL3Z/52qblB
Yp+dT7xU3OQNHVeNnTD4GVDRn2HN3CTH3aQRB0PU2zUX4sah4ybehM3j8TkkC2eMsKulrUnirkLU
pxMtC573hokq/grOfVFwWu7SYB6M93/kSBGIA2adLhya47zf51U/FnIGKMAApe039BM3grjNFsXM
mULaNk5YsKOoCIDdvXeqSEfyISCBST6AAHQLzFCiHNJsuZ+gBgTNkWWIwRv18ip4lHguDzwnsFfP
Wg3+n/kEgSp/7ScuP5NO2mKUF4Wc+1DPafj9O1CN7Z7e/55kgj551RWvDgktidcqfmmFMR8zYzIQ
+5S682xg349l48bFazTaf7yQJQr1thtifn4enlsfef7dobBZfvmhuaSwZ0n+ahUV0HSJ67UK/7Ym
s6fniaBwgp8M01/szcNiIpv6aRDqRacduLEAeTZs7DZuk3wtLeSAmJ7egrWLe7uSpFYaPZEAajYj
BMnL1hPVKyselq+ulRjtzuU13hOmEPVGWhkRYo9lQ3IOIObwdJAK6ZwZVA3blPt1I/8r246BxJrM
uGS6/puSThWSIxKU4NXg7KzlFdSs3q+I/FaKkUIuGu3g0/17VzYssGTlIO2+D0daMObmAhyUCTth
+J4GF720lYndZTmvEwpXOUoaM/stslSWPyVik57HM1SA6L80gyDLL5Q6ItKyK8dxvfrRfQK5efgV
KPbPyHVCd/A9ggwHo/XWhaTy7nmMsDD4kIpVdDTwLqSAjlhnEbWjxNFmcjXGyPT22MG59gbL72p6
oGXIe51qfFPrCvOW6z13wwYbEvFRJ30tci6voyEz6WQVKYdLx44a6yE8+2FU1Lkx3zRo8/cCkzZS
T7Qr3xioiW3ieBoWVqjUK0khedqxGYD34MxKMpuR7glsWoyKUBA34v1hUWgOa/1Pxhs+dg1YgXEP
kkRRUS98XhHN9phwXz3XH3SQC00knVzEiAP0xhUoH7OSN4yslv8E4iaCkIem0WdWgxDlxw4xnx5Q
XIvjFtqJPzThBNeSn5vyervgZ1bfLkgJSfC4RxEYcTQ6zSARQkQgN7LXDamcDivusCNc5LrZ++qr
3LrhffFiUz3OuhW/2qAbBqhAKS4ToW7GsQL3XxB17eGzKMvo048MjchdVQsoTQNqLY/g3DSu4t9+
sN89w171LTe6HHBWgZR5TQWDxL6Qpy/0S2tfIc9AH8zElPXhDfmNRE4f5WdlDBdS2nCl0uNj7vqR
49lWVfS9EKYxLSaPT/HTeFXj83aJ1F5EJrzVhjBKQ/Vh/8zlUuxb4rUV2VzaHAEwdDovnD/H/Aob
Ql71gvbKDs/dYHg+N7Go4UP3Qjp2ppIlbFhiByo6ZcRQR37AYOv+Q2AENHao2i/Wt6QojrFhRP1n
65SEZXJN1/X16GNJ3NAbWvqFwss1YaQbyCwnvipa81Jj/PcRel1dKOGY/3UcY1Q+RI/NZ80gpXnn
+lUiyStV+VvdcJPbXxGNg+PGlilfIWwqU/7yeG+POnqZgiAywE8eHdlCeBuU67ELHmKx8njTj71d
IOA/LCokARRjhT9esZABiD+koRROjY3kMvP1hnoRmxucKbdJoqT/GI9x9y8WryZu97dPCvdRdVHP
ngDaQXPQYqeoRJ7fLf7r0eaRdpW/P81SLaM3KyCwdvkGHzoUPWkREMAYWlgbpYMRAJ3gJzmdUCbs
wPygtvw4tXu0+4yxm/Uv8ad+LZuqhbz/K4AQQZJkguI7XdNMpJxNMFwmZ67liiTNYWVQKyHDWMX7
r/SjeY9KD+MKhUH2BKmXeozFnlzCyO5bgez/XNxJ4C94ed0so+DcnOAglFZqMj2hrSfRnZQDMfUA
cRGOcSyHaiujusevLRzQjX+mdwMCdlX+6JPfXlLBYsuF3CgEaBtmqMSiYkxgx6MmkSVoPOYOv7KJ
73atxwvK5loS6z83MAN6mS5WXnk3xNPlyddjCYNUqpfNZVYUrRgZ7QNNypc6tbjiplevE5yTRs6Y
MImxEWcu6AN8a63JKqBESOIO84wttgTafP+qHCoiDsEAePzk65fk+KcObBRgjgnKGrPhA16uje1H
3CZ7BRxP1ZNqPh9u67i4DgpF7ExneC3pw54qBTbacQf/Fs60konuX1wsPUlvUvQMdWB/QCX7cIs1
LZwvl2A2j/AAPLBW3Zr+ten4FBhk4XKCKlNjIJmvn9Xw9rPF1Tb6ia2t/obUMzkw2wj98O8t4S5+
ytV30VglZFh1uX+7J+ziI5mOKlCvUziKs+K4pkzs8eZurRC+MJyJ5Yra8a94yEWpQyERgVTTl16Q
TTKLEZe2R0h8rT3LiSQMite9Y4gecSU6l7krCXNvqv2I16lDAxERcsLr6YdklJO3hVccYhiY1utt
ROsMDXdNyDc1iLVBSd1h+EcTgo93/656vU1qovZIhAJlMwxvQ/yzS1ecaU5daLK3sir77X6CmXgd
Oosvdthx3oxr2E5eFDDZgj9JHRBk3YLzZTVdvXU6Sj/PpALGFbdhz2vBqecBklYYmbq8NZJxb8/o
JudyWH3ZyLnx+xXV7fpSJjFWMFzE8YNAAt+Stkm9HG9MHJ3b8rmGwNidruBSK+WB77frptjVTLPt
eDA9e10TnVk1AayVI0j8MtZZNjBGWhpECByiFiKnCo9is2PhM0hfWYI1AdQPz32lpfUGVbHeiWdx
+xxkQyErffbwGN+0wVzlkYeVcaMqDKgPdvZnYnViFEdhrIuhG5Xe3a8uSxrHzqP644G43jvH2hC9
OmQ44UgCDWb5Tvf+1uWuMVH2MzbXEUfPT4jS2oyyhg19LDx2f3DYnBVrqxnkIGhtZTCuTqM/8QYG
+U4pNPpZRLWlaopiIf4MCxl6khTCeZRqAm+z8w2hfmFCftQEDhWi/bmVFhQ5UN5hxKkpIU6sDOdm
W5Q8pjXkbq/FOd+rjZjf7h6yO6LLTzo0bqJcaAImM48g7wa28c83hsBMbcAR9IrJt5N9r5sCOR3R
scz+XBwah2YHejq62AeK2HH9Tj0wZfz9+DFD8IsWE0fWL5BGqy4T+XXYAI9S9NK4rj7GjxpbUqn6
6soI1StEQcfuVGfwtwvLZEokLodC+M/oTYR+qx8+fgZGNtm1RNjSgrp7dLtyh8frO6Pv2cQXkrk7
cTFhj2c1buQsAEQhoHM=
`protect end_protected
