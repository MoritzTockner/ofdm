-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xr7IL3YPNBpavxB+/U3plgeI8yYAVdAcwM86y25gvDjSuTvrp/ufTK5r9WoOc8FzTwTKZMOCqiQd
BuJmiZdOA3PoCSOYBJ7BVuoRbW2WkXNeYZ0k7yLjQaEbH1iS17CCvvAeAKkNWswmMo25npZsv6dh
kYel/XxkMjsu0Ol1ja1yddCgOw61ljGfVeqi5AmKLbzjf+3X1peRT5nKhTLrZam61a79upExwWl/
LMOM7nli4hIET1swYNdYAZxmcqLOeOf8P3Em/acoQSFiwdcO/2bDqRDhXj/uy0+JaTSXdWVfqZ8W
IMYkjJFSz3UkwVaIiK2QO53R36SWu8v9NaGPlg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
+ek0M/2JB4Zi+bLQV4Dp5jTquFGExc8Qd8SnhPw6qpVmhef9hFev1kat/szCN9P+eiiMDv/znukl
oLmYDKP4w1Ti2uvhYHhKbg1HkwZPrKGSoX0i0Y+zjAWJMOBNEjzfidXjVangKlMCFPvN8I17RVda
3ZmXqIpnda8CXukIHLIzlevFrb8aa/Ziy/s8uV+0aryvlGBS/GRE6j6p6547L8DSyt4WXjiLyrsy
N8O5VDP70px4dLcTwktgPJ2EtLve6btiMD1xWgsUocY6O35fJftkzFkDNtYHlG7T/g3d3R/yjBzZ
I+ym+AyIdSr1pUubXAZ84NHs/I2fva3Nh6GiXQZBfy8UGi2rPWvyFqHepUNla9qbxm9fXBzmcid6
3ixL/+JhlKi5XyrucmfGKLZulu2dwbia3Ukqe/MOmdixcLfpZUoAqRBUWiE7e5IcJB+l7U5UrLxa
i5ZfHc3EWv7+DbQoOj3UXgzLNvg5QRwJrfSe/DywX2+nTaMT7oAEoKHYV3VzOCG38FfWbpAiPyNx
+deQdNmMs6+dSgq4+Pm20Aw2myOZp/Yc24ksLbuz9RINcL32LyRnzCwXf3+m/z3sG/0nwu5wd/t3
YPYCVvmE+Gv8aQDXT+kh8ETKfgv1jpNW+auFTV81WjCHYcIKFeQXHZwWi19FbqJAvze3PUWZ1pfR
46M7IitAuwjMSroHlkvc3ITf4Cyy/8ETQHh6+B6vYrUcgIlmuAKWx1T3XE4jsBi3AOtnSkmN1Hv3
mcF/1wBm6ru0b97UHhk89oKYGX7F9vdgdLW6k19ChD5957KjdYrwSmnqnwfmDLu3hgmmZFV87p1D
MwAvzIoX4BFY6gtMb/tXt/d3nvAcGL64HUlpM9ztB+4IamUlAsFYdhEawt9xYrgdMFVEBUYqb+pd
+8YSBP4he6vmu5L/xzLrREPzXowczQE1HFWAJDWKqg42cd9AwRuS5/P1odrdOhaKkrtbJZiXJBMR
nnMysHqRzDzV5ojb4sWpbrmmkMKqPbjfLbAWXxmym4GJBP0M4YMBeG4KMn9i3fhdr9n4F8aO0sq8
isIpKxVk6EYutV1Qg4VWzdJjTeL1kelMLM1mWCm5Yfi0DMMz4chQjqLKm1fRbtKrtawsbuO1gAU3
NTOF1Mjt2rmJ1qBtaFlMxI82CaSlquY6NxlczPL9EMrlcBMvuIP1s/R++6KpFtuIT3nF5hVTnDeo
iqx2OAbPLOcjU6hW2MhQC3yDyJceK7Oc82HMZ46qXSsOR9Jr51/7mTiH892mZ1cT9y70qEPLv00P
z5NQ/4R/HMFD+p3mo5TYg1slUFlcwQ0KYyPQSr+xy1sFnI3fv6832ft5CkMgJwkHlSxDxtu5CfYN
UHOf8+a5Pq6o7eIBNINFGLU2vR7rWlqISM4Szfn75SKKnr0LXbx1Yn5qyrrYjQvkbjv0jA5tVHMY
s41zPaxp2SeMIwj0a0nZFh/M1RCRmYiw6pc5y4JDbfgrfBaxcIsIya+24PYiPFJHeyN62h4ZpYxg
BtaFwUghW3JJF2n6KX6P79cGmQ6AYnulSZ02VZhgvSEwJD4VOK+ZcjJV/+3QGocem8lORO52w9GR
+GfjwPxtFtFsRx8+epYcRo66qaHKe/IEbkB+mwzClPPjNU841818nxiKWZanOZjCmZiJNXH8qGs4
7j8zkB01gXp2i5xicoQ3MaO6XReLFjyRcg+SuQHhw3t0G1X/Sl6rAY9d9bZepvRShtpfdRoto0ru
Bw5uiWvAkbCLnQSrRv1RE2oQu7epQsIpiJcJQ5BCcs2vJ0YU7n0q3BS/jqdgStNUIpTMZjl8OX4u
5/GLupkKBwVydAV38pP/yInH00o/+SUKv9tkkK/6GJgtO+pxe8HDhuM2/I4xuXuh3lIZs/+s4LMr
wcCJyhpv7PhJSXG5VpNairAN3ZfpYqrj4XJDjQ3mWwFUqyBjiUl5Edo/P4/8XhmZ1q14NI4Spy24
8RqXXyX3pN+sUGR7tSOjyj++1Cejqp2vAuEWiLF6vMiRpWRn89k1/iIWGxDCcpTnCgHbEme30CWG
tv+9qLlGLJUUX3+fuVUXvGhAj1Ltevxe9l3BWSER9vAUvkCVdIt4dliDr/nCgBRdrXyg0XDfgwa8
LZa5XbsEv2Q+vZ9hgIyFlbOSJP2ZD3V09fG+MV0uF7e9JZUWzhzVXiOWBozyTaPNoFydnO/56ggM
K5cLzLe7smbskT2xe5ijDAGqLk1qJkhGXLMJLgJwjiaMBqxyq5Qs9NmDl87hIPvdz3D8rfvOv4G6
YWABUJQ/VtIF+vc9zmwjzkcBsPeC+eHEAeZKiZ8U2XW6i9R8hBxIRSzItmSi1vH9kfdpcsFVguyo
NfLAwV+dYmv2CTgpxj+fammSS1EDUZ7eBXboWq8rh8M8V3kvJjJb7oViV+8teFUj1oD/MbNdmxDO
MnvhOjbYHspewHbYKjNJTy1+dxy9tmVZPVp32BNsylJGlCj1H5OeImTFDBgaylNkRRDjJeASN7aL
blRYQu4z5ORVz6r5pf9CZz7J1HdqTX1NmV6l2OKEI7+ED6EtvSlUbUKVTbJzvnm4UaHdghcRHVgF
ON5X/LRwfF613nJmvRYd1ln7GhaaLR89pLalugMwDtTq6xjJzleSH/t5XOIEXmQspEK2NoA58YeD
aqjIwHyUyncYQI/TXuHkP1YTmp4CSFCVza8FlFrh/J5CQ2u9PrsrCSTdbUo9tAfQ8V6xe/xEYFYX
xpSHD3aEZPIGCD0aooCgHKyg+uLhUc2pIIVn5PItn2QnNEqmiml/m48jO6HHCnAZO0cIoMnWmZw5
2xXlY8gjOlxS2gDWx6DtDyFDyNwLlgaYygmofe9b4DFPZ5/3cn1fPWb+UHdcjCV1Z3Jccn6cQphl
YPl/qmdCpFquj4CV/n6wbnuwPoPjOn8TN5t0o6F5MBJm/og8KknhPqAWJji5kZ00sNi/9vwITbzz
FP/4qnAUMG8/t486rvKv21TE5E+GVcPShVK6VQzwtl50YViQ1BxcXZLHU41vLZ1zTTHH2w4eFLpn
3lUk8/jGHzFPXzlOOYNUEQMergecBGxMSYgG0AUxXluruf2aE58y2vtlmGu+/QmI6RS0+mWKPpaU
gyeE27OvPPmnXzpKQGBuuMx3GXSZ2ouTEQZMpHmko+1bAj71o1ueQH3Tsiw65cL1Ggg1TdCPavro
wfgeL2gJE6wDwxOgEnbQGII8OHxafFKdvUxT/jGIAihR0p7HQJf6lUc3+aBuqu2798EPHdfzTQXL
Yuh4/wtQx+VQ3/M/N49NYBwDDJpx1AXdqPCNQ8+K6bH6x9qRi2sdvRSY8f8b4tJOoi1UdKmR/SQc
xkgZ48T6NUPzLNyV0eq6Vpm51TedkEbxdsryLa/6Yzwbt2yKPwPgMZh7UXe3+4AKQrb4NQO4mCvR
aFl6QcRbaccMBorfZ5NVNJ9mV61PGV7gEngGXsI0NThixEZ1YsMSq33SfX5gL3Wt9BBItGZ90I+S
Lhir+qslLRWI+NGH20/MEUYGM82ELff0+FrsGWaRgyhzXO98AtR2OiOpIOC+10gLdIxZ9PtWP1vL
nHeyXER7fhyzTt6sXtjJ8z2jQSTxkyWaT5S1KwHTR+HYXdZvigYk8OCdqo+j0zn/bNJ20KyRcxcz
ctydAq0Ko4MB/xAIENTrphUZFUt97jTBp2+IxpUqYSNZ15r9rkRDYljcR5AqJSBVnJL3tslHZ9B2
/b19qSv8RAsxIwkClLZhQbuXLL1yfbjG9NBF84SGeVEgyIgU4gveec8bAovp+pblguCOGhFQS/NQ
qWqtcyRPfFzEPLG+PUG2FsJ7UCm7VX1cwufZL3KQqrRsu4IHVTF5+b0w1VJpo9MmiaFVlogrwfth
NpKB/TUirQ8NDlw0ZG+EdAwh4N8OAmtgf1LfvD9nDPVLh0mQd64mRElcY8t8WQFsNGTT5k/s4V/F
8k95ZhAYIVVgCd8twuleOjVZQZKOf+8XhZF0YeTxG1OQ+d3eTL96EZ9NSYm/t+9kWkK5/6761oa+
gQFrQjRq2DMBRSojwjkE4rbW8jzF9f742ucXq8g1pQt3IZ3qiTZBQohhRF2aOVH1Xl33OgLuSDMl
Qne+K2UWTCknJpktr09qjTnWJEsTWp9tZYPoGS47EEonbzgiIn9dvuhFsNM/3HdQr0o8dPi9sxtf
SU5ZXq5AY+TmnuVRsgDOGtdPlOvcQMCnI8okSaz6VIqVMJyiZadkurTmRG2AO3tOjXyNi3P7ernc
yW3LWiQRCxui0b/i5gzBs9ufh0hBQhXHzjGK3KSdrtgAak2CxBreOvNHcnSDnFBIJUtqegIHmxCO
j2f3wV4G2WtJTHZ8xQz4fraXM/Bb5YkwwCP4SJL4npQWLsNNDUQVhp44RzJb1Nvu/CQ6Wrp2tALQ
GQ3az4zkmlKCHriOEI1NaNZ/eFP+e07Yp1kvt0IYb5T/tNQhZk6TlgBbhH4EOHlcHn/+LJLWeniz
N3yQb+h7ubcbmOgnxrdZWg7r9wAd7hhO8tzrThXCbj918jVyFce9O6msPhe7dYGaL45o5WVLAPdc
fSkXGhOnmcTjAr9TWq8R6t+QCWQWj5B8kzA/jFSWmpvcjay2eLSIeC761uqAKK3GbuSeGTZhdJGW
ci3GXHPgNBDAej2wHszwaDtr2oUoOdEJDMB97W5UKk8hrc773wj5CWKIcAIhM7pJ56+Y4+3qwcLl
u2Qz1wvUPMZR9M2VmFYBGU9aoEotOSKji80/pFk3vj7RkQv+MUIsLkuiWt/zh0yMHIoItNZXByVN
6CN8O7sVPlU3dH60PlgrxJ8hdtQZGhqMnC7S1nPUNJT3y5ZdpaBIUScxvLxx24dry9FTzZwE2r6+
TFb4Syh8xFEj41AIU+9TBGPMvLwUrya4LobDtLRaHHP72/nrEU9nODJE5XUGx9y0x/WZl2mWAOcV
UI7UYt9gWPFuYkD/z4RmEt83AGsIBgx8NpkIH2h4e48jeNn1uifSmbSJ1kM8y/Q6PHPCZONHiEr3
yqwhGCP3P+KZqYZJxhuyBhGgxhyJjMud9VSx4eK3afroSvt11p4lunvKpu1U3xPV4DCPimn9Ac49
mEXysOV98XobdbJ3xGArS0BgU/YQ79EJu2jmgBw/QQuswDA+nMggqT8vjdA/cIsmaTBXoWay9TZV
O+sRtdWRc2fgnv/ml2NYcUZtM8ltlHqsPGSc+1NzfOTC2u/7GegSnd/lwW5bP9Bu3vpizYHH65UQ
kpy21kYXcrU1SHrghlMfw2aOjgzBsWFmp5TEWh+xrnQJa3hw2mVHEjZXaMABqgto5d5H0cqgE/rH
0Vp04NGwPEUoejSMMN03taUFnZU57X61LyQztw8GFtpEitqmvHJLnu783nmqd3xJyN76K+WgdR20
QkUyPINTvLN/BTs20rnDKoTGfMdIJIJWCJ5dFZe/4GMSWBleMM7f2FcKysNDKjIMJJnMj098YbGQ
9ZZIlW7Ydi9NSIhfJiVwD2zYp+93C4/52YwIDaXQTs8DCew+YRtz4kiiqUpCxOxABLFFjiwMWV4g
dhu5T53YSI4lEmI4/7LjfYbmJ1K9sJpIriLx8Lg5MZer3KHVaQk0n2+B/sr50BL7vy4tVcMGZpOR
a18D6Qb1OOSfksm1NyuPe8e2J9l1wUUAWn4mJ0JT+yhFKS/RW0b1+nW5pglrStQ+wl2ce6ZMLPmL
EvnYy8Mwd/AOEHMGbuNxTI9SOOOvpEbkVsBKsj+1DbKtajtuBtfVNVzbpMFaEjukRunAYa4LfRll
vutZcJZ+1tASBl34sCdlxk2BEefboAuVJy3eZzd/V0FxmOoY6bTyuxOw4uSlOTyqlITYZ+b4/PD3
aTNri0RRh6ickR2+j62vl671NLEMlVvygpQL41jDVuv57peWbvz21ix+u45JB7vWftiltd3oTFy0
g8mFnnFqBAtTxxWscDqm5Du3d8b+38QJh3RYNsI5b5jT3ywaEBxWWRZF15haBvlB8jZuF7a0EcTi
SzUlJWHaLz8Ld5lOVm1nDQp5dX0U3MVyDdrk6xE8PTzpy537Tu3gTVteWIJHDdZOtU1ruusQ9HIp
pMsvq/iTrrs6lRzct4nrvRIJaa8wD2Tb5Vxc+hyhWR+1mJE1rwaYw5DcMFtAFksN2QkMhn0Fok+m
y+Qofs5pjvekl6GJXHXmm8nmbtlWoZfx6KFQ4Hp7EQDEQ8ui4SWzVH7zqwDc6vKHgGqqZPtLqgYq
FQf/TXp/MYet8bzzDZyHIBhJWwevQRY5sziLChf4rl1LFpiuhM2unRcxb8eaTZDhnVrOTaIYdv0S
XnX+uB3O37g8gXJW9bi9L80BKGM3Npgbb23RdhXx+1VwnjdpR4/kjn/sfZfMyykAg6MjNy02lspK
7qU8D8hoYdLMBUfeMK4y7Fq5RQUOuSWZW/uKuqBzzKu9AChc0dF/9kP0GUe7Isc6w5PWuICA4Hjp
5zXuQrGIl+k9zdFo/js/UutXlSGWPAKIKjswScaRTe2/wZS0NzMFz6gjVmtXFnp+tB6Iaz3oNy88
05aol/XJLF7L0MxSg72nqhzkz66QaAbF1s6PyzvyLPV7RvxFuMWdTc9rqc9REnUVUTl++EZDUpte
kO80g+SScTrPtV6oLeui8sHDhzB+u+JeDlRxWF/5wqc9TdiYGhl/dO44y/WZF1jUS9IHIt0n4vI5
pCRQ0OI7DO+ucDU3ACTZVzbIhjSfclByz7EBE5/O9CnuILSJlmyqlb+d+snICqzlzJyFPSEfQaYQ
b9VDWZ9kbdbVgp6Tv+CAlVFGyPyc/gmgB/htZMYz0MH5AcwqrFu2o6CTqlkWGlyz2crgSwT3MkJl
pH9I1GB7RSXK8AuJGt+anM0aIOYCwkNvdZwjzeKTkewj5Q07EBxuwyaz1XvmdQvNRTLhY+FiXIE6
4yeIAue5BjUH8/+Ef2LLpmqLhLvv7DQphBTEhQLPKAE+/nOtYf+noYcHuiTnCbXoWlxheCO0/JNO
gPAERQaP4PCNpWxH3HfRa/x5sLjZST1jVNbSHKuA1D+Ah5Fje1OL76DWv+O9dQX5ZiyAHcy1ijdK
bxQdZmCbgnwO2bBUjADZqBFtUzAgxZSlIiHy4oIu4y0Q7bHp166yTwBIL22RzsBO86cPIqOVHJQ9
rpTSqSr3xgMDJKm3KG7heaRAmFCsuoMi7ihZyPTVGEUM+X+xM81xASDBEEevmopbYPGWPsj3YVwm
U4Zxx1AuZVyWATtpQN0iYksMbotpYi5hUisXH4fLnDOL1ua5G70T8MEgj9xplKspE4QckGm+6Xtp
xrkpqqyTDGlnkbprQIRIprgE3S4qHIPOcj6Vvm3ib4CVXSF+urpAIxJkSqiw1rmBgZN5pMYmy8WR
DqTv7a3gviqshyiTGHkOYMBWurKzf8EO8c9BuZefsLAY2rbF8RWf9QX86k8rc6N6FmA0NfMmgeZG
/TlcaSRDWHnAuca5Y9MBTZJWiPuLCIcAvUzX5QoEBTG7bhZ5DjvqeP89k7hce7QDxqY6UuuTkbBx
WmBCOHc/CJclOzKNbNhPyUCE7Pugf2dnK6SpZRjeYdG+L/exo4Dnvp6d/Zm3lJez9fJT61Exle4b
Oea2hDoBFB1D+pnBvER+dQl8pAGh/w6xoDGZ8TG6E19fgDitTVJRlr0kxJM9YnXgH5g+OPc3aAFR
Jwfj5jX2fD8jbmNDhtaEVBd2EjPlKpIhZcUn4FiYXcKR8Px/1vJEc4PJPM29cdXZSmZYP0/TdcOK
LzTqh3ayKO1t01YonM4Da7QwbaSzbojef2mBUclCxk3/vl2a9E4P0A+VspRK11awC65fT+dqD++k
HaaKcHuwIyQbvhs2skb5CHZ0k5gTez1idKyB1OdZ3hEMxsYropQ1zAkSmcIlD19FbE/c1ErfLIqZ
nGlrIyRZg6wJ93t324r+SGWv9kyZ+LkU9qkXH08nU8iCQ+mS0zk6xu58bUhaVdlOG29IOQcDjBCX
3DnS58pG1Ugr74utuFrR8powlb/QykRV2Is4sMW+kuW61Stmsr0soN4djJmE7/vppO+FHYCc72cR
ChkHjxtBOG+d3udENkK3gEvWaxfSW1IrdKFP0BKaGkKBRJWSE5XJQE4pY1J38/6lxVFnjQys4PUA
OqHuUqXwvr+q/knDXnDuxyozCRu2iku2USZtQ103gVCTtON+R+LFt8zZq+a66XsKBT547oOcPkZa
VhRYAmlC52TKXlwQ++PjURbG4Cdcq4+WdhiUZTARFxUo1/7uyUauRcfsriHdZ+9qrdDQU9/wS+ls
CuFDMoaMHtVtLfW3Ibwc5e1DM161k8see/TqOpHWmxLKWhB+PaeC3Z0A5IIyZXGfeSjyhLpEP855
Qm7JXYuqPA4v65ZSRqiaSSJTnfua4tswJCluyU1jAzJ9VO0jiKvggLtyqzLExOkqonPHXLXLWR5M
QjNWO6Xn71NJ37QdzAJcj8AZdOS4OzzRmTknPdBtP54D/MOIV7jQuU4QwHNVM7MwmRFXTMYEyium
SDRjmzQTAfMKXROrrlcPx6tQAst8QdOovJDlsLmSAbSI8fqQvbAAUG9UVjrfqTU13qgy1SRtDeXG
Yxt6/SNc57R0roc8R8MvNS/pXkyM6MOesSFsCaDeSJ1ggyGjZNkQGp/v46q/SMvLbZH67sYZ/WHT
SIX1+H+XBqEmi2e52M1b2BcfRJqWT4r57Jdc1+Q0P9MmRgBzdm5sHmOsqVVu5806FkCzaGFU7pjS
wBXSznlJXKhw4lccNni/Gh6EQF3UBKIUFSEqwgBqPwvYK6f2EQ9+dkEUQy53jCKpMkVpgIBSjWGS
6/RASQzy3+tSW62tZaVrduS74aq+8kw7XXBdsK7rBDR+yGnxqL6a0lCCUIIE518lCwgtwPA7pTPY
tl88T8N/m+lKDqkoa7W8sRyICDTnt9K5SDJqf+NnG9gncJHATb+oDHK8mwuSxDgaRf1idG3v2LZl
3LV3UZRjaRxRVywIPRsZX5IZEg4k/VoOTGPHCzxyaChDU0+2GUzeGBOoqQNJsHbNB8d089zMADnB
Zn/hvBeVfFTgY/j7K+LhQeqNQfNMimnElFIK0Hb0DlcV/aEUt7THZo+ZBDnEutxOckhA0SDuDgtZ
tX+/I85GCRFuIfBW7E4oAuFvwU/rqGZNmRSZHgpp65Z/z0bZvSx3ztFugmx4eSBWj/yWCzsqY0cB
+KxggoQ9eT16GSTrG23zZWUAOQsLLHTpYbXB5dXitFU7kTEstCB2o/xHUk8TFdF1fGGZvYNQjxOP
jc7OX+e+1WxtOLbLX0JiAuo6SLWH1iGQpMcEXuLzEFyzCX5fbw8IUyd8vp1WhYMVGf7bXJGcb1V+
b52LIWPJTz27l7KGj91VknYCPp8cAlYCbRBRivl9ReeIVfbM6XaZUQ+zXieuk4CjSko0mNL9HAqc
RYOGCgV3lXanRTxKCpTQ/B7FIJ7Mx/jyFMrQ6ZHxYBLam6izuD4CGr+JNPMm3RzngMR/iP7R4rql
Y28LhgCFIagrCqcxI8/Rxxs9xW9OW5vSJaLBZBu6QQVohqXJZwMGXYGuhEOMhrTNgeJB/LUE2bZ7
gVnLeH1T3sohKvcjyuzinOayPh1hPSuBd/LIeaaKHzLorVQ8+pB9EZTCOwnZ2O6uH/n+xU4hOHkz
bNN1swJ690AOQQxfINhFvYDIpzlTR+cnGNWzI6UEpkLQp7WaCXzDFn3a8sY5gVxlLoSczx4FPusy
uCdfU0tGCcGkjaIpiAD6RJMlICWlJI7pUMmxHA6SzWfH/PnNKs+NnFhKAE7L5JYimfrAQRQiDwtd
9C0Gmyvqe7dNmdg8TRg9d16SSU2WVnRtTXPWFSa8DTBMoV9Z7bEq3FSODamkW/XQPlgj5xv4bE2h
LBpnYB1dAIJWr8RhVUHe5sqFodVD+gn2ge1dm+6jHEQtxtQ9xrMVFDV69r1eshvOI4QdJhQTeMNm
yaxSACTUWNnYjXWlJlCHhbpCLn7oY13QKnUh/5MpFW3CAWl8CHkhHPt3xxLJxjSuVOwgwQqZtfGW
vutT5YCxqo2nLbLflT8gr8NftyDiFIA22KQ4Hq+PHITJ67SI9sKSv7UXyzCk50vOlnXEz3ErIhoi
uzpxcQfkxlL2f67pZjp7OQaL2Ax43OgkOjXGA/y3OF3Y0vgDHJWR/FtiH9dCXPIMqMa8508CSEW2
+fo1h9rQXmYPMlMNiPMka/jqAnWcdECXuzGk3BZPCvFkTEKErKRhz2dhMQ0ZUvcDkK1v1nLisU8Q
QxP2oFcRFfvrfPNBQdS5NWCt6tU3go5gnA2CNSw/UqyARnFlYKAQDUUgY0T8AL8NJmEIgnb+LaT6
dQOsbPg5j++H/X80zU9nwTXPCQtFVnzI5MBta15/t86MKLq5Z+m/1p/G8E1Jt19d7sbP0evtK9MV
Zl8z2RBhU15Qzo05FnecZg6mbS5QzRWm3PRxZvwGLYV9LHxLqubJI5QAcJSmMwyBA4/HmwF1REl3
vnOI7pS8SczfwOIWiN96PzT2yC4E6aMztjccez6SWMwjVrjs1ZoCZ7/aUcXBK53lYfkefQZ5I2L7
lOJSnO0/tR3OACxtqTyjaXjyg81LdLGTslHzL4JqsarZfJdXt5cuFwX9k/vLsf4Cg7UR/eWvCTO0
HWJj1aIpTH3QGKj7ZjKIRlCWSfFfn3AMPNieCtukFrZAh2CWjbKAfC2ZJFmcpEJEFZ7IbCISSu3J
36o1ARHyjt2iu5YWdsV+Nyvncsha0h+33LaPZvg1PBF6hNfrRo8B56mqpZeOnUuNxNEYOZLmXXFd
5078yXbEYAR+JfyU3cUtaiHFicXzVUEMpa4LmAzexlmSCLawSvcNGr07qfDY/1I67gxEVO+nhoUI
hOmo/Gig8SY3PMJ6+y8skqNQLdAiNS3uas7FmlRfOQVYcFwlcFr+KU1xx3aIHPRug3qspoHfPSKM
+zNrL5HAjlUUTpSWiZyNSBX6gtMlO8W/REXkcwTVy9iDJ1PehtLP8av8rsO/PkweooGrJKMZyJdc
sto55cK/R34SCbTvh9wsigZiiCUg6NIYtA5amKaSIUgwISkObWvmYIWCkmRBMzB7ycZnCVHgDIAb
rl3z+zBZIDoXdBpUEXQmLvhCxAM9pP25vmUc7nF7ufyAPy9i+uCKeAYNPbusVhFkrky5LKxbz/gk
g5He1/YJk+6k9gHLilBGAeQJCeAFJO9KOC4ZfI8QZi9ZevXViorBwYCDwZ6aJhaH1/Gp/ZScYBtO
uLhwC6cwbKgg8/h/th/kd6f6/4r9Tb8e3SWvBOQYUqf5yLYPYc8DcsmhBzsSlWxDCRlw0iNHnAI9
jLInbISFusqxDfKnsWFRoZx6Vdq3gtlTjjCnokAQsf7LgWPp5IqWqmqbg3pKdYt9zKxzU7l4pNUy
KN5ixXJDgr/mPRtxfxYdf589VW1Y/nNkh1XJVJUdXSGgr+y3JUwn/Xcgpnqf89E4QyzNqhNXcxTT
siXx/OLDiMYQDPYvziLLyphodPKnMvHIQnpenhAvWCJqpUGBHHLabw3GzXw/zEAVmVNd5L5Sn4Nv
RfyF+pdehQJS233GMWt/ejewiXxc+7TbwyYH90Jciuc0RpIJ75I5RrdGjKRvvA7HHfEcpLCe7B/v
jpls8P8+9KSce2pnNKvNv/hbPPkEogN5RrOzhblukGaPilakUqidLTd8/C+afdvtONkml/XcFdMT
upQOe74bIou3d/7tnFJfwtAULYNPLs5TYzt/qKk3bSOG/mwfGNyYI73c9U8jb+8bxF6sf+OKmWLB
PGS6sLgeCzve8s81L1pc/HFnFogCmQxs+RgDin9r5wfkZwXo+feLfrPnrXinkGYlWoChCtq5X8xw
yaswmtOXahyFuMoV6BmkKRC2JAoIiniSsH6g7xJ/hnfPI2FceKoviMkGVA0QgopwSQSvlqn9fRJq
JY0KUGE25ewrxk0YGdP+LUO1YMlo08DvdFJuucUzKJZL303B/WmKg6x/XHJ+prMxpLqPWokGXmBP
JwAMX1DldTDvS2NdpC1UQQoIZyZ4lsnZaeS6R3NhyrOwey7+e73hb8PoKFiHuhvdx1+JLxFn0cqy
tjByC8JUP2lK4YNcjBkuoCPIPCSBkHeeHnY9p6aTShZgVYkLy+90lXW1M857scBZvQlP5Q3jgL+I
1J3Bo2OOzUTRKG0GkRKHM8MzoQeb+s+5d4sN0uulM2vfps3sb57s3iYWwYUmhc6ieD6WpkfYKufh
+3HFew22VvXbQICqv4dxlMfVNxjJAEMpiMlmRZgHdUeqbBsp+w/FXLWLsX5H9BtUzgr6g6GwA04e
++m8M5QhzgRGRYZwEwWOcYTOtg5CajIjKY2q2yWakDWvdwKGu+fGRgyd0wvbGtUqR1AoJMwSFRSu
XApDPLlhXsyhYn1xf1w8PdG00m5x6gKoi5LtlyAqQH2FUxBVu+Q/N4Osf9kc2tHGs/12cyDfMDQO
ooMjp/CsR2g4UsQlOwToiFEyw9uJXGd/dPcEnYse/DafSQ/xbmcrff57ze8X/C5hY9J71bcLwGtD
XEG8eA6XHcTFXm8Q8cjPNBZ+NuLcry7oKOcyciCGdbyLJNwEk6918EIpKlkQvUEh2taJsphC6wGk
PsBC+zUBmEUFzjalyOfIXsjuUUMry5L74jiW8zOMmmbNlHo1vu3kkWvdvRu/O123Z4WFS6ASKRhJ
EPH/Ga13XJM+tJDlhB35zUqJrwO0BboeGU/JGXn1hHGeX8uV4DqY3WLHcyjvYakSLJPQHhXHZ2Vp
eO+4J5Zmq39Augo1jV2/pHhL8tN6z1aBm3L0WR7IdtZDwTBZOAtKTumt8mIFb62ySytvZ5TSNzkF
SvPNSULEmKAEVCEusJlGZhDkoIFdj0OJBwYx+TuOe5yOliKTSVZzg/gVpnwjKe9idZ/0FywidDMD
vR3IHm3mU0POewoM8CjD2El19TLjazMynbbd9oFPN2EGdOJsEhFZn+r1azPb3LJ19H/MEdv9gLSZ
N+iHYXsu7a25Wqk8dUfAoK9e/2gVC3GhCzoChjxaI3HLluWZUamvJpcdP+JHymIMsYFSta4f+BoC
vfGkrHWMPT3Bs0I7LbcIc1QdrvJX0GOJSoBMYtbMx3FCG7+w6B1AxVZrpNFlZ47H332EwCUHFW18
7u5m7KxVVKVlfMVkC7llw93IA+F1IUNMi8LQMkCvt1Yqab1+owC9wBjMrdi0wU++610OfxzDPvQn
s0bHBVwjVeRgQqdCQLrHhPUNZYBA7WchOkrzRFTJibe4zthRv7HhCZJ5TlT6e6E9OzduiuExqAjk
rMdc6Mc2kcnLMJMpQjiIim7DQlJh3K9aw4EeGrG+mH9jRVrcvgCUMWzbUlTmvyrpJVJJbeGFFbGW
p33kSbzM8v6Op53frFDuIpL3LE/xKiQFK0fSYXcRlekhs6eoYnkhl9vBcpV/tn0QKweUOmJJd69a
PNiplM0jWjJv95Y//4JDFFCUA5ifo4u9aAVDsLyqIhmb80X4vGRUk30SXP0x1TWWmnnHwJ3OgHVs
QplsZw09iD9B6+4UEnEnGcYjy7DjG7+fbdCub7iKbt+9QnOuDLv83OYaYYHzmegladvrJUOwDekH
zyYU+ZjVQ1KVHHaXFTc4+KoQ+o5EgGplPqGB7R+FhGj71EconqP5U1l5EzMa2dxgio1Gkf9iHPM7
rRqlY41Ua0Ft78xMrhZzfFDcki+tWIQOu7jjDREoNcLAsQ3SwwVweXF5ro2bGdN1akfBkcH3PO1Y
9+vCp9wIubfUbQaWPd0Wo3xG/T+N75sXb/ulcoE616qG2gB7Zu7rkC6qBtY1XEA0Mu82fm/hDvfp
T+OXpTg1jNbjKCWcgOcpE182CmpSfO8VTR13uVqXhpA+ik+oLUquBZLO50YGBFXsFwSKD+BmLyiR
tUnBSpPB2Z4LoAgs/CAHVUJhIBfbQapCwhwNLI5uahRnqDUx8OmlsJUskJ1oc3lrMSDqYnqg4oUN
JHMMIrXS61nzLDcc6FeETgDbE7zp7/hgWHxMpNaX+PliGuaQyvAUiHL/tGrLQanSaPSQnqncFt1A
PJu/nHHK56j5sXPgpQpZt9fq7VGyo8p56sbP6lLebzUhDBK+ImycpgXXBZ/FXT83ScUFOdjB9ZaW
Y7XAWzbr/knsrijA7CH1fhJmrLXXKpW7yU6V20YWyUMHKjcDJ2SkiJtKral9IQQOYNoDeiZOrwP6
I/jLpBjFHNNagoJQjnOIbk3FyU+Tq6pZ5GyFPMKfd1u/TdI6OGyFh5BWu2RhFUok3pRm72SYu7WQ
LcSfjA3q+UFVXGpfGVf5jVJVNQQ+RMj7qUIPu1wNppLQCj3yK0Od69WafI+tYLoxxYGAHheBfHiN
/Y2ueuaoz6V+Xld2ykzbrgvDPjnfa6tCflv9tjoPbU4y36FLiz9jpSZuhGHOZiXap3E5oSksgzT5
WO9+8TWkNzzWJ8YTdpcPRNhLKST7KjKVLMh0vg6LNYB5xzCyw6tK7WDlwioJCXy9psLhN2vqTgD8
gIuZOcW4z92YcJe+3yXpJO9sVHPhyzAHgfqL5ZO7bwOCVCT/zuTmwHzH5DmrJOJMCKsPszhpQa8Y
ighnrGTHokRy2QzMjJOj4N7jnUl99Pb0ed8YRLTF66S+6ydBAFXpWUM3wLYQQTpikiRZOEdFThJI
Y0nwAugssJ9QxtOFh1TO/h9wKOCUA82GhMUzJ3tD6NmVUlAB58I3QGaTGis2tJEiDj5Pzos8X0q7
T6Eepz5Vp+Bu9mT6+Yfenmjd4bYE+kb5Gwecn8zaw6gnAmBxUm6Jhxt7JwXyQDMdx14CWt2nbSU7
tvWbiD5jE+9e6WEtZsWXaqsi3f6B2E3k/+vBC+Yl95yu9Mxjj98a7CX2H5z75NSu/SRqkFTBAO+T
jAw19oFcGQ/xt5lzD4j62dKkKPchIVA4G9LwAoGVqOLS8gC/iHVFO++Q8NozWlIlVtKW6yw75ERS
J8pwe1ZPt9+7VE7tb9qVozDSlBUoRSB+MD9GJHy9ujLxJW7i/kIWiWPmqwhUq2tRPffB+gg568fY
wEOCzMfoNFS47DueLqKWHWfV3QBVbgXRIGuLixnCZ3eycE4+f4UFSvV8QIvQiyWCuykJ7qkioOn2
5vGn5eF3RG53t7kckJXYi0FZtJ1B36Oyw1jfQjtA+6zMPtsYoy5eU+RhUIjZ3RYNLoibup3atT8x
ASA8bk2wT9ipyqlcv9Bape/PsTQFPszY6MyWmI/2IVBZImTzQTTok5D5n/zmR2TkJ0sdR+mdqxFV
ZerDQBfWcEJgDbH9KNBW2Emnr2C+x1kj8kvDOWr+6G3VaHgLEPL8nIwNys2hf24sffDM3TxjxYsX
rMTTAgTAtbY+N5d9yeQnpgsYTccClYOCBwIWBS3L5OYhut+AxAscfdNCBFZWFKoNz7KRvmfhy9Rb
SUEew40DcKATZNegLTsf1t3HPJ+tTcfjELRG5Xgocu/IKbvdqU+ZxTb9YpwD3Lp00Y9GDULesl/h
Rl0PxFaHWbxY12j0X+3Rnmx1boBnWPswqVlTwZrNMQWxv7xdKEb/OiczyIDqCgToARVTduicIA69
kaHA4NgP1IdQ2V86fuMlsRpYb4q18bDvlZte/1zzUD6vf6xbMq979fZDQaKZgIwB9eHJSAB0J9HC
o60Tc8vw0q6ey9epUcwd1zaYoPcdKyExjnkZOwxFFAy7FTJ9HIFIu12RJu/sAJg2gE+x5wsmWsRt
s1An+PC70YfSR3N9tgt7RD3EnNG5ZGeMEV8SWZiRtzHaDm9MNXBYJkL/yebVHSESUkqSr8e7xBET
0flddmOaxmi2vGcSPcTZKSOe5sxk8CZkavVg6rIkycbeo7rinGcACe7axFV1n7zr7rC74RJ6UD7k
32USMaXgkwTQxPuqw8T/dqtWDMa9YxMX3OHKPnjPmCMcs4+8zJ5EYNkl5Rfo1ND1naerkYvTHO2s
vxszGE0Vrx9q/nwNsYJzL0bz3PCMx+42mb9RT7q/96VkvurNSn5wUM/DW6gCR0Am+hqF0yNsSds0
o0Bwumrm+dbeYhKDquKzSCWJYqBxl7gd2NMV8W/RZUdaAnLdnbfjZ43zqAfaNzmDLw/0306vtbQl
ZXjNmZxNFrBkrYq0SbJtpMo5AjIwlwGCh3IHZB5qiuWgy6VeFu92qk1fDkDHYGx9y1VR7xRAp/pI
O6YivPkFoXGrYoZq8U7hWuoEiRDupMaTxeh958Tb9wf7b3ZJTkeYjvQciigxv9ACVvl2TBQchMRr
Tmv4jqxXd8tlbGG2uEroZmz0ZqTJjrsUa7TVJWGRqOHvHb9MbY6Z7OgoS0Wq3R/VmN5ld4gQtXo5
R4LnAPh9F5Ct+lFVCxHLWs4fGCUodf1U3clToHFYkM5x3osqc6+K0RUApk/7UzR4AJKiFcNgs/VB
QD7mj96eMLDYClKuXE8uNkW+O242zx1zlIgVp+ylHxomFzuMe+hvOZqFpUYI/v6OVMb4m27eykvI
FEYsVVfQxqaMVRdZtjYUIpEtYF0t6kocqJM+uArKi4JLrtkvyLxp8BHkrHBrp7G9cv7/RGlcOrY5
NvdM4QARzRt3efusniUsjRKeOs6rnoHQLkg9aGoygKwBbgfBF5nmf1yRNJUtI67UDf/wk4ujtKkD
gMLBv5ihU1WeSmMmOBMISg4l8nOrVipsZgGhbMQXXQPLGrNpDYAbnNIG6sJ2Y7pOFc+R37Qpesu2
Eh3y+iM/ypz3QT8AogLmpTMlqGaGz+8HuCao4xN3kT4/mq9zNGgAFted0vXYizJki04wfmxt6oO0
AL4vYy2E0GAQkJYUpuPVYIKRK9/3MOKCqnp9i7I6v2InG8+2Kr/aqm4jil64Wz2wB+dHrE8f/Moz
qs9egUWez4AoqH91bJoi9rZEFgBHP8VWg68FUM8YowOzjHIQ09hp++gBrakixqpfNqeNUx4eirGG
x6N2V6O29m0uFxFHrcN9HjLKnDFawATDxLfKCKw8TFXusfKnwGjWVKpj9dDqQRwuWt+9/zBqtaQ2
+Zl4VnDkUK+Mm21DrhdoII886zLnJi4j5hXY8lHtX1iiIh3m0S3HMqhvZfLLzgbOkOY7KKYNiSmm
7b3jLObfVoER6OfeMIgQGd41eYPCVj5Zr0qOi4owuXQ/NmzWDBr/zYahg9ZVCFPtOVRlIgWQBzEP
jXZ2Okkv/XtVYVWwf2ZIwfEDCqMp0CSY3xWGyUeIrgpHfvv1CFavF59uYT/5d6tUClIfpFJTGHR4
rrL5MzbrC6jSsVuKsyI4fxbyZa2iJqExMMk5J2I6qTJPmtKDLP/xdksPH5bAp0fQyh84Xrd20e6E
6vw+H79rjPKrLvMCloFHMbZIgU8nbe/zpgBaeO0hHElR+WwC0eCx125gPCjsIATsBAv6W7R2B7Wp
mzPtg4tiPUdlYqdzJalBH0UdeYKTjLh5H0PmkIlvlIcizgat13h/VyIfF7mUgRPaHMK79iuOg2Ns
yzGLdyjE/TEUzWOl/eIJtLvTeR/K82M2HVyk24nS3kGnWDY/o7/iUtvZh8C8ViGJOR6PsVw2qorI
lWSETSZh5fZnTy5loKKzv2hHqRsigPSLx0CzY8lhfohu0bOB+pP1fRMCrRowzeibMRnvlSOrXa39
78Fvdq6bOq+AFp0EO3UdwFd1W6dAbUdXiwOuOXg65xOQGtWHieAfW0u0YejkbrsgNR+Eltvuw62U
Wnf98PqQMy2XOqn1sIUGdDVICn+bPv9aFzEuPg6TfRx93fneP9/d2a2r2qeQCqPrtphxM5eq3kmx
zApXFlHw7PTY1LKEt34TEuIMBVsjbsku9D+3umLfOk6TiWTz1eZi66LLrL/km5W/5Jn3T6usl2Et
B99/URM7v+Nr5b0A6d65wEeGepX5wGIdLHCFPW8KaeAjStPopo9klE1IGorJLjfGoJwnYuNAKTbH
sPLYNTAjUQGsjthPYmhgPav9vjmxSCbmESd22OdK0dugQyUMgArw5N3ednazxrDjlVTKcSS1oZrZ
RzNNmujN9wATTW0dqUlrIpCW1xWbs7sgDXsRxzwsu4+2wKT7F9uVCNfsKkSh0/bI4QTOcAi0MwoB
eACB7fZjlkpsH1t/uIQGivs4SFZCHeEwK7he9gdZBpUfeIsoUUDFM0gUOQENJiJDMWKQ5jPdjrSW
xziixDEktMZN9EWrYcAVLD9OcqTfHrJAJnF9AzkVQ4mHQzmKlUmDAp2gY1ti4yFAPr0GSstUof/F
zPYSwzkATGuGuk63ExJlSQGB3W+Sbm7VnjW3S8rOKb2nwOJC5pZDsqtLgEyYvaPyk2smOpuLbzb0
rHkpucncm64D2PwbFxWFiaJAK2ZNPjA1cyf/V96l69RbKh2etrNr4NK1xx19lRhNx8gzcFJBIm/f
wliyfmu/IRk4FTYWkDEJTamyU6QudX9at0s+rOZnmn5b9tCLqfY0WgXqPrD1eMEXqjqQ6eEzvDD+
8xEdYFwpEmIxTY0xkyOWTFKIdLeHPxlHNcaoKzW21W5HyfSp/GkB3D8NzRqkhNXKIWatc05AFaVT
8yNFjMGXWcGCK7et/OoIAkImILKJd6hlXRhXPtIWWqX4IKFpxweO5cyU9rXSbtUrdnM/48+CrW2V
vYwMLYl4tSiPhxXI6IigUKIRasVUS+HBaJCYePbktX+L8w6CHYRdaZcqxQoaf2SD5Nxh9X3mjdpj
oJEQioZbQNohspVIVfenCvZSd4fLeIYXzOV6SiWtTVfa4CEP9CKaHxKDA993ixjqNPb00PJybtZv
YIjb2KAQ3YBpCidLgUCKMJ9ooUzb9rjC3mbI/vwLdzS2CowMe0fCJYX8aw7CfZA4eG+bT7RVmU3j
/FFHhfGN65VZ2eIno2gWzSvyPQRVlH4Mr7Pd/U1XkV2SbbZT/dTS1dFem5cXiCoDxJZ2aCpkSFY2
UHQH+OpI2A8+UcnseH9YBj3AUJkIErY2R+XlHBkD4hb9pt/dK6uTmoAgyfqRWzARyeiBqxj2oS2l
UXRcpDau6o+H3e8hGjVB48OnDENsBvHQercwuomOR67eSRZSwZPFw1wbC+UfmCBN1+MrBCVC+IMZ
EidktYR7Pyc0fJnpc1c1zYZhL7kvNCQZDGe4y0aIovg6OM9idU0fvfL6U55870RtcUxSrJQ7Csfi
QyFTzbyIJ6SqZvYtbY8FGAB8kKjxOdMS7z9UhARssh5VprqV0Bj0XxVfvuI+RwNf3FebCR18vpjx
KBEKkV1TS1/zDx2x+CrtM8BE10IX37e1NLyZ7ungsuuGF1Wo8cqFbwlKAPzJC0Z3Z5nexfsGt4Ax
2ObcIpChu7BYyrqpQ+cO1oGVNEDXMiOZ6cwH8BQw9fn8CT9aHYeEdH+pJbhO++jX1rExpocz3C7+
1m0gJH/I4KhLohaWariOaeU5eM+B0AMYCd0TmLtL7vgeJzR/Hi9jsTuJ70X0+/2TA0W2OWyhwDKm
ydurnAfnaJwTl6+06tVYvWFfH+F/QZC0ekymdR5GIB9LHveYFe6DRS+huC1kPC8P7Sg1x6Jrh70t
7UjTlkRriQAPjQSy0amGZyauh8c3K5JzztK35OyEZbE+OB9f4XuMxHqxREzH6AyT1pMUixLxoB0h
/AbOERh+qfy2sAem73Q+Y4nAsotfA5XH2psnbPls5OnLrnG7RsrOVqYnrugO+fw6pnnRsXf9rcuY
UYuMFLdGxyFDbElLRk866+05pzez9UTydk58XpdsjvfEFXFZ3MS+IKybIoLDH6j8X2GxF0ef+jM9
63cLAayl2Ou8fxsaA8rEpWmn1fDe32px2y2srlP2nqGqQY7+889PPB2dT6AFSHKavtUyP8unl+au
ltrV8B7BwNynPsQt4l57w5Vsfafa39yISsxVeAp3w245CQj0hNeWF15WY1CvE84P+oYoZmGaMjas
0/Je0kJGGwhX66w/7v/klaxEOaqY+jFZPEphk1+lOnAn5FdKrucDYTaU8spc7eZrWsFbI55qx1i6
ZCccjBNXcbRpAZNdTXdOcYs3XuFMCcLkoZ2NcT4yvdFOOIxiiRKK/JkgvWPP5bCdkrLswHxqht8j
OlMQu6wfhNcfEZnz4vkW838xySKjhGKlYaz4cjy9SjZj6B+WM3g3G+ooyGcltbfX2LuAr+1oU3EH
EYFmvl2unrXIaQjmxwwMhpwmgmJNO41TIZpsqxlM10n5pA6z67yDZVDUEhEFP9r/ZP+Vgu43Cmu3
JmF82eN3BiT94PtpYxv6Xauh67PXQ9stIK1Kd/SMw3xpkNdYg0raxiaDThoQO+OPwpkW/cddHZAE
JyknH3Dz3Vh2OrnERLSdXbu0M734YRo01WdfXkz7zJ7rMmSdoDqmCGEeCunHqWqgiY7djxsJQ2T+
9rzJVJJW9HHErYDbvwWls8OAvV42D58n2fihQvVRvxkAC11rNOJYhx+NQ2RmudYfhBBFpe5hOo4Q
eCEgna05yHGSxYzhuTlNz3mWGN96sSQRV1h+22jHJPO7xB3PQxPuB9Ss0tKM1Q2OhsItiEOXQKsm
9NpfdrXxOaDG/fplxIgq8lb4iYmdIV4WYyylG5Lwa6tBe4xRx0wxfdSerRmwT2OGmKgfMgs94X6f
FdapxNUQr0oPtQDpn2lSgNxmIFlURllroPMsx6XpeDu9Xj39nQ/a8UXn7Zgx9MP+LweMZKyfTu6o
IoUM4RVCpcDxiPDkcQgva7BPd0Rh5tyu0F6yQ5IGEn0KWdW+6Gsc9SKxz4F5yYryPMyObvy5PGeC
J7ySMGO4lhTRKlKdbNE/H+itoVRm37iXTA8jUoePIqImeuH3+VcEiPQ161s2K6cGRkJXEauG/5Vr
ZbuOMHtBsKC5P29k89Tmn+fgxzsBxR5Ve4GA+R/eISCdd9hR5708lYmIpdunqn7aTaeBYzroK+PC
KrT3gA1TFwiMgrAxybCpRxwrzTmMCQdAACdWzFF4RDv+2uIO3+lKjYfGINXJX/nVoY1PtkT6BNne
lvrvEPSFQhW+eACRC13KCtFVQSaako/p/1UsQl+q2fE177mImb1SJBWwlSwM38ic1H9vervZbR8V
+N7SGG6dkT3TDSnP7eUvPzHzB1AvxIl0XzOmbxtHCn0ya+dvSa5pyqNi+lZjOPfUFg+Qft9X44qy
wVEy4avM80gfw7t3B8nzh6r3qf8UcnbABU7eMV63bQNfVJj5lZVkc0It2AASNlnDN8T8IWMqYx7U
o86MkUm55013yB/bRWgJzRMcCtKLAVb7mXF5GUixV/WyHg4kIQPHD+gtQVIZ8D2rSekexlEFv+qy
0Y0WHDDSE/HmTr9rYqPt8zFX3YD+sy4FgwQdvxbrK3B47n4/O+EeN1KWC0Y8XNuHXBTpHBJNFnb6
lRUFmrl02CgKmY/gTPbksbWrvxbVlwapmih1x9nyaO8Y87pH4UTfEYvYFFtT5OqP+6Q05lx6G08u
8JQy1SQ6q21iwwrn8Xbjs5vd88jVsbSOKQU2YFlBbea004cN+6YnMsXtfx8w3Uyp1Joq2NHLwKI0
mDDr0V20MVfFVbIXEhIZkUEoBoJ7Z8h0eEgw+QoKvBTIrmAFcqMWDDOvIuj3jy75pIm4YsBtYfm3
eVCFEXJQNXd/nB1ttiqtocn2UFQBpa8vvV1klCTG/8fXiCRDO63Q1grsdS14loPrkC3z8b0nrLLm
0+Mqx0SwC4WwRS04vY5R1ksK5ky+ReFkVC7/zjEJWgeRLuHgRVKPNyk5DiPkpnNuKnF1Zo+t5IvT
9+wGl5KFjU0rUKOJkNHK36XtPjtpvP/y8b/VGKpBxS8RRL6sKeiT5Ch6RroFeMsFFhwVS05iyenl
Su/93yn/sNyXJbawu0zjqSeQvR3aUUnGPBzOa0SIQObfXW0eFHLwIIcEz0yZhAb/lZX2GUs+o9TV
XodWr7a8LuiFoo7X4JctufzIPt1vhb3lAS584df63QfoVFT+rw3nUKUuj4yLnALmKXILAUpREdaM
xLaBFQo7YGjskenVV8rPuoLIC7LsbutLgY6vL5T0n6GKCVGL5f3G46KJo8hmr5VcagdrE8b5JXGG
sYIHCzbfj74lKK5RwU9TvQkTcd10JlQ60BPM8FTY509ADAmoPwKajMAR/E1Fz24SFOYQKVbaqubt
cfehAjshwyyQKnMgnkLS7xsKVLASSc2J+RNThpY+qgaKHccnB9Kq2S+1SNglh+tVelz8Q+OqCQFn
wc2RM6HFZ0n1Wn2F8Kr3dMiKb3qS7fu71TK8Pj58qo8OQ/lEtBV9CZxoiGX9G3MV6ACBzm+X3T7m
FabmL58nZsti8Kri1rPkANaFSFvZdbWc3UwgPQ5UPRK2R2/UVzF8K27aMOc5e5DJN/6+IQc+mV6H
n44eEqqgLxK+tSg+cCGGS0XTRxnH5LX/d8iauSlVSvNNJQlV/OghDPjne2t1K8ICaaZYks8+z9Uf
xRRlOQxadXe9xkxrBh1J3NExM82mw8497nKWKc5eAT+cCcUlZnmrP+XmD58Yk2jdhvOoHDOJvaWm
jnv7wLjeGa/dfrEmf/BtmJ5MlOG4M5BLtSjsU7vGLR86DVwMlEPGqbXPXHMeR+pQr/MZnc2EBAiI
soJ8zivIh1hlpnaz8RhkwZKtxKBH56J0QDN1hnymlCOcyKvOA3jF0ohlOZYbLIuguUijdgIaiira
CBLkFIfGDny2rzCzwpOVz3aDeFTeKXK7eNRr4yQI/liYQchmxa+e6qI5JZHfkZIg289qmMBkwqRe
QUTrCzx0jr928DV0iyBmRiOZuXvGyXBlbBxMl4maix0wxEYAY5qKV7Qdus+WeCrLnk5pBBQAlfC0
aAgLx+YWdK407bylovbG7DG2v+mzOrCYHRClu8uDtbuG3iMvlx5faAuBu3a7tu75Mg5VQa9Ekydk
6oCx9CSHdhX0VkR+JyXNLl1CZzaMmcT8YfYXrKVLRtyzJFJyA9F7UlO0AF3vYdZJK6DD9lCS97ra
hHhH0NpH1nlr463iCvVjWj+RdbD1AsPlPoFXF8yP603gn5lN41OYqp697POcZedizNj7AWz0Lk+N
5rXLoRjmc52fbOwIpqTR7tBuL2OIctibt5EGcd0yoypEvot/TxFsOXPSdOAlaES4Q4BBCyK/Y0Yq
jzIVGRbz99dUZQMhK5OlRkqGHpn8HZdlvcIbpDj6mXaUyhCIWpUtLMELzP/cgWLgKj4+02CtWiFp
DO0Xt2dw98a00aOrGGBhmXLG/JEa7b4pE7vvi2f1KfOW5AJXTb+0NuWjyIrxQxE8UPfJxB3mZkUo
gAY+qG+Y4zA7J40Ole47IYb7efXuFvnUuPDA8n01ywdG4kxqMRFlm6tKUGiNCEYw2/wRH14TdmaD
K1vp4Iseo4+J1VzlgE8fUr2oCQQO3wi9EpAeNsOKbDrjllAfTisnuMKt4AI7IBTHGDT2Wt44Ji+h
tlNHgs1OhlfZfiA1APfPErA43PAHJhcxgsRWVxCaE0yEOBh6LXLiW3IJvAlflfhZ+Yga+0s5IrL3
hDhRum5chOW+GyO+Nb/ba3UvpiCk+B7IE2sg3q+051lgfm/1+bqYSPcldAlZYwgef7mMjVnLau+a
+ijeFzpMz8aNX2vDF1w8LkLrfYjaME49dR2aIFBWrtGROLu+fon0NUBrFOqxuvfMJQnpzWkrVkQI
cIDj49x98sYSRsg8LkyAwXtACfp7odfUejQxo4zawz579AeQpTy2xZiCv11UW2vQ0rraeSdHPgNv
Dj73f97hUe+r4dqznRpHPv8OltZOM/Gac7YlzZ0OAfHUExljQCwBRlEcafCYEOEqDD52iuHm3AKI
jDEs7ADYTcYoj1qLheC6FgYOoP6B4oH6895Jor5pY8EtnG39OPb0+UrInx3EmRMYg+SnubJ6QuTr
gcI4eG5Nd0TQmwIgbHMl7wTeRaDCKMfyVDoiBINqhn+JGpu2HDnDZZJFdq/Q5FpbKWj798YzmpbM
mLzI6xkaIza39gHisswOrNomKRFCubVkhEScWinfnQobbMsePiGL/YNxZtboH8XGseZDOCq8Cx39
TPfg8n+SO1eqWj7Dhoq3GOQ+spINAEPd7yNMejLZ9loRLewDn/VLwHU3TLNM1uXq/SWJrLHjbxSY
Nb3A5xOr3cbO0L1qfx4O9Cq1HvxPWSYDNhm1GzX6vUdV1BrRBchBuWbyNvCsx7qCsHl/jxvo07ia
/5SQGqnMpJrsci73YXbRJBGCPXOyA6SCttU6CgGY7pYTMMRkNLkKFeB8VMm3vmuMBvtfmw1YGKEI
6qSmyXb/g5yWTAtWJ7F95h8s4wPwJ/9Uj62dSdBGsEV2UlNGf7r2UeMcTNrRSLn+Uaw53fmPEeHg
5nz1D+ivBlbyOAh76jWuYp7bH2qfQ4RA5bI+h8sQaVrNU7ikhvVToYFmUZdY9Pu0bn7G/sDNuxqS
kLrgW71GQChMVSlL5jDpUmXvUFBNGtG97qEdbuwmLl9L4BP8TG7jBfu0yG8Bd9o0m84gjS+/eFZv
YqM2IVqE+IHp13ExCJkeemyFIKg/T2j6KGkIU/8Uu7abXnzwMX8k3X4LMTDPkYHpPuxbLtOZjYmg
M9VahOhcOVIzwtmXLR2GSFgFgMKe/LYO2T5CgWLCLG3XND2RRCkyGKH/fMxTEhEYVRDa9a9ozjR0
SN/XJJoHo5wVB2xnRlJ6v9lAZ0/mSF6hrarobBqhuFy6EkQibE32674FIE/VIqbVoiIIspyykxGY
FjOfBTtjlKf4OKqW7v3+QNJITp1WCtrg/8APbgToUL1LUGuWTunXs5/P7m1pK/THp6ZF2nbl/GFk
EjgRZko1ddVDDDxsZRGyj+LHUN/mup7F3n+K1CN8C8uiR///T/5/W0ALI3X7uDNDRcGekfya72Id
beRfPwQuX9YMhWoEMK/I238A/bj1ch0SlI1JLFXsIK61DeSnlHXnZfy049WB40BZ2UfxWGMu6P/Q
e8i/KNaCa9c9ks92VJYaIXtn6E8k/IlK4PihRbHt/qalTY++oE13xuurP2GFMxOOri3thvMm7uzZ
Hgftv5KzM8qH9QtcM0IYG5N47vfF6gF6TV+CPkv0b94icQgXGuww4QyS4OF8z73JF546GS/BbvHU
v8gEH0F/zmm+ObY+YKzfwKoB+IYPP7EZZ0n+SWF4FyrASEmxbkFG++vasOQ2aVbXELgW1G+cNHVk
4EYgR9JPuIKf76GsKmYCCXDHCGR5fn3wwcniwipvdKuy/nqDrtFp7Dj8c7BSbX4sbMhJdXPPyN+7
ybO7miKiFBOqS7TwPSxWTj14K/XvHX/vF4W9c/+AilsiNGQ8DcUrWb1pe1l7wwLAmufcrBKe/zQW
J4MznPltx/G5xOzCNok/HyVlUITY2HxQhfqrv6tka82cQYAwwNXeTYehZwqkqrO+sgMObkR+I8LR
rTvEQ3Uwcf7RSdCx7sLVudJgLCEqHM/JSB1a19zz4grwdVJfZ393L25mW3gKWqlxLWRxOqgXoDsM
yzPhGGkAq6fwVUEoITTOgnaoEUZjFT2x2npkjLx4WgREKaf5BlYOW/l6RRSGzIkgfE/lKEOMD87o
gH4CEcGXMqj5mqFVHKJi3k4dqIdxUT2IoVvcKhFCYNG92oWI0Pxin6pdOM9EeuCC/L2O1MwoWiXt
Y3Dg0f8igz2OXuxbBcO8/Soaneipm0XSC1I2V51iz1U3jEbAEQKT0KB6/SIAbyE7Lkz2+IhIOlcf
yVEgimoQ1Z0+mga1XhF3DWIWq0VWfDKeqtwfO3aRoI1bkLF8Bvmf7RW80t8/3BGTOVXp38H1GfBA
F18/pPXM4M6KhdcUTfJF1k5NnePyNP37ZxL7lbVPFxNc2iwVMrnhR9Z6L+eDIdkC4oqOsLOW0+D9
SS1zlSClgA0nW9bIfzT90m6BSYV4OXJd5lys8MeFXoTZyNwOgtx2lgL7B/rdRhL0KSGPNhK0jJz9
yKKpiqf9/xYM3CkCS79X1I9Y6Y6KxtOqgUGiOX6ewfErrJ9u5cr9UPq9YpFLokFO30RbaZzeLfYE
BGNAPN+1OFP1W5PoBIqOZ/JAVU5bqSZUB7ftRW6qahQaK/B3JNyf5Mhhe4KvEOMWzbMZzD+PBYrL
Y/9CvCi2c/mhV3egWt/g+gr3vyGXZxi6hluilYdRK6Vi8BmUrTQbRCMP8alJ95tNtuNVODPh36eY
DKs/rSs49rlgBXMIoHP8a7ZCUFzHxYxmmUSyodqYLtpsyljR0YNgs2f0wMHOoB6qCmljKJeSWyLD
ms/T9S2JN6irti+V1q79zNAcS7qeL4jAgoZoWGDEH9gJ8yDX+DB3byi2FEYLk4fc8OtTH6Cb02Ny
wTN9HpFcRlLVjBq4naX+YEcPPWReCxgNrEATSJKN/CAzfQccNbH65WSvl5w3Ip47iHICFEzXn/Mo
XD3WEdb7q18Z/BnP00ONZtTiKwKWNUNlqAluLhnm6ebzJhKQF7PK3dYDlri3KGSnEYa7uFZ3O5jW
vJnuxMaaK64dAT8lJK28md5FlScdwibCx4Gd0ok9zs7NN/Rzg3LTDLP8K/5ksU3cwldya+4wdyv8
fflFVJmEUxs9M2+zMxnB0+ld3/fBNVGb0k6x0LlUFKvvakLgt6SiM0DDaKGLJKAtUhuAJAdJIl3e
bNC11dJvuD1Glthw26B0exOc1YefELgFOUEUNqLqYaxmxtumuGYInZoCaJiyZdfggxvhjZlxOnt1
loCQLNmy6fGZZdWXnlYezKG6lKJu08qd6WDlNjp9D/X4MvBr7jRvBi+xT1EodxgLPC3a3gkbQ6xx
I02f2vYJROuzZd5q9jeAKqd4LlELK2i3yuLSHCUqmK0dygDVradpUbDl85WG16XBHMkPhhw/O0/k
62CLkKxlAi3cVh/6FJ3FZD5PyFHOanCGrl02SukMYlOvIb6i+e5+itTfp6bHjbFUTkoAHMaa9pfS
h5LZl/yRVXXxuvOsEpLBx1Jb7noTPeWwrg2CekpzTlolGCOK/flyHiQuItcBRbjXr/X+QqNupDxa
gU3hl8pJhwwPHkzTmWwPSlEoysNth2BzproN08MjD4I8OzDWHUKtoo+WBjyz/e4LLdqJ3MZVESfy
8mtMMMKSJbyYv70ZAjuTHUrYEU5vxA0wuDEToSKKq+6D/v2WfDM/+Bh1XuhJxSBeSHPvLuEd68EU
cXVpb6z5wtAVHpoUgSQ7fjzqj1Ze9nz7lNfAT4He6fXy33RLVmWbwerUnN3bXsC0kWWDCVZQ99CM
i90xxFGyQutWTnmlthqm3IYZuD9Ub3UVQlVamcvnNzLN58mRAVjw4QBQ2k1ypOqFxtclFKGrt2Bz
NBP2xFRAV2Nk3a5Cc5em2vfsFh2/e8xHd3M1bp7yM+n8LOh8/74b/wZwNAVWbpoYzMr7Hz7/0xWh
f1s76zjK+ibMf7yThMGxCL+A6kbFlzQwNRkWvxyD/2d5bOLY+L5fwpINHHHJWNfFAzqLXuW4zOqX
q++kClQmMDaWtpM68TTY1rZhX7KY8QJsdajOIcIEtsupgXFafC6shhU8vMUf2qedDrMp9FYosv3z
nBT1XLzToC/qmpENKU67LXS53nwrDxL2RruYix9eZr0NOWPp7SAGg8v7Dncc10w/TaJl+9XqJLgO
+NPgWwRkPH2X6nZ3quofeZVv7rDYhCjI6qXW3bqlSElTnImzUjPi8uo4NqhYrUlRbUpQXtkdO5hu
sNtyu92ag7T1vgDAjbwTBe3g2y5Kz1m7ajb2UAPyJX3hg1nJEglmZX1VGPRSoDPjYE5ghr4BtQnv
7TTBd/EpTHUibg5uJEZhAIQK1+dbb09vqVvk5qvfki5hpOtQEZLpZGFu3kVbLMTkpGA0PhTbo9kj
scjusUBWbXnyS6aeC3v6gELfOhxPfWeL2YJQu34IVKK78fpErouSvNzc/iz2ixx9C5jBivPW1/Om
dnHNwAghm3vt+EOu2fViMUiGenKbcvxaXCHMzzHxNh2748krraOJRm8Ngd16VcUBTsOS9hEfDYvy
czi+gOlKQP6K7tDM8zyNbaTf3CUdYn1avGRNE5Ouaa18chlzZfmvIO9O6kR8uwGJRxRFBhiTjI5f
bd9ULVZkDdeQwLUi5dNWKXPe34uNmgCJs3+z4Tdf4Oujo5Pn9CMDivOYghYzrzlhvfNqU4BW7Qh3
e4lfDDK/pnHtLO3Kc64mrSg0yWuf8T+7sAoIHYoA27tL7rU5dWfM/M3L/0lokAY6hTEeyVigEhVR
JQtyfly9fqUKaql2UnynVGfR39QBrAZzMRmQaEDAtUzaDTQLzEek7r7cKKgW/rQYwCpqtXVR98Dj
hkYdipXqwMlx1sNJZyOXAQh3oAQP9Ff/1t+IKrFmc6zw3hBU7NuoGrDXPy4nlHaBsT8e0PjF6+VT
pbwUBlel1ZsZQHm/ONu9EzXGFlJdp8s7qLnFj2yhvwMZhHDBCNqNKXH2fZNXbvOKaJtVcbL9XuDI
w7wakScE2vymh4HazWtiGXZoSxdIHQJLBtbdotNCBmpL8BbccTGlQ/nDJEDL63LmfA4tG/Ph3UGI
QDuX5qBah8dVg4XO2u23Xk/ykbu6CRlP205Q2n8RXdBMvtCOsDlZwWBY2tIF40Q1vUbLxVaESgpN
Apu8dFUFcBp4dX/5S3GQFZ7aE+H4wUFZp+mq7qA+8274eAcOrHfuSuR54GK0FweriA8iZzTY1i+K
4BwYiTec7b42J0YnxHURrBkvSc9s6E6zJLnDfc4U/h0AvZNjOE0GDP+uqBHNYBaXE9syGT7k9eRy
GysjIEGgDon+jHth9+OvmdyAjjRZp8lnhrTRj3dKmrr0iV0nAvTIL8P+aPxycYQo4AsSseBBQg7i
hVNYrss5D9eXWWZQalAxwfLbEQx+IKevOySIb0gh12JTL/kYV1d7dsQOJJFLA8XENILTxFUWlcgw
g9mQ0f6JlMN0BWfQuOOpiCTGz9P8pUmbyUQ/idUZq2asL0xX1adEusr6t9j9XP7+98kiG6mTdcoh
okRJhmM9L8tfo0Tc9BN0dCrTx3Q1VNVfJqAlQedl42AX+NV5fsSVSeg3AtqNhD/hjfDB14M8U1Ye
dvlXJAxSvqB2nuX6jEdCh4AnFfJlUaqGTJ8SyJVDhq/pRTMEb8IT1modw5+mjjSpo7a55fJBzleM
UfJg+BbFEJdNT7GOfC1RCsicEAKaDHFaNL4hMoiiiCIAOVt/ZSi1krjAmYBJFJE+81uD1HH1xpnd
xzbj4jtet2vXZNxvNKHBLRMc3NtSJEEI9fG4cy4Umt58EpYeICiBYnENFEdVtw2qlO62DLGwGJcc
EST1/NjbhuXdE4EY5VOERvk4JbEPKahCc+itMwUZHJO918cQ2qSkIkm2djXSUnh6jv6uDPp6R2hi
h/3ccQjf0SR3HMCEL/E9j1RHdYQx2AcE5UmbPueMWkheYv2rNTDfXPs8EeQ+BliT8gFglKK/0BAW
WItBCBBu1Rh8tJR7/2e34fDMNdLkvM2WkbZkcNoA3DLT7tJaECrHWKeJdbyLgFbgkUbaAWhMM+kj
M+DCQYsmRBoFR6UGaDlPU0bmLx91cxxKF5cyOYSbelYBq8O7+YEmqeg6zkzkuq51FLbxBHzaFYFY
qH/Mmb9sJSBo+ifpTOMTgnCgTEwSFDd0fMV1jT7XmwAfgsKc2B0bPwzmWUGfw3JLGuvuAaUzhaZG
7QlFIkxyemnsvlrK0WnXvXeAZsY0VAG48jhC4OAi6XrzLFGh4F7IA2kssWAU6pm3Xju5j7TiSeYK
n7XP4lERbsdvqP/IYx3P2pHFF/+reXoeJLiSvIxvhlBXSNERTMgoIwW2wQi1wc1dYWSic031hRVy
O71jiny1wxhqzyANwGEKuujMQl2GS+6R7B9Btm6LxFw+2wM/UrszzXekLJ6uVD8EiqoZ5ynjHkgH
jL39AdTdysXoaTN6BmNYoOYC3Gqeu1Ff3oTecJCUAQxZ2V7A6MSKL+zeZP3EEUNaqNUNb26tkXLk
+lksos+ELmrRre4byBi9ZcfoRxYbvsceC6xmKVI+GSyKoYydFqnaNwh8H2ZeqtiR2vOaTqqaFeDa
qGCdAPaD2lvf8Y5WbMTclLJerrmPg1iAPjYLu/qW1U79ekVvTSLOOEDqUwd3YCMrBTK8C7iufodE
1lnTC5shXoyQ0hQvd1el//lOK9R7NED+whqUl6OT6eao3ga39PPxSMmc6CBVCRlUTuUN0TtrURkw
UjrogrO2VdCW0hb9BR73RCTQhW2nN/HoknQoonog4iWjLW41/8O966CRxosPNCD/OBEZcSrDZLaz
onKmtCnhcsUkbrdoQSARxCdDBASi4sN7cqL1sqOQmfDtf05bmsqrbDICEQTek+g2mmyUjxqOM8T3
BOH7ojKdQu46FijX/LNI06/P3gUK+L0ApYNf7Bzms0vKM8W/uX4/abeBaD58MYjT2KHiNUWfWUJT
Lg/0WSZckbFaRw/6IXsktLao6YdeWwt4YjtUhBg/DLgP8Yhi6OIoLmkQPzF+I4jx5R9GJHpJJI0E
8nGT+WaIAT9SsQTyXyc/K9Dp9EtdSCOBC26xp5x6mxn5fObWtDRGzP5Er5w2gvjr0IV+FrfrfTjb
vqJT3vq2LMAqc1xlIk8MG4tfCK3DO47xBMMVcVcdUoo1rl7Ue08HLCmnE2ZS8CeEZQ9wJhpiGQ8z
11CXKCkNkt1XglQ/fll/ADRtQD4o2r4ltRrCpwmNJthnSbsI7VLzFhP5uLp3IMHWHAHRhOobso1I
hegFYifzdoTuIeRGRGf5IHxGtTHZ6pZEbXsBevWXGJmf4WCpye+hQR4Kz0KfvJMybFZD4jI2tV4I
nrfzmRSRaRd7jxPXFqBILBbr1ZVcKbAlnrWYmcyRlXwa42ieIOcApxmzEG2j982jbuMj1caPZ69/
TPUMkxKfRnK9opkIyJhN6vevelM7ZhuwpbfP5o2ogGL6DrX96QO+7u7cj+OtjCrNAVZjh2wf5y/J
Xi0uwRP5LJVOsJyO72OybGcWRNmO+oHhmE8y1plZL7fP955Q1S3kResxZyHTSp7jH6R9yXvIjGVL
IUl3NetLzqbi/jkMKa/s9d2/maY3QYo84KNRUFfeWXxeSq7F7ezeyGgignN/YuN3mkqJgtyafEyN
AmeUI3N7cKAgVZUoC1jN5Mbzrhtpusvfk4qGmTtfEfAvYuR55vTSLIC7Ootp4fQF1DmUL4hsAVlN
0NbqcAM5BaJM5ZrMug283yhzVfgKpnimBDZSOcPKKsgrQzF2qZH7w7RFuqL5NPQDVwilz+kk0Wvo
/bDda4eOMBpoas7RBA4dTQKeBm/LP+ECw0Mm/xEcqGuzPFuGh4uduj6rocFtUvy5bK1nmjxVmV2k
8gVjxrhaK9NXO3LjvkjMcJFJjH1O3p7/R/tU5XnKwUpmD7xKU3OilCKIHFDc7W/XzQyq0auJ7WVZ
E7TXQO5pAkjWyIwxfDiux0xvBRncjno+codl4vldomMpNDW/ktlD6HFE3a44zRCG/ExobhwhcD3r
PEri7S3M/esy3SxYRoaD41YT15yirq6dloFkdZDu6gP5YaWhNdpvQlZncX+pwKLIB9ldLiZjSu0B
BploO+J/hDcfFkKGd63pJCeKb+jjomiw4v3ZD9ye5XLZrJyOXrzIx04RMMi2jwCZD8qH/2nyR+aB
JRlHa4VKTuNBdkMwblBR+8WR8x/g1JXJx9FojPQUFGwX0pRfXZCsTLRv7nMaQYj8E5vQhTiN8N1C
3MTg+nLakHKa1U75SIMDJjw6fxHTXvj67R94DexzeP7CUz1ZrFwhVqLYP3GxXWFS3V6J8qWw2LHB
8k4uRVohJaCxkSCZIfXVH9YphZgo/689IXLQ9pK2KVsklGKlfqqMZO/uSqyuy42eIMp+0gTRytqx
vYUc5rRhGBL0A5ITMLe95cbE7q3ELSsCMlCroW45uvHK3/MgrkZGRmsLboozSjsZ3kmxSdxDKTtW
2h89nrEgqsvvIXxCVE+0di4LJOxX94BGY4BNakLm4kk6pBIHeKKwptFMTnxWeZFnlsSTZzL9fiKt
l78pL7ZTMtAbNTfB/2FLQ1sb0VUH3fmWs2X+2QpgFKpg/i77rku2nUiDUwfUeJS4sf/HAaFqrC1B
U13oAFLLIxlj3onQOMDSdZe36uhhHchY9+VUj6F0ZWcg4KUWLNH9CVVg0do/rX+/GRpe4jF1QSOc
OHU/UCYc1GrYfQwg4qgQZOuvzdL9H8o8vhI7heQ3PQrrFfiQVry1Agi3cFCcHfzB1aYcz/uIvIpQ
99rs1O8pIeZI631Pe+V0EBXw+6qS/t6ZOprw1yHwzC8249eFrZBMmuUXHHua9F4SVEv0SWBC2Di/
qQLnmAWbSAoOI44RQ/NJIKZNYdNm2pq/BPXaVFUxuLiywdQq0+9UnHxIhifUM0iWoRhh7RyAEUVt
IhC2BWA4UUanguJfz60lODFQKNgczM9i1tbQyBGIK50tep5tLQyWLaL8/Is+t4I3/JXX9iUyN7SN
y1yxoLIvrwe9POmmLQaq1FRszpS/KuwRkz7lvE8F2jG6kEcbyAteNebh+XiRBkH6/kwSaH99DP+2
jY73fZUpEXzQpTXKyBbWokBuZZdv9OdyAop9bAc4povGa07PFsRf73OrrGfXV4dvWaM+f5nxsJVX
CWP75Oc9NXD2SV1Gn3BwaIpUmWdE2OBvjxceHfN5xGJ9Kpw27teCjxzS+COmi8Lch45GBLHa+DzB
cDNrD93GVlKXIdYoA56bBzjZFynbFBmxdgGBTRfyoYQMmHeIfR3cvq4azN2O3BLTXGGYlMIvsUiI
zbtSVk8RGpyf0X2ELguljf+ujEohrfS7lsJCoCEoQ7DlW8UfbH0uaTb8AHtDTGlt5hZAAFfABFo+
VISp+/7YDmVWw5CbRO0lbx/mHffCJmZJuGv6x91kDlFEMHd0hztWq9q81rlC7eqd6yQb7KQzJSZi
PV/8V0Y1vaz4EL8qGVFTN7bfiK2TaxhAhzAddHhqyyNfl4pewH6WYIKS4Bw4BofyszwLGILXak81
bFB6OIyxCN8yPFgHLpcWL7lAXmeWhe5izkXzkWVo9yMTp1NusUwUZhxfyPp9PmHAgaZrSWZHsVmm
ZVNcoWIzDW8gIUbCcPttjqqbVb/yu2M6lIASTWHZOJN0E0ZT+3foj/lYo+ThDODEqMWdMJqhHeQb
l62LAd/0TkeWgfu2aQ3NonZTzn+HFqsFsk5ica/5fBrCU81SXe35XG+GnLjTkvV/nkqCgH/KeoRS
hFYkKaiTcxVd+rA/O1OHiA3dXcNtVKLmp5cSRhDLMZ6n4EFs6XJ0Qx58niPHVufAuS+iiEd/2jyi
6bqtwqfsOb2ocVMr7tHwr1b2hAo9letIaM/uyAI9PEQFy3feYzClrN80grVuWhdXfxeuVI6ZzQ12
lsmrEQg9I0qBCdzOJWqu2leLAjBv+xmaOCk9pjPg1JFpHOYYi/BU9+9ZRoi5gzpnj0aa1Xn/nt5H
HXR3+7cTzgBiOQek6aamEk5rlV6PiUm9UZ0ODbvGV8DgyU79kgc/OHgwYrp9UzIO27/6mteLjhwP
4jNROGX7UV+gKKOYxg6+jW3vQmWLSW9/bUSSY1JSS/VJm5/l+XFOiU6HvDNXLYwYOKzF6wXt+XfE
c4wGvxtx0d8phImli9x72ArVcDx05h2/8eIIx4m/Zc/OlZDTRs53g8TEtn9+iiMqrXfbnPwJ4WJx
uMl6gB0TcqAv/6sXSmY/yQAypKevfPiobSDvtx84uY37PQswQXjNvYvpeb9vTyP/MvGd6+0bQhqd
ycmp0M1Idwmt3cCEXi3lATC4W+yJd1Y7hs9BrWIvV5Br2CwpjGLVsD4/HomTp7rkGXondW68YSVd
Jnjyx4Ef1icc0jGjUze080fXI/vmeYaS0G5tt8qLd1erHBm4+4JiA7dLQ2emHyQlXmDZLpC5LyST
nugbQISsduU3QrJsGPIC0XojtMChLor57wdK96FGTPJW7ksXk7MdLRe3d9KnIfy2z/qt21MSXIVY
BdXx1EGw2373rRaNyLRXT/sE3PHPo6g9ktqVyDKWha7n3crrJmikCouB2Gjt/yY1HCkbxVUhJKXf
naD81dEWubYVoEhbJ+Bp0LWl2K8gRuqUtFLxkxXFBOzKTOCbjOIxVp0OR013+jBBaQrUWqh8bW/i
iJyqFJs96Q8ROyTCopVcCshkknO+2aIe++QbSRkxqnbPPAMYmvmiyefnKh9nDBK12XqJGth+bSeU
2IAJBmQO246rgmdNTBOuHaPSYByA5lLJrz3x3xxylP89IkxXSzJjfBntFdx9t6TOYFftndvQ2CVr
cYIBcFqu5yNPHcWv0LCGzVeb5rl6ZoIAdHNtl6CFxsKAeR83TZQEYo8ohNmuHKn2WqErn/t+YirY
2hMiDy/sxK0z323wd7HoaUiOAi8FnNfM0wH2N8DhdeXExZH6lnRJABSOc20oSPEZjH6kCANbPFoG
UQlxzmxXN0VK8dWdMwM0SRMrrDFluu3305TY51YU7B681/Ia6btWeZ2pRT6pSV2YS9OTjTV63mvE
JuUVhyLtDtCQsvLZmA0sszvHthiwXj195JBrgC4ylymJj72PMhiPvVIgG0aqqX9bp8ycNSDSH2w7
IMykU+wXHJFWQkJeC21T7cRCOujqtunXT6iOirDHpR8NtNmubfwly4dzjD/B5wuQ/WP8KayKzvq7
mhkWQZB7REE23/E0W+OjNr0XvAWA6Xl0z+U7s7g/XpoHH0ynOcrULy7RAT+aB6fM22XBBqp1n+I1
ITEFTUlVa1YHrF8/Rdv700Q6nWG3HGbbWD5bamk3BPnEo1p0nkvLqy58e02ezkGx1ppXOFoIxU3G
rcGVn/oAmoOdf0QiL8Ju3bo086Ibp2OMYa6LKxNlZAeNuzjLg5XrL2z4wegCBTsc7szAwPz0aIPX
b4/Vpc6YW8zHG9V7fUvXdcWwm5d030ml2NQmOHwTA0x4tM2PPQieQqtgwfSapw4XbbbizHKtQR6B
MuuyLM+u90gDP5nakMV/CiYoOhyrU8HSvH5SYAAQQyESptow6/XC8RPimehHIEu0OKBCxd3b9SyZ
+hk/7wk1UrnYdN2EsHfVXHQhYksQj6mlxh4cMnOUN1n46ArwZ0qo6J8XoKZiBLbB1CCOoULgI/16
zmJpt/XrEEGtHKFJ8QCbO97PKHfWxUEgwdriBrNxpvTEuLKIpWq9N3yNtqHTGxD/d85WK+Tzy7j7
kP80hBtTLTuYDNCia/g/wRULAr9mmGOzEqw8Quqqh34T0Tomaef+qF0RBNMMhnlYtN3iJy7pCNGt
J+PDSoNuqKjFNBGrx8CIUd2yXxeKszUe7yvnLzK2I7nuHWqR8VgbO6n799AXp7DAlEZHP6Mhv4Qm
al8HbTwNAh3P5UEft/pGpL1zayQK1EIryGVgPadSfNE6dtoo2rq6ssY0qqws9LS7i/S8V3qkDoMQ
UgyqUp7mupcoF1cyEG/8GjnZoXx9ILEZ5S+bp7ZMcjiXWnzvbmajvOHknddC9/yWNBcC+tSN8gkx
ZN8nKk/dmk6ljcjr/Iqz36hkSkzBhgeNI/DGIEqxMcT865WKfdEIjA7Yb6R83/oUsEaf7pI3SqzY
li9o+OeTtrQoJl4/tdlindJWAPrrlH4h3eeroYJmk6tykuxV456+qscuvsoM4YYJR5f/gRPLbcCZ
YPEKXbO5xnQkrAQWlPep4DsnRGj0QibXZuQ11Ies95PkHdfDczVrOrs8syn0AazBvmPx5RQ1X8dg
TQAs428chvW8OocAwLh+507D7NsuTutt6y0oRFo9BUm3RTv89Jp7yCCHZeMGEwGznwElqGU69Te2
ZtZC8tSURrL813g36QBmWjD3vXqMup+/5Ui34VNYPo5RwR4dIzbYEHcQcumZMUXCxwrPRyTtxEf9
N16YRx9j1J+sLcIbci5MZwU98aJ6SDJdTEy3xv3ZiAfjJMANmGGWs1//o73XMYu5IoTZfeoev8sN
ZVV0ocuK4cCDnrZ/BZwYZk9uF3nWP7BHx60prcpRWXMjaCeEVltaCE2cYozUmr6kfgX6+osfazcz
c+jNdXI55nK7nMMt57uYysDeiQWQBX3IpXOhG241KbbLdv95mNzPIJywLYuuxkMkG0GTtKjxwyHQ
4TN0ihYmOJwcU8cPFOk6QAH6a8zb1hxzAh6wFznDJ1v3LbmJzLzFhC3cNyrtGL11g/PsceuLw3P5
wPHKNp0RxThAEITdkFZ8QE5/l8AM3wvIq40DnJjNJENUcgMVnvtXjTNu2yT42b9r7gRcTO5UJWem
6tWfST6NclPXwDf1EGRMKMu52ZrTrbaSe7LjFX/C2nSgpDlO2tXI6dgJ+k5vo3Hgo7ueCFM+EAJi
pEujosIr29Sygz8y9fNoBMqEDPp4jSGWXA1+KQbRIZOPhtsBNo9eX8zPWkR2/ieH4HpIA07qNvgs
oKyQB3cmslqX5FArYaRr24SRNpPZOafDaOb+hEy/PeOP1AiotE2C1I+1fSQt8SuUr/p0TYvPR7wU
IYJrIDH49d8RPIjMaHdH6xx/Inh3qkEKVzeEz1HoMMzuRPMdKIMNCgA4yjyotCgM5BJ28uPWcW7J
36G70580fn2/0eAhml6wZB+JdCtIRexC8+7RHDWrO9c4wtI9UPxxjXvbQ0nkFg2jtlNMESyIpBZG
85rI4uEMJXQPP9l6GlSaIiUFiJQnZR3iRgKAptlPwSm0KwE1yMB2h5x0KS5YAQKCb19fsVFTJEMF
aQK166rkjM1XugMoaAScDA3+z68EvjOibsmaiUkasgJ6xWfU3sEXX/ghjPfjfRVmJ3tMRBUoQpK4
NNn/1vkOyu2suIDUOchSZu/Mr5oHWQhjcgjG+uggxV8NMfU2lnnjEIwjWiNNql7VnO22wEisx2dX
K/8XVWBuFaIwOIRmt1W2NA/1r7rlDlXZ4jshPL/rvPQwcT53Mjsds5rDoYMUSY5N6frcrWtq+6pf
/7n/NIKhqKwarXvwTdfFZQmbAFf8SFjHxfYi6CnzTZIx0NOPDRv23YtD7V37r1WGZfY+e683hFR/
Wm/7aSU4Og8F0ZG6eYjyfcUIRzHi+Qq7QMSXeawtbJLWykzPy4N3EvdhbGKGOrcWT24WHlcU+095
9x+vLONtz6pOpTvn7M66sJ+fPWI4eO5CmPefo+KR26K3j7xlZSh8wWbpeAdMV6hHiu9SaO94SJ1t
9KZdyLYqL8V+7WiwBoUpeCL3lFFs5xWWqKng1FSuZgZ8uRPBzib2ljHaRIytRfoS6TK3mPLw1Inv
BkT4pRh23N3OPoW5t3a0IUxqoxO0FyebOxWWPhwLjhT8fIuxV4WzZv4d8Ma1SQkv2rShlS4GWeX2
k98qPzJpgLzbsqF7jYirfvCwUG4S9W7HH4ftARU+X5PrbqGKx934Q1V+JLaci+BSLVkbaOBcTTZs
fcWVuBkSG7bwIYRo5l0bm3pGa+gJTcP1BXIaEvvYxytYYQnJM3dSoosjy8LkGFA3HLKY/zFbF7Ro
k99qNuBL8PQ5AqVSaA83glG10lMvP5tgCOHEwxvdhDFawL6lVHuoR3csNPdSHbmtim42ccVpd0XN
Tyqk0bs/v68f05wLKt3mT00O3DWMRTq1nzDTNqIhTeYPfAER97qxNiCoubVB1xcP8OpE4dAVFk2a
Ukm3LozN0BtlRmerCOzAD+xFO3EzFpvkzcljxDDkcgigpT0h2dtSh7feWa4zGVwYUo6vyIozmA18
hA73wtgI5c4mMnM1sO4+tQwaAGeJjoA9+lZVv350xmufDQ3JYbTmDSpLmTDNGVr7Z4bZlkAbPom7
w5V9JVMu5Bgyp0gf/VAP6vpoL5U8h0v45OYyczwtZafhhoMbuwYVXGnPk7/Z0VFYOLCM8eJuhRiT
VxnbHpTkGjxWtW+73qB759xzIPATuWGDYPt0u59R9TAc8NF65k6Fb3XAsTHsgbdLbtu07IvUwlu4
sdWgFkLLsxULjijGVBpbdT2gDW7GwvS428OUAZZ1/UINCJWe2LG0bOEAQzZaCf0K8j5ZoBlSvDP/
mWZlYD1lxY/d42i7kkeRadL2oPUiK3mw/59H4RZlRKLxRiXf8MGBDDLio87QcnfLn2oPs8t22DEN
Z4VhlnOglF+pCxaxsgzLCwrhNUAApBudJorYx2lp+yFGfSYzo588CcjxqsRMsNw1iEWPJudweVBN
IZ60vKzHKJjWMOIZlNb7DcZwWgIXi7X8B4ethblrhkl38zocOz15fQVCuJT4I1S7zCnaj+CTVxKx
5GoLYbTTUbD3E5PtgBvOvB9mU4z03nYjsojEhPbG+bPuloS3elhkaoh/ybTdQ9KGnHAqglo+87hF
16KHD9ifw8/H6T7f9NBgPMgS1Dkt5Pi4mjfUnQPcqIwlsuALh2M3l7k84BpxPgxJCHoCxSzE1yet
QjFYg1nTL0cczc/aiXkAtLslwvoj6llwPHbMJEUp/jk5pOXlO5zxAwcdb6Ua6/C6tE19reocQIqL
ULYuNwfOuus02ImwvUhvagvpuKWvM6xtH5MUZPUODwJ+N/739rgF97Hw4tKoF/uADGx9SiGo79TN
IHqjz+kID5+FIinlse9/rFMJoZj0hh7R3AT0palukzdRNbG+cyTmdQtzOEVdIGGA3qca+oFqg7UD
LLjCDk+8YVX6+bxSCXms9+bJwwqTuxdEosQpZo4GTlNMI4gyGdyyScsNKHxRglRxQ4T1C8ixnTt2
xBO9J5eYs6Vz83kcZ0WkzIVNqMn7bVECnet/YMr6hjjq2Mr2q2qGegF27hD+NZ/Kgl9JIPHjjDl6
tHw03VualtwgHc0Q+CvIFbGpzD0vcox/Cp1ulL6DbnNoZulrlhjr0A9AH6UQnl98Yg9mgOQuDB4t
bI9n2sfQYl5kR1HqjgMTb+FlR5nY3M3OhGDVDZ5lmbWyIa/ndy1+5xL0Yr8vJ2Ek2HllEXjK4cJF
1Xb2c6WuwuSI95PPCc7baTtDDfvzP8oGLSIZkASJkCQ1k4JtG+Z5PfdbaRog4aIrAh2vPTMfXXxq
5UxGjgjPOzNpyiodqyt89cRdU2198pakwzGYG0uckv/FuPfW4zH8QlRlfavp12H+dNtv8IzjuVm0
3FQCDBxcrp3pBAxYlgzA22oxiD33qeNCBFnV8t/keAzXVLcg/O/2dpFkrOBNKYqf1XtcNWoVizDY
Iy5r/xnhXjORSMlWyU93SN/LERkmQCVL/jTBglaF1keidPBFSFRrRfQUhxcoQr5kADQAkmdg6iXV
f+DeUyoWXkDa3bBwTrnys9XeLaChAn6BUX/9BD36GFJ9OVEK8VVT8QM7qK8ZrHbHfpwFQzRetuNA
77+yg2Rrn3YF7C9tkRsTCwfYwGrx8KBnz3TS+de/kXC8cG5dugx2xR/B1AlUyHh67deY8C4FBO2C
JJRoGAqG/ZCEr7pZeOAdqyPq0V9XOOZHjodB80xV5jQiF56cha0+vjvHhxyQcY6y9Q7Z22BKB3+F
pMcEK3Ja2y35bFHqKX1mU/hW8PmbIt57ycSqEJj7RKQ3PPZ6wKQvN+fZD9jgK9AaD5gYcqMRRhuX
6YugeL23jbboBuDezuKgQEk25RYYR0wloctSgH7wuTs06+b/qfhy+VrdWg8p5EWgq/LGvgteV3sh
kU1XbP/LuhUF5qVsdb6Gc04Qj8r6GBuMRBX1mWwQtfK3d9+xk6Rzv2OCHjv7dWT7GrZ9J0Qokbhw
BJ/NhSULI6SXmR8xdfaN7DxuHg9nBwtYCL4UWozFKlIA3kcDn6aCT27Te7PqxesUUIUDmxQNWg8G
6mXjo09yvr29Eb453B1FllXrse70TgmFX6k3NNb5SYTGMv8WCev2F59tRjjmdSW8eroM4clrUXpW
d7C1+2aOlTQ8+P5OVPG62OKSqIqBXlPEZHHByIXbh7plLi8ltmoZ7ylX4K/P5GhJ5S1AfHTxa1Ly
cbdgh1zgWdpwI6NGZFqFKGonknYIB52sgZZzV/5alvoZ79ATNVKmv61o1HlYI2AE4XsWYDmreC37
cVMoWwC5hj/euphh7P5Dd1+vospIepdJIzok0KKJAiGB+tuQGLRCvmWu9im5gCpO6VzU10M5W5+L
BC5YXIOkje07CyVLuA4npybla6P9Ju0hgZJU+Jldwnt9AzX8LC6GTw/t6WKrA2eC5zgei47uw5SW
RRvEDa8MPpQVVaJeCjkkN8z9GuiIKheMK2gd/SAkHvw0MIXcrSY0kOpeSweAoMn76iBM8l5NJ5jx
v5UTH0lpFHngd8ZRBguPW7oXWzZ75Jq+ke9uzkuyyS38i6GReZFtBBaDvec9jTz+kYKiH3g8R9HW
Ib7ztnuiDmE41tOqgBNMTx6YqsWhsew9Ab7Gv0tTcCb8mn2MaPbdBHVRO7dFRZPccMtrXwJ0AnCL
RoN9dD/+m5RBmdhnEPiH8T71fXC14inWVgs2cIOhfko+wDiH9daSjY/vTYYMZUPooaTnFYBjcVSn
b7/zcllA6V7kWeEO+oxSTYH+twTsoZJPOVb+GkLhugLJYurp9gyLw96txbgoBcUhVgLKWqVsZT3c
XI2DSOE8D58hm5lBsRK41CJmrYHSYEdYxekaQFKHSczZfR4MZMV28+kfKMOav7RwI+2gtesdCAcY
A+14yWVXFdjB1GUo/uHELI9Q0joZqhscUDKMbQnFO0ApvZiuRIqN0o+6hu5MiSX1zvt1UyOkKFn3
/Q2PbYBR5MSALnKJShmQwzdsTawTtYWI3V/Rv7bAp2wXiZ5bojBLb8PB490mZrozragY2xnVB8J2
PjMKIUKDAP9ldK7EhLq1bdJqxSP0d6QE7u02H1++lPHo9FU35/JPLTkAk0wOj7vp8RurbvC7gVu/
n0d88DdeerH62dYzXttGGtYxXxZROFnK8HgxtLRT0EHlBzQWo6airAb0PaTFIRWAZQ6PjHPCJtpZ
5rIy3mcy6X4sXoHhwDu0AVxoSq3oqI6dlmJVSRFih+NJrfrFPU+bBlx+qPHIeLZ4JmMF4MwxkSFK
VqrLejPKYbv8Qm3WKQy23cKzn6AT+WhVtMrj9AsuKdbKKI35LU1jyBkpdK5zqo1bZE3gf6jfTbtO
96RjsewTyi7uz3C30WjG+4kfH3Z+dWev896aJ2123WyRQhYZpwUROEqBBF71bVQ+dsG5g0wS6iiA
PDiZj3O6HxDNUYajl5MOWbDLbs5IJ+H0Ng032nCugKYEAWVLDJlyHyOJuN49Woxqx054ZnFmgFrY
kZCDkd6RogJKxsbX/XhiU3S9Xr2u/JtW2p53uV3yGRWryP2NxKKdOONz/vAsv+NswEEFBTXgBuEs
mgrfSChNtpZGYmS83hCx5BRXS5sqDxXm5NZlDPpkO62Vg30C2r8nXDTCSWcsmoEbddMQtyDR9EZ2
tJYjUA1yJgHcnz3lBYLWofc6+G6e5hGFP9nuO6ECVXrL5XbUumg1p95y7N2ZcYQHO8mPhXP9/zpc
DmeLCwsW4nfbhuQYhSh7tMEwygHJ9Azf/U4lqRGqiJ8Ipa1Dbh+kD5UgT9caPi6tCYIhhdILMiTN
haUyM+zBo8SyXj4um4crBSZz8uMrg2PdGCxCTskuxkMDLkXp1vcPqz2ge86mWLXwMl2hVA53Xczp
fhv/LWP8hkAmwUKTt7CWU4XcZd4VunzhaSxS9sN0UvEFnjp4fjSIx35JpR0UVoHPXQEKBY96g91b
539Cn1IAYFGM5w5LLJpx1c5HggP64Sjx61CCxIIqsO4wx1WtcAMnrtHnnnJsQ7XWw6GQHbX5X/Tp
0DpP0PSqsTAZzyD+ORkllLfrRD2BOcMVZ+P24CJNSxc19PlJWhtpK1MngvSzDLTdZorFHNFKFsG8
BLVPN15sgbk46JB3mruB3R6iHvFBmhuXhPzRZwAz3LVrMycabLUHn0ymaUsozB7qLW5DTIUAJG4/
lOF7SPqhaLi0gHVYyqh1gZ/Tj8JRDR/SiJKkY/SARxemEj9L3+iiK4UkpNTYkgGoIctO77VlSGBy
LrK7gh+EvYp+H7Zy20+A0elIRZyEL9CLja2m8sslEkz+uKchjxCuMwdZDFFmllh0zhn1EoxpADI8
5j+pxCk9d9/Smd8BU32J+lMZzgTlZRDLIeTQWd+gWNsBa9rvxYu1yALg6aFqovqxcBgjI0PPMIUL
n9ybiYKl5kMKHr2cdGYGa+CBxFSJCfjUflzvSZQhVX6DtX1knG4lASb+bXLCW9iAcDuVvgLtw0cM
tsWdjfLNZUFVvS+yRPs7N+BQA/BjOSdIqo4WLKLyUpIjYubZHi7Q88NqpJEfCFc3XYhq/2CqcXvb
/NPeqFNE2CT0q4jZwXqUl1MUHJDVXA40AOqenjRKVgnzqy+z98aKj1kiY1k42xNET4cyVYNCC9kE
ssKnBeBhiaVfYYvl+xD+hfzI1nFn+iHO4Auf2U/a09RMXHz0EUKlrpFNMIpJ0cweq0Pds7TV2w2Z
12bzO6/fK09L3BaLsCvPESb83hb7SkAOf0+QOeuZqeqcALTpADKqkGIH4necpZoGQJ9TBRVVPwUA
0Nojj8M2O4SkH0zUsPGp8OQCSuCBEwasZTFBGZguedY1uhrKGh+QUooI3uTviU1msHH6Hkg1iFPF
1QKDXs7BLH/WsLWDH1hA3XeWiqtd8wJNmpYdThrry5Cl1uiVudb/fke/pqqNz+bI2fzKSwOLePAf
TNO4kjcgfbGVe0zM0ZgnvIbTU4XlXxLNOzaYdOewsoJXlKhkn7SWx6ljNGA7ApYtAiqalrkZDK/z
FY7jk9H6v/GdydaUEe6UafxQhobGjjWEeaqRe7RKbEY+aczdQpeSQlPZ/BR5EUkoFgMo5zpZC6y9
6kbf3ES21UgDTrtKM1ncozE3+KlE9Sn7oV7eV/l2Qe7fuEIpEmNbsQXeR66RWQDpO+iR47abp7ly
yMEu4siq86usZ/WWwHiGs93C1nOY8zTBuwPJoU+jRbezyD7VeThG9t4j0zuyh8ELrJ48mWH3giOi
g862li9W4A0KWu0nBH9jpy7AhsVdgA+IPhV7J7Iq3ENRpXINuat8G1W4Cj4Fr+gCl2KT9jqUwr7p
z/t7WYPQoVrNiwUVpYOB4asn66KL0HZmTwGd7lAbmL/FlWsa5Q4ph+886G090xbCbTp7eQKtAytD
7+Foo5t6T7eoXJFlUhsIAeexUB+9lHsUHK2gC9MBrrzV2Qd6SKXZ8s66j7Z6sum2PXc3COSmZn/X
10PNw9Vg4k5gBf7G7pP2X4DQDhwoOPgpfhwm9+QLVv4wKfnaTzxl9yT/M3aQg96EDffmE/5G1+dM
PBXg9ajwdq2lYcdqfg9GwHUwkTPTudPp72FjKvIq67QLXoudt8gnpMTr+Gcj6CP1r4k4KfEWQ26B
i5vNwL5SxEflqfGw6CNGyOUvp17k3ki+UaSDeLYseHMo4q63lum1x9gP6p9gH96NUXtoBLyLgQwX
Y56YOJyHwYPOTulleamOlS2/UhpoX8E/18Lm5UzK/6Q/9ZCCQ056pdHlfIm08xOB+Bw+WD1VR/WT
YAxpWOlzxfNI/hsnY3V6tVcGBk8dZjhOVwKtjb3czDHdaxo/oMnP0Kz33huo1F9PRmM18KApMlD8
VtgHTS1ac0ATWEGo3YOGUU/73+U7i1RI+WGVWhIGzNr+a2jXG0ep4CEBT1Jmp9IJ1lx7j8WOIYEe
Zi/b8RAudhOlK6ZIgaJ43Ny+lh1qddyJU22MqE7exxh1+DY9CPdqyje1fLYuZu8IdjOk1c3zBOeF
Bgl4wOxiMZo3DjiiBP8wLP5m9MBkwF4zQMr+oAOOwkL2rFQ92nOilKWSfMiVI6hkZYkUc58kpYhC
uj674WZZZvvsBL46nojUrekAdgJo8Y/b0aUmUbm3xjSrY/fTFKtMCnJLRZRWKoih0rH6yjf5QTAf
e8iHXNK2bxQInm35SSzaivazKsZGXFJIHoasqfRQmvzIC+VG4xqqf085it8344QLCk8whC8EA3Ph
/wFNh6hRSMPSTmb5Cxurda7l7GVq85jLHWlq837F6id9/VvTJlEU3Vt0G5/dhvpFI8F3B+zr4GyK
HqL4c/W1AEA0Hsn/PemJKZzIHALcLAgyAQFF8WLK7VuwxMVJpE6tcl/Tx/TZOzsFIvrSrBSQcKk1
BFgkQkAbj//vKKsanbzjHifgzUGlTK5ELxEJfakhFP3wV1Zus5UFRFqlx7Sl27cFkhx4DxXEL6y3
Z+zZYiWrFGigrZvtBO4nJ2z8H9+JRG+k4LoS35lVrdH3WqGKkr+NyMZ684b/FlQ0p3HIgMxR1Zzc
5vWvJawJ9W6Dw/dRl9E79OoVU0sWM4qaBJYF7+2gXDVIINhVtOh9KHiUl28/CTsvpAMcwEHjmkYM
uQ740mdZ3qo8ZskkMFSrfXwKb8HXSf/hYZIDrCWvtQ9YclBaPSPZ8s3AC+6v/gDGQh06mboJU6Rh
Qt/XYIv1wp8Ef+GYkNG1E3RT0T7pCL8yXbzIed1bJ7Ey2eQ/Z/pCTdD2BURVUJYKAkEskhwZ7BFx
9kaiD11GpLRwCvfeYTKNwLT1/wZXfF2jOzzZyFiz//hqC9RUjzTt5dN0h73icUo4hJjwxzXexSfA
lfR2hNwxA3XDBa87RW7sj9YUe8SjTh9O36YZyKtg/VwaRt+AeNd5rjwytcNC8GPy6pDYtR8PRpgI
JHyDspCaAbMK3HaLwwHKWxVd7GY2zclN30rIpvqHM/aIjE2QCaQ7PxZz7YgTMsHS4pOJgp8UjfwU
y+/iG4NDinBHy136lSXc5DpAq33dR2ULY7n+B4saV3ffzRlHZx/kbAp0idWow7sZ7Yc2qgVSDiEN
OgrDvCovHKkpj3b6/zaA/L5A+1C+pt4TOLuPMFXhlVNXuHaQYt3bme+tEUsh8oWsVFZ4gwlMjzrV
pT3KA0GpygBQmJJK4Itu5NmfX/XgoFXZJwmD3oPQxxAnC6ON/aa6M1tgLvp8Lj2P/bkm0w5sh16/
41f5C+0w3BQFwMWE6DO/xLSaDRibfn7CiFqORArXw7EmqqyhMSA8j5TwKbYN8JiCWEeihV8rGl6j
0tG9VZtiKxpUmTDH1y6wKFK7GbfOPync7zd3r4saqHYGC+KNmZJnixpDXxYV4veOPHpUM6MDX5zW
Cpt8SMxPlC6VpuNZZ6WXEiaHG5vBANPnSRHI3jsuJUwC9YgM7WLr+I7KQ45i+xlyGsiynqTWzvM6
/PLnVfJSx5oGYgNWxbkNAuTQKvn+6jjAI89I62AFwGzQ1CvkFMIF867z62MN4pIKICV0cLQ0Jg0W
CHm0BDWwDK3fFwOBzbyTMG88t+Lnl7CH9UsQQHbqbtJNNgQ2U2dU5P17zPD72eZBGRQEXUb2jjRi
EiMKncVqOvjYibEZxGS9SIgOUIbptOodhgJC1ge6tOtSZ0N223OkJ4MvGCwrFAmmek1tL/4OGASM
58JmhIe9Big4hDLwhg7J31XjJfRRNG6cW/MnzAQ/udPXNTem5u3XV/9d03pS5tIo4zbLNbUv8Ups
4vK98BxeTqJdBeyqjVUOE7pXY9jd90CzX0tL60wf1ZGGuoQ4EHkkqlelhHMkdjKn4XmhwgtHo/p7
uMyh3Ss4UOxh1bE2sJhvutqniJpOq/838fzZTF2vfyCL7yKTAKBQQZZv10JzXFc/2aASPsYandAU
7qZXwz7xM8JFjGsN7oVphpr19cySRUs6gYu1fo6jYO/BQbFBXAr6talxAynqLU0UUNcm945Ht7x4
cnORC/WJ8V154t2OnRz5f+9UEDrGpQ7S0DAUjD6YIjDdOAdqqhTsDY+UPKUk4FLNw1dIVQkn6BFW
Y1N8O9NQiS/pn+rQbYkT5QCzjeM6jkxfqBOrLqX3F6rKO/ACio6ZJiQqolS+fbUhhuXWnLn4hvKO
Q4n3yejvtqHl5/H9Zm2GT7UPePokJ99Q8FLEnz80oqZ82YM66X5oIDySq2ozDKoQiJlhITcqezw/
0Z/3s4YyBe9Zj8tp5tLmPg/8EOha+Stzi6ik+Keo9tT1GP+P+pN11SRXGg0PsGPME3MIlf3iwvj1
AApkqy38k4FLDKjqsQSc+NPwE5GX+9Ksn9LJ1bjatN7h5ZC1kRTqkfIWzjjjo3PpfMgDcJwcqhGG
DZm9msdBxAo+xsqMhdmYwfLuTHTbG1yhCNZPcsVuTj5AY3+VcvG8PlBuAsITjhGHrnDJTnPFxbho
nM7AKRsCEi4FexuNOCbXY2WX/66ZVooqSQ1tG5Rga6A4kBUapULUSUM4jQTIg/krrjlnT2lqmHMj
WVGWZeOKvXBxDgoKujnL1b+5u4175SNPqQfrb06BDomFpd5/kpUNTgACQoKdtWFboPynPkFUDNco
KLj2oCNMYDID2vCw2Ab6/NjSaMOGzjRe8w7R6L8sATV7zC4lgv9PhGfndWDu5Uy76tPL4JJ6XHya
UTcCxj8fDltnftbTMu+/adHtTLvemBJXFDKrbFK6+VNjyYkdkI7c1wH5m8dd4elgKkYOXovp8WQw
GngOC1m24tCRtAizF0EIViR9E8JjmiNaNJ1PiM2PXnOEzHnEx1hsZJeKFIzznpeUZjPMXM07DTvL
zqj4vAM42RduP88L3Eu3iK+qC8yuobzQh7oveyCtQ3FWgU4FKnir83d/hlfWaLWQsyNYqPyGjWr2
5uXS0QZd38Xt+PHHRZzsIhr+4zW8HBN5rZE6pF7Hc8aRxsryYnfOzvc3OKmhD1tV/i3Df96s46D4
UCBsf09Soln3YLxpUrTGMUcKmGBebp291cy+LCBRcTt8Kyal8ObeQTmejFtnj0GCrZ03ipqWoM6x
r68ZxcMxYg5YgFmzwX1XnWPxB0FLPXbk6bMi7rhlHBx++EHeVYvcagUdqDnBUFPk1gcvQs0db/p0
8jITWu2d+IrESkh78kcERw7MJNMNr1iyCP8w5H4RpoaUVVdfBYwyjZL+DRnwfudr5Ik5ohlfa7Zt
3ivKTYmxkFl6ci1HQGI58slSIbs/MBGwKkL+JqeAw7TKvmmr1G/mNyzjHcDSF+IRJJMaZsfHVuEt
oxWX+NioOJzB2x/LRnHr1vBoY0TV+6C3Zr1jpxak7sIC154GbXG/oLSN4FsVV3GfsOg8Hi3VU1UG
1A95bqeyRrmoVURbPSzM6hie99E0bKCIq1gPz66lP9s7ijjz71DU7eW03o/4Duqb31CsIxqvcO5t
mGM7L1g7r2uzoiwlS2lA9+0mCCLVtfu+xd5BobUdZ5WUgEHCeCd5dWd3jE1ZN12cp5bvbZFZceZ3
kb0uqS4QufQhF99vI8Jm9CBpgVGZwxgw8vIpfFh7GVb/6BoOa4gaoTYCeEIhnW/zN2M20GwrkMDe
37HnbnPq8lGDDBrRF8iAzhFHmN+R7T2GCnGKSUUdiMvr/wVhZwFTUkR7DewfZ5p5I1zZNwYMXmSW
G3wiBK4vKhzuK+lN83RfyXQwnJg0AtaN+Y3UMqI4i03wvXhyDPM54LuLOOhnUKnZ2VNn+olyBIfX
0ivW/rrEqy6mGnI6sj9DjUho/r8VtJQkrSWreRAYAtgiNQJ5H7k+vbi3O+aDjoezsBHW4dNB23CQ
1218ww1EGCtFHhenNVhIYHf8mD/9//6WOKSiGb0NBEwMXxZ8QCyB8J1iw1ox7x3gzIXlZWmykuJW
tS8BAR7l6zp76YuamKrMwCmdOCWwgcUOKou2BPQZ+hWAwhWoN3bbF4A/cvjopvkE2mLDqXcBLP3F
bz7BVABD0kPZTEtUT8D+7MdGIqGk5RkvR27iziLYjqyhNv92KaZjQE2kTOQ5ql5Sb+uqx6bjSLrG
2po/8PP3qgRGrjBAOkw9FTR//pflAIXsGurDZ685679Pa7NGy0Y9MTDwENaYNMWX5+m/M8Z7IRYM
fH/h0QPrMpfiNJwl4PwEkwh/zrsUNuNpepdaIX5YwBuu4dWEESUHv5qcU077oLbdYbyWgEgiAuBz
TnKuf5Bk6RwsY39NRS7MYYKnA7wopdVBoh9nzuNDKeS0Qv3XLILuAg8naV5dcyFVS3xoHPnUReik
0iQp3dUmOG1x81zeK9pPvuoJ1D3uwQdPK6TwOw1WcfRgCSWBgT0QQWwR9+270t0g3wHtLDz+Ui3J
taT7dsrzn3CVyLub4EXqgMmDL9BaLEBE2ygJvrF3dBwy+hURMRnoiUyDqp51Amv/oTYx+dphUNOK
7IQU0IcdaNOf0FLjOQgq85/jL8npyD67SPB0XVswjqhb7YcSY6Ofe+9lDPTQkUZdY64OJuZYHGBX
c0xy5GtAk4zD82nJ6bAi58kN37rUen0RTO37fjOI1AZHKc8FHTpOL6EHdPMVHdZYVSio13I887/I
o2u/JKMHPq+eGHSTo/XYF4jyGw6ezADoJ5Ga4/744ONj5UuM7bBE6mJljjsBWzum+wtlnJzvbnAk
PcPtbq6/pk8pRVysVFAGVX//OU/1s70JRfrGoVBhTw7D/QfK6Wk9InFwxf1oBtl0FjmSzqyHNg9T
0fVh5jtPPvsE6QxH5R4gjlZIxb6xSe0b1ouVOiVPQ+Ztwcupgl8zg87YlzuOXx9b6fWhXzgGET5L
bC6ez9+RUXF0IHzhYWmdGt01ALjByglBtLYHmhhFhekkGUmFTBKmsm2sf3WNXqOMS/S6OZkJHOTo
OZId760z7fKB5MwRa9M0DBnG3A+gPCi0pd8MANjv9iMMd5eFtLKvdNm0NgIv0ZlL1ml+VNF/lia0
J92F4jXelJ1YJNyjjfb9oq0VqTa+eg0OEX0+y/aYj9ymVVgt+xgrwyzJv2an5CeHkJbfRNVCp/ip
fAXjVjRpBg/ynPyimj2oZJFay2DD6VDZhRSw+8ue6eVvchNAlP8sr+U9A093j2hgM+vBJ9QJVi7o
JQIfJg6L9cDt7Kz3JI5LgzxWYRn9Rf2NARLR9bZnO8W4ZqaKfyWX9wFBwqwN0QKJ5RAD1tKK1wQ4
iFY/Ati3huxsBtJGCh1inOyHutjOAJ2MBQrYm5d/FEEiwaPtWTj5cEFIw2DWU75/6Vnz5mBtOaMO
pJN8tz1Fjc3pVE0YIZ4LcCQhH302arVv3wPlcbnxR7mr3B+e4ig5qlaG+i0LdepCT6nh1cA4+s3T
SVGBFcJNaIImFSkiad6b/M2YFM/o5DL29uNMr07haTDZl0SO0cMtdemU8x2xGWp9IJ3RQBR6OH38
20vSNq6RAITj4d4BW3/YUv42vcsfuianQt40i5a3GCBy8VBYxPhNIHWlb3Tc3OKVcwtf5tmB0OZ3
iWK2xlqpN4As2CDovJvBNkNYHujK2+IOJ5HceizCbYE7ki9PFbWSeM0+DIdZgsKVTa4pDg4Fb+Fn
ohmBiOLl5pYMvzrMJ/XhEq81WWKoOo/T+APjeKQrOxHFSBK37w9Pr2L3mWP6bwWk5M8gqxh6WuGa
+NaFofPT8DSl9pxu1CfZ6e0cun0pu+TmJG7NiZFEKq7JW+HF7IA/nnSAEqWVcmFqSW5yZ2es8kRm
PrMUF6iy9B3c3Tjzx4S31YgF3YqjgHJkpC/pnywAuMb5E4WG1KeQ3dMVzZ50ArSVXzZWjJiRp8bG
k2MhY8irkJBBryMCSYhAykv3TYHB4btFVnqQ5V993p4cPn500WNT2YbeFWuD9+lnZrucOqR2mKJz
33ps5UirVmmW3aVfdYXMx55qae3hc+l3JuoRUzZIzKbK8ZAMkHSTXVzzsg083j+iDfLDuXa4Ttlx
YbawTIEw7MbLf0Ig+v34lfax5kiCyuHoS22lYp1meVS/haERq3Fes9FNtZYKxpXRyKSnNV/SeDHv
xNeNARfVzez4Zir6Z2xXXzSq/T2hFgS1I7awQL9gKvGZQyG40IREwZKjddv2QBn8LpfF9i6+ufws
+ADXBy/f9ymsohIfTtGdn6mFvJ1UST1t7emMB8ykOH481Z/FnnjG53pPK7iQRUoD3oYjaWZwHH50
nEFv6Hm7qx4MrlIL/7M6tuMAY6z5bXlYX1M5YEhT6XfukTYjmpDde3wmceXRWM5YpxdoP7l1Nhvo
8JIyj8r+w8FvxeDoZwcRS24JRKinqqic20EF9STQqJyop5FxUZWfqlY+3jVvKDJIaGmJG0vsdkTR
Y0gEwpAo1ySp0Lb0/uEvznZbxrfUrB1wDA3mVlkqoaw51JBcdN2lzyWza3M7moGq88HbIkZdBuKv
zQe3bWvKGNgFXG4Leh84NRg5aR9o5nOdOV++3tsVXx/+k9opIQoe0HD+NhFUX1fFb9d0L9T7PVUi
exXeKq0Pe7vaXTIQGA6yfAp4igQTNjPL7upavZUn77/lrIVth8BpBq2vhwzOy7qRp/LqRVjpWAr5
Vlaq1khSL2jWHv8V3UbNfKmmK6MU39GaCJSyz3kUf73Slenpe2mrI457QEoTX0oiJsVz8PNa7PBV
aGfRN0nhvYZBYJ7t4OlVoykr+LG9+OJZgWhdEgohQ3hOIBcEewkIDmDKj696AnEIfi/8iAkkA0Vz
Efpv3nKZ5Nv288ZcMhwcjiw9r1ekWGFv17lbk2y9JhFJ8bdmAFHlcvyVBnOYab8sTIcSrfz31Vhp
+sQzhCgmFN2LVeZRc8DccAD3Rqdoe+qck5VyFvqLFxhjrV1Cm8ewV17F1ZfWqYHqe88UH0YPi7ZG
AfwiCxplz208z0pcpQavAftvgmqMk7eYp1Tqq7+PI9/cD+WMLIFF91R2R2p5bTosqoVpbXTltOnt
Xue69B9C2lLTmFQeJJFSIY301ovUVlVXysb9mJipgeuUGT2Z6yqRAqodDhfF7RFa/msRrB/Nadne
w3nXsSwbHoNBijL/ohBci7As6p2fljzf4l4qGSrIgmWFzEv9uohBXVS+3EHqFAVA1T6QnLLjawwo
JfunJWmz+p/1kHcU3CORJio1JO8Gyaje0zdey/8x6l0petGmm4bmWqzTMoWKe8zq+YhODTY54Dwk
9T1rjBq3aqS6hctpAZ3i7WO3d9ueeV7izB2203qUDp+3UXekOpz9hxlQ0N2/PTbKYvYmAhMuSRdz
iph+XlZaoVOjWpDUKk+Aba70J7ZXZl5MMjbj17CJ762zMhR1rTcljTa3Ti2u08zseKiB7A0kg9Ib
+wenQgflkqBAT+36oMP2bc4a1pztn1yU3QjctvJNbplHTqrVgQmOAmvZ/wbEdD5NBGFRKVk7J34R
ryEZtZngx4+HzOx5Qyd/UqxPYQVizyLh8gOsWTkqO30gLnrcRkDsxhXEYooN6twRV/nMHHe6SfE/
zYZDVu6SfJCnwc/6FZ9YvjEQb3LgkGd5i+9YlhcrWUqa+DCFPpW0NrKjVYNr2Esv/OAIdakJXZAK
rYdMYI59kWOD0DzaJSeG+IB/HTj4eJAHNMFfpMXL4MM+shptS7IS6iV8oL563mZTk0Aw28kC+wvb
/3baONMKfx5MKJmL3cVrMPcgP40VvdG0XpJlRp9AY3jfoEIGTdPbzN5IEEtqnoiLdokYVfm55dv7
8eUbsoE+KvliH/PeDYgcjpGz2k9IKFPbTcIoN19jmOTT9hnoqkvW2eqZIye5UPzvO2TED0wtjJAV
qtabgJGjchTvo5dOfblQxoXpeL3ZfoeBSGPyMYDmAfhDFHYQaadyw/75vKh1baubHm7rKpWE04RL
GCKULkyjBmwmLPEm72XH8bwhlN/0NkvWpjrfn2PQ8Bk27MhsKdSRLTl7BvsctHkWHx3JIQ0S+tFo
en+pkE29SAwrXSHKQjePrE+LvvoIf1Fizx6bKvdXEHh6doEn3kxyD3u6UAfny1Q3NXvHmNUKDPy0
CRWlJGJMeVG2+ZheJ9PVuh8+XyPohuFHwcBW3qoJtFVKVqVodzg0LggBObP1Ll5k/aUSuGc5M5a4
iGdpv5MYZR7W9We8EFlWxUKJ0nx1+mFJ2jbJGWBXJmvz5YMVvEsdlqkWWoThNLBlmtZjoSlcPfZy
ri1REzaqtzOZIue3DnFn6ZKuoHZcGSD+SvVhUtjQvoVsSifwKy3vE4s5a8RYZ0Hcbe+p0fEJ+x5Z
7cMy3yOgmQVlK0eXPpurs5ETzHBRhCoAh5qjXn98esWcMdrAZQvY65gIa5puezTM0X5d8d1Y/eri
Hx70eQ5DlltvsX9gJDJ6L6rKGNiMSHn2rGMHTTOhnhpwx0nCThdsnpYo71CzUjewscA5iFpVWj/5
qzqdQA16bm7i9wA/Xh1WHz9waodDpqZWVLbuWpErBhh1eLkot3wtMbGdwsffiSDvDqmBbJxS+eIe
dSLcH0WghM0NVOsNbEIl6kxeHHueHr5m0DQwr4CilYmDnF0BJsIVO3R6Y1q7H2py9n/Z4i3tKoKN
hUJFoc3O4+RyLrDWQWv99lr9wTiE3xT0bYC218QNlNBrhrTuCt6i016zh7+XXF23jr3nmBK96Lje
aAcDxwniOqPJmoWq8YcVRAQvqLm16JiMjpeawyonls5xoiPNhL5TQsy3kh82B9po0ZhhW9cJQpwk
ofAFt/9EhrAR7mu62O8VYBW3T7F3lazKYeaQz3vIVzmPPnMr0x8mVGY9QZQp9dNqxfLcfMHu4GtC
D3HIXRKHoOaUBsf6lpBnu5J6nu6uYUYfLvQPhEiSyM9lPdVmDPBYs6PUY8CAtpkYqk5vaVJfJ3NC
lbWAw2yNa9UeX2naJVkLJW/PXXl/afMNZvw8ROHEm3x2tY3R6Y4r6JFZ+DeJOpKkSowQZrb9CDH0
ttG7d/mBDAoqHRq57LJUluZnHYSZOLY+hgGAd/bHAvulHPRMW0jpmjzs39gDDK6eGB5qREvUyxi/
CSaZsiKtKR1D3XasZYEG4YuLiFPXyLumz/AYqLTAiVCheRFVG7sGzV+0mK/ApnVy0xq4uPciGbSF
pTY+FvaIqpbwcoDA5guwSnM62WlI8xacljctQc6VYbIFtngB/7BMDilT7u8DAZLXvKNwT+7oUqql
bVj2MiFy1md23gHlpKUhRvwfFS4po4m9HGc1XyTSHYkN5gwYmechv8Zxmk1SD6DiMtmqbLggcDAF
zoP2QZC4KNdcuquMdBFmSdTxKOwvkGMAm7ig5kyWHHhmrb47sMkYdA1yKV/wZlu6IkmKiDCJnPo5
uWS6PUaZ0wsMRWH3Bi2vJPxn6Yqf0lxZeHrempxHd7eUCa9ik8z6042jTmzRk8upFSE0CpuOUrmX
a3ReqkNZYNso3Ek+Duh5ULUp0YcfbRM5bdVMNaALs32aE7t81wMcv0k2vS/ytg4uIsUYxZrKWScK
PuJCZV7FZr8eZZSLMZxhac86xFcAQ6EqYyvewFpHsJgieAWpiwcxblSCT9xqGosbMwv8Znp9x3kJ
MNkHfdVUWeVqhQ/lltFJA48SAc4h9ObxApUs4quQPlnfCgpe0HDzp7HmzNqHyn0PcbYjpkTcHASZ
1z4kcofVwkfvv+k2qTNhn0GyZFr3KjRfL5ynwYToIo30BZDjG+Y887/WC2ZNmKVoxyNpfRZWFnLE
+xS46X4jQ7UVVARZWpZi1YopdVqlYq41qZP+k+vkAny8NxIbpNintMbjR7xezNFK8/3U7JOMMg1W
EF8U6zo1f5sa+At6mMpPKjmjKk2jGCi0/lkyEkltM2BDJm3K/gmOLsLpnmOz7MApWJYENla5uMXG
tGrCkJ1+s7TSomqPNT7J/BrSxSJjf9/pAxIlSNSjdhf24nR4rP5HRF4YHqLYi0kS3wlhhtcUZbmp
0irqhCFTd2g9JTDWGtvuv2qux6KHIcpE4AgMnf5IWw5HKha8T1jlF8X63DImgYTns1c/QVSRGQPW
H0htVgmGI9zDW8DUfzPl8n2slbGp3ekxp79PnxZckpY9akMdsOZx+ouYrfiC+Eq3cryuyMf+df0E
lm3o3aDx5HHxZSuP7tl97+ifJy5YFenRF0frTpe7THsq/L9DYVTvSUvLnpUTlpukUci8U7Ul4VfE
tGCbsLRQV5giqHvnGnevk5mlLqOy1d0eo/mxQ/iZ4VI9IZBIdP5PmpDvCToqk2LDhA7NrNQOYzcL
k8SYwuwqvCjaJdVpYxUH2/knNAyd2wpAlXu8VVemawBtMz5zFjc99VhX6Bq6hL4MTwN008/W+JVt
RpTo73+EzBRdUUsa5LITgbBJ/zxmrhMsqvKpXhqjV6CV7jPmkMyLQE34UthB5cPWXWEWb/UsV3k9
bE0jY1J1Nh6gbJ8gBWW9OSeOCMHZ5sR5HudDje/9HEWyvfjwFZpBzvxybvz6XZqYFTNFId9L2MNr
LILie9gmiVDVdLfkcRUWn52eXIDuiTVx/mPELmloPQobkGehiebU6m+qjKFp8+HhwVUsMUdzFIMi
xIsH147cpwC0GL3yd3v23ARdwT7h1B7OSjQv0xRVPlJcAwrjv0YOpytUPFcyNwpChiwv8Er7j1TB
vpe6itD4xQEEszuvXM+PO8fsEkYN2rqHXJ2iYkZUwVI3x2BGvtaS3AIhBgq5tFqodjPGT87Nkrqe
rUrvHVgP8KdlIas90s59jsLD3Y/riAb+MhDx1gqjXHxUXcDHfi/rXt/N5M55wUHT3UeBBRMc1qBV
4p4Cv6kIwBRlN7L7zPNH650Bg1m35xCCbVZ1fm3TBZkLp2iqFG2AcEBi/PJ5sYbau/VbRNM9k7W3
tK4Ihc3yxI9KzlgqJyuvdmY/HFIj9+nKnqjcGhX7+J+1E8rhrF1BtjBMhpmxkDI5hVWyXaqrI1PV
DyTmqrmQxQyEF98FHPVlbKKa0ZyATVNlEePiUcGEfH6zcMSv7vw0T1GCGxp6/icic7HItwSLu7a6
lJGF8I0DmCMik2IjX7q+BBMQ8nxYU1s4Mgm9XkSaIxHiNswkz0AnKL5hM5s2/gTbGuaIDskSx8ep
hNHpxU4e+ryspD5bGLTRCWVcczs3dx57wHp91Fkz1spRAvupy88kA6x69USIlZeiyDabBMOkOCow
oq1wdpkvmMoyrlJmYXSLnTmhNCYF981hUP1Ca2ewwl7cDXwVP7ROBhb8TimxFfmX7S1P8l7vM4w5
DlxHT0Fp6GdRVlw3A/Xv0euAysJIiQwEzPvqXMmJZqO0FQ6ngbEtLy8FVgkJ5GElmTh0Ai2Hrq4i
g9r+A2mit4BtrBKwPaGS9tr48ChkYDj06cjpOvNmrR2Nvmt4Q+DCSrF0nuIC4zWVW8ngZP+PWucT
AgcxFqt9vM8ftvBbx78tE6kTaSPd2+dqfauLWM+6BB/DKc/afLqkT7EL9bv/2ASeEmpHbh08mL5A
a3WBYBZZVCj926ahDxFfHO7BQSSfsC3zRQ9tS0Pvfq4T/OXX4R1bwYc+U/aubqwNA7QLv2u9odvc
KQFsbLdpSyURumfomf50BkEfwZkNxLsmnRCRuo+1XrnLRG+KotUIV3WEzlhl/PIiAaGTgjOjF55G
zTflTG6MaqJB6YWiSJCDRA0cFiwcmZkzW/f+X7xdfQvtUjSuQ04XaAqssTqqPPFoTBonD7O/LddB
KEHa6c71mqQQXd4Ejfbbd6HcBdJTJ0c6g6zdNdV+jogW8iBBHv4vAoI0B6aD0QnibU3NUdgvdUEu
M9t9AOwu5YGnsjCXgbp+9wLZG17leQv9qsk5onmmCtZJYVgeNEzNFxyg7Shk3y30n8sxipl/aUdV
v6ovn39CtR3xH3lD3LYjdauztLkbEoxnS5YfX/b7PB4W1O3kCm9HeP2RjisCBIYw0dXKXH6NKPBv
+cTayIerpuyb5O/wmSY6/qdUCaRCSmfhOnlUU5qoZup4MBJxlodhBR2SCpzVPpvm8MT9N8URjguw
i/bkyxkHEKF10KBM6zDfJ3QJqJ/k/WdZmrgUN+hwwVVxb+BT+TcEp3cFWqXDb136AgbAOsmk+VGC
Bp2tAPqwr0omiLDWPyyJHhsOC+QMAWQ3p6rd3jt8AUPsiz78ODw+Sah7um8DtjM+ngjuTfmKEL6N
9jlWrPJIcmKOJUvBmKtrCBoCfXZUcMcQnNa7HYvnngXrHG5L6NGL4dwwAfUJ/j3CRM7wy0zf3l9G
wmZcVEcQ+HUNPqMKqnvHrTLf9hYGE9rc8FfCscXM5VaieaiM5/xUVySBIzv4I7gsYl4IeV7NE46x
8VYdZC3k13dcvByITQGgOXNf+dx0S6lFdBCkCn9iKicKUQxbBh2VyM9j8ZfHoC2NBHQc6+ztHWPd
e4O2+RmZa3RkIa3APkmWhojjiPLVC7ZVfnHq5r4n61dh9/qiFoc5Rg5tqsao75ICn2DR1/SopO94
qnhdPy+Si2l15+QbQiSB62qmlF2ZihD1KQa2mjDcjXR2Ev1OoS/OP6Vzf7ZwKSLrEVf7CCNOdCd9
xWut2e35QB1/YbjJ35xOCrzj5A1UFcgo5QBuPpYwz+KWrQ25P420ifV/7QZYfj/av3uuD4vbYDoe
6cO8CKFAhG2eT+pHVcWLswXsYLnRkQ8V6q0sYu6aCdI2p46v2ZK3p3PUJUZlwVXhDkzik4eFlwLW
O1h+2Bkua7A1UU8S0j8DSvGofNf1eUuM24W/ER9vayTWR3kaC6XBsVSvKhDfWRlbswzsGJDmoheR
YPKMerfWwy/vWwJcFPnUmNjsBMketRhkzBTcPKiO0LGagXLk+nXKl5T2NDbI7i7PiQev3CKbStLv
cyoiGxhNPkQwnhvkiG1IeD55E/gDAOmDzqG5Xmf3h3t+4Hri6Fz/PJzAz2b5xqNV4eH+jFpGMyvN
bTnfDSbo6HolfSVNoYgIojXwb1FJQzIVE2XssW05py41HqfsGEN+o3EfCROJxCB9iNFCbrXktzaX
0492x1+9tjKXxErHOs8Hk7px7qiYTD1MWBuCW8zJcmMelroNpeP/27HW215PvCw4RyYqcWuzisr7
eEPq8tBUegYWNrIFmLXD1M/GsRl1VevkaUFsHD1Ar5If4w2QxkU0SkZHItqPrR5eSC9NukRYsNE5
NKHhjZ/f5/9annPAFQGDGSX8k6JaRf7vngTvg0dTYtkAhbThufYp2QMcFJyVBd0Ha96F0Ppy41b9
Z2fBouS9cn0dWhiflXLtw+FD3m1PFDF9nfVXDBktkVfl0TJcUurSd3fNb2iBSXe3Y21bY7Tba9tg
sjxBW2iej5YexPvBleeViw+Uu8g1xTps15eGwFHrj1DiZiNAOYfagZJ/7YP4+IgNLLXEVgnOV/yV
lPpP+TEP4i/LUywzAeX35h1E6xZ14Iiag6MsOn67QyGFj8Bgx6zxF7ASoR+dWy5DlEcpmEN6OXEG
7lRPX4e2GqCwL0g/cVcV+pdFm2aSsfHZnwPuqaUxVZNDy2ckdEZCYQE+6ot7Ctv67eC+5V8Ob2R0
9F65TIZgnZ9MPJG9Jku7AaYgglQ2VBOCf/rh7R/+i7jMUw0tO1MqKbUO83vIHg0Wf8d25fR6hmC8
n70bWrujn/2FQJQ129ZP/QQqs50bBFv3kzZl6Scquzhss9EXGqT3Fn/aBS0U5Zui1mbY+Y/uz98G
TqtnSfc82Rd+T3rHPMAcNAdw8aco6GnWOcYARjqfAsYHsTbe3ZOSzVjtZ5tojmK+TI2WqyZDjwwJ
pmFeZjtJP+DTAWLN4+DmJntISCs0gH4MXWyJsgyk5OCmvqmRIP7eTkTAChLet2RoaWUEJHbRzykf
TlMcozVOLATG+YsT9q8VwLtyl5ggMMcIGdlbxUjV2y1gAj+6vronC/odnevZ6vOdP/QhLpT0889+
Uo5DbaQiC5K1axvBGAKlWjK5YT0hJngfog5SJdKgBkSDsIdpJzIQsWN48OZMLriv5mopr+5BQ8p6
HbiP8l9eNQbMKntGeDHhp0Dqj93GMId9Lh5AXtDqFen8I94os7MdYUzpYNwS/WaBXMdQMcJrR/D8
oOAI3cUSM+4eYhbKvLV9UK2nhtqaCusyrDDLopNm/LfGZJrAtS5IK7973mwsud3R281LqvTnYa1k
qMs5WJFuIopL9jBtM+qa4tIqZ+HgRqe8emo/1NB4QEwwteb339JQlUi3nlu+aK7ZSv+6eXDCoDOw
pnxVSP6/ENbJRjF2DBwHQ2F+1JayJJmyXjsfA7Yqh2MAyYy2RwjC7UMfupO97U8gtTDUk6uk4ZBA
N4L2LwCRAuusNN2J+VcjxQA46CCBIzY/Ch0YCoeQK5D4Hz22DDsfxcRXYNWBkYeVSl0LIwnUeskh
BqvP/k3wGGG/JB4JdW8N15IPkIxfm8MKIVgBmiwH7U+8r+J5/Nv3Su0N3oPBQTgrWiM6aPAZ5qb+
rjcN4erhiqk9P3hBVz/ktJT2G2SZch3IdcmsExlC/qV/1HwYd7N2BvB/jFhLZa2aOpZp9AoywS/r
9cI6hhlhiJc7/Jk3fQeJGhqTOPQ8BGzadZFaZl5PAhFCpIfbJoc3D18VO3AZU8RJrDbg36OKTG3i
Sqp/qfMK9rOCRth51a9/Y6IIEYxWLYbi/S61HWkf7Eniu2Sne+TomFofGSwS+KhcxSrLJMBTeR2E
ZT9vn9NIY63Ff/ExGdE403Ut4swDXPP14c+KxwqC1BQTodDd3QoXH8sUzCIKag7Fl/0hJ/Cu4Uap
zbt6savmL+hZohk5oa9rTEJPcMGiLXl8DCXdnmp8FBXMPk7iwncuqWOnL3XsP/MZJCTIpLap/Xz/
FzrfGpXfhMx0ZG4XIl6dG/m4hggGmXDlpETdF3fdHAtDdJ0SP41BFQlv9pgO+zbkskOwDtrL7zl4
mgyCMl2qsXXDKexsQLS+mu/BoxnPbA0DNYPY8tmr5STjAVGIItL6fnQoMiQraW/j0qzWzRn+xIqp
LHDAmGAxnBPgBSPgdz+zD2g9j+30r21Zi8cQ3U5eS7IEt4XtHoOI6XlA4MKEwD0qR/TbVDulcbx3
G+Ytqekg1m87GEiYun3ltF3baFHgPwuWkgDJ81XLmdcz0QcEAE3uHQz0j/s932sc+bTOR5UpweTp
i84nNnyh1w2cePLVtW2jg0Y0zIgxmW+1SkjVF7TMxdvibycS6hHr6WJznnb/RKZIKlWmFo9mzmbA
bgwhN2OGKIuE2FzYY0DiooS1+qKQR7GB57FBhEhwSuhDV7nfMu6wke3IpcPFbYGYRAaHGGGI729h
GO9KP7ntO6hActIOOYGhyje26oYkFwuRtyQ7r/IpZbaDCuh6wkRp/vXa/rIVIQhDGS5qGiZlv2JB
hALqxCsYIP15VV6AUgRc/MQcM5FywUM7JmXKn1FIycnQla5XgF2I6bgT9s/+1AQAi40H1wJfmmFA
JuHJSe0jHfSUabpxj3cm3YUt8/001uQ8LOdM6JP6ANLDph0V9ynO3ClMKXD3gTV80ys379Xsm02v
eOMkNuYKIdvrA8A7GaFqRZTXXM/12jxbFSs3J8CP8A2FgxlKXz7jn7POaKKjQMZmhTzyZnk6dWa5
vCn6+YHQN3nB/j5qO7TCgLKpONGiw8ZJsDGwzCUR0NjglkelV8jCygO44i1p3DIidrrXZdiITuhU
sbHP9k7Np1eAQlNs8BtN4nJceH4QXNKMbOSMyJvMN0O1eNy0ISAPnw3jCsB6rB4j2mdipokT7XNH
3oVIfkYXfPwflNKsss5ZPGPRhsKUGzYWPBSRMRlDi4XLIwSBmp3MJ6YNx38dXHwneu6HZTrrMVwL
d7RhY2N4ArhsCgFx2zymJ1l/WtpJA/zz+2WNAJmtKiaRrOu72he4TRG5WXr6mkSzoo2KabDGhauq
4zWBm2vxwP/+y9uoaTPq+BlmJhY4TwLM5cbgmGa8lJbeJu/55wRYsVihDOmnN2P/XqEEiVDZ8t+k
LAKOwdC0Hrtw03crbXEk+ugvI6thbEqHa10P4TiIqaVavzeUy9+EkTweF7lldL+/Sw+4CaEuLrNQ
YuyiaJWJ0P8X72RE79hfPdj+C5FGTh3qeqpVRX1360yOqUOqSf0JYpVxHOJLhb3sb8PmkiwvrrNL
yLT9m/6n91CoN9jRYiIh3BLIfUMEIWu/enO0PAkB0qW22huyi11vBCdX2VM4xEtsMWnJuby8bSMR
Nwwc5QlmZCHY5r/+BTfLb7gRmRFYkkhoOw/I174ddRqkNwh1e8Yua5FnU+lP65IvcuwOVEss11Hf
uADD3+B6OuNeeQOrtCDJKlLPK01E5UUbMPwyJZ/c34KItB3jDFhz6T/OuEtISU9x6E4UtAmDZwUx
cN7SNIJlABZ6SRbAudvqMDZDVDDKTIHF70hltdJUZIkGpmmWiN0zZSy/qoSlJnH9+L4bgco+S7Bb
+GWMhCepGwNHFSztQRT4Z8PDDamvMkvCb0yxJLLqABHMXVaRWqGR6s2g72qsEmIxzJCBvQZSoemu
T2mEdsKK+Sq4xrIeODKyvJuSJyZXHHlzM1wlqtmVeoS56KmAhn6CjRJR14mvLaYH+yAynnBEG5Lg
XpILVYHzontd1pBHGMnINA6ryZ05Y9nqYgGbDyhBI5DaCwk87jbMcFfeNratY/npEli2hZvkme3c
E3T/NVbaP2LhYxz7CFCyn2zUDEA7/fEbeGjWjumIbOHG5Fq/6D4ageb0CTefYla9RpPBGcPgx2dk
0Rspu7S1EAHSAj8Dau6ZOGzJKYvcNNIwFBq5G24pVP5TIWEGBQaY1HnItyEyuttiadrBSwUJF4kd
5vhItV5OcGEIMsRXRBYZb8wP9WCB8bW5eI7wj9kSuTWXUBx2MfHwxCBC/S8Of0Kx5Mnco7B0m0zW
m1Bq239bXKz6icwg9CwdglCiZ9IsLLpi41nXC0kIqt6G5a1FUkMGKeu2z24vQwQ1gyNhIIIgD35+
8WwQHldS4g2ftnCma1xUcHmlfq8vvAPfkfrPYg5XywCYaqfnmHHH+AzC55AFUV2EDzfXoA++EeRR
8pVacaU6p+bDWkXJJ61ojqYdSRo8Y9Pzj78A11qXoLHFsXMR7iniH3LQiNS6oFH509y1bsqkHwR8
QSNdeR46qFEJ0WilJ4CqO4+9qSY47xC+NNmUN81o+iqVnQZHjVlYHjjiGjTJEn4n6mdqGwaWvULh
WgnS84Dar3WqZBRKpGtTMKQSI7Ey4mmoWR90NV20qU/4Qy7nmQqyop1MVPsHScE+2El1Z3Hy3yG5
gGW8rOags53/wLxyp2TBtNDUf7UZivV1cVC2rC2QJFdCuSiiy27WHEiZfLCx0ISeJ7cjNPMyMeig
tFdsZdwq4qUbOKUNeb01WMl3GXXOFF0vG0ge48OnA1Y6xi/vC43JuxDH5L1Ct7bMZw39Dm76hZ6k
m9owQ4h4hD+62xOt5eeIyRomvfowuNqYHpMtE7ve45tzSFdEbQkxy56cknKkVWMRH4XkDrvCGvwE
Q1tPOTfadsjcVVzQ7NTfQ+UnKw+cX+GL2gNFXd0faoqqehELIKb84pPawQbtQJgfPhtMgvnBKaP/
jZeAqoDsF2Mj+RkaI4GgoE71ArEjPBbY7vDsCBEhKuQV2teaXwe2oI0Fr/8uYVF23mOHCJM82ryX
yl7zyG5+9cGaGCVXiuNvsJbB6eR+r7ztyD87HhfFRTQxpjBGVRlYCVnNf/ifYg4+8S/YNhzD1t8q
pMSLjgVqVFHZWUqETDRorMUe40xBXOcOSv8lNG6fs85B86GQ8ei4ugO97B+MKXQl9mfqvitSQ8vx
d7NYEBPmALJWetQhhX/x9so+z3KjTHm2VLMlYE4t+hDPfYNmTqJ+vw2MgEj/guKtC0ZDcP9uQvFI
MQyPAywiukiUDg7Hmse3ZUY0ElxjMu6f0EJU0gFjJ+r/mcaKu7WeVaDwYfverifvn4Kz1ETfE5lY
cuAIAymGlMj4veqoiU5FnY6opfmnCLAgJVOBOZdx3rCMFdtbWoOH0brF9VMwJ+0LkVMkuHCgTPdJ
EMKzWphy74mpJoOqalmfI08YcqPOmLBtU8549jUjr3EZGvTfbq+f+HYUMWj4OITQhoPL06nkrnY3
DPVmMWVlgIHcXsrgUB0yhrvX19GdyPZavhbeLw2LGu1zIcySJ3KbtjVSH3hf/rDsGjOyX0B//a+9
qDzX82tqUzH+qLcEdE23QhoZGXZ+Yyr2wh2LjVIdyzeA+E+mbusYEOKkPnLEhEbyFNgD0JFjMlxi
jggM6z13n/+CDFNdsxETaLFDjqhnNTt1LDqD1g/KfuCRzL/uyTIXhpzhZWbm1VKtptonFybzQfKR
r2VE/nFmSSGkK7HM/k3irEdkEfjPFsS+w6kTPlzmnU5utaMnsnaBThYktDQUhMN7l7Vs3pb6hHEt
2rhvoZ6JjBdkWEQmhkD9no7LY4c8welgHEilFKTQlebPp5g0Ap7ORpby2X9hsTb1y7Fr0k2xpsOp
c+6Z2RX7xO1i+Uk1gDuqKqlnKS7lL5sWn1yR8CeNJKoluSmlFr/L6YhHkadR/dp5jniaG5Glt1X0
FXk1/3jlC49Y15uRpxzM6v00+ll4u9nAG/oswE3Y2O7pt5eRtsoiCkLxk9VvqAbBAu1fSriDz1Od
RNgtzA1WxAy/Bzpq3Ipd77gUoqdIvMrDhaxwZL9yJAxdtksvkb4RIjlq/ceksIRxnGG2Yyyg22op
soCCslV3xwPzVlCnFNGgCAdPfO+Vg1XwjCSyhsew/2EQW2CXvuRjB/9BF+ry5SA1B5M/EWQDbOVx
TBJDR0pHuByMbnbVTjhFGZLin2BROFiyJj4nkm2y8gPoIgLTLDGew0iYSag46tKNBPcU6o9wXu6j
Ap1Pvzwpj6BLk3CKdfcl+iUddLg9DN1RP41JMvOLdo1E+urqHiCe8Dy7fg6vRdI/3NUWDXWO8N2W
BbBunEM44RbfqjBCy6rBM5XNpiRqdJqfD304/FoelJLtHWDm+61LVUlAAZvHOLzazwm3XCj5IN38
5ecRUyOSgLcpe7R2p9n0L4LuUUnQ1FWNSn/7OhtmDb1CtjfaR5IUGueCyhzMVwzhBCC2S5AwbAzB
pWnUytGPIJ2OqHDVPQFsCqmzxVew9xgFvWHWKfH6IjpKb475QSFnc8Mx6P8leFd2gcWT1HisKKm+
Bk75fDqPzzfv+HZBLe9DVBDExwVqWc0QKSLObw++blqT0xwfEsFU+8qUby4n2qlGcjOI8iGBBvZr
p8IqNHL9fMhlEe9BuSTV4Vq8z7RPM/nxNjoiqxQO22uqP3qiDkqQ3ys2Z+TXyQ+bGj6EjxATA5Qv
WVFe3DLN55+akjGzMIFJHPh2Rtx5IqowaOiFObc6roBwGbCAcXXU37bwA1g0o+Yj02eXjomJaExe
lMTSTYW6MyiKU+f3nZrxk8U8xxyVqXeiiF3AVn9hYeJIltOk2bvN4WzJ5h9U/cZQSeoXmUQTOl+a
VkumxUdw7aR1xeVLIUmLpW1PoJr9H1LpdP4JYKPtS85B+KEA3KTojyF33MTjGye6FRyyxz8klUfQ
SU43E+VyZN7rBcQPrvx4E/CtqfmNeujDu4FUgf4iu1CE3AWhcbQo1K/0F280FKIwe+MAos8lyrRb
Png16C37lFgoxcp062HNuri4BhwJ+j0NzjwTPkaXfjUEDYVwClwhgi4eifoRBg+tRuWJsA1NyZod
8vNYjb3Jw3FldtRZgl64iVwFfz0lacpP7CZocHGbTyhAFNzRaq+ZLSIcSaDzRZH9aNPIQN+kAyDK
gLnQWuN+rxk2LXL2j9fJbxBBZVgQrIFEHsAGyIGMbpsZWfzjMXy/8cvwy4qw/ZBM1EYp6lvnmDax
FrnBm/RkXinupOOHWJSCWVbXh8iW7N0So7UWn+i8Sb3YPD1W7yvRRKukbPlOD6omQYv7DTmX5HJE
Z2mqUhmjpbfxH5RCvyxR8cLmUwJ/wTnXVgPYhXwBo22VU2aPxcxRNr4RfF00S9q/iaWFyAsGeA+D
LOJfa2LhhKE2j3BXJbXsgPr73sfZFTiELQgpV0VjZiMpJHCxZKGxHe2e5la4+SBfr+U2gvHJ5b9y
/tna1BWMkGY5Fj7//WxU158njROeHYfzJzXeIz7xVZ3BhaeINRziJgqRqn1BM7iA8EzeeuJzvZSJ
e9TJRK1cDzFur3RlHUS+ad6BKiPriqSQbN9JYDykaXl9MjbpXD5e//Qayy3y0LfOFQs11SFWYgxb
wI1qTcwoxWDY71xG64TkbqZFw+UBxsvFFLiuTvh8v5l+i0lK0OqApJF/+i8CWidShnD6ijoN3rL/
Sdp9NIW0CP9KsxD0zubjgTqhAhb72rOJIQ6Fo3SgGx3dzVLGGzK4aATyK/HYzbvfIKdjHZJsUxxD
6mseYFEDbWCVil4qPyLMK/LgJYMWP2u3Fn9/kQGPYuTAhRqbn0uu//P4TosGjd7uVAbdcFmkrLAr
ODhndR42T8OVU6hDFdBu6c3noH4U83QZntZ5aCi/+YkJ+HbOJ1RULLDlb44HiRQA2vbR10kvlagC
iZLZM96rF+SGRHSmKdHfla0wbc262LRa6QtM8GxS85quakgL3e78UAKLo9xTgOGLGHql7ZmL+mVt
+sxdxn2nkiYc5KzDpIbWf/56LE3OqhPfCVOO3d/yfe5q0Dj8rM+5OyzPGx6snMGg1tN9sXwGtLy3
Dr//QjWXfGlnayXfQiEqr509c1VK0LZWDNBcVYmz5lZkURnUaDqcbJoCdZQEoDHc/eXjcS3nUdCw
nxcOlGWhQnFBWVSwG/9t3netVvsbifyj2QmJY8jy1fmPjbfkTorRuZHaL8WGktj7KdbvM5jBnqy6
wbwtg5oftfT6S+UPFBLUSiW9r9EcF4NC3V+ZIyGDFhWeIVgrLI62KMmG3Tkw0mqrgCEfzIjbFeDK
ThVfShK2v9ej1nxWtUdnNxMT0dpnOncXEC73oEzHXoJS/gJKKMkr1Ao2rqUzPIcTJGln+3IDZm2w
PC0acc2IkVH0hHykpr+JQW/nmkShrqG4l4Hp4x5SpxnM98+XDOR9poSn2PoYhe1FzuHkQwpFNNsm
F8iDdnBeCFp9RD3/ukIOe7ksx853uS8mAizgu1/Q7knT68GOiD1Fs/7mrwxV6es/LnlGEI7ZwNlI
nx84wy1xDUydMfY8s/50+0THXXR7aTdEN3wVQJS/r8HvBRYK4htKKCn8j85JenUeLAG70qEKDeG0
4ymy0x+LuoF27xNNX/PFigUNk+QyrptkJK77apFSp31kysvejbVXX5Uq6RclitiqKVQ8jjk5VNjt
pshpD3z13cTTwZ4LPioxP5qjD2sdvurpwo1RU+Rqx0LQsFn75f6Brer1P0q0h5HXOeYeAt1FyKxC
knsC2PyF5C2WuJvlAr2HrSCCMS0IiSPI2ZKs452BUw1Uy7T32oCFWJs0YmE/o2onpnfsLM1FuZeL
AbKz//SSz0RZklEvOrax/idV0hJ6wq3+80qHIPmbRBiBYIA55P3Se+gUcQxGdz+b296exTd7av/B
BiLvo0egofW7B9x3/SHQM+y2bt5k4qMpGh11oZ5cFg2qfId7n8aJHahsLmTDEU3PVaXY4x+m+QPm
/l+TPZK3aarkavvfuR0sPIiN2fD4uQfSfIlhKEdqIbVuji9XDD9zF1vl+XD3ldRcYguxobRZDTzJ
tUJ8JadmtQLA8spp1vphNnn1y7Iv4eOu4nqZkXlOmNagOeIJMtH1frY+sEst7xKcxTie2zABesSS
wJkVPtJZbV88zig20IttxG9Ea0N5qQjCQ2/vCbLtWlu+uWcLQH6WL9GLUhkqty4/wEDFLT0k2eFL
ERQ+immV1n2k4IyjrY8PxPmPVz6MrwFcPJl5O7shgOHUmMK1BQMdVn8WgYgzFc0x6GHnPMqxaUJu
OqXJy+e7ccXY2UKAmK3zycyksBmOovW0unR1fHG6G9nXjYilS5T45wEIFlHyEkxlaGYh/fYnGC02
1Sme1R6RqlojF/X/pWP0MCRUZDPlqXC6tBockHHQ6h2RUwGDeZ2pTLK6w1gE8dUwaC5eUnElvV6p
rv3paLFdubf/wJbM+otRZL/OPxYck6bnXAPVyfxuu4SfVfr1HrbBdQzpcrgx8b+6PR4ZgORUvZdi
AhwQ8+9Fj9vTGYlLO0lLC5v2DG0cd9q4UN8BaWjkvOEkNP5NQZA2IlCRNn8nhJLE5dccrXXS8Ueh
tnUIjdR3LG0jIXlIpFDvvuX0fz+F/Y4TQVTaMIlQq4E/KXF/w8CS1rmpAIIgObTHqN/p4OJMrjt0
LoZkKxbL7SPZ2RA7g8RBzIFLCRZR4PAfpUt/6NZEd9KGqja7dHFQD90iJVYynAaEpzp1b5MoYufH
YCcOZtoV7hf7R2IRWmPicOvfAQMct+uQx5Rh9NTijxji2Vv+QAGt1qQ9pfoQa0uSP1TcEIjxcu44
OQzxDbEiQAPXbHfyVeovI0mbMvlCwHuAojBqHrIYDYsH9l6mI18kgcuDxaGo4ST2uKKZAUJpZGdh
Ea8bXktThQm6+TsxOkNUKNWoPPmSsEjVvTaUlsSD6I7K8E43FfOL1pvxX2txcxoZzmpWAiutt7JU
3Axa59Z0zdqPpz377a+rIihm0X+iGBRsCmzBytVXf1Zk/7IRxR2XAjn/8h3I1tvAXOLqpHkbSXIW
1bkD2wcGuxjIO1pZ028qHDm6fsAsQP6272Gl/mMVsaGzl8KrVQauVqU702YxGSVgBenwq9k6kB/k
1xp/rUrtvqoIkblvuIvRMFQZ2U+l5TwO6iDMxYXvV4iKz5JNZ7/MVXKr2stMAKQWqHWAqnVhn4YR
M0o8sqSUxM9hNz/c6PhtFoTMFJYcpEycvDdMR7ChVqTeo7WxmLlhLwXvr0pTDopeaPfYJ72EkS6g
5OzPbzpLFytRFiP2EMwriE33VHdWhRM6G4VyiGSwYKso3/SVwmug/388BTjht/TJoi6mIvn/aoc5
wvyhitKI8QkveC6Zg/LTDiCDGDXd6tqQBSfZm5FwfEz7DRG41DY9Xy+uUavn0Q9eUPjZaLMXx6k+
ilqopplPMkdxUiocJ7FbuxRJOXWDaUExrNbNHVzMMqRg69BrZz5w/edh3wFr4USqmmYm1S5LookO
v+iA1Sj8vG8zwAPF7+Z5EVfSB/tAe6Thd104OwhAoDAW6/7/Gu4uIPlE1SjxHQ9fCvtDsE3LmKi/
O1cHPGUaOYrXlS6r1FmjZK/WBTc29PCvL6LwE8BX2Yx5ZnXwH5EK0rGtrtl/vObkB/vdtgJaLrbH
CFBw20zktYq3aFfCPTJI3r3Mz6Zfi/7DCwEGxSm0pB52NKQS+tTjItGKj+QpQAhhc08lFXFqVNMB
YjijOF5i6TrcPeyC/I1rEgLKuqWL5ZfLnd+jb5hrTiE9hdUDwIprPD5zfi75/9sL1To06Ga20q5I
Sy2MPO8vvwLsH4N814vO61hKWxH9B4AXyLDv0+E0jSrZ1+Mmf8D6TfuTDQhSf632UjsOR+TbBu57
DfX8sJX8CoqqKvvYlJK34j0FsnN6jhas+lxv+y+ZF6dGtS4Z3Z/nTeL6KL7ToiVdEb/5B8qK6qj/
EvtVRAQiZZ08HdlJHlLhdzs864yw7kJg0uKHboubUaSC1cDq8YnfMpTEjndicpdjz+1CYaNacpwQ
dYyFwQyVx78O4cVinteEHqHJv+Bl00QY7c2KhMMfnHIDQ9icWoAyWnhkZOeNSfGTKhsahxBIJvMo
c0xvT1AO7qELHftTJbwHuQ6l+BusOuqNWjuxVgnbQAFJVh2x6jVHXM4DkmEWo588mdRBKmJ7GOnv
eivplpf9AD1m5D6G/eLsI98ywFBMdunoDU+ViK7nPpPNwW9BwGA9O6Xve8zmQzl/wvbGroKkGC/w
j1K3GuY8nQ3SU1lhsWUJAaFLAN7SDKK33KeCv6XQGlkRVKzvDi3WKaIiFIo0v6zTX9WnhE+h8jS/
4P4OQ2cYX8OYzaqmk50fEb75/7CvBd93C6HbzMeCeJl5JTRzraDxdBUgtAtTlSqkrIZ4lm3YpwAB
ucE1vmgcGFNoFonH1xziaYm76ltIy6Y+l11K3jItqYSrPin/ZoC49ew1O7qAdcFQCxGV67pIp+P/
7haivf9PN/bMcojCAticUy6WSFgeHX/jnA5C3a1JsOTshpP1jqsdBnizPAdDfZ/kE8cSOPF6pyGA
ZVvutao6OwKx5oukqHwhJb+3UcHazLRxlQdyVMzL0f+F0Vq0vy0wrLuCcq2eH0LxFgIeVUpjclOW
wD0QnwNvyd1IsvYFBz/bkrWdssGooIPFQsxHYmz1OBpiYzskNr7qUgMohSN2sLysQBRjaTCfkVHm
MAOw2vlaNkihEFMXT84NGyTjgthGKgV0BSBFFd98XRyVsKReQ67or4C3jDdseiAGeuIAzbiJv66n
5aFn2IQ41etr+2KIh1kCXffdnUuTnoFHCSJ0Hr/9PMl1v10gx6nyTwGSUsnsGL7a045axrOZR9Cy
FZSVOCp30lzu6z3RNoyECew2bAvauVZowpTFHRa4eKMuNS6h0bcaQuvm2xhGhgJaXm2/RDK/Ng1i
cS7oEEV43aj1xLhr+jzhynj8jOjPFFLTvuUEiNGEXj9AlAv+GvlgLipNfsIgs645RWiPNcy9LafX
mt+xYzcCDYFikPHNWGQXwI3E53QThruktvktcUuTK79u2oDug8JOtYiRAGeyuEJETl2jBFFl6uEy
ykr3HaZ2A7VtWBi6vlENrwQUylX/m2/YoFVhgOtjzzSFivbsq4SugCO+k0dblhc8Ou0zGXSF9WyD
pqxD5Iqj28oc6uGfKiPaJC7HFh/Am5v/aNN/ECjeGeFPO59+YMxbf6VXBhD5JEeM4i3M7J/+JMPh
of8V3d8s3jFzwckGLEMNt8ZT4Xyu/p7QsXERx0RkZm5bRSMricdo7jMhQzE/r3V6WduTwQPB1eAn
HJtToDdtVDuV5jjmVwWyhdQKZp6j/wzNKx7LU8k8Mr3g6Yivkoz/7nMlVP2PvMyW3hr38LeD2u+T
voqsEdAXQgb7Ey6ULhDMH52YWjgIUGo0qkvaeulzcN3a4Na9lsz8Dnj4aOZWyjOvjfD6DswS7VuM
0qFqQGZ1yxDljGH+tsO8G0zjiyujNyaHxE5lwp3gPLm2a6N8eMrkcjcLdUKJliKqriKUIvAXBDee
9SC/tkX6C6qcolCW18dLA2pAoyhVyODp0QHdtU2uJOqziFibR/C3m2PrQSmoOkjKrMm/+kKAfMjG
EQeHe4Sv8QUyHLru8L3QqCxIw0IuOzjwcr8uJjCZtz8GSGBRPNk4U3MTkj7HlcGw91gO9ImOht+y
E0PL0i5pXQG5zf4HaTQ9wRts2Pf5iZpPdC0ge7cHspOD4bPbA0mDp0Yoin0a9jVZ2VOj664mELz7
cev0WbSFcCq9/c/9X1YpwxVQYbFWp5VxuekTK0GzOqRwULkjZVMTXWwKVgbmtt9OgDlxWuKCyv1r
l1EMxuZvI1vyk98xaxxIh2G7nOjAxgT0G9UT9m6fl6SeORixOsjHY/HXBnmNqisLRA7y0ByNojEB
ClIL1wyNKvsTHrU6lxvhYaoS4jjgvydY2a/p0Cv34dEDuKUoWb9UdK/4qIJCZx5dm4rZZJELXTUh
dVXZaecdr+uQPteGxkUNPqiMeDWSFdnxiqzM2yPrb8cMXYCLDLuSVMTj5yIgfNrlYsyDaBqy2xtD
x8MnP66AvLhWIR5XFv4mw9Q/lGELSZTfHa74AxeJPVTCv8E8ZNrkXhlg26ezxyfJLT94qFDx/H+C
tdSDbuPlkVDVnJyKqDUNCMPYFXEJMHF3qKQf1rTtoSElWkOiclnMG7aZ+8mn0QvhIQIlgQVUSoLP
GlVfBR0H2LFFrp6x8IY/DsjYX7ViPPIW7EivV3IyAmuAta8G/FNBMfuXPLBqO/Ho1htBk0KNgXmr
N7GpnUh0EWDPPVyYNtBFztrxYHohviNJcxAlYc5JeeeoPOYeo3nbxK9hLzdQPUSL7ebrYjJ7GTkG
ueojz2BNJZaqxjrsHa8FhGPa++fTBrmB3XYSYAdV8NjioYxSEx/wY6KipA5HKGBI6TNcOvtBg+eP
Vf8wOvi/zp4jhuWCItIv4U3EBvZOJe35SfKCGfKMd8xEZ5tBv2xRU1eqzWqFyWde5Nk8RROqccyI
iNT1UqMguLLQ7xMwCVkp5am/4DujgyNSv+sz/DEk4kqvmo37gCBR5yBweIkDs3f6RBUNMUZ+IGiv
MsUjMoAVsWCK6lgenqUWtb/0NRIVezsGE5zMMkslgNu9oHVjRkaGQ3bvXK0twzdSgjXqERrD7gsc
zKdQTEJHKZPELh5Y6obZVBCvdQGjeG+FQyKZVgsg2XYNd6g27m95aEsXi4lNAHPJLCcyrz2/tcM6
VuStd+MWuIVz9/H1aUgKG8+vCMeaAImCwrQDq+guAKOGkQBlT1SIeB7svurh4ZeXu4fvXIREuQGx
/KiIAjDFegLZ0AYp+pw0kXx33CHDijCc9zrbrtsXod28XekXM+05UgFV8aKaco/NbeS4SsJ56OuG
IUbx4TsLa3jSb8zHaVhUcmrrTDWfRIC6xC99JnTi0OVF/Ydi0uOGbpyUPnHiW7EFhIJguT5Hc4zt
VQU/wNci6sn9B+uRBILspzZ0KqSDV0IFtCSBaiN9nN3m6GEKDcCgLNIldBl8B9NZU/tMnc7vQuI0
e2HTBq/SU1l+S63U6tIrK1sjMj5Vul7pUPVwFZqTm7V+JJp5dFwJKkB6JsREnfvXzMefvySsKmDB
xuhMgqEUck/mkaTD5Orn/3wOubai1d1OJL8Cn9zu18f5igCjFQOOVJEcmWXTYrOuZ0y5iKnZUjqo
igvYJ+0QbkKmp1Rg+yhIxn1DdtYlkZwDlkGk2Nqtskd4OfDVoksAQE2S1Jv9r1zhv6ST6UzQ92gP
mgoP/sWf6X3QdwjDKrn8hLlEAFr7WPSkdqa8m8bwA7M8Jgki+TnI6IPJeprtFCZxALZYWeHbU+fy
AkI7D4Jm7kiKnyBrlRugxzqhrrb/4QB7b7rP/JXGfWnATg/e0MNhOFp+GQkCpaty6YayDQn3lY2E
Igu+2poNitNQccoLL72WNZlHyYPla7J0wohgdYGfgDCXiR5uDwdadenVgsIEHg1gxjFm/toPh93o
kj8F0dvdMzQ9NtooSGBBHuFpwbKMhYtqAMY1Qv/aGtRO5eD21QQPQ7t91IwQ6bPdxiW2XVJXGoH5
UzpY8ywu+Yvy1/RECA3KCacsn4v+KzDkhk6cwZHmFty1IIvr7UpWXy4isVPe+lSWJVVRyqlYMJi1
XXSy1/ZH6iwgS/5iWmV5z7KsPnlTv93DAIFV1q3pW/WMDdnBAzVhhdz5okMDDg0m5SPLK80H5VdW
DIbv6+Dxpb4A8tEdVcLEwN2SypAmoWkWvlrB40SN0Ts/8dXnEDxYK2lmIPHHfP98OHj+o3osXYHh
MaIBN5dhQjE+V6Qdc/gJcPyDiggWM8x41+a7BW6yQW6tX7GsmQmqtYy0soxeryR9UDTnvcPkwWrk
pk5GWbL8Rca40spgOPiaWz8WkpGdCFlRsV9vVjG07UEEoofk7RJCOb0S6DKhs9cN/XbEv/vHASx2
kGhEueaXI7aKkY58GQVP7svx1kXe53yCq7wczvY66eIdGBsXntzsLt4Ud8VhpY9cQCydH5ybMT6u
fnvg/x5jC76/9ax6yv5pXRdiTTI/6ZULzjmfPI5A4wxOhQuX0vTCP3BA+hcZY0weCDaolYQXkDdE
Gli9Pq9Y31i/e8kkKYED2WLUFPqTt0dfsKrIscN7F5dYbPXSEvCy/xqwSP0SSvCKAHL+St9qfuqX
GU4FhhRMzztj2uqvbsn87/FpVG7YfTdkttcqW/jBH7PYmv6PCclgrsHygTWiOfbKtQ5bcbE8PBLj
pKlbZ99jqVHLGj0lgd/LQnWeRSAhJPxilKhaAl4esSHTHwc2AKXGczTb4+9Pt77JLXX0Td0mjT1a
WU3ncnUKiP9PECz5HYNpX/73Aow2etL1gyV5L0K1f7B7zpd7CXmOQj4t4jRSB7LcLqd8FjNl33Yu
UJ0l1wOJUSS1r5GGqkppYftUvpID/N3LFR6VOiQoIJ8zJ6FcjaiRs4eyEH4Rie6GLfCiy+X8mSF+
Osyk5IEcAGXsYcp5BAcZrHAmF9UkE2VtdBwhiVDy64xUi0EoFeqHUD0noVLcxD/GD/nLZHikOKPR
SzXmCuI1llVJlOKqg/eBFqA1RNQVX/GHbrosSXXlxpFeex2iy5mwvdWCkYNcOEHnIuZgEfLlMYGB
SLYuTr98EY7mm5QvZqVJrVQ6O7ZLI6yP/nFoh+37q/yYrN/dDE0HcWBHY5irwsLx1pkAZXR8ev/G
5P+J1HLVmGrmbX3CXKCJMZa6ht+dUz+ekBu1qyayzmvSJvXlIZpyujJDfUDtDdOcvDgu8vym17Dm
LPnNYPzxPeFtTg/vZ9GBMnV24W7C7kcHsyzlR4U+UH7TNYquNXSjE4S1LrqgMOsbhZYi9M1AYbk6
N7ytGhBr/oo8mPNpEsAQmrFsci1ZtJVYQ3GaMHt1yTDhF9spYmB6ocb5rJMd/xsxC8lMzrIpXyPe
mnwnVoZ92STtpc2YdydHNRqFGbsE6yWzL7cqv2bijQI4YVDwHGHQlquKk1FR+pyauyRfDVLLLxZ8
tNVqvPmQIpN+y6PAeOSAjy+VylmEUB0YZ8uDw95+yguGRC2/duqhnL2CzcYMKIFM+qVrtLEDLg+S
doZc6YOcDghyL8E3tQX4aKnVkq/BTqAe0+4Sbs459jh3KgqEEA6oFFyalC/nn5oAnTfAq0ALbj47
KJmo2D0Pe82tCnpAkRtmhQBZFKXtwoTBNtWSyXIus62vtp2WKuQcUtQj8Ym8f9zMXjr1lehLe5oP
hNrk1Lzzmf07qDXs49FLiW4x3cW9vPA+eIUm1CiTbnixVqEz/EJwkWt7TC54IbHVxth2m1Wsukar
nt262OHezTnNmEVTL36e7O/1Du2TXx8EPoO1s05hkVPUDS31WEv4KqQXjyBfOYxMNqEBCKf3LL1J
Zg4F09Si8fSoabO0xpIqa0nD9WoLILvah0rcda+HRLmzViSJ86CD5NMNkJ4rm1MzJkeZce8vyW1i
0Vo1CxgWlnEzmSZQWavayPhiYNFoozNzy2APD309fruI1Hzf+HTnofxbDchOUpYCWIXfXvHj0ZYS
TTiUigoFEDM79+UQXxwgZC/Hn4XOfcsP8WV3eUTw4JdKO7YIaE3cZWcCKf9bDsbSnKuRBl7C2Igr
K5nNG7VAVmtjtfuo3pITVOTnDBhiEMY0cKurUYkL2Uztu5PNL06TIdu2KpwKxpalT+DIYxZOGtoL
S7FhgAkc1cG1yeBRPK0f3JWtynACbEq2z70Srn/D6FQFUupbbdVDXXPun/RNnmN7xexLelwZpvKA
hzxm+5jvTQNbVM9Yqkn+YJgXlzhlbrroI5pOe+0SV6xvNmt5hTBtUd/HRkwV/ySe38n2trCnYGAF
vV1FWEoFeW72eGyAbu6InLivXuUauzFlBXbQ8czQy27OKlLj0XNQbo5L/6QKxkt4dALCFRIRJJuq
47YHIIA8aOAkiIZEwSXXFBSzrG0sSmsLoCTZtZX/LUvW/xFi8mvKhkxk3MX07vS3VLk9AUN5mjRI
YYZi3ReN7TtyiTLA27W3oiXa4IM4rx9hX6g/Dw0Knu1p21RYDsfYiMGJPYcotnp5Thj3yJfKU8yT
WeG1iuyfZsnJR87rGLuF6VimPgFjwpZOwUUHpuw5DGQX6ky4BAc3yRKoDMvav2m64i1u/hiJY16N
utoIXxyKBkwN0523o8aNCllTJz7oEJr2ceN7fXsbiGwdiD2PTzOXky1H9vSF66ubMxm1UT41mTWI
6mdL0jl9ncfvkNxlTBrk/2m/EX5eFGZbdXH1JEp/JpoWnrutRCQCgRrXV47Ct8Fp4pCeGDHS7pUG
hutXWS2/tAlW1SJXRRWbHe8zJDIWCBMoZTRZEqN2Va1jQQX1xjzyDaiyAsr3a+QICXpGUDIqrbwE
dA3IiPTdczwdhcx9yw7/LuEqVI6O/K67i0HO2n1rFcBdSkKaPflB6vEOzjFIhmkoUftj3BqzCMiR
XOyqiYFOnGk/3eh3F6nYyAtDbZXQBvEJXIzuVIBDJEgT52k33Rl1mX2NGJ2t7bLMkyK3IBlvDME/
htd0LBS6swAoA5KDpjZlP2seZ60BV2mshSp/UwTVY4LVhBMBN3jg89TcHix2jLuYNUjduMF7mRVt
QP3JLK/ykLGzVmiq4svxcKfXDQatuRAu9949F84oq0Xk8oogya3wH86LSVwpzvUAxbAAa8vC3BXT
plohqhqQFE4dsbohOXrXu4Vm5S67Npo9wnVqIe9hQQvmeEpIBLH+L9bDCBso4WD0MMFdSKmOM5O9
2WhKIj3r35NSsqjXQnutZKRAm2hNRRzfyFB+/grj5zcOwI3oGqmMYVNPnGkh1hNdEQtr93sArMhy
t5sDjyNtfBx1UKJYw9XpDcXITE496eb36UxFFCpLHj2ZzpA431aT2YM4cNq9jgZJMVd26XWVf/xP
NGhy/c73gtx1cD1bKZtYXh+Gjwywhw1Red2+YXwWHS8MEj/iew3beQnlmWpvUwI2ljXJwfgjQgM/
PXFc6/TN1AdoUlQvI82dAM4mA5xhmdpUd+pg552+y70RMHCXFNiY4eRrhnPmzijAzGsMJaN+1orX
vPCFD9jDk1BphBF+6Zo9pAqLqqJvUvJhXtli7tZ7MIxx6MIwcwwSxxGWshFKvr6pI1yxSbIHaN4V
xhu44Ui4T9nfRstnHsX+q3+ufdtZnJ8ip5GRjHXOKYhaUazhdbwMgfpBforhBiB37/QNDibGhZcV
BAokIdZwJ6BwDXyyUIxEzcPIQKS9GGwGoxmymy3+h3zDWyk8XmoWwjW0H03IejibU8S9Kp4i0rL7
zYVIzLYlQ8os6SOQ/FwHMYqpA8N0H7MosANXZ2Mc/5GBR1zwv79tRb5tkBw2nzi9q2cqDOMBRDQ4
2O1NE8s2Fc4B+/8iaF6iNzaFQfql5VPaJmov6G8JcdM//F7RahDW7ZHn1MGGtQBaiHjWR0tw3+hQ
tfYpF0zY9WtUujabYeGCfW7uad5angG02gJRqDxPAh7CwX/cShsWFqrwYjLg3ARU41Wr7g5vFahx
PyFMW+l7pZW+0Emj9IlEO7Kwe2Hd9ZLvBeq7HXNZ6n6HpW+XYBTbCf0m/533YlhMkqTp3fTVD0W5
0PM469RYIHq1yKi4xV6p95OfqE5dyEt0kalqHvcK3ntSIvB/YbeC2DM6aWl1zys6azef86si3bws
HZU3PT0hzlbJhmxPFtIYv1iZiVAMqVifHEeghW4FM4Ef69NBN/Eer00/KpnSLQDaZCmxTeviTT8t
a2ytJzLvBbhxBhOf8EPUnoBWhFWiEB1/2ERLUo5a6UeVcsXkXzo9P5MejWyWv5wrxxa3ComGSfy/
R1nGwS7RipQ4RUMlW33Wbir3+AqjlRX1SrScH6lY24qmd506n8ZBeI4OMvNi4SJWn9rmRgPToO6f
D3l8+Gbj3KadMWDBHDyjv8iYzAzP//JTTnTAwrs27zLxE17jOuHL1jINPq2TPjlm4VjPQCuLhB3Q
WL9XJ56Tf8pZsAR1hMZvFcXdZoAOWjbkl3XMPvueLaxrAg4r4D22v0KX3Ktuz//dohZjY6NYOu5U
xk71bU04kWOo7DWcEaJTygr69uzfoXYqPFx+kGHHAklYMVC19IdWCxjllh2Ienwc2qZhKoXhJwKv
JB+OYvu8uJWXUB1h1/f9ThDQ60XdjIzTy8TVdeSr+DnDSoPGx4Ri8hgZkkPBZnod6d0My6D34Ckl
jfqEUGaU3k5mr214cZs2DXzBLOoDtY4uZeEjIdT7OiUlzjHCfbYYOf585nQQFRIW5fNp3UJxtDDl
MhyOOFxv+Db/0LLO67jna7xjN+sZjGhwxwVEaFwxLKP5X/LaUrtOqt6yDxP9PM/UfHSf6uQ3mAZU
bDjc0yMQ73/vWrKZyKvY6Z3kVIlF14fAgO8Cj6/7gde2vJEPJSYJNUeb8zlrcHGt/YOY66JP0/Xq
25UjP+p6H7rJVAHObstMyUUk8AwGT3bp7idmv9cKMmLEm3rVcI6nAQFiFF+lMsA0Nu9a6/6FZJ/m
XXi9JbincPuXLV3xGk/yIhJ/UnAb3aNkhFXPDTdqKDd37tapWieqhdkb36ymxGotsLSQ8fpcWY8Z
/TWm0Wvh/SsE8IPLSsN/G1A+qo7lZco8YIdT6+B1o50sDUGmqT7H47/qa7shJmHd2PvQSBwSqMWM
McWGnb74i/ClL5WJsgUiLP123kiq1Ql+Ys5MRKcibOqom3U6+ZQ+Ec4PtyK9C/tjVM3IXx1QQ+RT
BmSVd6Y/SHGVGzKI2zUn5od1OBl4/mnbYMYiwS6T64+XXh6UxTzz32vbZpt21HkZ782iL48Sqs6s
0JuPstjAu+3S7nf8UQ14/IiKeN6VNkhQXyocOXKU07wN0GAYZlsWjNA/GNTLsR7H5DSsGlfQUzml
QTuPsuhCuX8qcxhy2x04fscxWKvYm2le5R49xbkVpGQLkRq4O5YkxxW68gCxucvCoirISVIC089B
FeCnA6cF4o1KYQTF/lkg0Zg4SKRfaK2mzKwy+QnCxGdDzDFxPUAaO4eFOqGQOPeqMuWHPodsTVEC
03ombRrVYjPdtjp/KoWvJAO0ZtYV+Tu+92OqsuiBNWu8s7b4BQe7ETIG1Fq4wmsJXm69MXu52pJ6
UNFbQFGvcAQ0O4SK0p7hNYJpmfowFZoiqyVyyChhr/NPruZCeYlvPwDL+Xoy41sOcuFuaJSOz+aP
Ac1yomb7cOZ+m8uysaqCERrKN/5mT4hQIMYBFNjawdAavZO/Y4+qyBPAceP5ipXwJzTIWyZmtX1P
pq+uKJDUWt3RSLtMIYzGBKi1SiFYQsnJdMepOrOVHjJe++hSd8WbCSoh3ZOcBXnYUGIREu29uj8a
ZGrr7/tDshGrMLnPevTQHr7vOOBIVBvNoTx6AdbU128mGnzWI02ADOc42Nguh/eDePxXNgYHFZLN
J/+bHP8/YTem0CECw0ybPbojPHuiChZpKP5v+bp0MdLqZ9s+FmDkJDf4G6//HTNWB0CKyF987xsx
m86pA2Kbbg/6HSC64iBab5EXy9HvcmBhYaFU2OAambjAWXXz74yLQbIntZS6i20Z/CyduN+YkZBs
yhBA91XikGaxlPIYPa24Mz7en/31NZyJmOxOdopSKgTyKB4ADThy65ElBPj5TlfUdsx/a3hrTnZr
NEpburN2D7zNu+R96tyII1lEKXfLe0BfVcgI409v21uqHFPD6N8FEQ6Skwl8E/g6WVYzZFPvSgEN
qE0QuQDv/x1pFTQnRo92SxAkYT7wmjKxvvIBF8D7zDafqOX/WX9HeorxjageGQNG/8VGeMn7wUeD
vejgcdpsXS3WCn2ErhnAsNTmDFpL+k52DQzWf1EHvTeHvQleLzfoJ3eh+bisnoq8GMtfrlSiOiR2
/7WBsLLV/WQw/gcKBFgtS6hrfFyaRzB1qEZFOjc0u6BsobdN0OYikYXbO+H/3fAKm2nBb80GiXQL
MydQf4v7cTTUVRR9PEF75Yf1hLf+OvcM2qZ2/cpYK7D9z2n+89IVP3U501smcENXOp4rEuvvHSX1
zPpOq+jQzSBLoTKdohOx29fOpKxUpOlMMVDW11NsdlF2xlLih/FFlfA8Tq7fiENxOZ48oC4MmFVo
s1Oy467g+3T4On8Ixa5h1FZbx3RfeSjRoFHltCec8txUA0rJojLdHbF1Qayly9ixL5wurP2eWYN/
UiFTNNGUkPuKvYxKowe8W2iHdtQi5ST8WbLtq4NeKEKC1bcFZdQgFMwO1WB7AYRvUwJNX19w/3k1
SmzhjDeDe4O+dU8ukLHTBgBZG54ZM0Vxusbu9voSw82TLcS1tjAe7wxow/xxU7FAnVK+gjZ3mSst
/agRW8QVT68O1mVivzUSzESyPzbuJt7KVrfKVqIRVzgUmSbW+3G/NVpxSw6KDfWf3nFtpapcSzod
Ffbu0rjvi3FcQLpzWR/FXZJ4338G7yYfs/nsAGkM5KVrBIrGsDnoXGx80wdFlNR3nTHs9yCu8e5z
q6MtKtAtyTyyWVIEi//Rcb5PmdOYG+aIHf5+6AoxUF1gFi+BfMV/pkj7FpenBQ17YSRI/osipBpD
tTHRJg0NreusLjOiV1xmWPHzUFYzbo2AKeA2JwYSGCVI5sJd+L/OeZiBDhjRn9Av67ccJJarm5aW
GJ/shdnmBaFYyVebVdPQ0ghP03Dzd5xGJOYlkmDwFpt5tOJBchhE1D+soxtn8/8aEs91oJt3Iu6U
Sb9LgajwVD/aSIk11NJAjJz59hK4Nmzu5FtnKjKhmyqA/rvm4Vt1Lqa2+vJ1IA7CIIbqP9rJPOIz
yaicDX7SQr9/WGFcnloeRqI4Pbk46rK3BsiqMsiiolJ7ghm0iU3ieTeB8qnO4uDJDNWwXHN43VpG
+0Uf/RiI+jecvNkNtiCnu3zsnu/tvlS/rhMhH6wu2UlcvtPThs8jfyAvRwWAHrjTN8XUuBbOkDVq
PAcoLG5eDgzBaxD7vTQ+Fi/N3Q6xIFBeaYmr3HeWz0G7v9m7Gzu0381qUgNO34jaZjeaI6/46CxR
KKFvpAMEKcyqCtPVJxOQLVKQ1FXDQLIPJxhDeXvcmczjakEqKL9vKt/5VPSaNeA8pGKl0leVG3wS
2fq8QTpjMQB5CweKxufGSdnSk0yAPiO8QTfGcGNBjCRva8/BgZDGCxuvyLABy9Fd42cgrICMatiT
rvt4z17HY+n0IwFboGYbfPMXZFkCwLO7U2vXUJtl5cxpdoKQPIu0BTvRHoQAed94sLgcZ4dD7MBo
zvdIw/MIT8+/YezYYWAolWuxiJ6xnad+Elf5mzstx/ysD8LK4qsGMDyWVuObGYjWuL3Ko0AY/ImL
ULKChvOLLGrWu0yh8e1fiYyEe+tlelZI4gLlOTSbVsCT26+DZ7qjw/Vo6ZBW7aawDvUY+QQ7F55C
ANP5SFBk7giUba+z17piNL5KWxEoCquPZRzO3NnoyzvwLi9ICXuamhG9N6BAk9abBLMTlcSdVaql
hVjv045ZXSXtovdkgI5GujSHzkRcUoKw/ls+rBIvi6emaiFJN4FEZ0NtWpFaEkMEIGwkfSzISEdd
W0bMGjlN0dSbN+2GjlcZRRn/BQaPmCyzCJgz9Q7ETxgS+Eq4iPHg4DLdQDECRnoU7i+ICX72j8Br
oWJpZV+vlbEx9TIQsinEVL0T9oy/G7qPWRq2T0bcPMnHS58300zZ1pfmtMPe5uVbwu5qQFwP6rQw
HBXp0dsXPfKeTlpa+Dk2jYZ6KgRxKONFNs2wp+my574ydDv4x+XcGsm+eoAUM19vKWruX591iqOk
1QsSPXRMwJ2Cwn3zFaIYw0e0yGmVElig08n9/RUsZN/u13Mv1M4wXoE2KxciCBf9h3wnl8D9AAqk
Yg4pWiXX74oR4FOEnTYNDdzYNlQtXS3UcUVFr3qyY216zzj6wGeRjVxg4pzH1WoFZBLZtZI4QL7q
R51fIcSQpy0w7yqUWWoULxe5kpkPnwi5IThUOP7TNQcywIZnSmSIoHpa+vOTTpzrbyBnbxycX8yt
gEkwWekxwKtF/5Qjordon9tEF5natqVtG+5uJAPLggmdppdziv9ZF+LY5oKsR5neQvHh8JOcfo98
HNXY/SC2ZISsjGJyKIh+f2wg/egtclQp22w2KAsJ/2f9tpAReQ+Y270tY5G4WMhWnfJT72oVKQYj
vzgn/r7VLgsXYvyFZPrTvpY+lk6TVv4KwrNJeaDNvfVJ6fWoqr98nttVjKA+XNsAPt0kt6Z+MVZZ
aj8idUIzDDBvo+/XCWo3vxi02NT+vnRnm/HNfYTkGZ1bAYVcbAPcFSUxsetRMqLqEXZhZUQvC5ic
TQi6iTrHx3gIW+Ezomio4gm74iVRGxPwmXZUajWDJSaKb5xOxv9YZFcLDJ0d4BF07HkwJmrjxhvW
+KOMNEbYcaQS4BqYoCVM0lesy9tY/oDQN1vqCynEXi8IUpAXI86nUYTTfBEv9mYr2WVfaHVGC845
YLywoPxIToXi5P2FuQgVGgPd4N0X03VYBRpfW9YlLU/aP9lDsDj65Cj1EBnHwb1RJIHBDbT+SK6B
xoG5UJ8cykvaDXiWf9D5KvVMY5Rgo8Ki045xIJwUvTw7aRh+UwddMIVlGyzeBfzSX5otPIKmvvX0
FFzQPUwmxcsV8ruAcHa1BtODJpdYg875LwvtmhrwAVA9wZrjO9AuPU85bQ7DGr6pqGT8kKDBjtA7
lIv5N/sneW9ypwpsG2LrxDBy6Lw/RmNvA946PEjLpoE4wCS1VaYARTVo29IOuB5Jd/2PFv3Tfy82
BVbj7/7HLJnSkp+vE4v4AUZxysK98h2y2Kygo6rRRj1n5eiDHx/t8DVoUwsiL5H1XfnSYLXt+e4o
ZVI+7lygnAOBK28WYJ1KFvf1oRbvgfHBYl2ZpF66gs7bPkvA0mVwBIQGA2kjOSWK+dVLiCRRfoGE
4SQRHP3iWRVPY8QGm+hwd7LwHnKviN3t40GcutQ9JQCQsOKUmN298zXkmakiD1bzWwU2Q/GFsJHp
P1WnKPpPN6PfLBeniDWMQsWXDPkJAzHfywJxJ+uDgoly89m71/9L1q3e8Olsz5vFdGdTBAR0B9JM
8GWbxb6U51vn/gGwoaxNpHaEs0JqRMwH1tnYFA0rZbrx2ikSAZeJQP02S8rrBImpNBEZb6Rqp+kd
kRot2c06OQJ4vgiWFnMTRIMa0HBsDDYvLtLwkTW8g5rdrKkkSYhrIpEW3TFuOMzk/g6e8AbGTyaV
9xskgxSmxBH1nYASxOgG13YxA/THxbDlN6T+LM0dnweuX7FsBPQ1kmmcHvDZQ3MPUZlv9rlrNGxD
MhAaylO+EcwHCxA83x0ahwQj6z9QeoKfJQ4dpUK1OUSVs+omsfrOUY+Uk2V+H80MK8xykLhq9o52
TxZwnrLafyzaVa3ynf+2EItHZ69i/pfeA2gTxE+SIOH9Jnq2bYps0ubHuUHcxvP3HpfW96/r0Ie/
bmb8QmBg4sL+q4t3PBb4NQmYkmNe8K45j1o5rOe+XNaDqV2xj4W+yKSzg7j9bf0MPXVw6tWZO1u0
uAcY1fPGfSCeAvVWb01wNKDhF7JH0ACEfacRcLXus1yHo88w4XP+0dEHhCBpvdrZmAiPfNFxu0b/
Y0jPzO/ZOssYGanoBpCe6kUd7/V50NDdRCCkF00SXILA5y642P/AnaQf4liXvaqIMIS+6IKxIl07
R7kMT9zzhWrr6ZfqsGhZPuO2rYZfLSWRU1gJ47DpVAzekGj4PoM8oWpcEeDDtTexTpWtbvirSejM
sXppDg4ZkEXAd0V3XRo9GTeZGsNX3CfQBsuXvKEGazeFLqFtJiOSXH08dbM5q4GsyaV8SwjOL/Gc
hZ/0GO6040fkjWOHAZzMEmCiwlx9Rbod9fD7Dj4q14Pb1fdorVtQGKBpRjHOPwKUyZar70Hib42A
sPHdBRNnNEbdxR2vQoIrQrFquq88eieRuJBdc+vURACsUXGOy/ZKymt0rKxj6+CYo2pmyjBp8u52
kf2at/R72q846FcCuZ+qYqxhi7QvS2gh+fjJXY2eKQ26qociKzF/da36RxQb0VceNXhaimt+Y6Mf
tw/y/esqpNPs+MJZJN1qH+Ozegw/7CB8UZ6iqxgyT4CI/M8N9TVmVIJUt50KMcNkH4pdDFkbaGSZ
UT6n++59/aA3QWP/zEPzxA0v89J+HEaU2YbVRp4+tS/A9U07OaQpYEu5uGrl5gWedIqxzhQ+mtKK
HffsrUNoe+EO0hd3Fm/s9ignjFr+U8QNHjkgyyAJwIA1eDEq1GhtWn99qgIcrYA0q6/m3LRib27a
To/zc19UOiIERtKmwI47Rjv4d8JBh0BnxY6IaxY7ktiY1zmFArOgCqVYk4ZGxXe68YSon2hA9tWj
heYbeS5HqBMat/+8Lal3j6CYC1hODIU2d0X8KkLQVrMXyAfDG+5vJFv6boKKd6QOHL0JHke/rAjQ
gBmgzI8N6epVJAArmhhOjV8oJigs+A5MTIGxTMYJwcM09jC2fimrpoFW+bCdbGL68UurCdB7hlyY
x0i8tTC4pa8ZopdzF40wEGM8yUQ+vBrce9insF6cD78Tb8cVSyAg7Qin95Si79CX0sQ9Mnbd0HYo
0bHYgnRaS9TQ8Vn/0/Pp+OV+L2lUK/h3hr8Xdr3sh8Df4HwQyuIu2zMGAUlwfCdLhY8pQQf5mkJf
YBpmQxSIUK7xpLWYeAHth7ScN7u5/K2Zjh5kYO+VsKsUZ03LeCArRmM+67UYTLIfRFDHWrvc5VU9
8sYrIteZ2zrWB2xQ61Hnm20Um64yqYPP/HZaSyJ82481jG5+vcZtoH2Pvwn51vT8Nz6ce0MYDERc
Ozjwo0Ya+zGkYfq+v1vJCypwM+zh+kO9DBNk+GRnzLHEcO5UROk1aj9zAenqBbW2GHzATHdSBIZj
92K8HYQehqfJOQI8TVilToFbIQep1sc0QJ4QvzNdT1Cld0cKUrrA6BH5MeVjBn2Hl7hYDT2w6EP+
laC3ZlafEVHHqNxVOmXjOimI0qqzmcmUwPy135OYXOcytshcHiu3oQi6M2O1O56jn6cGdZa4tC6O
hxclW1T6/ivlPxX5D43GVWz6KNm3pDk0ZS+yTRo1Q836IQVH9dkWAJkNUj8cj1zLnCW+hhu4mOpt
21Tg8RquR1M7O683o1uTJZfBLteRFAyi0a5e6VI9eUNF9Ek3p6Z3NwyN6oS7zhvhnZuAUxNgR5Wf
HNB8/EPq9C81vn6ZcM5xWcUsJIeslhBgteC1xhT7rnhE7M8JwPL5vCYycyirKtG4SxEE/mg4U+rO
8HKmw6FAbWpHMEbxmugt/eoaIbKeYntYVWm5RMN2jiITdf+xaBhx98+lwNUgiIFOgaEgqcUrJs2y
2Aca9Pj6cs+LkraZQo+slcmxul3gZfgcnuSB/vWIWepV3TCswU1hqTZu1GBP+CHZixKCuh2ZVKQY
oiDRIGlSWO+BVnNVTUUGBXj6sYlRZ5acaBbVjWPJiWd2opgBBFkPxn0EQ8isGEDNdm0Vfke55ZrF
H0paXQ3jTRC2byurKAf0p1E6/c3YSilujbc9vmR/xducnF7+qX0Th0Wb1Lwj+uBas8IUqo9fh2nb
+EHbzjt0F5KRGTNaiWwLwamr2ZPobwOThm3GhgyqT/guUnDPW8QcZZib1AStMI77l8Idx2H1KQSC
AQklAVUSMI8udY0JEPkls9JcsJKP4VKrmlIar24HFfLjXyi5tcFwOu7Wv987YidXML65gLk/siap
Dh6ZS2XjswrHOWuqiiqcPdkLT1XfR4Vz39RuczJQ6o1RffLijSh2emrlwWoIWDmktbzf+krK7Be7
OWGr5ekTI2chp4DUK5RNyxeLQo11HsiZ7NA5IoqAZkdMks8K9f+oYdzUgO25wOVvUcFU1s2e+7g0
4+awX2+H4nh4iQq8GeVhPaxpz8y2PUvZn42u5wBUG5TOtAldLU9VZ9encnEDv7JSMhcKdq/LAoBE
0E/vcqtP6qMpu4JUgJFEmp/4SHnbULMslTvd9P9aWzHyPd2LDsL651MghEbcI1cYbYCf+/Z3Ijhl
MdCWKCVDqk8mDY1RrMB+RwIuCRmlIoNL9DAHQLyvIZPKL3YXiIoZmmOCTAu4H2lIQk4d6SYgk4/G
BuPtynYV2+s1ssbYMVVohpFMgjI/icbBorSS7blrmS+CfaM6M+iKRzJwNKNtCDf6TStMdhV772Lh
0rukkEtMcQYbU7+lPsA9PaWeLgL/vJ/GO6cnIA7sfm6yRW9Ft+QL73iRt28HqsOdx/NRqtYU1p1g
hGeT/c7vk1V0xagkqTz1gq8/RjFYpP3OMorP3Cy//s2V4KB/bX2WDbOnnV8wTrVvytJDRHKpQB4R
Zr9IzTvT1y/JqosEZq+sB7VuaQ6RzbLKozwvEf1nc+k9WwHzpEaOGogJ0X/YSBjJkcvwSU/z1pTH
woq0cI2UV+gDQqPXlhN7v9BqJ37UhwISsoEkO/XhHL9hNsRVvmp7EGYM6sFcrlvjrMxX7tD0aBm1
08lTW0q7xCVcuW8C0WRJUvDt6tdAZWBpe7jc3eqQAyIP8v8p4stBlwGccqiW44SmQV5gfZt02Ua0
Z652sLTM+9zJu2VbX1eC/LIZyLuvcwt9tdfr/oIUTJYt3NquOEU1HCpwG4neV5AXmYX8UQrx+W4u
kh5nMAR1woHzPZzb3T3/kOtY5HwjdmVFkiaci8KvnsGqo6ORBeH/jrzzif7e4Hw+/FiEOW9sap75
gDOHYq3MLWtz5AUya0lDXOR3mJE1c2LA1Ari1jVj/Gr1BQD/z45DdAdk92YNfwgR+gQ7H+MUSzUu
3ZYtbeIr6M2L2LlksYTyWat/Zr4V0Z8n+yr1uIKrN9qsIiTriS62FsLzMoR9gYh0H//bMkQox7ex
oxz4mxgzHeHca4xkMqFvSEzg7yzBKtkTckO6NpXNR9we3OR1Zs0NTqRvWpZW93l9GL8gB584SbO9
ad5sja4nYsvKSvdh2Nn/5L6hWJEkutxEnXiH/Sht8cRCf1kREL4BuYhXkZSR+dxovFguFaKtlyO5
oiUuS7BSrfyorRYF3Q1y373b3uQu/JDX5hvV7rA+w9oi1DE5v4NOpC+2tR3LfBntFpfgY+KI4q77
94KL6yMiG0vOxhu9KQa9/IlIk9VWslRHmTUBPPgcvGtSSbac41+69egBLRZWh7kGE5VrLythm6PB
6S43EN44qV0zHg84BotDPoYw3k9Ib8g3o2coV/rqOebXE/rBnjLKu4Xa3p/W0rxBoi7EB7BomWR6
JOmvwt4FfSEA6ctpyaAMFlxgunakmCYDnBcCQJ2vEYd3xi1rHFgEEAZKb46XD0+hb2OwvGZT2zmf
U7ZETwlB8QBVAk5Ip4ao5M40NkM75b1auU3zMqVQMQMlCsq+8CmCd7C9dhaKlgK+rwXuVjBGYT81
gRL88ySp/QgArBSZ5xk2O5Xa+2vPNDVN4t6zZFPvbuGCFdFKNh75JsgoL6A9XFivtaGLPVhaYDtG
pMCe8TzTP/jduiaiyasVqBBbyEcz8OxgCIhWAVdgfvG/OCiyGS34CoX1PxhpWErwb9T3f64hLNmo
raWsxUU5B7icYusTWzEq/iSKNAqjiVUp/PJYBwzkrhcBq876OoPChT9erJoQ8VAq+nRcz2/Ty90/
KSC9d5H+bcomlhp3IyOO0qorKZ0t8czhmJvVbAtqrNzRGfYOBIjuXFAE7BzspXwzUcAhZhTbHqv2
boqQJw5sOG9KYz2PhO/SheOoVWi5irSPKp4RmS9KZHEv2s7IAldY6ifZ9NDXiIyNzFjTjDk+t/KZ
2uGGtkL8zXGlkThItgbYN7QrXi8GGi+UgKnE08SvoCapj1nyINzfLiP+GcKoygDUOKmql/uHE/GO
6XR92pMa0K+fRjuN/KwvTNmex84z0TTg2ZTsXJVTzb2dFLM6+RmrugY7/gbDiuHCnqrhf0zxK9OX
UXaIA/zXbJv+U5OdnrzoMxxUM7idYZXqL6gYIPllVLWaa+AOyLJMBHS4t1uR09TVNjKvIjTBjxFE
00io3mWE5er+jeFXldkiroFx1WcIgOgzBnrNjRESk2pJrLV0M9Vo60IHkNuwmNLdNWyX1xdEGMV6
NZXDggJS5bx2F/16is7Nraiwgxs4FjqXtdVqM1K28DXe3AR6SZXV0NQc/lD7johjKqPNTNonANdq
rx0frwBmHFTTkGcYeuhf60F/GLh6tjvps8y5Lcthue3RVk0JSEtJvlsWXs9QeSlf79tR+hpdB0tZ
jDgwvjEtiZ/GZ8ThP4kZ836lwIUQNIk37BM0EUQJ08qL2QQrGbncstWM2bM6pcpauJrmawAxLUdX
SCZl5C4HeOp4HclsvrQsAtWv507Wug1rrMX/szKsTen+F9f7BK/d76hzno5GyIwwH/xKmRuyLgyP
MmSrjcxZLogMXuasemKhe21E2hq2ozj9TMRYJesY9KaC5EMFT2rkpMyyVk21FZP0cjUMUwrpX+2o
Jse9+rnn5vYm59pXgqcrQOc6WIlrlfvnlFrbOMbYbhzXseGiB62Cnu3hXaAxCj97x/6Sg4e1secp
V74NEFIT5UJhgy7+9dtJ2Ix6apsDyhJirsT/JOFwzD+niX9jSoMWioylmQfBwt7jj//E3K3pv5By
yZhwr6U9+W/22B/sIkKzUb7coH1BSR3C6rzTNIfZtj/OYk4HoRZB0A8vUyMhH1tJs8SSftHhCvdP
krcb7F1ct98PT48GsXqnarF6b0hhUsw7EU2OTd3ksVqkqfHX4ElI4CZ7ygFXm3ItNH8TbiGgro4I
z5xpRNNOqo02UVtr1o/29FZFnjXW8IFHAhjnWezitaSB3W5jbB363AYGMo22lQULTJTRdAEvcIWP
t1Xpo+dWUv7lTl+slpyhWCFDz76Zg6nQerJ+t3F8e3eLQ+tM2gfD+aGLkuTa1u3o8Y6ecoe6lzbo
5YlRjaoEIBRr0UJppt1WhCg/zYY19je6o/8YUv0WjOfAlDJnD0vcEpqZ5RptD/6j3x95pIYY/VHd
c2sDmTZU9kbL45NS/S1GtSyWHxhYwybSdT1hm9Wxql+36omV27YyMyXFlYcPRQ0f45kTNbcZmyoW
CzbWfg0hjDqTxcQca7tQ24i7iT8canjleR9At75yh9HIGA10zkc+scDfztkimvxGculUI88WnQxL
QDpTWalyO8RHW10CiWOY+gzVx6yS9UAMLpNm/yWPUqHvjTWTWh4G8KkA7c7dVmpiWsic3EKJB0HJ
UvloV0xKEpUTe6fRreQ/HzuYtJu+wBDSpsZ+LKflsuHLuLPXjuwCVC0sOaT8UxSKPpC67lRq1BUc
R7LFcyUBhXXL49xzYPymC9PecKqYGRQEU9bxSghJBsdS1BI96sr+I1gEgzUNArvAj3QpHyZYafi2
/DoYEu0VlSsOhmuoyvGdUZ6Io7fqB6a6Amzr8rwIa/Wdl8kvcvwtNip9l0lJ6j9kbH5/LHBzICOa
YM1fa5+v/rVi7F0lbVxsZVnRQdyLPLLSO39qdNYxSAths+BP65otOteaw8caWiBbD2azf9Qj6FNH
7+2+pmsPVEnlArQ8/PU7DXcwuCpXhjtvN34ujnH4mHpNwuHWLEZ5ycvAhg6yFXYQ+67RNsyPE+cl
C5XXweswQQEY4R62EgDWGvd3cKEsL/i29DMlKqSrCeYSAVR2+Y16/QWkQ+dHaSeWXl7LltNpZnLO
zMkJGnd6QPYozXOfRRczjSa5jPG6/9QLBqDcWd2lX7Q9a7yyyA7UJgsLKu40mxebqzTW4RV0nW8o
QsBPkW1qOqKBWYW4quSk4/YiF1VHdX6yk+Hkul0bPvmFCt0/mYlcxIPbc3qkIhTB3BUGx05iQAVD
dysUALIlLl/uV3hZVWWMxkZyGcU7A+2lYTFB8GHuGdpyt+o+MpXVzrqrESVrBSR6hkQCYf+3rV7o
0HSBYhhVzH0XjEK0uXVHOa7fVx4OXlsRM/fmJs/tx30Lj9fVjcKnemgLwP2QcjTcNrxmbEsu+rhY
nqhC44MYFS7DpUwOzFk9fis4P/cTHhNUO1mraA5FyEZI2J8ywfOuEdvzVWEp8wl+GZKYnLw9rpy5
erCwJ1MdROu5XpBLHgO91S9BiZawVls4cnos2Wh5nGaQt0TzrQ7poL6NZk8nFO1o/VG1gcfSCGCl
459J8R7x0ANnE8KhNF4NOUEMWXm1RVnGVqnsGcluN9/aPXpQa15w2JCHDf7ZNA7Pr8ZYM4ODRgLB
mVoyds3Qv0YFVG0mcJaa0FOXN56Djn+4qN4mB2HtZuCH6PGDzMGU8fkUfPDEjm4fI+5QDpcA54By
syFe/U3MBKjUs4Slx1fNN62ga2W87A30HqfhaozU14fq1wnyNlcev5lEJOUkHl6I4emkg4yoVSNz
NoZDt+lzOpuorVshXeJBEO7PgDGmlCs5zBwSCPLx51Xs36HDRUQa+ZAOiPppjKjbYGci9LYPA7ZY
NSuN2rCrNtdWjJO2vxuedr06EdeC7Ml5jXw0i3NtayMoUyaaj4yO9jKBc8snMUpTvN1ybFH68M/O
9qwKpSPogjdmkBeB0sh6yllKFbY2CZmxW9VwS0PnP7oI1XJmzOxGMUUAJd++1fPX5HeOQPRqkpxU
Iob+uFr0hKo6s1FbrRxSM4MsVEy88l2AMj3hCRjpK4w1FjUMgKD54S4d3bCpd9xVYFBGG/TJeE7p
MjAr/kCMxUjlBJJ2gKLq+pqfMtvZtBlGogZRDLy7kydhr5cHWjUui+1Oj2CkyRxMDeQBLnVPsVqz
dwOX+/EvJlNMnuompQ8IuLmXFLfLyI9zZOVISYAWcEzOR09YEVNb4fNWOyAIB8vmmPgFI3sUhnB1
SqrGxB61uJls/qAegDGnrXNkWkIKmmPjWXIduwkbsN4oyJpj2aeJw8ETt3gHMcn+eP8fbEb5mUQY
zwJtz84ujq/riIvTtO5phR/IWLD9RNWaSo4+KVSeRwZ3Z5u73dkYorCW0J19veVcxh1oeF34Nra5
8t0HH0YcGgn5/hOOjsyhCjBfgPhOQOhvUDXRBKpstiysvVmzUb5ZvOOneeWoYIgepCR1XZgVD7mO
98lx3oDQhRpmtdG7rUFycBOKWqKop+1qTdYv1/9M3P0gUPOPtfAG4aGC1SRN5IcWk4oz0Cx6Bw36
55YUjXqTwZ9eUyn61Z7uUXVSysM4uYEVHktn9Y8Oqhl9yedWgtibvpQb5qJaTUmi10tb5YYdctki
Nnu2CrIYd2Ki7ZgL1jMk4LcbIjCrVerbxACwbqFPOpK277XIvy3m+nbGm+9TbGMtiztvnyAEx985
4t9NYBpXB7KFrO/YmBkZZUkmHDobh/vCZXiepXwYSykaV7WrTgYkpj3Y8zlbovBnkMS2Pa1i8d9f
63JtD239Gz2vMtD13iISgYBicwlCk1yB2xU1BDVwfVpFAQ1s/g1pK/38yyOCCFe0BtOZ0Id9BqMu
I6eO6tMPVxCjWEwfSzTuiToI9I8cvXyvLF+cGGoy9x8gPuGdSLZmaVqDjm+8d+ApZT/iDIQaJg7D
DZKGlwphQIPMhBIZ5tTdxnlQrnycW7+xWR046bUtRE+L+S0dOpT1n54eiwwqDJtlaEqAH2EMKKUN
dB8CsEjapQJiZhWvoRtaxIXFxQS1jslbEJl+qoLdNBEmff3CdnzRLxiTXrOrKEYgxfzCNbe/yKho
4fGLHzzn+vZJanJV6qPvnITiVmZaz1reMGkTMTfJmDPA0fVxHcgXg5VneDHgi2VDxRwUxFWsdC4O
VmjcAhIJ6s1fil1t3Er8daR7nk0mSq0o8raU98eF5x2bp+y2rxEYt9JhE6mBV1cFxCVR0u6Jwqsn
Bj1tX7daSlC2rtInyDe+FOMaGV4ee1qmZVwRVSeDS9sHGepqqWLIWhBP0jW8yxCWP15IJ1/eMv5G
m70VzAOVbSCqpDrkdl9HxY7jZUnETGk5woPatogBJGeeYmlerVRTYnefQcgYh68ennQxtYRIR41j
Z7EH55rxMjRqDl8C9y+EfxuPGJ/pmpAa21EmxLVB6YwH0T81FdhUAfp3ml6VeXrKOwHMG0WfkM1T
t+lQxZjYmwe+W70AU+Pm5ahQ6j6sXXz/bjbJhNLgxMykFOHX22hVs9CKK2VTtZJw1EzyUGJmqEfu
EP2ZGAqa2e00C3OOiP5ho7WzmsMpN4F++PnKo4TvaB0dtp8/t08uGHCG3KicFTB2JgyInLAgaoAH
rFuqyRWDGPppTJmy5o5eIAFK0gncH2E6oPoF6AgLqI9r8YXqum4vWqgBb9b1LTFVIelVxkAZkS8O
6IHnHzIjaIdEotEulHMJKVwHBkuwqzk8Ydsc7H/N6IkjG8Ejhv4KP9K3zj46XZmIYDPpwhl+yaVt
OKiU5L6kgIBZgWlh67nLMYVp0F+jMVTKcJh/76LrafNVygzuneU+6FTDtU1omwukFWOFrW4qVntp
xe8Gtr3pfhnZ6DbU0bKYllyo2adaad7gk47cSBsn1s2ePBlez2TdQmN1GkWdXadvBeE9HsIXR6Qv
LZGClcUq4HzANPnYtupZ8+bZLZJkcW5eJtYcZD9hEBdDymXTm680JcFojKSg2zpz8txVjkqz6tfp
tEfttQ9WGxx8uZbMHcp3Fouq8Yf3hE/81bcsifGJwiuTUZvdY6fOCQccuuiFVgi1OTjqqJk1LS0b
LbrQdb0e+jM4u96s38hDLfSVfYWuXc6B4BnWomknmpAQb4nRrfYo2HihsBoa4jAdODRJDVtYkVDl
TzIajeeLzdQ7EI1rRNnAyAXjvO8t+psD8jxgjwlUJRlJfykRZheKsai3+gXIjLBxwbgw0t/WTCfc
gdvGDyi1PFjgPx2ZzEkuafP77A7Y/vgeWjoXNcmaG5n+U1aBT1ubEvR1RDWsosoqkoCcJl0GbGwQ
DldgNc/lbignapfhhg2MCNVO5fPhOjPPz2dmGQQ2Ybv+7nI8mYl0qhYYTfFIe522hSKtnM1jOBKr
nPuvg3PSR32YEfrZZIO/p+lJlxl+XaZ6CTJcJ1Usk7VbestGaaaz0wjNpMhyE2xxCmufGgb3yZIp
iagwJg36HgSIbL6mFbyi6WrjSWWVjbYC+JimAdOHjb8bVZC4sleYyeEKVhl7aioYq/LVZkn+VM1T
MTCLbTJRo2aPhsgVLC5sfencoOCleIXV/1/cdvR0O+rJ9amZm3q1LXtasIvg6Hz9GwIBMwgw+HOS
nuIxxHFOjTziZb8jfuC+OpeRiOAoqf1yWdLAGo/aKwqrYk6Vr6LZzP6cSAEeCVmuLyQHucXlUou3
vTadmhh0HKZ9GwYX/qE0xeoxcZH+Dlzd51IANw+mW6AN9K3pXdIO00OmKsIHDy8xTgNclI3fVIUZ
dE71O1pDFjacLOqtNYzBDu3BI4DiZv8fEuTrdPMmegh4pqnXyL2Cf29wVtMZgf6i3apKU3QXJbmR
q1TOg8QePWoLiYPE+0bO4IiS6F5D5f5smTp8nLC98UtYliDvhVpcoA03Sbf6vUNPOwu46Ioc7127
6yYOQ5dr8BM1Vugz9e1kfMQVKFUmigto2s16FSP8G9m1TaF5BxXQlAGXvJrDgIdd6LGmFysi3gmy
sVNGPfCOAeNhXt5VZz1bQqfiCZ0NLAM/U04VKiQcPyVgFm8pGkBasECL1ehSnv8/BxlvCScKN1Gf
4i5WZNoCSh8HitHv6F8I8y9iK2ZNbubdLMqQNYmr/j0Ohgx1/RW7lwFPQkfkjcbZUx3p1MDS5Oby
Fwb7i1w8XEbLOVgfv2e+73mFzj9jwmyZlE5Pj6i6MbCUdCis0XadVlFVuMF13HnqRodeuhhIpoh5
yro2vJbzLSsedcPu5nicKsIqA2mRcp6j0u/RR6rC7M0jY7IqiIKChVqFeURdSeKDlpcLE32hQnWV
mwP2OCRgY7RbyE+adzMNF6M32esX+7TbIMqUaFt0v8hnAbfSW+oSuJPD+YKYm2hPBklywx3x5jXG
NRsoU2otjzWF1Ei4cA83lOnoU386WcpDIYfY4WNDspv4rz5rd/OJlPj/QlJukYPe8tQG69RcoRb3
AvSD2Hy2yRMNwuTbKVEz/KE50Z5ncns3cY7jLUdCkUsAsHZQx39mXXtKBB+BKQBJTAA5krPFjMxa
lHredGnC9UV91xQf75hGsyD2RpzoAj7ItBHvCkYpXQz5FgBDBqofUN8aCz+aDieVNXEiqNL4MWJu
rvIw0tdQbrcRkLpRjdUbg/IwOiiBLP4yEYGoGRlRrqs0jgpp+vy8w9yH1c3Lm8j+zW1qoiJSsC7z
0S6ripD50sHjOm+lEQg6+WFawFgE0vst6ZPTPlB8CiguvRU3y7sWXcWTyfxdU4Y8MDpbJY3tpBTa
/L/ta7Dv0SzCmI3GNi8QcBqJqnmEr848+uwU16/9zh0cd1z1U6Vuu5Ex+AgAs88j+0BbmIJg+dJj
NRWgZf+M8gSHhJhDBi9h05gvpEdiltRCMCc0SQjAUKMKDQuNcy3j9sQPLfqqfYTM10uJr1kcTycv
UBfEd81REXeoH2Xc+xNZP2nV4chu5VMM07un6/vNC1267ZFdV/SCrqf2FNh57eQ6nD7Es4k9SDoV
xn44tf0pPcTIQbKYtG+0L/YI1W/j2SHz1DVNNBwGdg35Xicy2p9gphgRLuuYQ3T2p9KfioQDF8sa
ogVFSLGKMMsK+f/Iq4CljgkxdN7wFtrZQvjEtBl9BTk+TvTUu2cNR+O4Ot+Pwrne3MJCxOOs3P6b
cRooigIvb0G594ecbfEruyEaVFEwHYpSEMBRxpreun4uYSM88h1e+BCnxugtE+ZFkeY4IYrZJZpl
VEta8AvgQtLzUhvXVzBwaKP/vNgtyFfh3aVCCLfbqbUcb+dVuAzUKUoJ3bFXYHFBWXKhQ+P3GYmH
uJ6XvDF6Q2b4ePu6O23ZQ+BtS3NTJVYpCnk6YIWMjaqT5TruuXxrNad/8f/3OcuxKmfYhwgIgYPL
K2S/zbeSSwoSke3rFzBQssUKFqda8RRH/mjPoHiqc+69G3ivOrLFp0Fv1Pg6qSK+kUHQZRpWDrTz
M7O6CFVKJ0c3o5RMcWRKPZuEOy8zY6AvgF3RzqXGniUqEvX6FXaGCL/9ev9sdmt8LpXkGHBe+Kz9
g0J2xmqvfwaFqvqVLN9hBlCEppIPkLXNCcJRpBsBlRrHk5HA/b/xffD61szPRjW/QlZENCzBHZsG
ytDCLSZPEctArXnL1MySr+xrTW9crl2E22O9sW15Ii58+q8+lPTbX3U1y4ReBxs9gVJM63Rl00bK
YXkHaOK6DhShAB8jUrQYPQ0a9tXre01LlYL/dcVBqtBjm5CmYeIp40sU1hlHNiF1RcnXbkVoyccZ
ZIwhkUksAl6jzT3Q2/L3HqC8n1DjWzhW5S6QRKm3ZyLULmANaKhHS6GNP7F65I7gDO036a/txpIT
fCZJmN5YdgHRnRsraCZxoiG0PIUGdVOik8hrTLoB/AsmetjzCpvA5e5ZOBHeNVqReICR5z/vjsNG
dPBGd92Hv7aIWLq0DnSLrkcOzhBAzhOGmj22GKkocElJk+T78UVzC+oHKzKuBV1dbOP7DSX6xJkd
0FxGqv5Rdg4O8pNoCXm2h9M+erEyjJzsceh9yfPp8PV8/gDfhFcv92T1QcaA+XJcckZigbzV3D8i
OMYceWXYzvDxczz9ZQaihWiNh1vlqQ/mF0pS+DkSKTBTq0SQJNqVAszz59dfE0AkdMkql2tI5kWq
+b/i8bwT0TVzx0F/BKUsqjDsEFt6CFIEA7ytaqg42g3imMrep/D38jYpqdPe9+1bshEtaYP25RzD
VtaoJk+WoiGtg+/Z6atE/0DhGUk2WfervxOIJ/tx0Ikf0lNBebKfMkuPc9N2HF12DgzJJ3rAwTv1
SpXe50HwX9BejPO7Npw9vfmEdRJ/J+4AKPBZ/KO4I9OUQCLy1M6X0MIOqA76ohVHwVMUbGYWVNHg
VtKMdPNFrsxyPfN18x0IbtfJ+wMbBFJJ5dEAYl/yajilNagByYdRkQS4n8pcTmHh4DeVeeRntrn9
SmgwXiU5YaNvEHVejNPL90WoSWGJ1w7lQ2+j60dlsNud0k9f54ng+kPR8Y89A6BVWn374snq2+aS
//+Gll4exTYSQkdQI22RI8d+Kt2K/wDYF6dtFcVfTSIJEyJHQYHAcHbp6kVo5VB1IijRckGRTcWA
Id5/vYH9T57iGvXV3y/bNyXuwj55vVmhAZJGACcwmOcY+gjm2OpzqBT/TJXyRzY/9ZIZAozQV+Mx
upG8GdPgUVEOBkVPJLvl/jDIfYaiQ4FAcg2DV8IXJ7J5zAG178AhrzGZ1jysYimz+wx2A6BmwT/c
yN5wHlNtIzgJ+NYkQ7P3Uz4dnuGg2HxRdeOnIspR6OjZkstOkdWurMEOEuJ6Ica1FttIzTuJ6IKD
QJIg4anwQWN023T+Cy5KOh2X79MdBadMqX1t9HWT1ItftZyZ3QPOo7O0+n8IQuvdzNVCJg7eQeFl
Pgdz31xADkslbZ5oeAlWZPUVNVpTAFRnK0WHvpRm3bJnXwOwEqX9Vk3P19Ohq2QsMcvjLaax2DhM
KvTtYQrdkG1ektGyu1iTpFZKN8LL9GcpH8KDpo2MwZwZtIcZwz4433FIlaIbXnFWu3IK/qAFJMrH
diWbIj/znKWo62jywwTRNicg/DO2BaLtp9GIdyyFwvwHH2PJJee0d9bBgpoT9O3UgwEPXK6obIxB
LSE7eMm+4zdwGwz/VWEkzzBrhFYbhy/0B5kTjS9cv2n2YWxFqPsu3mf0cMfA9q6d3YL5GY8f9qFp
a7wNtQpTHIZVhY9H3Goou1nScoe/AwuIGRaaOvRRZg9cEHdT6Gc5umd0Gpv2tJ6PPlT1Wdl3Ex+H
4sOr3o1LGLi3f3h1mWWhe8e1LaOGLOm1nn8Evt7JRvFRUDBcbHmFu7oUMRUm1YvK3RdrscjgRfcP
4ogLXIATwa5dZp4TgCkW7nv1fmjSCi7Ynpa7Bv4nJWuT7YR+zRZUwpvw2OAyy86y8G15fdQB8gvU
4wzlqYCh6SccwJcAx96KzHiTD8UXjm/kswSea/Kk3pQj0KjWASwhx5qK5xU8AyBUrUDTu602KrvU
mL5Bn+6YvKzW/RuQu0V2bkBmgdPwEMv8S4ZrS5RX4uKSBnrM9XAh0JN8NyvqjLMKBvoYav+MGB2z
2f8wDdhuIaisrGgpYOQFZ64bblKGxXBQZZpR5AssBo7wIk3LhIhU8kUmVvk3kTRPLzCfCrZmkCpU
28uKUL9JUoqvKaYjU+GiYVX8Wk21GPOgqTx+PHDhpTjMAoqgzs19eQFZeWSejYnSKUzyYYclJv9t
85/OqE74m5s+NoG96g8ZIumx0RuldMmo5vr9beDzP6B12ThaWNOimv+wfWmqUSxMNcoU/B/v6gPK
zLkXpoJ/6LS8nGFPkdLR1JuwPebC1Vnye+d00mR1fwAGTHRh0s5A5JChIk/53E//dmIUuOSzLcjV
BOdPhUjhiYYsA8a0R1EikQ/dYjpTSUu7vGOoPzq2bv4Ur6u263JQDHXB65/t4uYj1y01uc91g0NO
pwIdpkfA3Jf9azfMZcC9+VZdWuHbrzS5dbnVVvCpTJOXCISK1MOgmquDEQB0Mg5PHC3R1Il6QR7c
2e+A1ritJ7JX3gwpuBLH9rQCrAO0kWpjxnxEtmsoKGJaIgxk8ZnnvSmA/MjXhsxbhM3O2en9wp8L
U1wvvKZJjhYqUdYWH+bAbuALK97UVLicbCrTdb0CsialfgfpTA4ryMU52z+Dv3MPFgGHe2KVCW88
qgjId0WH/R2q/Oq7ZuMu5hgk3EmegzwTrQkbQ7yIHfG7XCj3qQMdloU1DuGG4Ej4zMCJG00F1cBv
crC4Zl6A/LWrofa3vg0Zij6HqmCpZ9RalAh6O2E99gC8jWldqPEYEUVKju4Rx8h9YM/EYRzRqERD
sJ+6P7SpzGwIFggCiqWMNNygGA4pDQ+Jg9M1c3QI4b/64g5BPPI25e3mogqEViPERmTzjDBLcxUQ
Hz5tkL/VArCjOMPhVnBPk3ylQEzGNJ/OtcNNL3IFOgxsxkOHkDlDoo1ukDaENMuHoqXLBsvx63Ah
MTXzbT9rM3BZvMRnLqfMOueA844uXdIFjAiN3lGfEsWrZR3LDTkFVZRrWc31RnFkH5GyxKrl4Xdr
E/fYLetZiqN+MQFYZ6w9oynxe6UezSnjf6RYpW+tGE9DLFs7n0WcD0nPpPUuIpJxLTo/J9eFha3w
XjsSt3IN2c2j3UB38CIkx1E02AhvQBC0MJV95bu6nm0daomE/cf//xPkisqRCA1Oj4wfH7TAUVwa
Os3Njhiopw83YQYCdVujHzdVzKbqaUjIPLX1GHihargXzf3iRMWTsGVqZuj55LWW76ArYLyma1+n
OsA7GJlYurWGkppCPoJMRQvafyqhkyKig0lGmJmeZFYF/VaHVXIHawmC6yJ689J8tIfe+/K7i1zb
qThQzi29J1z3vx31OJtann4WnZVeqJjLWkJCHSqSGnH1sZ9d9lRxMme/VLkmZuOtGvOGqQszy5UN
mCx5abSrojoQAxFbPy3GxYW4xGpYKjMmYxmOBZ2WNEEoaU864TSltbGul6rF3tFmMbxRwTeTI/HS
tpZMVWsXLqb0ukjD3kX23k40BblDLb7HwQBJY5pRknDgZGXAxorkeki2hdc1b8V2jkBKYZnLIJwf
UAjpZoCiIMR1mODMv5L69XRGOGzzMAPmAcoRscx0hw32cWS/A7MKBhDRDfWZlW/enLZ/688OERGf
JewtLPF6BArl1T6BszXGYS9PJL01XpECo0CZZmb/zICVE/1JczlumpgPDIGkMmMdiffu+qRNx2ty
3Pz+ETUa6AuewyicNgI5b6qRAi6HrmU8P/TkjNaZtdXbhEHpjNkiSekVYHWZxXi6m719jyabm6xM
7Tg15UjkTV6A/f1RxJ4/qdeuMtRJAkS31kaWvFHfmvo0x/ciN7LItyPgrY2YoXwRQBGN790FTqFc
lxUjD5T2l5/VahxEkolwQXM10vpGaY+ojJZCQrWpv/jaBGe9D9giJOyXEhNAhevDzj2BAzemDga7
KkQbz4c8k5kKoDKNombJ5wNfHpEvc3oQS5dwysVhblOhXcTgw8Z/hy+D1h61qE51aBt99wIldmi2
mWgFw+kQnevU6VQyyDXSWhpXHOqzuiXZ5Lo4DK60fzyp4VUUcQA4BoUmfvFqvCQrR2ukKQB+Jkrz
XVvJiTsvFfBF0q6MzKd8ZZAHlqDp84E+mbhBsRaQhCjobZV+QFmuqdpqULEgYX25cNbM/H+Vuu3c
vwkynfNxQ4i299OxSnolyR3n64f0YDD1GskWhgOgFxaj2lTSgKbsEhZJ77sd8pjIT1ZcycF05M/J
RU6Uczf98g7A8HRqgAtQM4XjtaqY5U6TMy3YGoaxp9dOJ1nVHqY1yP1sWc8tXmvJG8/rGAtWzk5R
uh9P/olrdv4ZmIDf1A4qjGH+GviibJscPEmcS9RCr2Mh65BeiL8/37BRBR2Ukk8HEepi+71wXIvY
WgZJW/ZCZnAmvGoX8XoLriTGdW4w3uHNt2NDjZQJuBWYgUJ363v0AZgKyGF1t6LGLuyuJbvtYfk0
DgcbPQkQG8oU5h4gsdjAM1tBUs7MZ8WmHp7JJCkkjAs7xlNoo/hsSWXhfq2igtDXnFp/3IC98kqq
+zj+4vn3rN55t5CGWdt6IY3O+ZN7DkZmNH1jMchXzcFyjlY/ONmlK/jN0J2mlUFCSpNdizG9OqK1
K5puR63PMi1/56qf5oXBPQhsEa7Z9BCUHc+EzEbRdnBwxU5qCQzcVgq+bb7LilUsCboJxvGbTvKY
E50fKq7e3+xNI2Tbt0OkbwCigU0x85nvdZXIg1R/pOhPtPjJczPf6ZJgRpcY+kpi2H/r1fxDVttZ
r74LaW7DNGFpnPD6vTimaPG4gxcGdlFrsqmVqtWDJ6zqdRVQrVnQuTP9LIou0UolpoHFBv8YI4bY
CMuf4grxHPvMeH3swoa+rZ2Smvv8snJ8oeLNdoGrcJz5qRPz7xYbhHe2EQsokfudk4J3RGMHXN4l
CtDjyQho4VExrUZy+b5u8kLZ2L8NisQM1d7k2dD2GKbe6ubDr5gBUzP3D/HjdlwCXYLuLHLB5uwJ
FIIbaYZ4zr9USjAUePMMYXcEQldL0WNOh9NskWIuv3pjWVbT9SiJmXwhUt0RVRSydvm/m3SGSr+v
8cVhFNDfGbKyIq3BZgdZksFf5GUu5H1DTrB64v3MiZrXpihbfAcRE+/LcdV7PN9sTC7JHBT4QDAn
Fi9ke5aee0vN4Da5yeJdioFoCd/s+akRjKo5Ys6764+H32uYwG399GobtG9zvLkqGy+LxDSkYQPn
0WJtkjW4FNw/FVNleqTbzPuiyGIy8lQqT0veIJc32wuuS73NyNssGUhBcGDGgXZkOoFQtdbAlTa8
pWILyaWN6gWag7i219FDJqVE91oRGINlmqurI6AqtC1jsTloh0K6MAk/+9WpngQ/Jn3/OVy3W14I
8OHwWvo3eDm/Mraj9syBEFmatBdbK0qGkkUyVEk+Ff1ipOGdmQXdcL54GlfDzdQ28VSvfD2MEyTz
sKn4d7aVQOU49B++0N47KMOkPtnm62eGk5HZmRbZF1C4qzt2M00O1Ikz8VTC0iW5gkZC629Y/MEt
+X3eDAI76EaXOZ87H4ONB45CbOjZQu8EIcm7ICiK2RqOA0/ktQC+jPbYpGza8rohrhvglRxNB5cp
EtRrVkE9+TEPsi06dIyybXLRenU2sW8mKbyPfEYPRIe9esgyKzQ1Aru77ybFnfO26qO6CnnXZkRt
RNwvXLQREhSx1nMNyZx6+XAfwYrAsGDuV1rRGIk6unXJJwjLlClmSxiHUuqXiggy6P5qxZzs79PE
j+9wl0uf1a3WJEOgDIdgjjFtrI/ZeQpu21VHBpOBV9swOOv+G+cTCpso2Ai/Z7RYs7j+pXl/M42f
67wdYTqlLtv5Cgx9NG/h6JG6NoFL+VzE/zCRN9IZmrskCjKTbjdi3a7lIbG3LOU0OEeAn/cZfxss
t5NvM/Lhy0RtaawLoB/icuQr15ukEAxnzbIfxYwR0RogWwLqY15pyJ7v8b9KGJu2ILyWLS0uU+EM
PtyiMQExS05s8m+wcmxJdL6N3v+UbbiX4F0GBDaF1L0NXd5Kc0XGPq1FSxGuT5XU2oFiSsgRsohK
anFnBGzVgS+GBKf+oOn81snJxxDJqY9n7meab0wDHJtbeNuSa/yvIvl0qLEpQI5JStwwfDe2DtKM
X2hW8OzdmIqMB4fMAfucCBUvLGUlSf2O1Q4nFp6XwS+cH+vPjuB2KHnaDelHbhHHNc4G0MTmJUt4
e1fjAoeSh4fR67SHuYGwdJAVVFHkjQaqpOo2paM+wUSoUve9V4XfwPBpZROneX3IMm11iWPCeaAH
ZltCMAKEEIn0ZfTl7ovjIyasY/1+MD1UaUE5uZCN1LDvuhPDpw2QHorGya6uy5eAeLgduOq6K3ly
HQnPlvE+6VUvi4gGo/VxhKzain3GjgFtxZ4BIKZiU39R4YzGvtxRnjKHaQpKsj42Qsrioe2GLFQX
VYGKuRySPflfiCl7+wpI1FHhz/Lk6xRDY7oBEVQNYBCUO0j8nkQzdpKhTY6bHnLTM/phuqAm48+P
Zem+iH78dhM7Ru8XovhHNGwM/LVoe5RgS0L6+/b7lxzm8kqhTJbhcMuZx3mOoEMTw1TGZBDN3iGM
IFZYSlNVI6tJphBhYzClo78PbTOXHiOCT9nUpuFXWuYmSlb638fMPhSmXT2U5PXDiPJvP0Dy53yj
FEUq5osUM/FRiKpRd517DKUpJMRkgtojjNHlb/qJg4gdHKyO6s9SEZcbeKY8RLUDpcdzBhBvlfdN
2kobsNx1ZPefAH5nQZGjUDciB3/eiHi/oZQ8gSoOk8Sq50Nm+2AikFka8CoOYN9JC2xiYLq6BsYi
VWTXzMPH4ggWMetGkLhiKyK/sIUlmCZ8vk6OqUAwRvfclXGEbcqKVH8lwJKGaq5piApINnEeqo8U
CEcDZ8tKOA59BdgHsIebFEsdN1IJZU4XeNJDxWt8/Uw+CiLkC1/O1A7NXdAJsD6Lc/URgLZ8NdCz
CtghetHDMYS68r+IAQsFzz5UqqDaSfSnTLANUzCfnHrZwprykNsLa+OxkvIsRwFMpo/1lQCBph/6
Od1X4pXPdT9Vtdd3aI1mvQKxBNh8XEXVJ+0+i0fOgCQ+YUuiNRh1GLu8/lol7V5h+Unn3tj6WvYV
3PNSTJHoMTQiTR2BF4fZZ22fADCkF4Xj+JyBsOMP+P++iMDo6USiKEpZgR4tS6ehe71W2Sp7EUH8
WNRW4u/tASbeUAIFFp0SvV5mUmE00Z20YLSXTxkzCsIjQ9YxkloIiK85PPsu6yA7pis5xCFtU7WO
cJsKru2sIr/ixb3GDOAb43467pFekmpggu/IkdypXI4qGJaJ2TxELclqDbwx2QtfWjwjTZdfyKlg
khiLPKMBjJ+Y4Jk4YEyKtGT+jfJzmK7zAWPQCCnPflmsIYYEnrtYjhsdG6KMknSnuStFP+979cOd
ZN78F5+iOMCt3IgjbC2+z1t1yjLER2XEOnu28gagI77vPkAt4+xMqFpJz2uDte2JnFoVPq2g5kwj
6fnjkGDcOWWOJfvRXrl83gjgtQ7OZV25+pGEZ1549HivDRmKM6TqubIB0nuWiULEYxJ0vZmaKSnd
hf1C25qblD0IT3IpLT9wAJAyB6vr+JpZbbYC4dES5vRIET87pCCAtHnKcPJYsfxmTIzdlSNk51DL
/qgpQ4VDJtMpRU9ypX4DdchCYhgt4PAGexH95U3626DnUNhmUprxIkJzM6HhzWjGN9vWNF8yZBU7
0xKnCdtEpTK00A8h07KyjoR4LhcEP6esmHEPDLsV2HxmxAPr0io9zaDbWJQalcThzCv1BLGSiMYW
wBYUvs6m5lesq2URGZy+MDs8pNDrV2j4pfhyX82ip3SV6vEPsIkVkfZGfuduMvHYWAMuSIXdT8nD
1YVlrHiBA033Mw8Ppc1RelVa7m9PBf5zwkVpHprvkuS3uW75n4tDD9ml31Sxoo+H8bIsPQEWcM1O
Np7Mf41XY1L6i25cxzp9nfCtB0X49/au+fyGdCOc2E2LwP3PNew6OjnWLzIQlfmJJm2Yfp0vgxdl
7QLikvX7d4py73DtWQ3M8RUFFHiu3VNDZGkW0DFvnXIR0OEc8FyTFi2T8nN6WANXGYztwjuM211z
yRjx/+1szJv+hEjSIhvm/bYeR6gB9SOTMGkzmu7KlwrulEHee9qqBbZzsyY3nyLVE+LV3GhgRi45
Ju6UX/SR3TC4lWBV09Fxb82ZXbOpGLTE/VJukt4slhmBsF5A7mlK8vGG8c0iLseY8aJPi0VDJGiP
ftawc/2dzdjMmFr61ymF8l+5hYGMZI1rAmvEfQz2lsyO6Eelux6DJi8j2c5sjk1YaE1J2fWxQ0+O
9DPOeeslLADI3JPyjiiaGl3cznrK9EAFW3/LoMelJN4RIZlk6waYT1UgWrPaieInDcSINQxueF49
XYVOnfovYavZNS4xJLdaIufDbXVZobPc7+ofjMGIG2N7Z8qh2WvAJaOnafSfK7Eqa+YnNzo8osE+
O9eHW4vUduUzbbb5JIADUn9A6DINL9kmuCjm6lOchs7FYVI8JRGswnT8S2DV65gQ1VozfrSETDoa
mqw/WSvFaz/xkPYmvSjE8oEYQ4XxWLY3Jr2wAdRj5OftuLDX25MJ+VnPN036GqkQ5RN0xg+XFgeh
8mhjEs24vHimCWnX3RPkvmX/ZJIGkOO0M32Y67HozEh3Z98kCQ6sNVGEaFeCPtGSW4WR48cO8BSg
ak7oPzqhXBVM0My1zorjaigQeUDJW/IlvQR/hdoW/dtnS6bNfmmHxMLW5RGDfFZxszXuDJ/zulkw
x3Jk8v37NkhhgNmDzdbeBwnLmFIxJwoEWTAmcMwqA7YiN8kALowcX9VprqciYavW5nWNd/A459HE
XARqh/ywu8ECj2w+hXn0AYmb9CvvvbUqu+8rVv3OHLORuMVBJIExhLESR0suZ8b/ksjm1KYCTrRr
sOnUNKFLvRUE7JAfz2zto2++8NN0EPbhgG7G2iFtLY0M5oWVh3e9vrVJ3oLFB6LMoUxiePZ0Kvae
Nx4zeYu/Lg9wEUDIcT8gpLAAsyZo8kjw/EvAeuuBSYaXQw/lSyJ3+BRr2lnNvuRsM5Hg70o2jOaF
o1aeoFdRY8em6CN5OX+ndzQ+UDpDoXwbTX+tvTYZ+r6nldl+2sQHY+LP0XsXBf8Lty7FDPX7jbb3
+xlR/lwz05CW+PLb/CHezccIQAJszpKVG3oHW9XrjKGNnplWhV5dxd/K91ZEU+RNMH2lZUknN+0B
3zje0Y8mf2r116soz9Wem4p4s9AhkDiAD7AyQH32MSvjboZZq2vUm4A5HzOxriexQmXD5pxhUhYz
Nn/t7/zOAfhiKTLLvGaeDjHMGnztfUCOyf0FuD/mrICSRgJR2aNdF8ftPdNgphjLd4fUpnobBg9q
nI3c4rzQHLgduaiR71NdUNCo9BIcwHE+pbc9lfPD9Tc8gyIiKvZH55kuGzwKZ43HRFllg9e5YC6/
B9od1Zu9ecbj6Vt1BXIqOVKSuBzXD8e4hpnPH88ktPlxvXjfCNuCTRJnVPIYbUtD2tcJJ/DgfIYD
4+cPidS7h5U+8Lx3prkf0TDerS2lgtAOHldLnq9m6jT14M09VJBFqaD7FLv9iISED6oRoQCo+v1W
LP1KmmbX49IlSnBVJMfyAFMxd5fa2iFRaBWg9y4rkhPcP0820x0M6F/RLLwLcKCSebPWNKj5ir0N
nBXLUuKfhrmYUJLstdwzYJ0UIaI/5uhsotuU0uxt0V/L5RYu0SAo7BTunG5P1BkMRfiFZrf1M85d
cgZxndUoCRM/shI/JoBNXUpUkE6gKivrOTDRjLfW6XGlNcjvlGzMyQyln4t9dTe5IXHv9YZZTaQy
hBDLUVzuFXZ6rmCfh/6RNX/F+csIwUwPbYm8VAP81MPdv9QyAcTUaAuitEcaJjsFCrE6HPQpwi6q
Zgukf2f4IWl4X9AoONfLlIasbHwAbmp2dGpU/gIMCw6kKWpL7EE7c5Vso+R6FCSbk3rW5My4gjnp
tZTRElkhegeN1zDY9LF6dMz8znyueOWO+dZMGucWOZtYWh0HsFFhk+Yz7KFFHKJd91w5So2OeGUt
FSZDgnO2Lafhb/o+Y3DgvHekT1s5a0g0eaireGkPtcCrb59P+Hlb4g9J4vjM2Zn+IyVE3NAdLZms
ix6emIIbBQlT9X0CLzwI+SUBsuMH0RyHtYNQwBCuPltXchXbaUZ1/sppk7yVhoHwdqj7Ijv3DxVo
AAqhWcMfCPcMgAVnolV+Jc2ZkVWdP7yuEn1tzk3a2aN5Eg8AbKB4Hb2vKEo2rQZfPmzOwBs1z8UP
PNQP2jUPcwPmoPofZ7YtbS6SShPQMOVn2FkJR0RyJCtlb8v0P4XGJpGU8wiRr+6+uA+sgOdPa5/G
kkgKM+b5zgaRcSubsII80axqD5OO3sK+nSUH93BTQqr+nlvN87FbWQcy6gIq88Yxj4itX+slLCnq
X07MTF1bmPWk9VpxCKx/gVnEcKxJ2bKS91T1ygYu7wQjM+l3H+gJIcH8a3QeCcBlicHKLdxLWHQg
I7Ly6oh+yqWU1wHRl8SseNNAaAiyuQrtOheT496FwUfqv3DOOkcBhMfMJqUzBQQKT3agzKs6HD0p
WZb/m8HDui0yIuKkaek6XIHZa0ukrwz1c5/eIvUrUEA/LhXw2jWSK2tvizbYn9pkadCvrmkRsTH0
ZkyPHbLD8nid27LoVgMkFLcIvhx2Vr2cxqxF8xjO4GbwW19it2CI4yBTJghdukohnPp89HmEfcuQ
Fn8o31qPb+iT3bmifzb09wqBp4xhj2KRUuh1auyZAr/l7YJFZsfu/AmEfYK60PwDvAcYck2ISEQ/
/0F9xHdXLOXErMK9uUdrUrJkD7mariAj1SkWmD5mzbDY1jpZwjPVTF/CeYpIuMkIWHya9eyMPW13
jVF8I47GkZR7DQK4Dvg35fetXbkn9HVz6FygPah9VlKab/qJNVR+EJe8CjtrElV0Jh+xdIaqwD2p
pd06BFdbVAciIjL3Hs9AdgHINgPWh2aHfTv5dQsxSAeGrd1L264vI5QyvN1sbCqnXFuhq6G4JLxP
N5ovtvXdJXU1MfDsSs71D7dwhPco9d8Y6rEm4MpXXLDm0fEyyTi+nHBnbblmrwWJiJDyF61LDtz1
BEJr7D4kK01eTaUpVmEVNTnjt/h5O/9cWWtfhkDnK08RoLWflmdQQ4yx5+PQ4Fs7mdfYDWOETAEK
sRoJcBSi8uY0zacXnrI9m4jiX2xEaBXWEzJMQPbf0QlIMXXFO+YWRSE90M5ckRD4utCsqtunG+Xa
KH8llG6L+BRkLnn2vbm9HzuMlZuY5JH6pCEdtzzDk7llJ98O2ACa9Cb6Zi6L4wnX26ulB4MSlYOz
RPeGzj8Gor4AlSO4YfFzlNhDrkD5ki8Uomgxt/9VYRilGMsg1a0UZ4GfG+MToI7d5azaMUfvWmL8
yuNgZn2BM/U5FOzpSURAGjmHW3pZ1QHbvqIDvaQoQQcZYRDaWcaX7KC/fDjfMIKsQ74vw6BTUD+5
gzHPkC9K+Jxd9F33slzi9JrkPWrLgaxlaHEacn5BBePnRQTtgJhSZHhQQLPMS8P3B42kp9k0awJ6
rkmHbB5oSbJLXo+f/nR8xd/g5Ef2TF+674XUbnRaiFV0rIJlhumJxS3VdcKXtGNNj+Rg4HcWQyyM
AcLlTvZ/UGn7sjUJ+KGSc/vPme8twMv9vKhgKvVW7ou274c67MHx4BqP7RR5f1iyt8tfPGNYyKP4
XuL8SMG/w9GYt/PI+S8dWQw5DzjbA/4W+OHc3ikz0HCccG0sLFGgMDSMw1f3YIT9+5mjwd2c8NGE
0o397WvEVoocuHpZiY4XMntcRrEp8fTqiZsOmW+UZPiCp4aTHYoZrZm9Jl9tEdpJpCsTMqxepQjl
12GqZ2XVuVo0rhx1sVB1kAkhgdf6YRJuEthIj222I1lk0JmlODfKNRldJtAiVwfKTIpM5xcys6Gh
oEnXRzgW27uiLj+Ok4qNRdtUcE4r7ShCMGQbt+Y+62avKMYuDiAVb15SBb5tld2FnPfEpepVvvdn
8zA0kL8FBEVqHj+oKYiBwjecfJlPdpSEvFNuiVgow2BmQ6dgbP4gXmIw3+2dQclMouAOvVlq/FmQ
D6oWkyPLrLci1E4hYeBmAUjUwBEYxWEBm0NVBtpVpUFrFFA/4y/1+iNTnAtJIqL3FOQerL/8uGGQ
kkvmN2/8YefGh9SCBgO3OsQY7TuR0HxThk8U164j1SGertztoir3DQ24rJbJaqy6oubBfVylsO9y
dAWasxaCyXzDVvXB2m9eZuvl1Nj54PXYeyVQWRLxcozCQPgefcbFcLp7ukGOPx00sVx9ggpWFv4Q
Wrlym42N6FWfbkpLPfsyDRkEAsI3WWnw6j/aHMzZSsWJo866nQOl3s2XLAB4kuA4wiYsepYqNDNx
GRp3Jz8WHnCdjioY/C16Nh1lr7pLnplz9dpzJVdjg9rM7UxVaI60suC0CwcHnRvSCOvCt7DcQXub
btN1iP5867crF17hzGbQVbqB/ELo2hsKOS/jhMg7bgdOCbxeKI1A1T/2eAFn+GNyhgXK6Weqi7Ad
y11XgLQDn9Rysc3cxS/Xf0N6pyvT/M0V3FzMW5IhSHTMqvQEqMhfuspk/9Bt+rGwuzuRF65LnO+s
s/GEPaTT/LxZ7Aic4wlzR+HZj5NLE8vCZt6Ny2Wv734B4KhBH5KKqZORYm8+DUMIzgkLFOtSOgrZ
eFReyHDl2L/KmfcdBH4YfL2wKjd83wamEDXOH4Ly5tRmMk1/QUXi23bTrlLMIBzICewC/+8BtBd+
UEB6ZhRpk8gACklE4Q4U8ak6SEfcCBd1tSd5/KZUvWOkMTy18AYaNiBGTWYHW/IpWRuaepgeYHyQ
0GDzMbba/DYjA6AMjf9cvP7ENO7FAvMQccHs7C9c6/c9wyAuETlRKKBCeXjHYUB6OYNwUH/BDMBU
0E59HuXFK+XAlSeiHFhOyEG5DwT8NrFnOzHRmwLmZH94dmN1aeepuiO822+Dg8KVpMZ/Qq+sNDWo
GdGDXxQEShpOXZcqcDxFgI/yDbY4Tmn2Zwe7VhvK81H2NL3HTrqg9pg93/EVJ22eKUvPZUf+uUHs
yiTCgupcdXg6UKQbqobDmLZ28erqXeFaCeL/T+OgXO2nJxzaAmIutPWP9OLCGVqUT1QUmFTayiIt
71NBfGSxRQELvJn3ojxktdbBlJT1J11PAG0tsG0XbDVw/7p2qrc9fy4XQpquYhuD2LjEC0DSgM3A
H1Z9yk3KoY8nYGnhcp2gvHZXf//mg+X140qgMujEnNnm+9S6dtpuCjy0I0vu4NFipOkTFq65OKCw
2qmX0ZoWYOoZA0i3zwx9yGUAGaTMu8wbfnRX4Pijr8J5ni0zqLDhsXTXFm7LPcG6VE4h7NVWCm26
XZ8flhMe45wJVt6mbM4sfQT7A7tx1en1+iJ9S6Jh7IA++RosrLWGhERx9VdF+fciXNAPm/B2oWvw
MHbT4doyo7SD6q/l2FdFvm08Shp6IrvMuMVhQZwg9T7GgHMreU5kA/OdHeOvrfAFD1E8aRzfPx6I
QKBFvHSlBqc9OEvUit6kjh+Xwu1JfB3kGRmZDJlQhW7sD0eGvWnT03ow3wYNTqc9spD6S4KRmou6
bh9DT5QhgSzidG8I70Z84SvNwRIwVDcvAuO5OrMvq4WxhQQp/4bp8tjbu6gOGofmFIL6LSM8SKUI
xM0rpSk6OoyIgquBaxwLPY+AoATaRMa7KprWeoIB18qmgUl63PP6n8aVEXPlTHHvlWWkoQ1cEjVE
WyCAVSz3icfLeIjCgcj8bZxL19QzU9qb2CWkwcRMcDmx+T5K17621MeYKazb2fQPrRW64IJwnwpf
xM7cucWFzJ2EDOIQCkFJ32NDgN5A1c0/QDs4nWJGg5HAQ8mByX59eqPB+5WUNw2b2l9TBbMz2lSO
Gwy4ngPACrjtj/VLS+wcxLCi1e/HEJ9GwOOq1JM4g3DreIeEwJYrevxJvaVM/2diNQv7zw1XSEG5
sdI3ArmjnF0NyU42so3o3+gPbLxAARalHZeP8XZm6KDN/GB6tLhEEA7TwjywehpYtgSeF9SYqgtt
Eb6rRtizeYAQrTpcN8NLBc+g390xCUwAJKhxvllVKpV9uIYFtoRo6dSa35ih2cIQu/m6Ifx8pUNg
QrfTGE/PLvFW8US3RoyDghqVvtupDzLG0EczWqQiuoXI7/ciP3d5JaOjN6B+peeHUgOBgr2lwdGe
evrwJUaMgXcYnQVzgCPoVuEwNhA8q+9i6ow7ATzqQ4xCyHMpPIn8VRFpRlbX06LmG/tiEaKsfNvE
oK3xIpI7BOnE1j80iXT2rqOvKCJDQvLrKt6EvbKeKH5u19CGt0uAeUwRZmJDEkJ7nwaal3G53Kih
rRMDu+9Yry9nVllGir5F1y2oN0NwKeptoVwDiit4dy3eHHmeofqDAOgP5+tcyLf4AqThdl8W/DI4
ZttfVVL3uWrEoQm6oCtQISDURizfr9mUnUmoB75wIto5fPyBD3ItdZz+6VVvPwnvtoZ1Kwoz3kEn
HpR4gHBBU0Cvtsyk85akmewJDCHBMYxoVNFvAHNN7hXDgyxoNyNXEXxb3VioAtT5Gd8mWMIKRpKq
IktrNpIA5CUVRkvoaF8gpc0FkGTTStX/Td4ERFfXNYdwgv9tes/KIFjpTOsN1sbq49AHNscACp+O
KDShutCOtXUJ0cSEgH2+6ZQXAsNpU5OAdxT14245iUwYKl3rrHiLd1hT9SZ8edhu6RH9lAzWDckM
aJ7JT/kby+XDR2VNvQEV8ng/KuYDAWuagzz9THilTbwj/hYfnJYYfOIuIWzEblZ+hzZrKVEq1Nyl
wXBlO0xcl03ZvwLffG+12JzPHGmt6aP+O/S6qr+2T3nCvEH6uU/dU9havOA8g0VqNeXrcE2Xuh/7
IrH95LUemaDS/J1GJXIN4i3chSQ2TYg+mEdMegbIM+AJsJ4uMSukdurlHHk5lfSUEgy7JHkzd/c3
YrYDBhm/LtOrWpj6PUaAd1lxIG060cPUlYGsLhMtV+t4ILsUIXOESJyoVzDXU/XhZ++unlaGFMPV
THMK5RSLsdX7hSBtAkvHtDW3o0n6awTrY0pvVUAnTzC3Ymndm3HXdoZkcrM+GOtbJ3yOQOn0nzN2
maZbZhYJSPdPmXIpYJh/jBe4desP/awR5BrkbIuicqgWT7ahdjkyUj9BA5o0oWDyBaRTUI7MGNH/
mxjYl8TrCMn3I2t1egk9rPYb9pUbvBVDA1muzYh4a1xv5Wgk33cmR2l20VhLXS8UvZkJQ6RgiO6z
VfPm48htUBODkISxEEBdYvSrY//bViD74wND3FPS9mB+ABO2qaDGhaVojNGqmXTIuGSvoWGNkJ6O
voUXsn5l4szCrLYBG3f2nadSXdCUsRFTXLGRrFcBCC8WlIrnSmAiUdbIuUiAa8Kwqkkt/ChFeMpH
G3auprmq07NttGhk2fTwItjZLWhVLL/qlbVHB4aeeZmDadFRi1mT9HHvj21S3GBQLOObnEOjdW7F
fTpR76KVqYZT/SX2Gq6uO6YYXu/8EsV/39fY3F/DC9+7n+feyjVKIYcXQH1HLntalFONLt3pEHYn
J3cpwYOenDDaRsV0/va+8FzIIfgk+U1ff5H40Evh9LS9Ew1vT80HOChLmVhnhCuFtJTL6ez6WoY3
Ip9297SUWJvfkjUQcHcFgPA3VIqecqcpJvCtNjXUVhcITsX5RLVu3+CDDOk+pIPQy7NBirP3k2Ws
/qvl11WUQKRfgfTAQ0A5j/eUIL3bViabHLptqcncjSzyvdCFKoVMY16gjts6kTL9rYpmylnBbA87
R482SLBtxb4KVR4skHj+VcKEaxL61+ETkdpVEKL8SW3w7nAywdbCuGiQlFOrU+Sq29PvWHyRFzB8
I6u9+1SHaceJZL+nU6Nt9g8rueAM/hXQaaVvKcOJfzOhvnnCupOTa+KGXUd5H0/Ps9h2JiYgz0V+
7zd/+0+pr3gpPb0paecZ2b0eQxYiIe37hALNcbJNr9GVXM4cZ5bazq+CjlxdB6JUT2UwplTq2uaF
7PDQl1tK7DeDOslXQfvljOVmYaihHpyOl1aMSH2PM73thjwKCkCBEgONOwEGGB9k854j3kwG3LeB
k50/maYbDmeVqi7rudiyUhKigWlPs1D5oOuZ9nKHpnbwRq0jy0M0Q3F1DmF4B8deYxwyZyO9MUfk
3t7yTusGoTNwu2pRp19tBdeDYuTnHxplZ30doNniMKpnmuNbLTdtoIb7hepMcVpPDSsndzjRvne0
SCCnz20h5cl4PCQT6lM8lRkV6rbhxzb7zprgyZTkGfAcb5epIrlrgDq4QlPA88tFwOuO+PdOKdz6
TWtdJildr/ZxSWuDRPMFJTDI4/cLMJ7/V3POZb/7E5hMNrIRkVkszDls2finxJatD0kFukh/oQnb
x0ue4oGHrg7lRCY8i/KTvWwJAyb1uYjprgbegON2xVhN5b1JPFcd1/ojhm5StLI9BPbYOVH7p5Y7
zLe4C0x7sEHDHNIGgwsCGh2b4k1zAkrUR9KccDy/x9Rd0b/3b+kbVDzh2UG32oHbJUdAdnBH4dMQ
wFAzW0pZXz48cIW54t2M7I0AGqRb9ijMZ/DHOKanIK9TQVVxGINm8/Awk0+1f7R+Xo6gxS5QQ7yE
A1gzTblGtIPN29633yyZt8beIHwepeUKDe8ANJ9De3/Vvl+DoL66iuIAO4Blhu5CXDAKpKOlc0hG
bC/3d2k4XGuXS4Y/ii1n34YOvxYsM/XPnDQqLQmNatLUOc2XW0nreh6o52D2NcSQ4iks8ivYW9lU
JoiI13LFB6YWnC1WuvWHEtakOHhbMOxvdN7poMpnEZwdjtCFak5B2I9KFMcvvtAwhUP5pxrw4ajd
PggUi5Nw0iKvvg+bRM9N0Dn2JT57tyC943C1EOtvcj7DIuWOkuJ5Hh1un99ZQs6MUtSYnQWDTvbk
+6QTIcucFBrwrK9S3Uqz3JICDgF/eZRr4nD+mSSVjl8Ikl0nxgFzPjvbbjuH65j7Wf9/1hzRSShL
8aLz3Sqe+ba5cxcnpD/Mue2vzbWvOAd41W5O7HemHl3PEV0vtdgrtT67zUkqLWVr2KziBtlJK4W3
M8mjUi4MCuP+dPrW3KXE5rRWeS3tNa+uXpeG8zsCyPshO+8aRVz3j13PCYS9jyTfEMkCbpvOvtL8
BKk0nKEWLv+NqzOeW0BdD11Cm6Uc6yf3BHKEtjD+5cA7IM5fU4uzxHDkdjTp/mBh4uZDf4+kGWir
FuoHg29JdV4/EJJGgl47xDeiw/FJoHCsBfhqSPnj0+J9WjezdSXg6Bh9GCmwf3OA9hFNnLfs3SSv
asXAUbXl2Gzf94k0EXTw96wX3AO0h3Vx5QP3Nq20JiFsP4SweILpDc967Txt5VKLC+64qyPBfeWe
01zysMDUyHEv9fsV3o3qrl2PoZpErTGKkLWtOhefuEEYIrwBslwL5GC6l1cA3es5QKT8jXDZhysP
VW3FYrGhHqocQrzUKlQhMkhxzSy3A7hP2QgpIQxiiSPfnHuYOWp59t9xa/F3vXcs3LR/7+blgR+b
Cuih9mHUXQNixdFgyl2/H8JXpq2uxN2wmQtZLvf9EiUYU2EEMbsTmllUG8o3G0kfoNE34QSLmWio
kc8Se1f5IK0wgWcO7Y+xnrGf20V0A5ng92G8/Ioy997f1iuJhGc+kV4OrLlp+sy6zBcAtT4jcOUT
OwmTzgfAhyr2qy4kZFe/7sAGNYBJR8Efl1vkIT7dDYHOR3a4A0Na70RVeWYSNMXKBpJbO7FAvYDs
rlnQ8va7O9qeyNd4XPRa2sLGK4OwbzeRl4KGlZpW4qCs7XwlVQVJNZQH+8Cjh///WC54V9FpqFDV
YFejCaT3UzBJjHOkdSBCPdfrX4AarMNXWaDXql3MBD7YkgHC/XkqmsIVGUxhMWkEqAAOdSPsIwbq
p6J6i9Z6ADBd1Z1TWOhjJirmn/gTxlLw/Iz23pd05L0gNfQxjuuHCDNFPWhIIpXFKUeLxscaR1uN
9bMeo+qduydulpxB47EO4Gba97C0WfD7E0RiK7dkXF3uGOulV7UojlGLv8si+Q+hFoP6prEblNdp
zbWj8hDMZiJLISPs9tdX79sc1PeuncWy8bSTBkZgW+R5R7yzW2uW6JjIsnFNR6/e3+tA83ffR3n1
nO/DvfPl2afY8klUiSO4uiHwaXrY8+iyKos2oG4RRlk0wEOD0S0thHSJZSZkas1vh4Ho6+ImAEdM
mQJt9jDUN6eTfwMytt2BspwdH3GM0MIGAqnzsHEsE+657K/eejsGI6054O5e4OCkfXlMwcz8ROq6
FFPSav0hDmEGdpE/lBteTPH7xsoAGZDhDcd8tLuOdskka2KHjF6IEsovztSs0Ys9s4SqJ04uNz5Q
/rpPbH18OGlSWoCJq8pMpwg2UR9zVKoE8l0MXphcHWTUVzYIg+CQEp+T51b9SoGVeZW4xm3rJrQj
/1xspKi0v+XMRU1SJVmFAM65uozK+FCr9X6/PEESdYs4UOxPI+mao4s1f+BvkVir7oIJx5Omxsj7
sbQ1peirQIBQV3zX/lXtCDLKU5wRizuqF3/Z5ZlEZjseYmHWUCR3v1Fn5HMf1k5Vaz7uQ5x4pQ6r
m77xsyKb/mwTpH9itGxYVsfN/uvIVMvIX7Oie5auDy+KMiAJALBvyzf5xaVQru89wsAkFP9hskMH
ue83kLQnw3tJNpwkk0N3vvc50S6K+cdK07AUUdIwhkLRQ43rHhxw5PSgTKSQ6A8+DeL2ztxUny54
IRCXFZVXi2rlzk3lL4aVqgmF5VGhx47Uyb/nG/ygNporLIWIc0xyn79XHImBImjv26T3HsONJqgE
pBwlvH7ZJGCv30yNe0gMRuF7951tR5iPC/jFGJzpOfDq/DueZAia51G9y/VT+znDxfy47BO5wfca
cVJfiTGLtNdIrndPMqkqM15hA+zulsCYpBEbx/ELCT4r+Mn4X0tWHNx1sm2TmLIDhVZrO2vi5Wmf
IxU3dpPsJrSCXl10wAHpRPZI9g/jfSq0TQ8V5iEGXJdMweJPJT/PdOCisDUALcC0+4qGQgPqFN2t
7GqDYJzHHYAn4e0fS9Gp6Iv/H2IPCcc9uS5M+aXZggnf4NBUxCh9YzTQlDDALLxE2Dgbhb2KMxFG
RSzwy8kvhhsHIzxAceUXDpFL5f1MigoKpybTYOkjAI10HCstwBzq+WiKiRr19vpLvWO4/eM9jEFM
vjYXIDwrQz/N9SLJaYKYLYkLp/K6YX+CTmdY3kOxq+HV423AuTKvfQaefVzAUoQfu9RZNni67kg4
EGN02LlJnJSBoH15Who8vxfsygTKv9P2d1NKuIDiovm5rax+2aSW//lAOIfv/7tAXdyU4F1dnPPQ
/mWdN3UlO0P6C/3Mv2XbmK4iMIO9ThIr5bZU7g2IxafOvTFblhJrjN50xxwDkNjSri2c5DvU2E+X
njjmW5/KPmyRuZ5UOlCCSK48bjRBM6XvfWiYrY2cdtcKphN6nRkT7ALu+NghPa1Dlweq+3GLw/BO
go/p818yfLV1taTFBlBzAeSsTYHc/pzq8cu492jzUbLdxho1i2SeivtIS+R8KX0kEkeSXTG0EFdf
gtqBJPgWtnlspjlhkM26m174G/sArXH56JxLIIrjw5yZj8PBWDN12Smd39EMtBTVYZy/9WQSG56f
BtXvQar6YqgbpdPBAK6a+xgVOY8RuuBo/baCuteN9TkOIOONJLNMnJQobTHRmD0uNmf3XriOO+Lj
6z2inW3LC92Fbi6S0znZ5V2wHlmckgY3IkS2bA5+A0euSiVEa8c819Yhk5XS9OGlXC/Mu5UFHmS+
C2abf1zBdLlKeh1EjSWOE7SSbo02wRjTUbyeEtLUl9P7ZsHPiTq2LW7ocv6PA2pWMDiq0czY/KLD
J+e1a22HVa2NtyzOW90rF/wLz5P61NiN9DbEBsckrXTwJBHyUbcYXtNbfFmgRXWLfXMuDKoNIP61
iErnxGYQFFHE0/uljwwfOlwqzgWQPoKMQSR9o8UH0lrIXA65pkSSHg9LzEvO3OUGG1+4F6dwwV6u
06/BtqofM6sLrPt1A+Q01mEwodFG7u8ADfpd4BJ2zPS5YrzCenwgKzDbb7Mic7+tuT8EHWFFXy01
MWV6qzsPTD3PhioBSHoDX2qIsOCldLuofcy/77eS38UH38r7tX6ka5dSeF5HVVTqptgrBX3OvuKg
yui0BNmb1Epz+mCBcEMQmV5R1xZkJVow0hGjJJMxwa4Ty0c9KmwzyCByZAQe/Aa41VbU7kjOeI5C
APvZDTIpyT5WEjRYgEg/1FEo4JEQqA5AvOXeUm8DTrZKKERLxYhD/kzd7B7/CqyvoDhsb++JYFWe
Ag9vdjqyo96F40nb99JXYmN+ATOBZSI6Jrc14UUQvBv76WINemBPN+MJIQ8RahgPHQAxmhtiuFEH
D4u6gR27Fm7uKRxSJWkFdqFdKRQgDj7yQR3lZwULIUTzM7swwAqcWVJaVAfL19sccXCbBErosGVj
sf2t3XR9+UPZ5BTenNJ+w9GngKoBKqh4A/pTV9mWog3iYRRhJSH99lxPhbJKbSSQ4wqn5aOAX2Ih
OoD298MuoFdB8AJ0vFlkA12YFAbEDWSufwwHiBXRTclpw7Gm6DfQOL11RtOpWnaCfQkL2ntYb5sT
emtf1IjaD0AiZxoSL3bTID3BkTuATqNgQo0Sh0L1xuh8HTg6N6USwffdQZrA2MEp2wKrJjn+ibM3
f8yUIYSk+0yepczNq3WARV2GoZf/yTWjkHLAGrare7obb+gnCfzoRIwfG7WTiKW5UdEjseATjP1i
8+H17GYtP4r03DsFhqz7RFm/sDz3LDM4BJhBD2vfB23p6dXebw+FFW/S/m0RRZyTxi7Z5Z8mp1Rh
jWQCfJxdTXs/pNa7ZO+mm6uneBMokf+4r9raG+VARz+u0+qX9uKcExWsvZVL0NWRuyUxdozAyvkV
KYIb8NdTr3BMV3gZ00KFd7xnw9aze8lAHYrSC0MxAcJ/ZB22a0GuPirnMR0Wb7GSbMDdId3SllQp
C9CedN4K06Et7M8mwQWvR96WsdcBAxQh/ihyAnw0FgYS5dsjD1CfLTLpJQE/Pw92UZ75H/i3Iu+k
yk5G3SFgiUEX9BSV7PNHi5+Lwu9VJA88aRF/lHlmRxfjqDwlP0ND1rvXITSQRmw4mbtylHr6DKqs
pmEUI3WTCiRfmJ4DNT49HMf97rH3gjcqyadfrYusaWMN/JEUrblHn6zPtzl8BRwu1xaFVr6UDo6S
4Ff3M9FdhFXqLWB44gdAebMmITvuEDx++1kykV9rpSsm9U5oUkENKD7SfuiWlxgo09E4Tf8kNNJZ
vLwknSzFM96by/15mt9CQtXGe49yItjgrE7aNt5mISXkbvJMlN8M+6ePUtUACM53ad3G500KKSaU
1LIL1619l+ZkDRTew453txmypb5Owa2d+wyGMhdWRdUKe/jlWNqPRQtoPMLlMdSGPeWEDs26BgPo
MSWVo5QXke3rcmNyzz+CX2vvD45Q4wD5y69MINnc1q01QdSSGxHZdpZ05w9oS5ZU2YXvbr7ofqW3
Yd4d8YZrGwsuDIkoNh/k7/3Wa8vAGxelmZhTcjW6veLF88yoLW1VpUCNzu6kx3jYVoBIk8NaBme5
f7qa69F9PkmG1j0UnnWnPtyuzLzGFQIZTFEqmh93tdbrzBiVfiaqv8OdXykNJpUtVO0O/90x6gLm
essZtfFedzoAqh4CRzm2EG96apvAqIlZoByVxVQP15ai2aRN9f8Ek9jfUUFLYqHwekJCpzycBSyV
GwVoHigvOR+5OqXBSL9fPOpQIc40rz7TPw1evEQNAvZyYue00ch7vnBiWMzl6gK/Ku5g9cN+KhFo
U/1YC+TT6DFd+FOBiKZz5h4jHn1trhmJTWL2IBw7Arxx4iuuNSJr6DGZ3eLYOBtvJTu7Y/JSPQsC
NvOURSZrKbRZ7O1fBcGmqvnyMAPCxOF2AoJldO5CL6JlKy4bX/n0pXa6qu9GAL/rHGFQRtUvSDfN
vNp9NM/jwM+NoKbh3+N2G0/PAOd7lbdxLNOvbFdxAQVky3ffHETBXZvVKuv+htqRq2S7ibwn6b66
JbOyarJaaMDPLvNIaeUWr59gR1k+kfwtxH2OtXHaO2BWD+kZ0ldCgQzsu2cRZ5E9++nIZlSZU8ol
vAD9bEV0Hjo8ul2pLBwXTq6LC9nfmyFSJmRm36GS0VBJug+CXIBkO18po3smxIpthr/xdguM/9It
w9/daPWHCY+JxHuuyODZlsV4LEoaEjCe0+aBZ86QV0D/iKJ9UyiQJwH8yg4DMduX9iiGc2d/nrOd
VBeszt0NeFlyyHkRZWNvP2RpMpVesZZTgLK+axXRURZw5bMQ4isRxiUsSt8Sy6ISAfhc6SKX8Ad0
5lwe/xPDMv9zXjapO4TWaHYbu5TrL+400fNcPfLlXjcTm0W/BCkZN0gEgoQ1LRhh9yUTKC/f8pFK
SuNSIWdzBtyHr8uQxzDotjNeVeqP0P7rcNtypjDRssS8+cDYWP+KPb0rM0D3xm5xEbKQWwqAhzMu
a4fqglL+F/YVr436zDJkmX1hXUBOjG/ShHAa6ml+UUIsbWWERqia+z6p6Ye8RZPYJc/q9hwuiG/L
HHs98Mf2hQQPcS5PX0tpjN6WWCOdsUBdtHUJeovV+8HvTqDk8d2OnAi2eirWFGiEb34iF/KJRGg5
/QOZjpmXb919RPuUrrhQmru4ydQbwcvv+9Hrv8AgS1DeNoBB0uwjVfG6YQw6UMc2nD2FRcUNrfu+
ozTbmOlxM3lUT5EyzrmhL8i1PGusqxITvcXRUGzlQYjzEYwZr+yHmtv8m01/2dJwzj4i00nyQXmi
fwpLpW7NEo70t2qWXnWzRA7FKiUtAMR/JQT9EAkLpyLQJcDtkDX/wjeaIEjEH6TtwFf7ECprtShm
RpCQUkFt6nUATOA6XyNZIcMC0VR4TTmqtFfwNog6IWaHHmEL0uv8Xlsr2c90hNAXQ3l5aloh/Rn4
DBfbdo06byGjPaJdDnQuz/iwq5LHbZKLjR5q+IWTVB2TTQD7/PsWenUL0I5cKgWWxD9B/HVV6HNN
JRD5/D1BWUn+F+Fk4rsnQfxnOSwBRqFso8mdVKDlbadZ4S7dUUzt5jZez7xISD/bS06uITpyHPW2
YaOCIxvHLZ9Bbdb6Hf8cvUgYEPGHvCYQj6bNFp3D2z2pCzan+m+w2T5KSw1ReHgLUtOjgVKGkyYH
qUkW4toPMzIZMIoYGf8znz0bLQO7qcAkaNeSBnuB6xB1WVb6kZFzOshVqStUA36NP3nMMqWu7du7
Bq/AgWPUuyD1KrYBeraVkFv8Iap5V8AakORAXI8fswgw3ByU9ExESEtn60YjI6c3kC72cTT8eCJY
OtgjBEKjv0U/WSfXGKiq491EeN9aCojctozpuozqA52UPQpQyNRt5xc5aMqhZ0TrIGwyP8oI2IVe
6Z2CqiPC+77mOMtnix26fsxhEotzkpDwyGbZmcd/9PACLJZhrGZEsTXOHiHqZ1tS3/7EhlRYK2/9
xgLsJWBSC7/WT8s9NPzRPnpr33Rc1CCt157oa2Ku9XNE5eIg4hzKo8AJhTaVlACju1z6TrniW29b
jutQIifNhw7+bVCvlyM/lKPa1UWRioq6oRYFBW0wxYOgH66Hyd10m3lcaUVMGLSAzVMlh4XEF3Zm
7HQ/uL9UXhf12BoECajICq6pVUrBNiMjBYpmqZW9ulYNQBuzX/KHfB0jodxzxTJVFpci8ce4TPbJ
fE62KJqYSKnckpAMP5oZhCDU1nZynKbfNeLzfd0EcZ+++0pvgqrO7oQVnto4Bb2csNm88HDMXz6f
N89TRpn27msheg1lg/Ht6oG3JueVCsopccKlnzXKvC6sD/c+E2eIZKp+f7uLQkaxwBWJxwC4Pi/Z
hkpa6d6+5mtYDcPn55AcsROLcHyvBspPDYNqktvxFQWE344qpQF5J6m9JK5mOc+SjP891/DQEWR6
DhR0nSSkDj0Bd+i9RNMxeMEjQ6HsAP78IvBVYs8MrpWg9gX069uUqQwv6LBF4232RGHOfWYM+SJF
TXjle/StCBBprb3nOFTcNo0B12CHinMckwKI714rxZMcp83yAnHaldztcaIXdSD1Pu2zNqNkjp04
p9eEBcfDbDg9HOkeKDo9kap531/MvSf77znQ3xALWR0/INq3USbtZZS/nMworo89g4orfZvuRSI8
5PxdTZd6DjRvD0+Bx+sisaH4w0TqBvJ091J7AMXRN9xa74Gxke6Iv10Id4rgOp+ifGB+SIz/ksXb
rVDzaa37cplMqSmFMk5cW+gkzbBP71FqCN+a14AYXf/cZ5PVbrg3/Ci5UAr7mn+RKmLlMPH+57CA
AqIvrZUrqpfuoEB2DbpwzGBhirl1FfrHR5XSyXDFiRagkla9PwMGtAcwDqdaXkFE3VH+vQk/pXWN
KqWD5k9Bh36Ui0aLlgZCej9BVC3UhaToNU59VYbVJ7zZFz6L91d3rs+SbrjZwadt+VAypK3ZJVuL
9vcgjGkaE7AHYahXp1ecZVYLeYc4h9dOKWMkJhmvh7Hh8llS9DHXWu74Gr2GBNAKdeKrx04xZswU
oMM5sTpDYynk1XOAvQ+fov3A7B3FUI81+3Hdi25qUT5BJfm2e2lZXRKXY+7IyoQRL9a5zT8ejUFA
hAoHGHK8MuIDBiZTzaPOTdTdzGJ37mYInsESky/c1LH9zHAxjuq8pUk0sj8sTDfN5AZNR6KKZuzS
1rbZz825tXJUGzxjR2iEkVzXKs/NI4fT1Xmxhdwf++yA/GAlImqgyr8bxrio8Xs2j/ZbrkrwcMiA
62YCfSVpQgtvDzWQVAxhRJAfzSfjZPcLn6SbtSF1LaHgSKE/w1LmV+yt1M2HsuG5Lvp1r+mS4cBP
KJKgKlY2/D0SW5UmOCPz/I3XQ6W/OzizW3ZhIWLO2bLh9lYFBdTDisoJuqmqMbrc2bprIln0GBA1
mOk3xHPD2b2MDvxJ+rhTzY3ILJoeGhgBboLD1mdoW+D0OLTxyBJk+p9nT4TdR3WUuo7Ksxf3zmxa
1D4yNYyieG/8V+PfKL7pV10Td9fDOrkUJ6WLfLrjcjYCnCO+WWKKSO09BBwkCufuVvOJduA7EI2/
Ft6+dmsLAOdgr9Hg2VEavfcdilOTtR0ake83oijr051HfdOb1NPG+sQrnl08xkWF8Qo7Bsiw68RU
qixZ+PD8GDT/Bm3nJuwtSlIZqG49WDfXcJO8W8GsDp2RGEmrQ+gtttccfAQKfbuCtyCQ4b4CKacW
xTQdBPUwtAtjMNDWBsA8GC+15Nt+ebtqD7TxNK5mbhDhphtiY5y+cw/P3jbYRrcrVOWk1A4LbH+E
Fm4D85atJbRerWWOxtS0UEsG0GMbE8YRrbKAnvjXnl2P3lQq8o+s6iJikOcTun9ma4P8+YtgKd4L
m48IE0kdQJQKPHe9zftmXxa41Em85Go1AHzg7vKsTswvKqK0MzIojXk+0C99sQPy10DicxVkBPro
Y8d8Ohw+eqXWEZ6+tfr5SB++fQczjYergjua3dalKIb9548DuI1L6mODXcEeAOHIUnoAP2bvH98p
jlY2+LFOItfPbQg67ewu6o1Q7tALO6GFNs/2ka6VqPEobYmCFgPD1rpSyPjITYD44Kx2IG+dwixD
XZrwJOXVrKjaKBJoVmpBElfgApBBOAa4N4NVkbu0me+R9wId9tKm4f3cvUbO3AePBhRd8xpUIeSL
1BgGPheTHkUiOti5AYuqi1D1Ne+BIjWahtxRp9u2XV+uYJqKigwED2DTjhhoE86PRTeygAoJuWdW
vb9yzE6ohMHslJBPFxuVQ+ZOzvfxa/1Lr4KnxZxaQUt4E8/yrug/F9Oj2Qon/esYO2PS9zamGg04
08qe/Hgh1OPKAzTYcmphQH/vD0dadmJ7cQauiTt8OJA9tD4aZZL+b+8xsehMm1yVSz8gZUk+DWjR
OWU8o4DqEkAqkAXTBIoicwvMzNTpvLTrFrzXcJJoZcSFTg9QPNZeZ/P9+eTh0WCs2wwdsHAzTGrc
nwol8pDD4MgCDMuRpGDjhlIiqvpGG2uVHqKc9tEw6fKqvwTCm/eDVRaGokBJ0JQj2pYMlt6YWcNH
GovYFlbunXJt7Cl5K/JDQsOUqGEODsmzT78n8rvUfomM1U5WDazeiTzU0WDnJL6tvTuA9trqQYAm
ybVNrFX0LI7kavfgqrDZwb9PivUmgTk0EuypfYkA94OqjFqhWRSPuVk54nOAFkO0GlLi0+1SExzQ
nhW1zhiQgJcTIqo6EgniDjSiUgK0ffkAps/peSaFgBsBq/E3FAfXxXl67SJkOPv3p1VcnBE3fgYP
knsLZswY5e9dpFMWB33TqR4T5TcA9yXjxQuJSDmeJ118RD4yopZPXboImus6gCWq9VH9iH7PSri5
Zt2vXc5/Mudlj+pyTPSoRhwCFlMm/n2C7r0Upv3ADyVNH7fq8Mc0m2hNgYiMVGDzuE4tc47oArOe
2ZZh+Iw4+ElZECAANBJVYEb4Zg+i0CxKVOXEXIYoPz5nPn9OHGc4fIp7dLbP4O69OTveCb5xO10l
ZoIZjmghRnwG3lqYBDj+cc1/pnY2AXZRSc/j/3stx96AICWxsDXkBufLlF+gCSrlaIu7Gpnb2crw
Sa7mCEoiaZfvTmE8GipnLK1f+4WQXC+Q5UjPp04P9pro7fwLdAN60ONDkgk+QvbX0gQQbOJIly7J
tGLXZjxkk4w55P46zRDqBNJqNcN051KUdp08MpdCz451ByMqwfOPUDD+0B/SaiWb3HGyBr7Duzmb
r0MqahEbDyb6ZwQS0lARFHVQfBRkvcjIzyybIrD7vjh4jR8OmbLl1vfnJpxcaKJAuolELW/8NtDN
8cu5FjvLNz+QFLl9JsVYhsPi13pzyqA/M7ZVLCLrzKmoy4wGT/OUwjjQn828y5CLGdUFuQcEceKU
GJQYEtBWcOVrPyweV3QiU593f6hFxHTKBi5w/ORwJPZ/S7KJNobEjtKUDG/fL9THMHxhoqR19RU1
dZ3fcaHGX+2yYVn1Mmzx/aY+03K4yML697GCAUCGHIQjcaTJYp4iDgiaP7nxc1Xesl4eKcgNFiq9
LvTplvzYUCuC07h+P+tRKLbBnJ0phW1LpVUBM8wU0sRqJo0zyiyOR0UeIY+hTzR5Zosu6A6KnVL0
oz/HUGhYIWIISkQJbCW6+XHos1By+62aquuj6cuCX5SLO57eDkTzJixpj/AWjeNc/NkgsdVzV1oW
GdomWf6LC3h7DDDV7+JuoaPuZe5e5FgtA45MRrpP0SPVWBU+ZzlJIvKqfNeBpt+KCwqY6bXTuyHm
i11MViG9CFOV5oKI9LyJg/ZK6MggVk0YjPDKkLex6Q8DTwAqMUXmn99OClUS0YxUoprDJvL/RIow
+gQSK4dAuuy0SD9+TA9kenQQsphdHylzdqaqaUdNhHtiKuRA+K8DB/gEUjiWHJMczFO0qdTZbQq4
T6sn1w59Tua8R9l/XiadWFW1Q9TdD9/xZgmOzFILeL0k/1jRz+2EuMuvGDEirMPQDqcLT7wqOZI/
utQ/gbhjxzCGHM+E0+tg40g/gOnQeCUo7tI9RemKCaCQQSNYHlY6NZXeTnrSJUwPZDO21j86xEfT
I3IKFg3QMjuj9RNybZk7blz4ggGINTIt0I/AsjGVZJfqrbC+4TKXVjWaE4PB9eg0nmuhJu/NdspE
HjREtDGuxM0chjCkjcnLUFGRleKRcGHUySfeJy1ANT/TMthqRuUqEphayZq57rVKudl8y5rDpRnx
CTvzYLDAltcodtxNFvjxHXWT2XBErTNPCcBx6TCNL0VmSKhoLxZsL6ZyB/3FIwofy5FW8lN+RsH9
u9gyCivtjWPhyi5aFseYSHhGSEahM31zrHhUT9vptwYXOYp9JD9riLpZgbxSJfxXawbzk7zeJ67m
7yyEgDNac+3VGN0L6ScLcZOfhjmFq0d5o8jg5z8hh9cQE8EL5QdM46vUVRpMsA/mCzzd8i4AvhSC
4pMl7+WShtnOEz804o41yr2UWIq0/1chR72BZru0nW6OJ7tfLwS78cpaKgfgFBDvRHpXG+RUnbPi
IfL+WklNCkFXAbaWwL1Wt8qusFTuDPCL2GOycqfvLf9idaF3WCB2cHjyG7CoB/0o4krhfW+gAFm1
udIE5acHQMsIZ12q0jnMW0c3d2H5aCai1c+et4ffYUlCD5E/s2EF1dfj8thgn5BxHup0BETUs9fZ
FeQVmd0/78RBgoIeNIfMmrb5iP6dOXO1tOgWGJxdV1GDIrN4VApB/2yhRV4nineVZDtpD/CENKNj
hKEI3g5gDmiV8oN8lhahz86AlPN9ZwogrsHa+IYYlqsAryw2GZ2injeXTO7FAVkbR3O7
`protect end_protected
