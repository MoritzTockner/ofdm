-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FJxGOeRg1LTLCncdH3PRb6VjZ0hBnyD37hqLJcJerYDcgP8vGbM9oEbXg2tWRq0SlScDcmhzxN/H
hM7GY5+YENUGnnlxoD8//urcPFpCQA82Rl2bNrcWkI0zfQSi5MGVg4CUyaI/fCTdR3mN569y8E+9
INEGvOLqM1Rcdub5CX2tA123l4cru2vhubBRiKWxk0kyKVOun4ifx2xlXiL4MrdGRysGmWB7XtIb
qoSRIuzF0pDfSfIFlIgNlD+Ow5hkBjaaikVqLndKhEfcOZIhYJFvL0JjXqX9o5FMbGZExqJkNWLq
7/EOBMdu5ZvBseX0WqV5nyPvPymce99IusZNZQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
e5uoUSoZjLXc3FStzgJtRUFn1GswZw3Dx3nn1+//FZrqZgRwUgVF25umjghlC904S1A1eqC8qgkQ
NGJphDDTvx3kP0T2O8dbRDDv1dOsC+9bG08EAY0C3Ht3CJSU2HdAJU8/ctbOZKvzf3IlL2malB7r
KuHIltW5+CMxa5Ni6pODTWZHjRCh0jaI3WH1aJIg0z5wSRngdTKcBeubodBKcIymb2onut3QPgwT
yBaeU9+9YQoRGVS5CfaLvUQF7pn0+PL3uCbONr/A3kB9c9WtlTPcbvh3iPVBmZ4C1EKX5CXa5C3k
eG24E3AdoZsvg64XMPKndj7X5FI9+PpNYFcmUoPTKi538W2UpwH8nCdhtCTsPBxThXNRTdLkNDA1
iJf98NCTZ4+ScxCk9C7fVGWUz9q87GWORZlowbazKtK3WJrM/263Eao/3fpZpZ4iZRWPjRuRmfE+
vErKIdwFt3+HO7RLBIzfsgBXzXGVzN8y/uYT8aIt+QCzTJYnfu53SS2ix+O6DcjJXqPTBIeMrVvY
yvWaD9nqKzQzNBRH1YRmIvprMWJdq9hz9RXvd7OTiwQUK/FBUIFxF1ZPyI0kcXs9pW8ImU+VWYgJ
EFuueEXYNkYVPvnWbgMfQEqeaQEepcl5pVQNYR7jHryYu9za+czy4Ix+7A4vofRUgLRQgzRM3IhJ
TkogEd3+903fGkNE6NFxybRhSUgcaoIJxO40xG7w4szAN7wQaNCHdFNXgu390yTMzaDSYxtQw5I5
tDTB1DfSl3g8S+TVMlsqweMQRqMCuehWS6yDjP+ORj+6ri2XtVbS68YFRu6v9dJ8DXqfM9CNBl1g
sT8MIK8zF01fL4h2IdU/zZ9lCJuty8254X64aH8pJQz80NyCqA50uTwR6qfMZ2RvT+8Egopa6iC/
L3o4PT1Csapv3xXuCI0CnSFFoAb7/SbogKwWnLsZF5on4A81QJDPcPep6kXEeC9yMD9sSQMD0wp2
SynFzoGshMHfygbh1lnjnxaVpel21+pIyi+iDq3prD8S1D5BFvoUrDqV3wrynI4nnaKoY0gKGdlh
zmSPLRKdqBb9EuB1x8o2UYLbvNZgHfTzwZ32vWNwHFnWz2M904ZeNzi+vpf7kVs4C02x5tVUbzPS
wUOtlBE8dzsFPnk3Xq2myZ121zuvwGwUkSLZiCD8T/HKHEw93Y82JpkvaxF1LVsyUAYqL/K19SHf
U/I75dgh5hjLvi9TODYgWRUjcoLDk+ryOYL9jEsoyMY6qvbdtkjIhfOo86KQBvrXKKPQT4XAO1VW
XgXL9yTULTXGb6k79UArWT0Yd3Aeq3/7R31rxgRi7ewtjeUt+1R+heDN9V3DULBkqaVjwTi7OoFo
RaoUFcI/H1qoXfabufqDXtwlHNxwgZ8MB/lc8K5MezorXadA8EiStPZXN3HfNEF95AP2SMTZR1kH
GlumRBWIsL59Ebi69YlOqwa5VGTQJX6DgReGn3riA5zZrykGxzLqeN4q10E9V3Ec1Bin4ROnUU1O
BzQrwfkcvmrkENVusDL7NOh7lAH2bGeE9Pdp2VRULRGboZKrMslv1M7HwA9WLqIfBIBbi+k7FqpM
HCKC22DYmbT1ouL2Qih+yoj/Fl6i6L/jZgfFt0sD3Mgmq3DUnN9iMZz9hGB0DN7oFteX4Pjto9XJ
O/BK+HwiV/WsuJs+T5V/BJz8VyB7YzFDd+ZS/NTnH72YfEIfoOgcLZPHAtNpT1cCRv6hPhOOl6lf
4G2OfQ+QmgPJjcdoegiZu4vrcPGyCo5fPa7dGUOeiea+g7PgG5KluC2q/KpA4/vFYrUNhT07Rdhn
kovejbecH3a8OfKVkLG//OaEwgICQvgxKHzMvlQ2q7Aw8Qls8G6dv8PyrMXxjUoU3bND0g0p/6YU
OonBGqADdd2eLP0t+u8WyQI4wSPAO8WwDAABUdZVuN7ksiiYw2/bfOScMZiC2MFjCKY2xbHF+o30
WzrubqqB28XhgkE2604AT7PCqwUUa9IriWPXrCAXfm68nrD0WQxnJ4hNIpUGvDsYWiigfRvYHtxv
LPZbTt+4F01YbRPVkX54i7iiaDWQb0n2xd1SO+KBphwvnImYojMFCMy3WTiRzALKGmOmAGRnnmVN
SSiambpyb3SV+RWsfGAsE7kfBrdffOuW+mm4RflMHvAyFs4vs3uW6IpJFdOolW3Axwdb+mHpik4K
ewkqIG2n79+QZKIBPPmyRrmbhF/5h1PaC3IZwTpH7m4F3sKOaRUtpcV8LtivbFXazbBfnn40IyiQ
tQs2Ior9ZqUDO4U0oK8byr0O6BtGZdUlUz/Z8Y6a3ciVHWoVfQjAYQdeTB+4b0YTRICeuCoNLQYJ
mZymsJYXHzG6e72Ckthw9sy5oYOqVLo2w6aHvje91lTrbqq3FeBF+e5BV72FIptwq0ccb7XJAyUu
eyv1mLMYy2v23gUk2G2t/XUC2GZOQerArqr332FUlrhRWJJzhdA9akLd5HeZZPthcUD06grKl1GL
gsdjz3gKyJGUufThuSdpA5ctrXS8nwk3L20zNDagSHNQIVQeJ5PJVQSreTUDq6MnT9XWHNBME218
uHvLCKHZUWP399ZZwoer8yPmzuvtlN0i1CeoNkUC0hKbu6S2upsvV/z7Qr5YXzdZ/uik/f0ELsGt
tjNuDVvsUSiI0v/JOG88ek3zRNpUPgAtoR20bNaEjt4LOGRubKLvJT5sa/H+txkCdCLqGyx7b5kV
P7N0AICNqo6JUSwSkFRiP6MxCT+o09pKfZ0zcT2N7OJTRk11Y0mhcVxZXSlZj+fMcAvQC3gIednN
bTF3O3lLQUVemBo+rHVlEepjr0gx6tO/jmv+GJV69xVVYNduUnoVf/6t/IJcWsBlHYE4Cx6ntTy7
ZdeGobEA5bll/Rf0I6FJfLzjQNaCgYT/0mfntYPkuOfSpWH7Ao2QS1vzD2GcxXzSClSrzkPnpHuC
qYqcWIPrInri5T8ayeV6ClxIGY/w7if5Dh2y4CC3VFzgSV7+H8CPJKLpZvNuxYXflCQ9ZVGB0fAN
s9POgK1HZrnpj6hXVAqZEQjtw151vfsNjbsCsKA0+2NB5KkHA+jxz5Ffkc5iRYjNLjNYSp6ZuorE
es26lUxodwP/szqg/3hpHmiGgtMRG3fO6BCF5ZFaLvysQuVtK4hkYZJL+MZdUSDGubL7fjlpg1ir
8WeF9OjXzffmt8bZdSjBZ5xT19Ixj6TBlQGGBvYIPQw1nVk7yGL/jMXo8n8Nd0rkhWBWrbO6Y9LP
h309dmvvGoqSt68yGBKTczHDuo2Y4eg1ZNNtBDqydgZNxMpPVO3enTZ20ARqvgEhFPHkX/9tV3pF
8MM0giHtvQMt7SIK8KiDZYiL2djpYxPP9CXWKoOdiaGMvXwW7b+Y/LclsguHD2kC0kuhjROPH1gH
0+HCduOcb9GmjmwCufh30vdxFeC8X/ZuDXPtjWgZRE3EatrJCnAyyc6TBcb66waBGv3K23a2R6GL
BhWWxvtwtO5pUb2DygccOM5ILYnfWjVh1TyMldxsXXWclEWLsoXKyOYebsiGoNBsZO5hb/CVRBe5
iWuYYf+jwb5rGDV+A6ObgMOpW2d1ucBhgQC6AQBsiic9JoMbXe9k/BV3U928OWawLXAofbbB2U8K
30oNUHV7+X2U5mhdID/Bpyot8Y3/SIsFX7wU1hpVMgFNa+tc7qB4DGIAtFC0DEAazIHSpyccONIB
YVvufS9m9E5F/N+x8sIl9cPa0wXlUbR7PtjHYHFz4oT0/XSjS7YNon7nxtEFPO1mR1epTTcWQSpl
/VyuF1JTZ60g2ANfq5S8ibM6o5gzEuFW7SlnvmivHNbsgE1HdiEiGtheVjvTz9mdN/cgLsnxTkLH
Ac5zy8F3rRjGyDWkCNXM6Ai5XapSwHAkrwMzQOR9BwrNvlYvVczW+eFewupnKDqFIpKL17u3QiAG
sf2k1Y+x+GqQdlTsOnsHVqjL5poTaO8Pe6awWU3Xto/jpEmMMSzwKZJnzgdHj45DIaXetiwQGabx
/wDlbmSFe5tfGSftkHoPKF9qdpviqqUFBAL/VsK/G3EoT2ri3jUt7Ny/wWBxMyyrYTclvGlUAPnN
C8Ewm8oY/e1/XJRGY/ZypEHesfwNaVaFTOPgOKysLzuFNVR9yXeSJZjvyw7Ccv5m7H7PjJdqp3ii
6t18sfPhXFPakrYazyxSEcFRNWSCjiOUKm8W0DUw7dB/N4f089/33xje862Wf96VSDm1gTcpIm4h
3ozpI+syA+H4+hRXG0zLU2GMpIM0tY9Ka+eZSNzaw0ZFoPkiWRzOFPgrgKCdDQP1KDiqyNl5bEDP
igYhv/uMq0p5UPLEz2W4MYX3G9f4yNCHUwaiTBlp4fWU2PdxoKWnGj9DSbvOopgUeRCho15GbaV8
o3nyzH5VOfipilFtzhuG63BjGqnwc1T0x1jQgICP5r62cpnw7hFPe0kOAoyIiB8EtG3IJQCFuQ2C
ejK/TPavftQ2aI+ZlzlTELnU2q8bYyfqnlZCvujDIpf+DyIu2LLSPQe2f5yNVsH90AbU2rh4NIsX
uGN9q/ZKfnEiYeR/14VgjhnDYLqLQ6BUjj/P/ocsGJ9TTYWD8F4ZBhaZLATDF+NxJ5FGfOAAzmjN
LlTD0E/SNlFMDp2LLJDlrw7evfBmaKpQlv+w16RFNFRmzq8Cvf8QrfueHav1uOLTTgbQ350pUS0N
61pH3IokO+BNqA2HQ3InTZSQKZDVzMwTIK/C0Nr4KfMVKdRjRhDql36G0ZI4T32123pDR/iDAMx6
Mf+0NhbsJqFv3PNKQE+rQSe22ae3AANUgf5e2CK8yWikdCIKZoBelwpxhdhiY5snGtm7tE/Vj20B
vdQaWonaQNYANI1XBPUeaO7Rnu/N1UZyLBRfxkUNYiQ4hjsXH8DEiqO7j2XNHa+0bend8glVe1Hc
aP6dVgapwC06LFZqcHdYOs8delsA/yV8WvNqL+mTbUy/Ufh03POhPQw+RyUW0QE7QiUR2N+ncRqb
YndFYH3JyXlm/NkKDOWoRPUdQOZfeLFVOVxRf4oHtUepyDni2GbFEJcGg488+GyYYfWCKts334Hq
1rYCs60W/bk4oljQcp047FRormnQqFE8nn4zhHC7sO10t3/Xyjm+BztF03zLq9paKADDfAeJHpAf
R/beYHOWxdRIvameRiuJLBWe6mphE1XrcTBg8AQd9OIXepr2ZguWr4k0TvaPz/UkjiCEEgmoNVeP
cRCYkRsFaxQkYFPDTczozArH5iaGGVpEF6Q6gOiGG33R+hICr+hPJIvlaAeWNodGO8YHvg7DcySN
RiTghdrqPCQ7SgSdMP7Xtl5c5YGZ7WDmmOXBbOwcetAMwwJbN7RrRf+8EeHAsIQmTLLX+C337ISI
sDHI7MOMxAxMB3Dwis3trXZsZUiKwkANfaCRob1E7mUryNJrS80tLsf31S81Sfc5YMrpb9luBv3X
MFtPIi0filUvzaZjNDb9bZcr6/hC0A09VCV97553IIcNj0uDmkmPqJcYaW+hXSDc5gY8OG2XaAEQ
DApU6g4Xhd6CCi8QZooVhvo/B1OpAVvX4Jsr7xZmVnknShnWofPVJPkfRuCdzZgyYODLeIL+LkYV
tdwdaN2c3zWO4a8IyfanXF4gBYpTRkMA0tP0FFzlWPLCX+IVnxcyLV5EEI7okG7gvqaW8LV0cdNT
ysxH2hlDM6NKYLHKh9T219wswQjamV+ZP0zL+JVHwiSszPHGBxxofBDqtP+n/xCBcY049HjcJJt5
nuNqK71jPqMvTq5PTU7ffjsmZenOF1HY6BAOD7WWOM3U0CYWtunogRBQBls/zZXC0FFsSTZPRTKu
txFhy1RbrFt2ZIF3gS/+mMSTj4JhUCDjanDs2VOvlOX9kViIOYFOf4iCKZvsUfQk2zcbX+TLDW35
fy+S0sQIFN2uankaiHRFupTSPaZ68uGcPw2ZL5qDWjmQP+hXoAEFDGZzXYloXHvwctmzZ1SMFAkG
+YBBcUHysv6K928xCX47DKeOw1xLGmyUZwPwG5amUXPpgOXCKrXz02aXMdkpXKVMzQLqIpmrYEhe
neVKJIZNm7a0A1SMU2FDdSwd+GpG1URS/u2JZkyjLYsPtB7/Z6dRwovoTtnZVCGoV79fiYeKDXLX
G42JthOFggJR71UTjbJ+2XYR/X3R2ape0SwTA8ofs+n57nZf1sHtYSmN/MPZntHtSQJB6GtL4RFd
gKM20HVVyzaiNx8XuD+5bRAeqGDy72iey9sIyNrHVhLQTj2sfTq/k4OianUqoGaQmUx4WxHP6yzt
9ifH9memZNWjC+mtVGVrCL85/4DyVX/eKGB43w49F85/Zr45dsVBY17lrxSw//2tuL8zndp/CcfE
vCKS98YcgzLfdDMYOlQG5egrVuvv7VNh5Z/RlHOsN99XU2wRGIPMysdsAfackxUbSQ9Lx/5gHEF6
TGIQLAv1glS6jv/g8utq3JyCRSJCgRSq8bdPfeY09cR6ERPim35dP4uf2Gi5XkXNsOOx6dx+q8hy
TtCSuTRavvy12aMgdphYSKZmWYXwxY68CmCsAOchOxc4921bI1WVejEUS+stV5p62YxSK+qz7vid
oMwLbJbx5V3tJINqWTM4MV0yMHcQZgJHmIMTE5/jaRE/cwa/6dZ7Sz0yYaVkYTAhjP0aG9Xm15RB
cjKQWEVjRw2qltUB1aMqFn1a6JQPcHHYXS3ugFvr52sBOUviqYi7Z27KkRxzdu49LXlQqnhpbfu/
bc/4c8eBxcbQP5Eb1HXhFe/Z+04cgOysGSN0fdwwiktzxiNPyOpY3CDHnJICWcxVKR72fPGBu653
lONRp4GEQLRCMBnoT+XTY09VxJ+PEA3tCxLEgi5iVwRHlmpLXdQEpvoUwF7kpq6c0CoAnntFjjvy
2BfVEN9LR3dF5xUA+XB8AtQu20XjpBousmK5EyjhyDWmVW8iQs7KvuWjY6i+mg+mv9EriHDPxW2P
6Hc6bd4Jfh7Q302EEiv2O72XlersQkcZ3WmSlLw+m2UDqjQv4UyQYwtTDRlu0+smhVPaL/8oqhOd
13J0CvMmuqHT1TvC31rf18acUr/sQmnN4ax5GPNrnaJRj0WUfdG7VgYnW7b5aMSff5tMsX37vIDj
/zB79UUkSQKRKBwIzTg/mnPFOOAFHaaRP6Fy5shOP9Gg5oMIFnO6R04fJnwYTfq7k7bTZ54mk63T
G5rvrM9yepbKCNcHpz2Ax11kDf2PUlgIH5gyhu6Eo6PKq//v8xgLEQ2aIYjBj2S8FNw9l033t4h2
hYP4xBGvs+2gZwzn4xHpUBzF7kXojpR/s6+YvCmiZqA5+tt40p9MN6WDuc5aZ9Sbfvve/j4t9wxH
XODY5w/JQ5xJ/xx+IMIwCeWA91lbQC9kwZ9viobyxXJAAYY0dvF8YfW9d7R6/E3zyP0Yuwo2EV8u
7kQqfVjYoc/MoaGFWQ5D19Hx7zbLNBSTN1apvtLVXTNDwB9WIBYsNPBCcV4gN48uODjcey0y8F5m
XrvsI0X8cUXDymzB21DeRDKtsCyNK2vmCQOFcKwHzv9pJx1lDOngVuNJR84Ts4gc65qXgAfFHwfs
7DhIxQ2AE2orR39X6PVhg/2TDWmR+cEZMoVhn0qt3ZRA6ZLgf1aAq2hGc+RicUPqrqMSzu+khx0U
lcdlA09wC+47dso46yowmB9089RiPNh9fk25nKpbXMng88BnltLQcKRvbUBD6Np+Z9S8wj41NE2L
FarKOMD4sct7B5q1XNDxnX8LaIvzEm5QEuEQvkwDcGzyY8UyygkE3ygHTuwGLSe5ZHiUd0bVHSgL
Xeihv51pWFccIq7F4Lt19rDwwjX7Pcdj16KRqYUTB+GdytfiVXSmPUBtY+No6xHwzgkE8B0gRsly
2MwUai8e9BLRijxSXYxTBbABEhXP+wlyWAp1GoD1rjiq/Zgpr2jxgPYKU0epkf8XxOlOtbzdZ7PH
pQQPlL58a1lM7u4FsxrEfZEzNwAojb5mEzrUpvzuebZ/On4AnzZ/4LOeqysidJq7f5Nlee1SrLS1
rM4WaLovldwYR4Im/3r9e4UNEtU2Z47VSLxPr6JvMIl0Ff9CLAJ5C0IeM2mrs7wwGWN428SxYP5o
c2bX+BiwF4ZQMBF7KSw03rxFvSKN917X6NPW437mF6Uem3fs6KqtctTTI43ZoKz9vF8Q2kuCTBhM
jky6lxQJGPHPwnPOQ630IoQkttUssJ2+E+U/N/zb0qMfO85oefScb1ra39ywCuhf+ONU/xUhi1Bs
00Sqfxp9ZJNB24U8C19riB6rsE2qybPlNdNuZrggJs2BDKiZNYMRRq85XLAcSUHsGRmap5kRdEys
T3eczCX3nGW9+WuJxz0l9o+1p2zETga6kzuyScD7677T6ehiFEK/DOFAETZs4LhFxRt1rATdNaSf
zQHT+Z6gYbANzsE6+HNHsY1b442lLRgjv9aVjWyk5LhhKB7l6oCOPjMnRK8asJf6AmD8hQD53tNT
v4DPf0CnwNMidN9NcSkeZuRu92omGFuyy7vT/4Kf6sLbUajXG63n9RwcmKnm9qyLFjCMDut9gkFR
coz8htfqlWMJGuq8OgaD1lsUUUhdN35g4AaE4YcPTye1BiS4vLkn6p7sYJgETweDvwU1gxxoBcu+
Hd1e3VC/jQuIjdOe3T0aD1+SnLSvDuxb08wAiJK6Veye1QxfVzdMtwcCeogY1jaMesvSUOICklNB
8ESgTyqheFhPbkSvjWXDmVOX2KsSsk2T98Cl0BydC6UvZhI1JhMmMIystSqDXAuJSBTxMnY4amYE
5qs+OWeehWK+Tamq9gFML7nUQLno9gBvJ3iGkHas2dwBRKgu83AGPeYA8UQ0ci8F8MgXB0bsiV6q
2NDDB6kr1h987nf+PxGcbE1mx2egaT9zV9+hyLCDJsJh2hsd/IBvFJXXZjV3WLVeAomNFBCdLYAq
+znFntlVi4NGRpMNEgGIUav3EKCTVPCFCoRPInIHYUQudhHiM+F0Wug2+dyPIVll7qy89rpZHaPM
22qO9UIQY/8t8IOdKarJhny/kkJmPBJXd9FOqAxpxurv8hrdxQlPn9wJHrRMxcGjI4zNNhfzC5K3
n9vLE8tfVgEaz9SuIsdF7BL+xVgK5EYa2MHHSOq691GH2HqP7p2M6qg9attY9xHk3o6MnLDtfrIv
Lynde6EbtVvnnkoyfG1lqgm+Nz3IKww/5PX3LKE2fZ1ap8sjbig7P03mvbnbBvuyFDocJ++TGOln
Yhp2Gqa0ON1ndaPc5SqvMvt7xFwN2iJnGV/F30bt/+lqrbN37z9QdDwWDxDw2ahWV4LpN08GuvMy
U1CcfNeXnbOlKI9Tx6Kl9QOMBxYLUY8613OW9Sg4BvpIv3OhgKZEw98nEO4Lq0k6CxfzFF4ME1yE
g12HQzCPsihBkr4NvSgblogHhu58EyQKHpe/7MOOPqxfiFn6eQIQyTCuZTSg91iLze27Nr6KI6VO
WoXACBrQVq6Y3IUlObpE1vkSG3uC4FiNrwa5bcHrqOQ33qs7NlbIjw7rrS2DsVV/WGQCqbB9Zj2R
Adf0rIt3tHr2c+F6mzfZq37dNSWSJ9lByaSU+8oiSZRe2uDam8MZ75Hlsj+9V//4J+Yrs2zEBiQa
qIqaGxRORAjn/GVJvPOoyUj122y12keqdEN4VxZp0EqEspKBXdmsfKzFjSwaIb4gUjy6vvsJTCl5
FAUUtniqt+AR2JA3YFVU5g0LkTSmpUoiSFkEQ1fmOhPn1OvARVRKStUkGoWDOKoDQ9MFHuDLJr5w
VVD5uzFCYUakPkH/SKEsRDQDc7wo9OYlmFNoA0xLFgf4GcQpFmCT3Q3tpDjVmFZgxLZrWvLwNOaq
QWzf0ZxFzyzfPJ7Q2bYInj2t6fFFvC2F47FHtyJU7vG1q+VbbL4JXDZOBd8Mt49ICFgZlWWJBO4L
ZqafoLnmW1LJkInREjqkd52hhaRbCxwVDHwvxgiP7Bqyr+vvfP4eXqXrwRj8VB1K345aET2eQZWf
kSCzqfQoKiJtnY1nZXzg7ArxH3LH2312sLebY+WrqyreRj7PJBVp0iAKIQ5MVI7QIrJvKvWvK6kc
hvIQyWojy4V+XWIbkRCJzEvEvviIA9F1vqBlYTtgimPz/mxsbJ6XMCcFYGpuHCPIS//Wqslxs++f
fpt6cUecDlBltK9l0uKOdCEFVebC9tiy91/XYYRnqPXkTHfVcZBSQFZZ6+w/8k9Eabzwo5Gsv9SG
6n8hF6jQYfO39ulviOVHFxuKBnjUOpIfdtaBREpWsK7JxeL34S7ybHWK6nvVMXW0fJrS3dRp+Q+H
MBtkuod2wJr3rVko3bLTScM6Wlmc/SUiJC150CeNtQMorQFSP0kilsqv/BxGSbXOpijXjRnCwTpX
s3oPRC/VhuAllCNml1y24A9+tAAGPNcZHzAV1VBGwDR04UEyY0VHu48TH4Lnm5PH6KNr2jzmxSxd
G5gg6dA8TFD+5S6isKHo+VE8qdSX0zOXYOZqjW8XZR4DzSZB9iWfXlRKJ+8ft9zNfoAj4cSUalWj
ybKLktSrtWxHUfEJkoNydM0/+X32bdSUT1nU1x/goOlsAYHTtvcdFfjsfovJbUa5WCB4lM+pI0z/
4GdppLgjw/ZoV2CQc6vKKBytP8Gc7wFIXvfMkFQe2wiJXWkcFwFremDKqYnUOM2InixEX9+EJTd6
6yODyL/HKN2TbiGiMrJiu2Qx6jZy8Ni7QBgXH+Gbp2VyWZH6udWEOSnJ5ya2MMZNx9HatlaASW1p
/60jFcbQ20tHnlK1hBD8oTNgWGYY1wDiGtcxLAtrWfMWqeaZ6ms60p+WFStX0MOBh3mclNzYc9PV
c1ngkULtK+7ie8pfWGKpL99tNeFJgOWsRoojD+knoNzK3N45/cf++XjJMeui+bKGhU41PGo7dC85
78hK9+0HpDAS6g8udTPfbwar6/plamDTeJ3MrruwHnA8zHlCiALXD3NNzoWzDelCLW+iz+6Jrcqv
ta6GQZsfiBWXDiK9KKqOV8X2IYQmzzSaQOamVo4HigDTOeSmewpSif3C1uL1X8iFAgAi6pf/oVfp
Ms1bvQI74SnMEvMsimms+1fGsaCkzKOPXsItmSR3
`protect end_protected
