-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RV1qKlFyhP63HRK3RALWLe5h4OaP57tR1M/UdxiP3moceud0Jyjl7cOqWjlVgVOv9LEdR/vpEsGk
DoQS/K7uJpw2Y5FttLQbDp2FLFqodeEZ9xhsoJHK0NQWIYycfHkntY15D6kic5iQgqBEdH6bnRt1
txXROyIxBIPb3Y0qbex16NjigJ0PjK5W3ibdvBSQGSeOio4xbjuKWdLf8UZFXka5N+LF+qOX0+BZ
d+cZ4vQdXy7DFdRSwGtetEY26+BSOrtvXRf1MBC9hc1gCIKesXxDsmHpp9+bBFjwXt93A1BkdKH3
V0p6inzPgkFhv3nqXGQZXGsqQt59KLDn12pATA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
A2hh/Jvnrpq2arPWEvYRCirnFOAI7jR0dRfTG0pBmesI8VWG9+Z5VQNQw32OouS0xE+m1wPcqdI7
7WrE/rVO+I5ou8iHoBNcf1/DneKHjeQjejPlerqfZmtnKR0dP2pYSLo0522/W+j8mwUKgXL0sKoN
Aik5qpONNS2aznTbVInTbwJBTsiWut3SDEo0tXD6A+rv4eB0mUkOi26gJuSz687vqe7DzUeVw9zW
qxF3iyAy5qWx+spNk4GmyTibjz/yeePCcHZxdYOBmLdp8N0VzcDLMts7Gm6h0CxA2mb+e/ljovuu
C7AAHG7oWmnU/GHWb4cwSIfu4aZlHIZPxF6TBspLJFv6mTu/KU8kYNNfysdL8S7xtINURTjGSsYK
kdMLIZ941xRjkvtmsv5UWNW5+9ZNVw+22D+XZZPsEYzRQsXXlyFd4f1euNYdwZZv8mdvV+FNqAyg
1FLv3k05biwwhxYA36xjORrnmzi6kxiukLfirbglIxSBlHR3Nhl3xOaweULBfYrW/JMkbq6V82BA
XO4te0zNP1qRzkQn79eYO8FqG07abcvXy9Nbg1St66UO4ymxgi5nGESTwQlR0InR4LJq4RbRUliJ
hMntlkr+RQsK+d+c9xRg0e8UgUGsm8sk9kP8NXKLDhKt55k4X/IG3YvUmrOrJ8736SUdYgEM2fAZ
Xrhzo2wJmPjah5QTddP5Cgsx3A38JrYSQ++16L/I+X8xu73S8rK7sfoW1n8KZkFWWobj3geGqltE
bRk2L447kGdA6cVYiFCpaqC8+koSLlxfWNjo+wbuHgkZt77hsn5Bva2aFxa8eESUtAa+z9kvYzgl
Xm02x1qql1ujuR2VsYn68i9Ag58Zq/51VkX5UNEm0/sWEbPz1euDUztXib9CGWiAYFfCVSUvW46C
jdNnVoB3GMYxxFsYaOrRM9nBBajZrTd6S22Z/cNaRqsPwKnZA3gEqgJl+GGmYbxJYRfBFRUmIs5T
LPjBEd4QxPcC7I78sMGy2crLgo6ID8cnDInGbzJB5y7Y6Apce4E/y5inhAbvnS36qxS5p7wZtIDs
JoB+YvjsbHWOLMlrBQRVw5qA01CQ6U+7qZEtPs/Mc7gi/tOXXgbVCxy5PpVwYuHQYa3hDyX7waqi
G2aRr1MoP0F4rexrLNoU21s5clNKgd5VQXxypW9vBrtNszaDnjk1+32Tb/ywGzfWHdLLA9nAwa/v
hw/3M8ThWFjVNinLFZv4iidOPEEtOCY+sVPc4xQFYPFjjXIpBc20Pqj0nhPg8aJT110QW/1J1INX
UP3XTu/XdwFecKsOFePx664QDwRSqEHCeR77f8G2yGYCxcB91Ie8LauxITknVE+K0uzFQv0o5qe/
hBdKeI8Bhqmv21Pnlj5MTl95hqNhXMI0YwDoEbi9JzgSIb4DvlGFtYY6AhCdXK41kU4h9fyYs2de
Ja6IlS8qW+VmSNhxs+EXf3pePgJdWpc8mK/4h6pg/fU2ePtBWuLLeOtRfCFSnK6Q1tpy2M9zqg1l
rANgLfTe6JAjTUu2kqSGzWhgAoz7nSJ9xMoKGHAODbf8tqJQajycWWLCg0m2C0+4toNGFNV83fGf
woXZJWM2jvFrQZ6t0gMa18AI0VMNo2M3FI4XNfFGa/FkXh0kWCwIL56uekQ6yyS50ekXoJIFwidt
B8st0n6cAqKYsrxv8StdkT95STfysG0d2JzLwuh8iTIIDpZF++G09EataXRZayfJzzZ9oz38BBg/
qrPDY4rhzKPYUpFBllBrdJYG1QwYxQcXFiSE67hrj+FIrz9LDTWAQw9QUA8TovTBCOsG4Wq3eT2E
GnlGH7zxy7TCcuCeBe7OOe4WjlB5F6Vq7RLs3BUFtQOVdiEY/F+juyqmiofN6EEtgq6uAefhDOCR
RpiPhOdMZumqOVrf9irLLJrK5LbZtVIeQl35/sEqW/eOIgUgjl0UTAHmPeciR+0Hbq4R/IIVDTFk
UfyfsQh7DDjPkVqlSDmTSIl3PASH9R1DPUI2O+n0AmrbyvbNNykSvJjcc1pMYgjsr6DYpeQzN1ip
oVkbSg69ToDXqEk5ZlvUEnTtX4UYW9v3c3T+qMQ7EBMFQ6cneJ8tdMuq1pGfyNl/FKgxo1jO8qii
xIdtrALhFolS9t943oK3rZGMuHEfJWSzSkihS3145BlDzQu6luHSYKfmRg/nwU/heKG1bbtFFSP/
M2olcmfYgLjK+GB5BjDyBYJ+pTYgegtn/YHxgXMmfSh68hy7g6qxe6u3j5L1SLgLzR8H5+glnBQK
eNS0xt8Clkh77mHvriXg4MX0o7eDsU84WbK0IWJU+AkA1Iw3hOQSvw2e6lRo0at+sBQACcgHVh/e
getU7iEDK52a/OI/hw1P1vJ55PAAtGoOAfDS3WqcAcVpVByVuc5obGq9/et9wNTA7b/i7ZVTuuzt
Q/VkrZLIWeTHbocZxQzwyegR11JMVt261/fPyB0D/5bVxbKgSNZ5ysDBpOLVcTrw78DCsjAfvy6e
RwHAqjVVyd6E0qmeB+O2HMyQbueu6zTVc/Ht9ciyXi3U8mtunALhvTrhrE7refYS1huSHYMbgtha
1F2YftZYak54CisNbwDiPPkZPGCvs8bPdHRcD6lI/savCFUpLLu+csWXYEgdNrx/s2PwB8WqsG7K
qhL5cKX4DZHkLhSZnPtfN+c70lwhUBe/9wwtuDHbG6TRG3778vtqy51b9aEj6uctzGvDRVQ4bRhy
EfY0lwVlpVIUuRq0tfORTmq4EpiYorL4xT8G0hXqp1fQe7BI89R7axw2GP7zSNWhRnY+u/Yl12zu
uXlit+i1Y+ZDpnqiFST+5lgIs8HqwvUkK4DwEqLixO+Vt+efjvqbYSTMiW/sp6YeZqx4bA2zpfYv
z3QYOBjDWXHJ3k25Rh4TlsJTztGmBNSGr6wXHGX06id89HOYyC2DjfmOgGg2S7IC6vmIiiHAq0jK
FhMCbjieD3F9MrL+/wsfBePyUU3NXlV+QDSznfochurWP27L1mRtJ1M9ugbRtQRr/4TWju8rBQLd
3Q94e8Gx4Rs0SIB4/Fq/hniy22yKlqwvgIlVQ51VaQvbJFmhSyjkgyRqqFz9TtguoILc2vT+2PhZ
+l3euie0JESIXM6yEiSvzPdVTRZA5lZkHkj09KY3JmHb5NXvtctCiYQGEUzuOOxGTOfeziMWSMal
m+DaJjTbqXdCC/PY4YOETMs7XwiwJGema9/mgoQDbrcgdQQ5d+3urHiVPqBD/g6EvaU1YDgWHY7y
3s/GP+ZKVTVF2mFuEk15WZODWqa+O1p7tgKHjHAdhsh+/RdB1NRCc4d/Km6bYXfPX9GAMvBbaLjO
SWbudpgWnzZ9lCXUhNr8O6oFVznsDQ2IHCbf2ZWci0GJLvHRKfbZqdBOQ6m6HZ4YVXyPMbHKlYlV
00+UJZocC+T6ciKnczVVhurDjnK7AkZ6HJApyPo9kSQeTodMCLsROYcwcUG4MXSpLHyuFtdhxSim
7K4OVzq1zVJIcVTJvD0hph6WfILBXlzfE53uaS7Gx7l3skD9ofvO+32CNiHi9wwyQ7xKDQn6yq1/
91Nqq7z9ptqyrD90NMfzQoBNZhTcnTKtOnglab5Xnyos3hV6hh10cN3rLiwl88HS1HLrRvWegQu4
EseU5m3t8aWLfL7lmoIFyIzeTJ8Cf0vdLBlELwweXh+6LlYC/4/+vUMYTprNz84GDJQ9tyG6H/28
AAPf6X+/FTj2t7d9k1CGfFfhC7QqbAT8Vsv8rR7OYj4T1tW6u3l1zVmU0CdU6SW6TYXeKfFe8Ljh
Mm/d8JJIfrowbJdnRbE4N3cAJn6LNcEUALuBu+q8EONfAEOMYTmlMfMtWbGg9ruu2pBRQZcZbF+Q
AM6bOWh6nR7oZenM2vDsBKHCfSAABDY+wRogt4kTU6vmUlysVBoYhzppxWN/1pjMnI3RrHB9ojSU
PPq6enCh91eH5I8XLcLXyg92GfVOK4n0SHnvyn0BQEJddlkmC4I8YPMCHAQJbzHD5yBCSTpiFBC4
NbJeF2MRZpVe0MEMyReUr/ECGdLR+WWD5mvUqJQspBp/0l+zHT1dtgi6DU6vLaWoSOogD585ym4y
mAhQJdjlqXZ+3MdMiEtO9xWrdlrmuQyhgIQKzPTPxbyF8WVElbRdweMFqkKbhROCBICrkZAgn255
Moy25015IGxJeP02Ny5/l6ZDiOlqREo8mPPF7k45ECNzOWgtpsCOyX9no+PN0LPLiEWMS9gxSSge
OUBBmeQcl9l2iMFSZCejBgjvhnt6Tg8578x/3exWOADkIF+a84N2J2fHWE+nZmx3uAcXSO4L0OYA
33UMFMbZSBhDR4f4Mt+5d9mwIdrqE1H+d0R9iW1+1pCsTyKglFNmYt9OJ1RFvOY3YSg8HMLF06yH
Zcf8YsJHHzRoUlVU0TxwqAoRmU3a8Exy1UnNdJc/rET9voR39UJ52geOK2MJpIno91N31dDLomQJ
hhDPsfwTz86irh0p1VvvbhSi3431MKB43OcwmUD4z79+w7jGx71/l6hobobcVaRX9lpghQc/4/Wh
KQFvfqAs51o/iLSuyEI2RgKf4JvkPuWFvChLHBL9xcV/H+DvS/EXIwrVrdr4mUtJbyasJVvw0L3H
ZJ195Gkc6ZLk7ksiQNiqVFZltB07GI1T4CF0fUQ1MLqsk8UK7C1hkTTOHEC1jWILiR7L+JIi1D9r
ZWN7N5qT9idHA2qborCA1NtoAKH0YFjJo/m+ri9Lh2HZ+pmsnNiKBFLIzEe7AxYZ5fllLrwP46xu
8a+jFerBnD3OztBKOiuTfgfjrn/j1qqFwWmCwkeLtiqTSSDJSpSIQUZiV+AEdCNnr8mmTEKwATW8
vN/5EmjQ5CvxtebKFD1SiC0B263HvBJrvQpT4UYCcEzzVt+MxveXXExiwZ3qQPpJ5u4E/ut56rgj
gYKh4PK5sd0h5x1K3nKu2QBAhzn0qaO+68cnDc+L1RZwWs1ZLI0gGCsKQ6jA/RFxzSh8kz/Pkoyx
8xOqilp5rbkGzoNZXxXwRBg58RpbBZ5lEYfLXxjW/TMyYQXol1mjeOROyK7nVvUVtviAzGdgL57/
aNRaFUFsGCuJqwGb7RbusuhmSQUMNiSn5tYYzr1R6Bx75NzZ9uqqnfHKrPj8X3p9wCTc7ism63ts
0LgD1AFRz+g2ac2Pt4MMiC5rI77AEoHRH5ZeAcQAD0N3l6JWngWCVgvGVkZ7fxtCI8N/LRKtDw7U
uLAsV426lFAhXIOCp7MUz66iOi+44GTfor8YriR34rN7dBcNVzomElrRyGyWtEd86MrDF/UY34Wr
mzRfYyHB4QdkvYmqaY63Hb1Z6RigO9GcgJogYc+npkoeXMqOS4IUa9X0u+pk6kaJt6fKGvMq9DOr
UL/DdAi++533QxYelygRnumhmMIdfD19XhOOCF0KTRthRHE347mq6wZtsmLc6hqyieSQkXX4VluS
EyUD/MqB38dKz/ZJma/Pr+8nrfXDzZgW6opCQ3vq1AO7nK1qaTQdvVdPNpGbe56GdXIyGMUGxzSS
u14wPCGnzBUevJCnuL4CkKqJ1IghjI4/NFJ/2seChCiDR3KgNCPjedHv37ZNy47VdeLzgW8KLetH
xGkGwRuQes0UMYUpRD3Klb1O6uAjjWAnuFOVqw3IAU2+A4dU8Nj8B+eV9KaRMRNWcmZegQ6BXxxS
PCttCMDs1VyEFBk/uAy7T5D74d5S8TEsGYQxQFVpNcA7xHttdvQi+OzVhPZ4wP/2XOUl0vk6s4ON
SRlDaUjmgcwL9qCAAaeYszTQwSpxQVYKS2pZpQmU29gSFL86EJGTSn9St2qdEYfW+QMxls5cZEHR
+Ji6NPIt5m34gos3V+gdzbtCSB5rXah5mNaxcdIJfExYZpfwJjHdT3o+QJ+A31Y4Al6YQ++xgRpZ
PSt8BJn73a8Mc12dz+HN6qVqr/6hH7j/CkM55p2W2F82tXYFJBDY+noIGZ6JpVCz3FK04OrGUYU1
eNSJb2k/2Rgb7T3k9+XDxSYch0ugw+rYW9VF0gVe4SsqC4V1T8wxM6nRDMpvaqL/JUgy7GeSV1WL
KAO6eWXx7jvm0yxNE7gS1WU4bk2TdAjhWyxoj3w3IUZUVfn+JM4EJ7PJJK59UnM2Q/ECHg6khGwH
1zszC2NU4WDTvZVT08v+vVyQOHntNgjRoPZ1fL4jM9/Mlzb3nNJPo9ukShQm5Bwv4+kyPxhTRyGB
5/ygTGUif9bTMd39N+WSHh9ldVqEgwBy3ae/7wEdiIHP2hoHDSAkhGcimrkrRIVghmjk5VNEH16K
KYat/7hsLUIDS4kNwcRMK6OMKtPKf+0CWJ1/DbS7MEuF8WVKaYTfTtPtCyKTtN27NzNGc4txqE9N
jBtM0uKUp8Vjk3U3x9fffBfNJ4A8Gy/JMUPPFFcOuBrK52alCKWrIo193Ps8EEkym47MStNy/Cr4
u15RqFRpReH+m8bpcSW0MaY7YEGd2fjdyJSnzI17Fz2x1EWfwdg1LecgOIw7L3v09tc9h1/5myLd
n8+wMvIgdsDsSXKNi9tS07Yevh6rAWsGUJdMc+co26v6axMhqFpy70sK32xw66e+pkHMG3nWH2gI
DZDaq5Jt+254P0dPBptaymmrTHqTR99QgPPGdkvhXbjZOowztQraVQ6g1PWJd21MBLpyQrl1Q2A3
kdeeSRUvk1jMVjhLCogjs/PW/IahDozf3J0MB72Fiyi5JdisOp7lLQFFbRs+pZ1BZvkB6RU4mP7e
z/Z2QRX3h6TTciHuUIWVZotiZtGOHXqcqNi2s9V8xxKBcOXk7FCdD4gEOHmPJEpADuj0F79zJ4YU
FYmr0UMWNU4NMY6Zz1TfLMCbFtXmWdePneovffjPpCOYiNY4mrbZLb1FdQ60YiOEirUbuQ5e4cZt
OFsJTZmpXHdg3M6NmdY2HRRhAC0+dsb9tGPb1di2LARfu+PBlKDz8wgw6wWj4dtRfmnf/DAv8sbx
QxbcTdp3YyQGo2Xi/KBDTrenmLuYiJ+V4mYc1qWedbu2rgvGPz3MJ6uIwdjv3RDIbKtvMWOFz6jj
XVVNDd2v+nIwNjafMzOuMQ3iT7Sb/IhdDvNzMKxgw6b21iwGqB5YXZrhO6ekzx1b5gyFuku4rpKS
Qc1zFLdFL99qmz5EOKkzEUr7ktVuLIZ1FB1R7jShrtf+MI3YV8hXDQ7yZekaoB4vaZdtMBTw+/6p
egt8P+HHhl1fgRD7nMxW19mip0lbeS0wyUD24QpreJG2mNm64rwyznbVmT6dVC3m6nglSsHiOeeb
TKPg70QVFjO5e14TycrjEDuU3X5rSx3LRqhmJHbpmLoSGMShMlyZeh3NEwk1kslf1h686dxZW8Mp
Qv9l9DY3PfAXfppauyizGh5pJhOP3VZGNk8weL3bH3HRQgxBhbgwmxULfIpnCpBMJh2y4iJedSVl
1elKCIfGXe8hGlzcp1GRTmvxBGaZ2RGTI2hCsmni25PBmG958HoqvoJ1qRAZe3pX5RuO7S16bDkB
8p/r70M6zmlS6NqErbWgB4Yz2WV9USZm65huVW9tQkFi3fbhqrxiMYYnmfHCZ9kVGB8JOPUmScQR
bLQwt34ZWb8hV7jHu2iipXzl31qYM+bEkzOyupjZSFbqcJ4J4oBGKZq+OwcC6TOFGtPF3wo5SdWO
IE/kgnASgHI5xDetIcR6b++D9At2js2LnlIhf8WyPvlakBs6Lxy2pWGrORp25B/varFlFJibc/mi
ug1TPoBy7l6FY7iDSsePJab84wpe+1bQRdC7DdeeaCvgFF9Xq2ZO3K0IRoBJBiYFsjDRyCh/GuSB
bpAzL4caDO6U0d6rhmCLOV7q0Lthv1vy1MKl/GFgzrgZ6DYpcPwCVlR8KdFxIb+RyYi8qMNZtDRL
v0whdCuO04qrUj+RiN9px12Vvhye+t91DxFgh3wF8abOZXWPzqoYTFNwJCCRoln8ePjGMvQ/4r+y
UJNnQp2lmPr8/ksHYjK0lSgQyFttbd6WcxxwR2NcuR4lTnm/Xq2Iuddquk0gXuZKWzNPo0fRZnnT
ypAEXZNDcjK+WcmNx2nJEB/U+fAmsttbNC/HqDFaQklqPKpDEflKyzlKJdf3sue3WzgQNPq6rpXp
ExfdHW8FY1kLTrPlAVa/s0cglv/Ryo0ljmqcLiBw6r6dZkUvcWU/7C7O0aagEtjRpWlySCmL2fdb
+y7X6HvK3hypzljxI+d6gMZrsU6Afk50nchFWyu+C/CaEcVCanzX70tF3qu0RV4O9SKbNIqxV74S
4aMYSDSOplivmXdmn3IHeR830x5vTSEh0MG6YxoxsaP/W1C3l5S1YTyDIZEW6lRQzboGfmIf5V7K
eeQAnqGvOQwmj+Ig5vDPTipAszTSq0LcrXyY8WZkOcPTTJeKMKK9TfQL+BX4L3sWEZA8Ws5kZ0KT
2OU1Fr6DtKJQXJU4rtG+8Bebf5ikxlrmj+TlwlxDEkzgyeuDCnbDl8qJOHar+jV0A/DUHvYU2O7J
Rb1sChOOde/4A8K5nYuPYxilrXXCg8MdCCUBonqCemoUgmLAwahy4qmyC7xQwSkH4iWIM691pziZ
Yp6Yx98lHBuqmB8iC5lr0G/RqAHlriDfzWzriPoldyvd+DuU9oIKGEa5wCPYeah+E3gVVHQw4eOf
zYI3CGdBrfkbpHP9RogkYH0ccrjxu4Oe+3VpW6wmcdPhppJv5EeJE6tUM4PsbBUTM+UALJ1F4ccE
jMfOpGqgu6a5mOewwW9Ou81zBuWpAkBnN9V8bMDMdC4xejI60t0I3y4QzH9UQdhDte0KxOybVo/y
FKXokB9WA7H5lBTpV6mOAAyXKqKPjqEdHsewgjLblJ+ufnUourAA0/T6QJXAC++VTYZtsNNiE0aD
nPoZ+xhfdskdwHVgppzQSliBUECNZOuMt4xdvxRcPcINtDITUas+97Jrj7zJnCFrKugTmrmouSus
hIDcnuHYfZZ1Hrw+qGCG6iuX6gtd6Pf5ADw7v9K16MB/t4NKrZQMR1V2JU+MPWbMgYCCJ/YLeSI1
2X2IP0dq3oJtnFaYelgfqIrQ83tZglsaQkQiEo04AQsnYvwqFXxSbW+ZJTx/1CnX1nFgfTNxSw82
wFcasmfco5itOGwWDZ7JNFR4yUeQUkjX1XtdLLGwjr2IkXPDhXQSpt72cZTwJMfkuunZxFrY7QyJ
zYZ3MHvsyRQoH2suAN4RIM7ZXG/Wix7Pw41pzzWkSP23EL+inBS5oroOlwaEQiKVPgT3CViB6GaF
uN/e4T/m+YRGsjBMq6e0c574+fNEjhB984nI78mgatFPbfb/8pLrYuZupgUNPovvYVN0hT9kdKWj
FyubH5gNDxgGdUIGwr0lemZNFBnlycpVzqoTOsJ0lwSBGFrNDR5rak66L0NUP/Aw9jwU5pvMzC3a
zdwNtf7suPTsNK0HESwfDZEXv/gLZZfIH3N9BSqZu2cNK+Dm6wY6rIdJepn8NIq/EswIZ6j6ViQD
RJPE0NGVmkZg2MEM/k7fEyfRPystHp3F2zrxdWnVXMQ054HzOzhpagin7dTRgLUKQMj/39RkLj94
ByCAMh+5nQlG+fuZKxshyviYwyquUum/VlsG1DLzKxz3Iq+H0rpDIuBwlqSvbI3XCRfNiBwlZVfu
BGzvV0lUjYoi5Vik2gPGkZ6ki7FbN1hAHxqQ8mRSf9Iz6w/1VCvUXMWp25inlz5C6SuSgo2FxBJa
FPxzMwFaLqkp9t0KEXaCTiOBl3NIdgHxlGaqM6uQiXtzZytv6Uk2BxOatEoefXWljHdk6zU0XbKB
p9PzpvbhnUg08J/kPwqyaic6O3qb5GM7poLmFy9n6odpGgp3vITbBbYJGtf3E9Res2qD4H7TOC30
Y5WT596Dp1xhl71MmTSwzT2eoBS3EqLktABLs5rPF9q6nOGmE4WUHw16DSj9ifd6XZJ+sH10HA1U
9M9rRZUW7Q+iGuQnhmng2I/8A3GrprjlUGv0hBtFcWEFnu+sQAllwyY7SsHkXNf/sC8ycH0wTY6Y
MmtbmaqGEdcwy3qBe0swu9Yxf207YwcliOXYv5jb/kbRCQHay+CGvbMJ/Zz9ScevS6yPj1jmJEft
e/ME+eHdWg72wo87pS3c5T1AP1ENu9hWqMeVsLVytGzHzMdtcJfvStbssS6OEHcXJDupvvHBt95Z
eV2QF4X9RlQpmUsTh1RCO7rVVvPzhKmW7K4TxD1z7IKQWLCW1LPAxvIKevdsINDmUK57yog4evRh
HRt55YFhNaErDp3TSHkV86zKGfj30UddVZvjLBFhV2+/AuhDYPaQDpc4BpxQ4Kxp8xkuktxVWlVH
kd3uUxO51QjTEYEIXSJJkOBt4MXTESJISpq000HsrLzOd6HXLz6lk1EbO8JqbtH0cKooRKickvlr
nGixLO7gL04lxG8h7HFzFy06VtPKcxWfSz4KWT6IfAmId+vakNOCklzJImA//lrC2yTb+CsnwNAo
d97cWhlrFSn/d3odcQecwvZOdEDud4QccbBp4KEN+g3/rT/jkEgMtYf+Oqo4Wd4l4q2HVPr0OMDJ
IYs753mhkyPPbiDaxwqOrRDl3mBZNTuwGQhjrOCXhC3Ehvx69rIn1EZfhJh40pto075n5Fc5GeGX
Udu17Ie34Od5w+bIJuK4Ok1v1w7erGPQ8nL1fJpZiZtdenEPNlDkp8TWBv6zCNMtDIaHzPgDt+Os
wTp1xCGGLmVV02ES2FK7gzQky3eZQIbP0v9nUplLHF5xxS7kuQ/GVAcbvdW0kS0rlAsMJShd4PLV
M+nkHNyh+XKPYd+XbHy7Sh7zqbv8xfJFhA7xHXWu2kH5I62FeVk4FfPrfEM5RsOgSG037hZNh+Lj
MHaf7v2zudIus6zaFlzIzMnnFQch+06isbMhzM+hk3mfj9RiyDmYTV6CYIsMPcoldaNH8lLYobI8
1s+R+Uo0KDDiwaDM5jw+g9SWzNuUNv38ujsuEgaIP3K+5rhL/7mqqsIB+RBpQwpQewoNiDLhNpc0
XOIii6bQUoFKCvccg7pnxNQ9gIysirR6CeCkRkX6+/eOxq/oqQlVWgtob/d7CjXUSWESJ8HoneDc
ZdyonGZqeMlCp+oOgsn/4w6pRk5v6mJdK8Q1wleYG9ysWKsq7i0TJ/qKjR4f7YmIlR2uXL74fgCZ
lDq+KY6G/qDO1/jhkGoVMvceDrPEqfC0nt91p3Es33jBE5+PEPzKa7dU2h7I1R8rezAtiRHvqxH3
9Xg1j6QmTTu5gcwuo/MBLf6jQo5YW2m8TGnx9/UVRHnP68GvQ7lWJp9AzIvG1xANcXRVcDLY4Npk
iyx+UufXRb/nfi2sIq41DWEGBn0eeLBAHf0B3DbaRSCYbgs9X90ejAQTfwkT3ucmfiO2QeFplT2X
aDFDsfTI1idXuOc2ayussh7ugcKNIymzny2gHnsQwhy/wFdQCEQf/pt3VBFcoizk2SUqnReHp9fJ
Y5IcLbEph+iqpxgOZ4vVXWEa6qmRCmVTaxRhIeaPmZp9lPPBkJfO3AynJzkRi9PLxopJ3fI4SL1a
IXNbad2NsjmKBBjeXW1/LG1fU+fdA4X/Px3Y6KOR+brGoDctk6QsO5xlQpsgPK3ZK1IPonYwBMEc
229XZdsbeQ9dK+bHyWElIdSLfItB7BUPhyvr1Z8n0fBmNSg2SS1xrlVBOGK6TidyC8O6O4v6qbFA
hPwMdN4tJelRquoZYZAArJa9w0DFJDzxo7EaYNytgpL99mAJ09j3OPi6Z8PKKrPGyfo94Zhja3so
hGu3dzxbVuRdvHCOwSJfd0nUXr6+3XzjZvnUv2wIlOat8GUeFLPwPbal7vr30A/QtLOwtsGRP9WZ
8uiRpy1F08diZ/xnjrlMgwzn0QsvXR5orjGuzPRHo10V/w7mIM6KgfKhfWZiJepx5kYffBi0ZPie
EUUZoQ0up95ifNiLRiR2tODhNHRcomeU1hVJD1cG7Ff1cZE5itMwrZVPuU7JHK2AvB0xJHykw8/r
WOulbPSjdgw5HVFzFp+RhmJHmtfdbS41ukIQ61Ryo0qytHAFGrPZu1pDpVNpHyXajX9K2f4BZH9M
PlDMLRVP2KX5u+TzKclhPSUIhmCsQ3ir7GJEDDHPMAEwKobJkKV3eA/aPvvEg/YO/Q9nYPrLmw/O
3n7p5XoQmRI9bJzjdgokji7Ejh+cjecqxxFC/Q9ZoxGMk+3ITEdbBwS6pXh4atkAngVOnjb+BGRN
g4n37jmBOjqKjLp+k6EQ7efzswoK6JjHnosZz/cNXGfL+83VPQt/UAIqN1ZYTTRL4YtqrAzCrtH3
bDcEKOulXxeO7iJ0uyNqoceLUI4jKIZ/7gJsbRfTTWkJaDPIoD8S1+ZjFLk/wqWW+s0FIFcU4fhu
CKc54IvSo2XVZLxiTjMAbp6pCIisFJfrI2bIM7MB40gZ3N75i701pbytonFAjKb94p/++QP4mf8Q
blE/JuTVVFdmGzVaLqkofONYxQyUbCkbDplPgyJKlHEkf3KI000ZA4Goc9ax1jJD5uyMepcnB3Aa
ygaH9SpxIHdyMCQM5ZAa64+5JGvUki8tLEBO/oW1+N7lhXlOtY3VR7JN4QOicoz1W+lmk34MIsnq
S08TE+0xMHSZy0AS5w74XjCcohQJRofXdYoGcYPpbOb2fM8GlIUoW7F9lCDU5Sp9cGHBlSRP98nY
wH6N7MXMaKSeKBjOWubcMiPoBebqfD6qw7bXmNl7ESdbRlTVLMry1CHd/5I7nhUBe/KyZR6pz+kn
KQF+4ExYx9qIu61Le//+eIOm3nDiCWp6RSgpv9fws5VELJj4aJdk/20UpMaB4EQmPMf5qRAoUHtq
/bRFrUxwt141t7JmGOZgvUp+POe2WM9HJyDtJ1AcHSVR8dTvHmoLqSgPePaZGw0ywGlTbpswx8yn
2zlc88yEzTUgCOTO85KsrfKpok+uJkwdOH5vI6NepHNtXGvJXcxBxMGRx8gpkbB8FYNYbQp5VzcK
lbmzptHiZgBjwMqaCHSEKjKHnIleFVCnhnCVcY3Yr+KbtDwdyC3IsifLNgZ5Hn0jC3Y8ctRd4KVe
RSNN3wtPuXIpVAJqQYNrkUcxcnB361cwJMiM35Z6IRT9yuiDcYSZyRksqE3xJBruaoueoe/F+oOU
sYBN1uDZhSH0DX6ox4A0t6TVR1tJxguQXT2eVuT7V947AmjmxP8x6PwwlenrEz877R+rQ8Jh7A6C
BwOxFRFERwxaDfSJkrt0aKXWfypFHcBTe907Yf97lfko2U6WjZ1jOATPUn+EDqUAdS2493oratJ/
rTB+Zatbhh3c873Diia0TKPRPU0QyS/hGw6nPUp2LEK8JLfDV2lj6VdPaeS1u3pgyOKWl7eBu+zW
GQXfS9IvwbCXYD5RSSocB7M+ikVOTYUxNzFuafoujb6AIWII0g3jD/Lcuzag2MNsrYjTKeyuQjQS
d/a6UJySsuIf0+nU37wSsec/EeNbSUscgbcEBOJvfM361BwhJ4/tN0BAB1QVxxFEL6L6O+yGScPG
0UM8hNDwZYe+c4Gbm2OGKcxrvOjr1rHMePTXxGtUPuiFHqSzbbkte77EoRWuHIeVcduSltq7CbU5
anmwoy5n6uHAO7hSEwV2EUd7A0+V+CZmz2KeOFeAbznwgaqixbbdXQL7YYudl9N99bBFAi93geVb
zLayUfsfPXgBMdgVVJ3bcNiDAaN0y5dC8uWnnMNQXCj0P2/RtT/SQDb4M+LC5rmA8HSzpcs7Nh+T
7zTISawNsiYJgTXq8lFBztxbMQVMBgoy8i2F5e22UKyS/D0rKasD+8TviEz9exDfMcNZpKnB9C47
ZWB8jQsrNaQ/yLaHaD0W5Q3NoH81D14LBw/grrUTh5kdapczheyrJMrO1DyFU+GuO2i+wa8ZXwHr
8n5JX9wwIwrpJHEJUBG3GkpIkRPT4FETbdjUFMUn/Ib8iuGMDdOEKnZeZToiE/9lkeYcvDsIVDvp
AxnPVdBz0TRDSA2aWoySLVy9r5Er1gy2na4MnxG9P/8ZxuST4c3NBzGAmWNgIZ3JCNR/Bidtq/kr
38Gke1oykDpRcuE2mDJLf1EHkvINiBVEKhOBxZWqrV1gfb3eM+OwFVYh0jw2m8jNPnLCCHeSnvep
68hzjVZxJzCF+vmudxa/zGqB29CIbORG9y9rpK6QIo/ndbDZgEum0baAXoChJJl3uVwQCVd54iNL
EkSU4BDBC8WGMX0sBwvEjKbGm1u7mJe2RbrP0m2OTvbohqia9+QYbjsa8JyqR/qPageHUlYWrgw8
Rbcl6YVl4bh8iaDewurMWgzPX16rcHShwTbBCnFv0B8Oe1GfR+e25yiuSSxG3jMjCsyC0pXvavOz
jTFGYU34u7/H3ywI+mplO+wMStPmT+wD0fxvEGGsPECfl9hmK0o/4rNkNSZmzkBKaHYKSYbEIOSh
Agki/mqOGExK8Ai8WLRu+N99qc4Uv5TjSioEnVfyfBHTngTcVV1dMLeUNpKysV1zwzaSWXzci3hN
kQO1arkrIDgafnDgKFz8DdRrY3R/j7ZadMXub9xStoBs2SgQRhqxmL2QvAtOeJ/uFE3K71HVAnGL
SmsK5Pho5iCQg2JnVWacPhpfSVaw+3f7fbQQkLVjI63Ceo1MK04nxUdkPZr43M7HghhKywiXAEXg
NiOGl7ohkkG9/Hax4U7wsvYXvFS2aEaDoNe/YJNXIHivyLM5y6apGItPncKfCrHRYCONgyRvcl5+
Mosiw8UFxq2YXzUGzvw7pI2aVTuPvBQePzb5iuulNsxEU8F9SM3Fw8No3Lolu+jO1FiJS0nJPtpw
fZHmOuSnKLLmCMPxCrBS05HDJOYO6msudu3tFEdnq9qhAjzOYoJgYbXqdI7TRj9Ps9/XKcnz486o
v2m0KYT6gahWpcFLGSiP/K/+hwhfDPVD6y+goHub8AeeQx9t0yz5chqwYenzh4O+HOBRMKsa05xL
lEb88ugAe/oH1JwupnhCM3X8ugkgv6iLaBsH/6wIx2wUNl10OBNnElU0TFpFREWwuR2xSxOs1Y3t
gS2oj4ZpTgfJvyO/1F3Fxq9lqKWqUGrqLCb9H3bFvkliY9HcF14+ZqTqM8Hi37N8KDYoGcgCjoyR
avighyDOCvMJRZPnZ+swXkwkH7VPIX60zQyCmjAic2vAEck4jb1udxzSoW8XysWjNuFXasJrn3dB
67k/nMT4XYSkSNSL2ySdU2TURVkK28J5hS7REY9T92ZXoy5lF43naocWhlZF2sIQ2mQGoEQSlhu8
qLYDTfsx2CdTmsWiAGRqKPVGkOzCB6iuXxO5KXZ+elyw5VGQztGu8pHkKZL6B0oD+s+0PSLNqCiz
MfjlD0H6OhByFsfI5r/t3BsKFEjOQhF+acXhWCOpGh3I0/YB6P3MlR9qbsmL/PM/ChZGKdlSTrXy
IgRgoztuzGbPKziGgFiSCfphNFRzm7wwoTAnsO/n4EZh62rv5KFjl8v9uPhOy05qtiHuf1/8Oewd
HLXmSKsAPfoJuS9aDuq2O6M7oJL8+sG7z2NmE771RAKxEAdFKy8YZRwXTeBBrtn0L/ByNMbUV3oa
ULVeZHlgMhiUGCm5NMraZBGQ31VeaDxyGnn6uMvyfN2aAEzzvTwe51I+ZBmokZSuHXZeyHzWsHv3
+oCSj6CR870Fl3uSNA1xzvO3KcS62GeRqEaQwN1jqBVSmH9+1vYEvt7lIm58pfT12aaX4ORATLm7
v4OVgKps+X31+cRypELQhEmo/TkQ7ZFRu8hwyWKLK/ZxJpNWHayZ0oM0PgveYPzlEJVY64738wRg
eMEKKHaud1Po5ss/NAjtAN48L6l3RB1tpfaqhdc0U9YOwDFHKVKS54bRenWSfMxxO6XhAOSqntUA
aIhMm3uWeEtIM+Y+oklQMHUWXSVPb2fDR5ksRuNiplNZVlkkQ0tG2HEtfdj/kqq8/DnykUY0BdqD
5YythPPfti7vuJPaE8aHJEF6TABPb8S4VbOygx9szjJ7bOhyEN9pVYlqM8F9aIC7nf1zqcDk5Fcc
kyo0uZ7WN2DO1Qf1sdvKDNOjqEb4s4ByVqKrK6EiMMxwihBQq9xRJUBwpCQDlbGB0Fvu6EbzkI0W
jKe4CjFYpX4MSUe/Fjx5K4dgqebthqDDCEUJRXrqQ/B/N5OUOrsnYrnOSgRAZGyNVivDGMMZ6sFV
5jPRlWNmNT+/MfIUPFzBw/VX91T1i9U4CpFyVAXtGi2LwZHM9nEiooCBcafOFAmCunlsm2m581I1
FHbsGQW3+C2eDxcFbP+fG7HNlzIZ+jXQF6OY1uzxG5j6N4P7tb18o4EaeAEw5+mfeHRErdx5sBsM
IMrz5quI+7ttb/1zzK0ZzW/wjtxKc5moRO3uhfPRZSDzKoO0kGm+0ayYQ9cdpphsx1n3n7w/yUpd
xYL8CxFTEK9K9R0wz3YiVTfM4YB1K9IYEunidhNRpz94KYHsIX/AYQ7HpoHVpXGEEB1KDWPpwExT
KXlBd3Y/ad5Ok0HAC0P5tefy47wHX8c5Div0XR5NyQmugh6Y+QKmacnG1L2SVllSxCKxI5PK2oJ9
uDcZwwIsWaLsmW5BHhhATcD0Xc6ocK9tnYXEcTa9HVvOlnERhUgdJaNELqXYlUVrgb+BJQfotb25
TDZgYpZ5X1XqzWlm+MbsSYDeN68lwtGOGXRRmyNS0LUlAGTZ0yqd8kHuhlNDvErnAe7jM8hFMd23
WGYou9Wek+H9QKwPj5wTdlUYjy6ayhHM6rneSb168w8to2cu0KH2FrwPybvQDrmFnkm7uLyzqw1k
1zOHmPAXzFbgVnChckYgwlXUT6t/TrVHzP9YnbIQwDj/2KxFD+loynq14gHMAXaqW8n7iIM2mCCY
vcHlRUMn4nPXByi7zGkqoSAsgb/TWhPdNCKPX/y2LB3H8JxFdFoP2RL/JyZOLx+SBVH2sY07UozN
TzuySVnbLayaKi33xjtR26htQ8S/3/2cZaJRKDA46P+KKbrgJO/oc8nbngtMLMXA5Xu0bleQtwf6
yVk/SnKQ7V/Kd11/DcrypbopmdJ1HKq+7gIaa3RDzDiRt/eGUBMR2mzz2A5bFHMREJmU2GRAh/zv
7P2sjVmUKoit7pnR0FwPqw6jYs9DfE5yBOlhIyo2vaK/YqwijXU/7+Wb10IvCFmmh74Ho562SSQG
TAp15HpmaRTIC8/EqVPcpeh9L9XzG/IRtN3izgkFcsEWWWlBftxW0EZdtggq19G7pf6UOeHvK+ED
RanBUfyAWYjmITu+N8JhGtndZdZjJ0e8MsTzR9z6W7WZMvOD2gbtV/yq6cdjx6Pe0sPPxOUVJlTu
FESBnxs9kLGA3dcV62JDoVg7cfQK/K3sEooGItxjH1veoYN7NPFxx5skwpnTCfSovdH7XTAGiTPj
tkRgdSt8ASSK0ahcIpHS9rLxbEwgkQap0M55J2JJdsL++rP92bzjipDvtR/Zzk5wziq34S8FDNr/
73VAJK3/2zKrvKMTOjWQjrhOp2RyuKvwDRQjaDnIOkIdZQXFEDJ0Ls0U+japHDQHGoMkEks9OJxr
Is6OSO2UKpikzSCvhNi5q2yOqz/2NpBpvZhYLRtqvcRf20Q+T3g+GB0QcLENKT1uiT5jDVN+2TSa
ZfDGdE3Gofb7j1goAOQmrvtdix8tTHkhQVll/mNZ+ERrwPsyTv2kBuFB4y9i2NixveuHHYzMbftC
A07wY2Eg+lmiFa7ZTsFWlyNfBQ8BoNcB34QfrhW8WEe6L37cQXft89kiIhQuuFU50kEO/l9IcdjB
UolXQdaY5uNyrfGaopzQMpmo5q8E2e9ePILduzj2Wn/eFKp34piCo4uktxUl8SYuorCpw/r3zxGP
Gf4Bopjcy63BziWNjLqIH8OiFobqrWy2vAOegqy52O7pOn0u/AVeW9WvaZMs94V7C3u2RuL4ugts
21UI+7nkuHu2/rjb3qTYK2gru3MfMbxq8fsPeRzwMceZHhqEm1Rmdnji00A6kfSCPFZyhG4KiRz7
KaAl8pq/PkYZtvNMLPOjGpQJFi2GXhBBoBAe99LaHCIkTRJutx0EzWkpH7dU2a6Ts5ydWP3PDU5E
mEgaWsT/xPpvOt31cVQ6633nJ7H3apIppjoNA1VEv2hbGp6RSTKbH16kZ39MX1mSar+kOPvxX83d
DXgHxYYBaDEwdZGfYo3wuHh7WtfPVEvTFx8m5WVwqj0r/4390aWfQ80w+8ypRZpv8DAS+zHWPov0
EecfZAbFyeP0B66QzeNK8KZSfd+3L/VyDrmA73gArBzS1DyYpABN9JhA4HQcPDTVDFok45sDkN/E
uq2vwX0zhCKEQOF4uM9sUPy0hJ/X4zCjL/vCyIV7bzhO+j6erzj23ASySo4bUp2ai452LkT7iNUt
BziiE9T2pJetU0J3GIw3al1gArVLNs4lBmb9E7xYVQyoqqd7iUGD3nCveHVOtvEeNr/b6KGy4aVG
4iL3pKJ0zyOYl3pSNvO/OCkGpZuKzdaOiytCoUysKQqMjNg0AMCBEpE5DV7Tbo8adkKdL3KizuBE
ZD41eYr3BPscyHXso53b/IDMk0g+Pun5t+8+NObUS5dcL+5jvl0WuhldevhzHF72qwSku8LFaCOm
ymST934k2XhZCxsq+m6H1pGG6JZTUwEKYu7fFyUcT74bfkaqT6EEyFq/BA1I1Tu/b7kYe+hoXV3Q
MJEYu18bGbsXbeoY3o29I5NI7l5DQ4DezJHE6NyR06iBZpZQuyqV8To/HCzeqNIKQJOLRRpI+A9h
6hjkZ1f8S8+dMgwIWG1MzEIG7M1SIj0u7P+TG9ddOMBWjRMgZhUK75WM6kcRMZWVuwAnG5QW9+A4
3Ptzb74b/xi2VAYmQiGFrHeSSg2WuNs4HFpWkXLzE+NMLnKS/6IpHReucftR0CWobC+lV4N7Ap7O
bldKp5mrXEAIbjpmgG/QFdRD9/oq+V0FRhQm0/S30+c2biSKa+UYLAxXPkORUzRafNUvuhq4of+o
232SaQ4OKbnOCxLEpMr1AZ5XRpE3ytbB5Tmgifut4GjGd6uQZo7zEd7HX1JPq/eUXGNZ9UvD0ZI6
Y7kIzQVaIHWesOE66VEzTEh4ox5Rusmikgon42POARPXHF1spXvmmUIFP73+AHayV0+SKK2LsNPr
eZj4ZTfDpqiRTR2RqXi2lZ80flFDaqO6ZeltuWE88Q/lzjfolYUzNIkyTJdMTbFfqXUGOXQMtHRo
wiRrDaUDLdqeg5tvmBD+m9lZyc+rye+HewEKxauMCwL8BrhU+G/VSOkHVCARmXk4Vs4rcKLlPl+j
KpRxeV6YJ29qeavAGleI0Ed9i3ZFTtc4/TLckft48FI5mV8R3SMVDOKy4N32X7ybLmEEPHOJNmmw
yixyfC+jg7vK9k3TEo4sC262P3Sl3j1FW3hH9jlMrTynfqnYWritAaafPUyLhHPaUmRtbBCMuLLI
yGo4TmBmY/h+C8lnbWUlyNeFv8/eQpFR4AfzvAcsPxH7wxBA+KYqa7qYcfgXIktW8xumT0bFEsrL
UL64WrTtQGOmIF31b3fEGSg/TUG+AaUMHAJvcjZ3d89XpEXmq16xvdYwXg6eQsnWwOLesNOpRv/m
sVjZLi2wR1G7Loix28FxP65S6pvg+3wvwxrjp4jndSIoI6cTyvk1mr3mrca9WDIEqYGBI+5EcWzI
2HVL2mHlscdQo+Uf7eeKTWzDT5wKFu48eWRE5HgFDqJB1v1kPLlkCi4id4z2s6RdSsc0bi5sTOy2
qYSAp7eGhz7ymxpk+8oUQDxWkBWOVJuIznClqIlRBMWvPbXQsykLkSUNdgduutplihdosg9/eN92
43/MfUynDPyjcepdK3Tye+5RTTDlVsVE6z9yNMlhusuNV6g6YXmyRWWCOHR8c9ffDfqp35m0YHAl
OC9TK1HM6NiAyDHHDMhn4YpmdlJQ8+tqYSub+KM/hutMacC1fH81Cb0KZBhuhqSZU2TTx2wAfskw
+MNeZezeJ0zyINaE8JfFkbblVt9WjjCCcSm0RN40hPMpajaod5f3Oq5Tsj+muBavsHxRAnFQTDOB
PN/SrpzP96O+NxFlgZHnSQM5W8o/m7NvYpBmo5B1AkSpTghw+PzHgyInI2O3ubwj3/oWBMUm7iD3
PC6cDSmRJWrPxh0ADQMD3SY1y/piHUTZxEM+myPULugQ6flo+ofipMmNgItvDX7J0UyiR9TMXoUM
mmgOBaoXkTp+Q/gI7B0Kf9CZinnMA95e6k1Uq/icY+FrQzSzfyzxQMDEKWhH7NU5O8qlPpVGXi89
6HzajFIpStoLSQ7XnXECmNV1o0PXSy7uZfup+bkUVFiVKVwdeOaNu2Zbkb6enu3DuQCsFI7x93+F
/0w6bDD4JSvG7B8A4tlYm9nNNu0ijlLWDiEVP2l0GA4lltyHkkxOiZHGz6pDxJ7w5B/25YdpZ/ml
a88+G0o4Fy73Zg2zDqg6g2Ds0N7UP8ZzLnLvuOo6NxN4WAn6ds+YhNey+yq2PPqCyaBTuaW3k2MI
uU2OI3RF9BqQN3Nvy0CLlq7e8damoZbMeR4EP2eAqE7oUEfceNnB0abpDYVpAymHDxZvfgHi9xPP
RIqbXn1jYtpbOthPTQ6xrHX+QqIHKaCeXUdMaBi5wd744G04xFqho1cnpUUr77d7aBx8t3g3dQU8
m8/3A7M6ykC/pthq+BC0medHAix/eve7reh+7kjG6+QralmUZMuKl3rmRuZst1wV08CF9GOPTV1M
YgK/XPBj5f+bCe3ZswsmCILYHwr5+EZB+ZoSqf+7VUBUSkh2hiGRm31/eaplPNsIaH6SDtT9WaZy
/Q/KkX4MrD3qb9D9iNkdOk59HKDdAsgE12U42b5elRPQXq+a6pJARCn0RWYZWCZRHRDoeEbsaF0p
VskaindQR8XkHZjOBtV7tX7lCT7nmLhmoW+wZuZerIwa1nzyz+TRa+Cs/2wwCL9MQlx4st96F5sn
6czBzb6rbO+hDDIiWA69aPKHoG0pFtvfdvKzyvWTRz44zdqgVeknD0tLuvSWuMuiOksfNCAgNXD/
kReOrlL7cTIbH8lowRNsX6sYbwEhjhbnFplF4qkm2lLTGpg2oEgHwko6fdaJh1b0rGU9SckIl3Rr
xPSoyR5cmic6/a2hvdWGDKFlHQC31N/n2pV3pqWjB9R7f/30Y2QXZV3ECW5O3r1zGZbA93v5+5jq
GfcFsccDYkIsohYn/Bz+IwUPSxP2ZgEnsysWaRi5nWjh45CS30GxuhHFQW12QSBQOGjIJ+Cw2TL8
rOIDBpvMVgCbjA6pBcRFS7VFeqccW6ETfoIr6JMhyRxllx58x/ChLpRzGiVCfMAxNIrG0FUg2V3+
G9BhpP+FCCcUtRkwValsuoRifFfZCclGMwgpjKWe931JXUDmwtfiAJTfUrZfSPzjCHnVHZ1zCRN5
jlk4MkDtRnUMxuShzVx5/RCur9/kBzBG+YAKC/GEAdSmXp9LvNEcUnmcwRDwFKaOGRu6cfsfbQ/D
NWsW6BHBeBUby2FPKtVGqBKiXl38gxtaNRUtcx8pFQpJ5xS7q11YRWCwibTZN+LmDYTWaDJxE1RL
TN1iBSDE1jo23pEocTmC0bPPx7Hp0oJS8uExSeatk5W9Xj08fRxzkzNVxTotaotVNi/3fpe3JDF3
7SkP8sinKiof0w92vYV6s1MTaXckKq3auzZdOIrK3AHpZnbAGrMCaxmrJIwz346kgBgyTcJZvVUD
W3nnnAMaP69ynwE3/+bW9U2BdR/f8pEXgSyQWEJbXVGoA3BtUKfcmuvrytrjkwHt2sDAVmSin8zx
iirpQBDZxoIuAKnWsf6bxcDMiLrx3jk/Pqmy7WyFLULrc3EowfbCOkzclOipqdee8zqAM1f+lVn3
j7cs/QNXNx3nizLYynywbbMG3f6WeJncLVkeVUWSLwYXp0+KZxFavmF6iTgOy9A74tTUhAmUpNn9
THp9ATstlxlfeVQCGOGGwpiKEwu1rQNHDcyoRroLfGh3EiBKjZPCrKhZtebxBDuRA5tzEYqr2cDW
PjH86EBvC5EiuIfOeuITPfm0X5c3YJaZ7FUdaX/sR6psYAbA6qTMtKbj/iXHJxDgoRFU6bTE5Fbn
D4a3oEqiFP59iTfo2aYk3xgE4lJ9h9IXwXTimkiN4L2seO67/6Q7Q4p1MQk9zSxF3evz17740xyX
z5WRkIgvK9k5/MICWmY+2D/rlvR+8z3z7vCKHzBr9xm0fy2ZHJ7kG6508j8B17Wj6+gwqEIT1nE3
N8ApXdBgiqAKsWucabU/Kre25WSgAZgzCSv9pSvBDWRcqY87RbU7ApX7yLOucgJiZCnVL9JLpwS0
v0AvagZ8d/lp9Phd2KbjIpqD9mLiBNcrFYoi2lbF1qrsmnji0tAtOozDwFOyxyvfJzisM8lqUr5g
s4GjPsvUZtrVjeYgglZ3Kz8khbMyOMgOV7UEP1oSoHG90XvYMdptrvfuCiSHzB4PDzuSOkKC/jgj
8k3nAuGjM4qGx2gAe90m9kGTLMwMRD9lnydZY6c3mluYYvPWANq3k6nm3Ai3EYygyycoPhjw5PBf
29/SvLU0fzl8k4105qlcD02YKBlwRaIUBp+C6HDxQVQJqOYwB/763kOWYxhfej79l3taKdFAb2kR
drFKPGtxS8JcixUI3O/LJG5ro7o4z+z9WLYwW72QPhSrf7WMz483Dtvxw6rUBLCyW6YwcVKlFXuR
XlwKl4Gqup83+ibxKBxytl5iSWgZKYLIxu9g9gtPuytv5gblReSe4e9Yab6Kun7A3VPB3eyie/MU
TLoXgVuDcuR+uTiOLFryFtUKeLS+i4thcplOpgLpCP0ETRg44m5XUdCXhPxu31ID59eqr0XL0dMY
m+8Hr0WWsN9tYdY+C5TO1iLELX9o8NSyMw9STUQxGwGRKgKMIKvaWHU8H6hdquiuRxXTGiRf5hjQ
IMVZxt+czX71fSpmkwrp6sa6aRPa2enGGzV9hNO+lcj1/4y9AS4ThhHaKxTSBxvTgx5lTgaryDfA
FycbL8zEWfyhGJZ/k68cnpWk9kVKx5s3mScIE53iNgFQQQBLu1YqCfIdLJO2RrSff+74OoS8Jd53
FAiIgZPQNN8kGuE2Yzlzi/56J2py8YlufP7MpPr3iOQEeywGs6vD3o4rLjsFK3BfkJnHBTPWlDMC
wYlfLajeNtaw3fwnTTJx5bf1SAhOO/omHlDtuR5+eeY69jaSNwM2LbsHELky7WbWmsMngJ37ST7K
kFcJmXsilA1VabMu5QAbEiDl8NV7hb8ktHzsu0gJoiSTDdsAgLqHY93aOQ1QahG3DygX+1IZOnKZ
fc//bVRQbNaL/N3nOtrVWRjGyglmfijsAFhfnt/neIwApTjHVg33pDfCnzlagPHkboaZNHeHhmB6
My4bRamsVuTxHTRBpMT2i19oDiu4tnzgcm/vprDH4fNJEqoYOEy5cnfJv3CLOqLc7t1965qrTa5g
FX++U4UhTgsDHYEdPh4mUdGkeq2EqySQCoCSjYYwYbx2t0z/udV5inUfdUvFM7PndXS4hWGAE/gQ
yEMiZEjh9AS23PmIGBfSZ/EKUMnsk+tubWG4x54tKx+LgyAtpKWP0APddjexEy4T+qi/uMk9t3Yo
gzcd5ovvgdZ/ftR+coTorsbpkCjZIKQxE6Y+qReCEDYZrnxhhFlCHnXdH9vvLHaflHHEbZm/Y/5S
zEoF/5MbpUXDKA3PPl/6ydH4sDoTKvaMdb3MQqSGshJi+MiSV/2nhg2Ftl3TjeZfhjOeGzHEL9JA
hek2Wmqp/OqTMnf9bQcLnl6RBXt6IxjZvuMjNCG+Xk1hGrrR9y+xD2gXS2mzFZWruo50+/YmLrDI
8xI9ROR/ucTfedSvPxiTY8SertPTi6sDXnsiMsLsDKdOB5dZZiPa3fvUlNDOfACtgnuru5FCEurk
lOR1Ir6TXYXG98bHaHr3eaLBGjt1ktBXLNxAWRurJy2eCROFIV0Bb8YaiIXBGM0ZDDr0zFC1FGfQ
n8FRi/Vy8jWpXNcMVv+CXWF0LYtN5Er/DqrRBE9oDJ8r2kXiA1w7Ke7g79SjRKfcVJBVrYZEYShx
96Q//oks8Z0/H8z+RU2yT/eR2/tqUJ7LaxnYp3hkvnereqbGf2WbpaTtuQ8qgeMnuyHZ8r0W3hjh
rNXmEKgfkqqqoyjCHgnhmcocAhSTmcbo2MJ6ncGSGw9s4XvgO3Lf5gxtRR73tAVWfwehRWYc5NNP
R3VBdLEaFpja1u7+gwb5K0N2LpZBS2kTaqOeCuCVQnucdh5p0W5DNFgyzcwAlCK4PPZOZ+RPikaY
oE6xwwW2MoCTq8QFcDpl5eb0wCXsoQPP7KDEvu6GWQlmhmjzs9+Ft6zlLYtfOj0bQ5B3N3CUwkDu
Q04DGkGJ5ltfAfjYnrS0aQXfipdPJSz+S5DtmSt8h+rFaEYUfDpiQE9ADZN5miJl8nG78viVkm0E
Kc1wRrxwAdCvO7ZIfY9gr1z+smConJbrFPa1W+KLo/O8Bf/lEyi9OEyfJnv54BORhG7okeiprlIE
2cH4z1m4Czbwue0zCIVwBb8I42CkHBNqHtAPP9fmF0KDjB1biwsr1uDdzSNnWiS/EaqxJNh3MsyB
tbh9vfUl2+gb2fGcPZjSD+DhzAXhGceNQNN68udsil4G6FPb8uOIFR5NeSi5D+jYW3xr0TvwFT1Y
TYFe9+FEVw0Lwqt5UlikdJeQ6f8ElC7zagRov4IH1jFjCALT2jA9hkjj6qGDlz2p+ZhSvFiTMMtF
L16N0lnc/mI3huR3QM0mY7XKEmpuOJVe5TC9l3MCix9Q/0H0RnZKK2ASmgGyZ5En4kAeAmsPRHfW
a1hOWPgSF6BnwVclcQUvYO4Q+YLuRCXmvcXgnq8wuwSQUM/gxSfPh2DR8bGRXqqJZrefLfdrmhLN
SqBkw5/zJfORWdSKyYN43wMgqgpUQuB80U6jmYy/BrI+AOeX+z9p2s+fST+yhBH9tTwQjTyZm8Xa
4PFFswWSv9FUwYWPlujJDQV4DZ0v4/Ep58tdLu+wil8sm5solSIgY6ZBGWuGeoE=
`protect end_protected
