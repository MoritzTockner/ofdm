-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
IH8P+4x9SMM9GJFI1/dfNE83HzEAIO/7WbCcDOZ77JRyeXRfojH7UjPWHD/U1qk/EYbDy6iw4g79
xASBHEKPDzDOmvKnVUHo4aJio9MQk7AS3Acj5utbkBVmhUgz4GjBZj6NLhqDuRiDqRRItRUXy2pA
cCqF5sedSbRyFwrrI8sDd6T/d3feZkKJMYDw89Eq8sz5Fb/oTAoK4FQSgFDKY7QUKHYL3Ssy2h2p
y9krL8nqnlqZE5mJe2iiSRZbvOnrWTS1x7vnQXXGoFXpC76qvP64T1drWXNZU+vMDkDmRjMER79b
L8x9xWcTx5MSk2dHieIkMrIHW9nzKW7YEH8xiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9472)
`protect data_block
D8RLDFDvWkOL6yFkhCRRl9Y9FYBnA6nKAqym1n1KUMNxJkklcVN+fcbHViW4OnRQSGb8x313fY+q
tx5tQwfsY17BeLbH5w6xbTqdtJp3C7kZcjJ+i5m9g+Zt9FFlY4ZEAChEjgfTsKsWR/fijcdHdtW3
qdX674CyMzYisqCZsvu+MAU4VGEWrEF1BVaSY1Me3F5fOMSDkNLkmOLZDrddCc+lTXvqGlwmahDh
Mjv1hwlnuKqLFSvKCHfaR2+O6V+te8106mkL/LVd+Xkie/Wm325Gc5tGQ355ITmScsFCZ92fYprg
Yde+NWE5ML80Ed3NpFBKf0+GVd9xmj2A8Y6doQ6pjv6LzX27GD5lpPLc6yif8eSlcKsARrQAVTGQ
xmmApL6Z1WoGf3ywEzkd1kRiMwLI9oRO72pWtEGDxaCRJ4YxhhCjpd+fiUedXDeFHUxU0X8ZW3L6
NWnCoJ6MiAw7UgW2+21KttT1ivFYvQWHqhBpc79eJtca/VX/RU0bw0LixJIEdTuETxDvIXpWR4vY
PT37ObSgESWAXZqe2gaaBDZI+8O+0AMr0LqyRURonOpMVpWvgyms49mClnAQgKVJtm6HOvQOkI6V
DRM+1hWSE+UVSZTpmsNotiv+HfKB/W5iaf7yucqij77UmKMP8UK5prNxrySXvP0PZH33JE0CGkQ/
PLhugkaWergOAugeTZzAz829M/9UOxpmhaAj0sF/S3ixF7Ih26KJb8JzXYX/V7jY4UXNGaQQxSAD
kg0BcYJ3BjC2khHRM9+MGcpfwrwD8RLHelbGSeus5AotxfRqR7nVKEIirKH8TaTQNDdhpP2mBRJq
SGaWOgJ690iwG4oxTKABhvR8+ftUydMhfyzuKrneQZUe1o69Qv3BFIST1dc1HE6QlDSgxojV85Cn
yNFCS+kQlJp4/4fe5l7vUmYKun6p4wSXOO9nvQdxx5t/2YqRV5seWlcKlqEhm4cUnDsEyor/g2hB
vuMzK7Wj6XpMTNmFDc/khvoHFTzLsIfKgblDdp5mkRy/y/OgXZZh1hfSHNC+IWlo9B55QPie5See
7nnjLHjtkcu1Ena3lF5dqn38wc5pKD58PTitASpd0QE6nv9hoUDYiYy0CZ/OSzOEKxPhakFgjSuJ
8sqgEK/DVKspj0RdgJWB+NSWpINlVbPecj80XN+Ah2dQcNzHBjG1RNzpyIVK+nTQesjo7nGz0NME
U/TUA0VnxeEYmC366p4GfEVzfjxOVCJCN1kvQGHH2kHuGnhr1ldiZwPDGNnnmg5/K49iNcped7Yr
PGUGRjuObACn0AeFh/3gXEscd9wyKzXO5A0NFcExUWRXLvj65JLTGNkXG2jLHFzbpQOUdHQBodTF
jc3LCROPj9Wvip11PEaih99DkQdYTaWamfelgqXVn2OY8SCd3bqyg+GPGeofcxkLSWQweJaz9LjW
plHITNYQWsFlLrXVgINATM7EGdZtjjh4zRS2+TborrF5khotyVLnqr01eOfMj1UhVXIFd+8mJI0c
JDo75Yei0On+Fq9hcnCLznAQxS8fz2idaLaNCi8SPMi6puKIw8jkz0RfetsIe3FMfh9WVoCxmDT3
IaAMwGyi+mf7Zf8aluHQtbgwW9+qH1hJWA084MzI5CZrbGe3gzGHKYBxGN2vri2XlfA5GwkSQCjn
T0PhdTthOouISbpiLggx7qUOFeCFDjSqrUCiRNW6Fz9AJWOSHV4tB699yi3r0UgJoEk96+97RNPT
uAUt8NAPm4BDjcmMqog3r2zZOEpIG8gGNE/UG+XFIKVlhFMSQN+AEI9j4x0G9KqgrMMCrsxCatf3
ftEGrDZM5PA4OzSo5H0ONbwntOmFy09wYOlxCmHl1EP65wTFrauoR3JHi/6snO9uDE7IdvpSJMsU
N/IN2nDXlfdL1xhzov0z91Qx9h5GGV2D1bOo2lO2HUBQHrVCmdMPZaCqvY02NJKo2FufCRJe+FbI
8GmOkvsxRNfHSDOS8mKzg8woBXXH0B2YD+fH+Bq+eX1qWfqHlmf6KSIIUb2FvnJptA84CPQUnkw5
eXUoBWb3YF1M9K6ayG72qgv9ozwJ1RyukN4TGo4l17nNdlBnCBUp0aeasZACZ/gzCjzEbn7kQR6y
dASWktqypscLCAmbX7iNSB7uImzWYZyKcg/v4Lw3/Tjc5wraziwbrkg4oahfCLY/kY8Q6OtA/efL
FfiMxnTMEiCit0zJ1GNYw1G7d4VO+ggjFwJ7suCexbrR7NTNq8nNi6dkOcWLepwKu5nzD/dQ9iLz
8nu8BwmjlOjybnPUO0qPmg3+8KoPQb4CpYIc687pcy1DCTZ5Nz/kHNMkpMXxGe2wVGhYJYyiun67
4qFok1FKrjiRgPFifGXClp0l8AIrLbguRh0O5p9yczMiz6tvKwwJa34QdRsJC8O2O8l48s044sv8
REfLQEAcAKNxICI4eoO6FDqC4lB39RkA26TVjF5+g1r7bu/hRYoEpObegTp8G+t732bwSmlxUA1o
tmuKnrSOyNmi3IT4Vq0iN7wOFUpvdVTOLQtEHs5AjccybT61ygUjHUZ2zTIgdCCElkbrD9mMt/mX
01fnAhXay8A3PCDxNcC2kCRGN19X5ap9heqYlAGa7cHc2Ni0OQpdyK7fR5zUQ40fMomAugPuAP7X
rCtzenipgAF+KZua7UcKZpNqS1P7vfvdmOa+jWsK4wHOsbsW7flXagegbzuGefyKBqu6YGBpw0nR
hR5eK6oyJeSRpDHDdyPRLdGM4j4gvxkmUhafSqZcy7Vpd5+V3RVerz8o5let5edwXu+uxM2brb3t
+dxHSpxKjQURazF1FaDP7J0CXrrFPtQspmaWlUasDS8hAx5qOaoqEb20uvtRR9BgxGFybjI5x6nD
RjwAeEqvaXNh5PakyWdFMjx+sMV6OmOfYOSBjNYARD93gkUpBtyItMIuHfH8bfDiUyfk6+f5qXME
oY00LZmLHH0AO3wRopDfiMpYbzmfq6KjKKuWuwLAapEM0BdVsGCvG+EdssACnw8jUPh1qZootlly
8Kdc/vOWRBI+JYOXFlppe/wRYNWY5b7MxV6/Z55q/sPHMzNx35NLjbY+qv5jTSbQGIj0BuLFI2Up
UjnRahygs5fM/qrHhW4RYY/t424ykH5xB2MIHhQtZ/7xXlJ70DG61F024VaED5I2EgRyWRxGLCFq
jNwi3UEV+/52HqT1NJSvkzq1dCzDFd5fqCbKkNYCsp4QCFXBRT8SvTt/aXhm8fXytTPhdKBioVpc
FPwDgXaDOWmIKcQd/7KjlkAtXhoIYm2ldGSZ7x5nJ18uyMX19uK1atSpY3tbrE+/ghViGktw/JjM
lBM3oVCdX+0ZhJgqEyr2DKDhNwptCEtIixfPQf+MCjbrDcWzluhfkS0GM2vqpsu9oT8H9VYJ0atF
sPNwLnuU0L8oSD59SJ/dU0nccaj/ricHZavxOOCH+78j0Ra74njCFq1+DGctEzHH2oeculrE0wM4
dEcbeEtQk/N2MiRkp+I+5Qhw5vcKkv1LQUHjHODaeqX/BMHsxmXb8aw3wntus/ATvZxjX/WBDH3A
ItE4JVG0850CJi3d3ATXxJONXKYqKJZmPXcYAjtLGz1LBmXY8cY9IxjdIB7WXzJCletddGvnnjLM
YvSYhm9nS356oqrtH57pITfaRYbeBuARoZrzHZxuOpJ6fu0ifHIR1r6RWbpYGeBaML0FWHUaUpT/
tGxP0WYEAjxEOR+NgjKmx2LLmRtaJOaNqykE+2E1+WIGzEzf8V2N3R5DlOEX3vTJMym55x06FKuC
rNSaUH9f7XNi7xBEwDguNSMS3BG06y7D6aqUMDJ4mtEElyiKfVYs3FI7yM1qftDHQmyjURFoccvh
ZGYG6qYxNyAoXiTTbU2zpdlvOq9Kq9uOZwcqOJebBYC1Ye5k86l/FnZ92dqVshHz6Z9uDOzjq3wk
V5LFiGOfXHvurACY67S2wJ0TuyktjirZTe4fH6qa9/5UYBpfwQdajuYSZ/0TApGdMZ8YxqEH3uBB
Up80pM+wjVDXq92zD/FT2VQGRrKGFqIqa+vhZrXqEJo7YA2+u653XG+zSzVCpriQwQtX8dlK71xF
akwlP75NIBQW09sY4KvIuweX6KcJBAx4txh0SohwfEAU9CGGdb9sjA0gt3zI0Xgy5WrcBcHygeHn
rXDFEcLROZwi8E2mSnEZXeYW13W1Rm3rCtCzHiKkG4pN3p7lSw7FDkuuU0/jPKZN2mHLtNv7WKxV
x8Zqlr9iVUU0NaG7mGyMenkkskbsIc4xsKJRkXnBaTev3O/m9czwSGJWKGuR1vIQ/fKgFwoYGh+E
/Onjl9aSwgi9eyTW6mVhlQ2m/c/QfbuZKE5ery0JM54v+5/bV3AbV8mve/sZCQIOAxKRmmAolrs+
bMhYT3bfrq/yDJ64Nu72NbwymXTi6cYcSgFKJ+B31K2PuvetrWGWck2HO8CGHvF/Cge4+PhxVBcF
8Kc00oKFgkk8EDRKSi55ncE4xSVdD6KUgdQ1cRjxhTG85Q2omZ088s/nXGBFKS45SMqK8NOE7C7c
2JUvHPUenuXiYuNKf+Ex7bfE7I1UtTiHysAbYcNhfcX5BUOveali9UxUTIW44FqHwsHHOtPrHKlq
W7uMnDO/cOie4Y4NtDt4fZPZxuWWXfGCme3AQf9LRwMm5JLgUEhdvGEp1BkDPRxupRTNmplC2AfB
7PENlsUR/56XduKppfGDuW6YgMuY7mASyTIX4io2kWAYiDah+W7lGZO2u2EPldry6gAJH1wf6d3M
wOS6N+SrZlmYnPo+ReB9l/FowH9+oefzmBeokOqmphTYcRL0PKTuf0keZF988LDdV5ENlc4gilO0
NkZj8SjcL0g9M6W/CDY9XLkPRLRYD/p3dCPEf0cH8nKDoEDJzUA3/l1a6jAS2Qcq4DmZWU06dgfa
KciVQ+Lw3/w8jx1TgFdDhvhNOyFQ8vsWO6vC2UA8Esw18JL3G+RolAB+VQMydym1Cr4Bx+tdAyds
MN8+CU8Ni++OYePmEm6+wAsTsIfzgVMsK0GFBzuOW6vP5ZUPFp1k9uzQP6bqhmZBl8fs3Uxku1ET
fGuF4IHV2/ninfyy6b7SeR5fK5xGR68cwOfzhssEtUbS8Pgqr/gSIqpbNoFPxNs62dEAP+kQJFj/
YaZuxyku0Vf2xVr2MYKYgUO6BlP2sA6avmK9bIdRyEY2aLRZwy5LBr4OTv3LV8nP2nD/6ClklHuT
/7BgAQbKmgVmJNrcUFMGcG4IlNn9MX+PIW3cpynjG3SwOA6NlksaYhdSX4xDmTmyudjbast75cSj
O85nW14mNwU/Roe+o77xfpOC8fB66TuHYJeSQQjTX0kFe3ECaIDW+mxuO8FFouLTnw9DdnVZgdq/
EBN3CQ31ythjJ/vO9c2UM4J7wu1A5O8s8VL2hgmd1KKQRetxBOcqkfYH0UL8DUUoeexPSxyoP0PL
DANkb8fNKF413+smNV24QMToaSskeVKiD/deK7MtorAInV760X1boxqrrZK9lsHJ7kuVdZ1uw61Q
W4HC13LNnSCtBPDfWWO+BiI6mpjiRoxao4QfVqA3nbXbNElo6mQHTEKTpYB2jIXvHgYUQ3q3XJPL
Trrpi3dWsKHPczbV2DRB/r6IuRjqi6YgpyLfthUH8PjmVy+Py4ErbauxmrqIg+GTPciY6JDUe0Do
n6Zik7LYzKUbojZWRzT8RLyvcFEeVCc6qhN/G9Mi9kf0bsMTWiMF/7a6uchn5YzezB3Mu52xCqWF
WX6Es9JO98qdbU/LZT6kLoW3PL5s0q0ncEliJ/mKmporRXvpLsGNk4f3pHE/I3ntXmAOU1b1NtX9
1ygLJoNGNx82pUv7Lj/ayFImLYlgyvlnqelEygU7Kybr/vcqC9PpfqEsq/CpY/5f0ZJ7fAf2dwfN
0hhWMU9j8z7S3/tdP3nszqh+VTRskc+9vNdUhfmDqOWoyqLx/hDiPgiIKQVnZ0MZ5m4ZcZeIW2p6
5GkLzwynJ0n4K0yj3OKeNAKIWzw5VHiiWJtskSG/0x5TQqcnq/lgpDHl1Si7X+hf4zaHiXNPDzo+
Tm3mlAXUio69MnWVdWb5KUe+cfjk8Tl9pgPgibGI8hZd8ou2G7hpV6ZYvkK93Ayu2iYwKlsOQLbu
UL28L/4F5lhuaGKm16hgjQQe7HGhkKyNRlY80w4z+7y2R2L5yCPwIwqWJmYS43VbhbGlWdztj67F
o4hbowRNVzV+SdbiLcx31xlPCJRw31ujS+reT6mHFts+2n3FI0zpiLK820eRBV7f3EdAFakMog50
iLpFS+CL4OPluubqDV0L3L1nkWwtGg2W9r/CYZR1jvXvI9WKlnwyB8/llaYH4zxQFXvErdy73Ucs
CEzrlcgQe0kLW2kiV19USvu6LdrqVRQ1JEGj3vn4BfGNHLiBcxAZHR9YIBaFR+aobJo/F/EMM22c
fnAL5+YkPk1/Zyn2F0WWTWxIFFVCLRhIXfFJtNXgcQPJEx781416DtSPoVSUIUNY8z0BT8g7/Wsr
vNFhL/yZ2manNJCNX81736NCHIVnDvVGR446iFyu7kgruoMgEFKZbJa2rbxaGjFWfrTt4I3SGV4e
MLWsWWxAt/3W1iMIGnNu56vnoKt4rzyBJEmx55oNHkOuNRRo0V3hRXBqRmsRyh8q9vD2Gv6tN63k
783W1dmhMBVXiTFWlmAexCP3/xCpJd9nW+qVmSMymec4+lSTaOwUWDvezHpwO10PvIrtItGAFNXo
9wlC9IdPgiRYMAU4IS/o3YX9S3H3hRiWWdjnRbY9ZFARodn1ELNxoXkBMlSy3jTDEOqEnVaLP6GN
8lPpxAOEIUv1iPx3wbPcJJuhX1j2BVdz7DFB2DasSCP+tp5xFljhfy/1kRfBJfXYeZLdIFgCzMnK
tOhyv3/8vyjfr6wn8cNZmnge+4h7xowkjLrX25h77+EOT+WRonF52vgrwSyuqUlfEzu18Nf0kpxf
zVvenOuqIwj1w6j9YijE23r8rYh7pahG8h8KxdauGviH0vlEhB4qbdOAI/A+St1vtZY/OxvknPab
2wBq6eQuQO3wWsGO4X6Lf6mxmED/UINUv7BqsxPjKbKd5DIidSpfcB2LhFHzxUDYCZ3W+BEGDcRd
LlZElCw7okMWkPY/UYQvcBOwO0Y9tUHX557pPRI9pZrtENxatzsLoymhX1x/UjHGLsx9LpO9G7Rs
BtILb6FHeaXwPwAqTJhmECIQzfsBQZjxV1z4oIRfdnYYGB7ArOAdoqqkW6q2ESVHhEEdX9RjfYkE
tSwCF1IMkR2RwnFtbXfZjGQ0DAKMmLn++mbmFDyEmzj/DmfLVLT7EzN5le8h9NQr7q3tRfE0vL0C
6AfPTxqw3Rbqt5FBJJTDKcT8jiubiKbxrs7SrZhL+AMIvEQ0c2YoTrJQIlm/pt6/xSMF+q7kFqTX
u86lOTUmx1NxDDJhu6Y9RtFX1392ymRMlSkIPpnC1RQTLSVad2ybIZdiiLgNffm23qLJEW4Jh6kw
hvl/pgaBV06ZUIXXdcQmO9C55ZOy1mbQp4D+BsEUB+wB4AivfXV6mYfVRoKQ9mgnlX3zH3xPFFni
Nwjuj6ISfvcMWPV5sJ5nkqPv3jJlIyd1W/Sw6dTprs6FIUHPRnWzcJ8DnPR6r2yDV2NtwRdSjb2e
rN00qzJlvPU+oFUnt/Bgv4prUSTCECkJyUnbEb90BoMclwh0CFw0wUk4JLscA9oC59AEQHiIFVQ4
aXJFWoegTQf+8jeKy8pl3gpagU+/KrapwpN7ITJix3HvjzFH6bNcd6CGjnLucym4Ee6YMGuD2lOI
HG3DDvm7ZLRJ36DOwqyjQeR0EktaMADRSHnWx5j0E7Aevk4RnjMf1aijBLayZR2PcdJnZa3nWalk
IJEypbLP6efFFjtWSzfak3SVxj+viWzabBhN827O40gRn9OmeYKJeE2/fWOC98X00YxTyGclBtiI
uZFFO9C2ijg1a3v3SyxbsRoJ80+LGjK2UC+ut4mBAXod+xD8v+TkBfzoTuOdXMQhKKpDrKstHZiv
42TnEcA1buqefWACf2DNOn/U2D3LsYotPBdsW+Z6+IiwT4MKzsZBRzI646NR8C5EVWJBNbnZzGJ+
iNIKT90q7SQ+p5ptW10O2cEZhAF2TcDQMUMx6WS8YFHIDfk7J0ZwwqBXiSlp2I5LGZbi6JFQOvGQ
hjcw9n3/sGTKkbWzTvVSznQu6RpmCyNI6C8Qti6MWJAOFzqPNHAgqrnS6Gr2HRBgFrd4G15WldWm
TILPJp0Dg/qpGBubIAhluLhvFRuwyCpiRSXqxAbt5mFF4M6P0GOKUGMZ5i5fd7RAhaIZs7v2wUDD
D0c9A0zzRLBYz2KyYOwUmecSnhtURycYhrSugWr6stYHY1OGlPKQ/Kl6x2Gv8MKp6RX/3M6DOPHD
gnOeSGzM1kvCRGhDJB/K1wWuwK8B2kcIA4XK6PgCjY4tIAzCOEgS6KY2uKDMszIEP4ierzAhWDgT
aA2f/OdbARVsMDO6NBeM5ph0EqbG8HqonSrfuT7i9bkcAnz/TxJEu+P+NBvNXOtmWcXPmCkdZNGJ
gFmjFU1LjSXEDzyOl4Be95aacDW2qfQS0o/o6a3iwlOTV08ZK0ofQwrfQCWtd1hE+d6kWgmpI+f0
fIoQdORzN42LL5K99HANqny9Yq18EU4z92VuARfE8Yz+PeK1gkXLpFWMYI+sC+c2P0OgPBZyqkMe
RhYxw5mRbp35BlceFOFlT77aql6UfEFPPHpGy5reM09dd4CUDUG6f5GqFLp1ZJ282qPAHlAqulrY
HoP0iOz55rH4eHpYlVlsT6/DA8ae6o2XDvUNqARQLYbaJ5C2ml68mAI8lkRSXWpbLQM8sThLlg3i
j3tXJBykBWiEIVD1YK2l+bmlZD83VJ5Hv+1rPogQ79+nwB32FxtR3nUDStR7qOYprcxi8zeoLuWY
s+GYAPeRNXA5LNMyj6+CefT801Hc7lDmEj1vsJRqEOv5uQkQ+/cYvTJXOScZIRvMuBymMIp0/Qy+
iYYYwQwy5mKZbCAtHGyafUv97H/zsiqB4cHrIpZd8dPjZOwMe3HF5L2nFqoFnEtNy25v6UANKB8D
5OxU0iIep7UyEvWIF/iDTz92Q4xfwqGL56xm2pbjBZsy2HfhhscJ8Tm/+pOOcT/kXP6i0KyJ5Pti
p1Vz61F1q7HbWu6LYnSef100gQDx4B/evgwDGzx6jdaPXPXi3NgR/WxJudykZI2c6dZxmFZW9jD9
ehpWfnujC9qgPu00neldll27knZ3B3bX/1pNjiPro3TPbF2y1lPmj7SlC7gf+SuhpW5lfKucKF53
9Lj+3a7ra8BE4ujUBYbmWjIeeYuszy/hc0Yq9C0VrnvZr+yc5e8sQfdHBvSUk8utz1caBocRhz4P
KIiFPZzHUK+i7bT86nGN1AvTNC2+NSO3spcZIvstQj8QTISPB5bL35GbMR3Ov1j5GDgKaeaQdyQw
o/a9yjErbdukFtRlQt/zOdVQk/R6Cv+mQu1M79BaBifI0umXuP0p0Mep9M5JISaJbixuYsC+VF6m
3DKUGGwU6+NFWVWi5LomD09W4dkl3QYVfOqhM4SbeEogl7auBMaSuiFlZRshC5rJrZHwKKHc7S1f
i18WZu2z6cCv3qQRQ6PNDShqMPp3KLrBYpHbRTiOM9NJlV3/vJyYQCMnQtKMeiCusbbtKXrLJbU1
bWesk0wJI45db3GzpkUMnY9eeYubrM6JNvHAqT+H1QjRZ6s5C8MhN3xgiMgWAv8RFbCdo7lO1giz
3xCglPHvFsE8JU4Lnq3P8ff71w/NCut94yuqCXEiK939IVxssRP8cWZ+Oafw4D6GkLbsnR6ZGY9J
EMLwMMdqr5KP8olvWeRL2LNQqXLr3fQ65i+hiMyytp+tFlu67+IQ7KMTzqBL0lDKJx5UGGIBX0lC
VuA+gY1gA7kGdbysHn57qsxhul3n++a1alOtwZmICYqWN4BzxS3xRICnaWmtB7NtaxeRAqGOAk2x
4awtt0s5muwXvry3cG6i395LCdIQhOWvUPLu3IH/MBxmWgsCHxNjeo4nw9hbFRrpS08h8OnOHgGL
9d1o78rkFFbCxFyndbLixRweb0+Axv5YAxGnjwhPU/q1NZG1SyzCfojSMf7EbY/rGlyU7H+jqt62
L2KQ0wyy0o1uL9nw9N6PF6AhXsfYalHi2d3RTWAL7QxM+fIB4GGMaDizk1GzyOZ7I0GplXHe7NgA
TFx6JdS2SluUbFQjIz1xqSuR7rdsOZycd4LwnkbGvchDA4b0263LVZEK4PYPUfE0JVXNf3cdeHGc
fGPyxGn1pFvHfKkfsNUO8cWikNuRmuAPci/TkNY7MwBC0LQC42vursiKwLf8gi4l8JNXsF75qhbC
Grg8Ou7F9Crv0o7iQ8EYvxWssmHSRhJcDvMig7sRqIK9xQW4aCDMZdsWS8/Oa2F+alYw1k08/J4Z
O0Vb0ZbtWtG8Ig7bxH4ys6QSGUdHLWx0vZLqxvG5PzRfepJIYrBxwnoj18fodbnxcTQxjMox8KKz
nOWAPlOS82bi8ORupKc4dMPKF6FNGXB4A5B9jh/Ed8dtATDARuMHxh35bSemi0VsvrvOSZEIMBcw
zfTxs3oiioiY0ibT3+5j6SgmhiQ7uh87GXLcPza1Qw0kvXq+dlKD0/Opge133+cEjlzE8+QKbRuO
7uXjwdWd0U/6ETkPMye6guXr4UbRCYNQMR23TgPlk/T6UKpl0KP3tXbIYLjyfFEKEcX7WC8WWLOg
iDcUJDDKxz6eW7+ZH9HXI5Wu1CexBRjEf+Na7rLlih9DdaGQyNvjyCPrAub8LPH3800lPEotyEcU
064CDXW1cXbfNWM9+Dvov0BNtNqEU3sic4EU69A4KokgLP7Ox3Ked2CEMwCZhHXI+aVZA8daHxJW
T39+/Okz5MhmL8GK5ZsFfDWpWoE/4Dy6uC2O01N9XQ3h8pjOazr7ju16d6wR426Wu8YzZfpISPfj
s34I64rXpbxsWO8BXZwoFNAotLcMYJzRu95B72Y+yF+wkROTgjTtXkFqbrugKEfDv0WIquKTh/N7
3Cy6s5XHoGh3HDtqv3AMnx12IlX2eQHIE0a+sDMDLR1QBBiLv+blLMG3KQrFDBXWAm5/OyTci7oi
NwKgKy3sHDsDUAfuutPPcECXmxqVQmZeSil36DA0sa8QhJ3yycc6XXv1XdQoFiXqMNzt2ezR+myn
z2mZirO7yLkveE/pl3kqk0Or54wXPv9Jo1BquQ9uw/BsHZVx85d1VJK7VnC+9H3UY7mzUezLh2iy
T7BGAkYx26syGjTKtQw+K3RiD/MGXjfGQGvx7AgjjimxL4iPdFM/KvxHj6zXGHPxNs6W/cTv+cjQ
VftjqkplfJkXZn77m5PvMYEeIxrjqJjPXX3I0PD9/W68gjLAC71j9xinuw9cS/HPiM8Fl/2pBTO+
W5Nu8kMhrXGXJuv/DZrUkyMdjG4D06ao4OqqyGeu9p+Q9z31HtdcX5tnH0zKQCzc6DZf4XdsBLhG
C7beetAf8GobLTLKr2T272nPLhQeAjWpEpOkWh2H7+nmpGYSDFUQjtO8Gfsbm39fORkn4OBdeh1s
2xRrUKrgHSKVAXtXw5XJjDRdP/m1uB6GGBoqIySUUozBc9xb857HPr0trLfjiqsOSFEZQv9nxEx3
EhMl9P+PHrm8GPQZcdbug7TVToyu9cNh+lmNXTDkZShv1zp7iXeUvwHMgeWx3kokJyfEGd6WAqUt
sLeH0znYJgT1AQO1ihPtspL4Exwui9pq+NO+pS2NqMfy/8Q758iieeOpN8WaFVp3lgTj8gi0/hNC
HACFM5vHb7zZ7sJYl66tWEsotSOrDIxH1sTxCQu3JZECnEZADFSytuO/H3XzrUja3DMuC3NtqcCb
g+8yVf9h8hpr3PDErB0sEkefhxKeUTd28/RJSawazemFdPUPZN+WBoqvtIFMUIHYMSQ51M8jp+Y0
1u2hweX9rO2YpXKLhLbUQ9VaSdqaW3PgnKVXQX7+l9WQKypsWc21GeAvBTAAIgWR/t0/g+cHk8Ii
vdsl84rq98/DB/vaYL9GIdkM7TEhIEUg3moX/kHoCqtJjMIMJMxdO0QWsIigksSNqUZo+Ls6vXVc
6Og2E3dqGWBs+WP/oNyRcLZr/deXCzenYCLsCwqoQM+Z4pIrze5sNdRV8gq6rohG3zHN0/xCyrBk
REZwMNm5CuDg16l2glKFy2c6YRTVQFyvB+pISLWJvFmMwx5Izb5j5Z/4Ho1NKJQDV2B/d+QWNvI6
JTsa5mcZy8jKQnd3yaOcIgInxhaDDtVFwMDxGSWq2EI9qcArlTWjRgOqz1pGCPrRRovLW45capK+
zSh2fMSTOHDdqljCY0JUnyoD32FkHInwNhIPPR6pTObnxaOrDf2gbquXbG7B1vqYHmMPrwzC4gvg
B9Eo4MxCTbobdJtnqzhQfuzMqSByG03syG7+wiqPu1nKRRSK/l+w5Tn1c/1xkVmvwvBM6rPoSNr+
T6dfm3sogql9enlsESX9DlM0BQ+dPa5ffsQ2IiIATRIhIY3MlZW1kr/+PsU1wAli641KIDL6JJOB
k7ttFZDQxIJabQ==
`protect end_protected
