-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o9vZgYAaJ972TVO4N3VQ1Z+z2zHbC3Ee33ylx/BotPOLtoAC7FdD3VuSKPTIVON02YctOn1vbT9u
Lu5nrIjKaBUaYJfUHUsQC6+57npDkRnvLPRqwmiKXBtdMskuRoxFmE/4Vts04ibyZPdIz+M6Eai8
Xsx/IATmn1jDfQbZcs1XZUURNAPfTKx5wtOD92FCs+EK+c7enqIqqMEfos1gxlrR4keOQ0Q9NnsS
b92Lz5FbPh+sZRBfZPUsi/x0PN6jQGoPYhpbytQpxnw3fse84ZUsO173cLEffyy3FNSQwYC2hQEW
52eASotPS78EO3OTJ/EJlY1XqaW/uUT5v+bqoQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
SSEYNFUH4DzbHymqGtiv2CHTI8YSFFMu0Wc7v2aiFwQ+31m52iJDXkJu++y/U7mq9QBLozGCig60
+vwDEyXxINgQDp1250ttvIzuoj0YKTBudzOD2Xw1jveeB2wNQjb+7WT4c/yxFTR/luCDQ0nRD8Oh
mWUUOeHA7+SU36tpEyFeVTNwiTdMPJGW4cnwFUzQCU+HauXch4p4/kz50VPX2c00ulsn7qXtiKgB
YMi7of32VRoUDXBP+8AnLSZQzgREPOQSL0UNY7xDdS4X8CdP/UuNmEIbWOP/5mv8ppGgFyt5VXSu
OPDMaXfl1qx12av45vzpcnJv/Er5w6aR4otkOLENRZBMnPDswOHkGAEm9yyC/nnIs6oL9+QcOk0l
IKPoYvsKUS5HGeXon5nqH8t/J2tfssmZmBOwOHKWhbd3xZzP1mDcQWv7KvVJ+I1E7MaOR474rMBY
9kcbRtaEsPypcSEpFOhoSGQFpHCB6jJEomdA60GgBh2bpeHWrtRaq02YXkCYJ20UQC+2vCWW50e0
xvShC+zeJ49jQVDbFxlXS48P8Y0PBV7fIPr00XwSWJRuiX60vAj7qWfj9Uf511uraZO2ffKHVXQb
9mCoE4pyeC7xlZ0MS3xFeKy4yFyoSjUZWzL0YyHvoRxUZrOR6yFf1CRcjg9R7RxDVMh8ZHIweil9
76oplukHL8XHM/ZnKciaoc+cd3r4VPDQ2MQDKEConsE6tpqQWwdL9bUqU43hsGCd4afNA/EjngOw
Jbc/o2M2pZjggiQOjzifvFqj3AWA5L0d5CIPI4PcVaArpFUbs2v+laa1c4KqrzKtlMBZGzgeciac
17rM8ShDCtbMKDpwFKMU0E5rV4qZHtGjlb3JaKxdyuKANconhxahGDy2zS+OuoFsY1ufnPCATmdP
Mh42ySNmZ8+sFAddnC+b097ZWhXqzS3em8qYuD6CBIOUKf0cGYx9Ai9w9x397mmwcUDd+JEe7clO
1KGtNJsLHBQPBhsAn31VED/3cnaS5HvR0+4BQaoQMuatq7GTmP+X1Uc4eblpeArZQ2YEBVT5B5Mm
u8Da5z2+AAGjFdiVwOlbd05wV6XoBMDj0RMMklsC7WmNXWAU5vVu6AruBdjdGMcNttkOf6UFlG1C
ow/p1S5W6NvuBQuVcgCkbmClNp6PIaadGD8/JdLjZEpdAN68cN9fy5H5AvWxO5D9wi5eU/I2ROsa
S5r2ZyNRYURtZ03WMp0A0veKG71skDDf9MYElNhFeIdgXLbmsCcFxc0jgzVVq49ElKQPhhXKki32
2Kjg1gPOxRqZOaqEl35OTKoucihfuotSdyDrSn+22TWo2/q1AHQvGtcrFypmAm8dVxXAqDiYqMoR
mnN2qT71d6DtoTlvWY6DPeuN7WFzxR/OY8tDxEa6kkCUZLKQfOXi/HL2BCIKChokrp3t18qjB9Zj
OwDSF4zfqmeVlCbEmTm7n5Fl5+pBDTQnml2djPHo4BFjXx/aAxCuD4Hdk0NuqWvc8I9l9yLbbQuE
dFV1zsbrX/07avnLTXkY66VRIUzjTkC+YdATTUY9LpPSd5JKP4M4Kcimnk26F781JpCnV/0ntpQO
u8Z/yny7g4p6ZAESEsIG8y8bG3Qc3E+UdD0kiXb0CpF4Dah3f6xdotcDlV3Ixc6moSgykVp/LQhQ
ZItX0Hju9Srgyym8N1TsDQfJAC7HEUCHYtJHCvTjDK6HR64Tm5VOkK8OlG/Fuj/BCekHh3Pc9EDV
CaNXzmFpISiBOr/4dMAS31GKFcNJbtB5kUMebWaLXdB5xpBchpVHrkewuRzWQDES9ahRf+nB9Uu0
nxNehb1zIfoGguV2kspo0tHx7SIkZJ4+j3JsYBN8DR30yZN/zoAcMPeQWZzbLOBAoTedvgdeYj3G
lBjBMum5CYblcg+xnl1PNxQmOKPldqwIeO2GnuD3PxU3Lm4kqdrnaJSpyqs4Kqkus4uY9qaKRnBJ
SY/oTmIwCJD6DA1X+47bNliWVcFi0s4FywRs1r8YpMW1NHoZwQYH+tUrrNM8dRJeNZsQo7EwyzuV
Qmtmebg5PwOoTdJGZ+N6PQoVRFsc22FZhiQnUf0/t/UIwcxRu06IGo9MDqg0kN1fysAcTRN4xq9E
+KuV/H1siSneo3hvgHBSsv7vtGTG0irutunO32NiJqoxHmTJb2r6ddp+t+10eXvJXNIeiQm+iiuA
i7aj8WtDpH1FqpeDYZA7sYk06GEZMRx6WxVH7iIEfnH54eHvM1DsSdIfmbiaEyOFn3VPkql1B6+z
Utb8rH+aAzFlwO/JcRL8JbrWnrgzV5LBvVN2nr6/OJA+E1wfdUCmSZDq0Q3AWtkUkWMdo5Y1VHtE
jhQdRnjCeL4nUfCfkjQ6AsJC8gH8h9BtEARHSLcX5Mt2BAFOc45TuqGfBSTEsDQFe0cFCU4XSh51
C7R5qROLBgRGQ9yHy0wp7rA/PxrR+BIJdSGZgSEzbvo9o03nybLtdPUQnOKcn2/qDp3IrlFvrUFw
rJXf8QauDVKwBnLg3tGbEctKPDDBeCCXe/DO4IeEeM4i3BrhdXX3nnH0P5sfEqzFa0ApWfbxkFHG
c5bb0XG5v7MJr9Oi+orLFUZbu9WzCNXwI5ZI8z80DbBXBbLTDl44XmSVr6bXDsFZYbQXNZt09LlZ
sNJgd1+4PR3o8KO93Bmjqkx6TxcGjbYvsENrKtVx4jlTD8PQRk4/9OoI9Xz1S+dLTdQR8/aZkQCQ
0sPRDMV/DZDyM+ugl64hc94M8+3UwLEtjixgAsT0YrIND6MzZYxJR0/UiGqBzZMYXAraQIdPBSQq
qkHGlik3XC0osb/2A9aIpPkuxbpvDuJStFbsORi0inVHu0h7EKrCt7+LTzDLflwyuE25TEj4zDaX
Ym4poyyz6i/I1ESmGbjHrLnHewfX6k/wWVCKsR76i7SFJd0kPhv9iLo0qB4+tg0ZDuV3NFLY41tw
K/lBZJwv9CRLSXluCZvd5bxNkdyfiA4w7GNfxN/X/8+M+7XkRhif3g3OllovsScai4f3wt6u1Fi+
qGugiqav57s4+9GrkF3Zwb0E1bznAMlFWBv7dZaS9nlE7n/aSJsW6EmhDCGBcxjyhMtlvxnoRy9T
DrH7y/k9hEXig/jmTMlO34COa3Tyswt7lSgzFBD7b64TmrfZkL91a5ODiViJyj3WI/P/lHFgqRt+
mIchU79oWwzblAVrdELmgD5a+LdzYCRfu47e1Ffn3yk6iccZc2JBqHp8OzkoP5NnFmQFCWk4RB2c
kUt07awZMxtqkxIJHYCTs7DPnNsqfUbQ4pCIcvvyT79wTqNiqxuo2zTkaC+QdxHQrROexPymAPeO
hxopIrVz/UIM6LiW86jS2RkbteDYOJd3cGr8DfxN8JjNlovdcy1jCpF18VQLnbCBpbxlUbDpvKUI
q8jDJgaSgBjwSpnMyYGKJ1wn8L2G6UYVRbBujY3gIeFzcYopMQTDVEtb7LQlpz7YO2LuWKp0O6xe
HVxXF6HPxTppzxOntW4C7jwBwNW2/3kpfvC4vrdgmLMDuZeR78yODjygWtv3vVgZHD9H1eM7+A2E
MHeK9iagk4ygyNerDkEZ3G3r81CWodHfHuNoRqA5jg/f9A4CXHLMWuBYiGss+2QxDleGBAP+eS16
nqZsiAlzYAcstp8uGXnq7AC/cmCZFg46O/AggCslYkJwJ66TagFBwZpYwavXc7ZpkysHM9qjJyhl
iQx+QAenaGX3v1vlaLes1Uz+R7lCQFCUT6FWdf7fVX2lUsGDWLUgjHPww3bEPY5nFc/ow+hYYjr9
m7OJAmpUARTHwsevCralRuzEOLxxbu22enLfG1s0jkMwp9GUzg5uqBGK/ksLYyMiEv5n4gi8+9bC
ASlMStrA1pAaBlfqCuP6g6aWFKJrk5jn7zyeqCtIvBwK/f6MIWR5HbRGi7kRVthJFyrwFEuJGutc
acr63121ZUxld5rI+7LtBfvCMrFk9sAnxpgcek3oP4oUxjIVv7ESccbFAnOLA//J02a1I81TwMPZ
mhoPsI+Frl3Mm51Pbdms1/6VYLzP1xe2TYcqJFZpxNX3F0oPq4vhwaEpkCJuL6wNp3g6rMkjr2yD
rpG1XcNlSGfzm3ey9LJv98yP81QYfMuNrMpPHKbQmGBQAMHs+pKMJpEJEJbJb2H3l6b8ljEauPyp
oHJAjMKsNViWDN5v2PPg+v17t9FgIIkJa5H3a1XkosARzauvI7mODf6PvA3Jb6XIRb4y2k2rm26S
wOj9MnzuBos5ueu0CCcNU1RboaDOakCkYdWNzy0PugL0NJnYWW8wwqH0aQI9Z3jEkIXQyxwiyvgd
dtp1/uOd7Cgmihvxfg5E5gnsbEeJfCKCUIPNYv5P1kIlpJfBFm47hYUKr5W3+LWsMpsFhpABTxhi
DS9/r7p6ZSo4GvVJrpuLyrHT6rYPaNsCCJxed9whp1OBPiaSuvH9UXV+X004TglYjkurkP/1uNzo
LCrTA2Gvv/YXwZ+OKQP022q1tjts3sut5HajfgPRL+5at3tnndSn7WWZcQTzJ1Bmmbo670eSle+s
VtJZX6IfISCnBPvY1p7d8WZTNJ/mmaYsnAOt57kHziy/DpVjLiZAAuzh7oGoIqR5PUmEDLTcpEvF
94Uiv9il6giPnAXlTvX+x5ydZpC/Dp2IV5gJ0i5/IFs4bBeUGuJRbMkTTgJfUbymu++fXU8O8LhH
J8eu9WQxoViW4FCyndn/fzvngtUWLilq1BhaJdQjkN6SsmoK+6feqB1soYr9NUDuYS2bD05f2etA
+pY/FN/qorzM9vBKpyAtwq2wrbr4QMPW9M676oQsfa6JvAorwSoG4YJ/JnDzdN4hFccPVRFHsuVu
WdTlhaZpUblcWbOiu5MDJSr3McgIW2odD0JczwfnnLxN1zunARrW+4/fXRye9UUDjc6/oAfXjCXW
Rj4fmAaRJ2zIssMivlAZN4LiDXWhv/zVtzOIPdxM7LtZrw0B6nUZ3Ak/g2U3vPBegSRyY10qljqW
aW2duHJZZH/UrCA0hA0ewRXAxPXsiuIkx3LmCMr653Wbqjd96GJr7+5aCQi0BedGKtA5TbMYuuOt
0l5DtK8Bx94DOa4WSw4nnQTRFzjk73SthOpzeEeSuvaMsaFwjlDH/LCuagHCWb7Nzqe+Nd26oUix
aO8r0M11bmUa6rINlf7LDz0NVM4ZNx3V26W4BA7x62KDJIrn44oiPzm2sNsl/SLY+e1eZgqQxoP1
gzZTbClW1fUM12iXLMMhpS/MAvpZV6DvAyX4nPbjcaInn4q0SUz+VagNWYrXkTbIWaNDeuY164Kg
UAEWr8fgaqRRpA3C1hYneqAmSikYnnPNb8HwmUIHSy9FOH5uD56FeGYVsgV3TuW0DQumisK2UegV
j24m2FpY2X7WdCt/NcMVUFo1L+TZke6oEUtfxgrlnNs2LeVoBHci30f3vVfqDGDv+KXtjmr7dXLb
bnbo2gOjo+/WJPFWFUlK65tGH4OYx06Ez57OaRylHAWBeUdJ362nuIAj/GWw+EoNw462Z97l7bRw
1+pq+89WiY1G5z6Sk6qMWNTLCnVItPJPi7Tvlnx5ALCs7mpGGQ9n6P3yNlA/CbiCI3GmsPzSK2wF
u/OpV6SqFrFxM+kJqp2CXMNZuBgzJUlnA4X72jdWpxa/xJqrfVU4eIvfr/1+mGXmUIZTwjhc5DxR
E6kl049qHVr6+KrMzzTZx4tHyUvS8A21Le22RxD7q1HCZApOe9D+355abwmHnAh1X/o27sZb1hXq
4tBG6E5hilTn+bwVA1wDu/Lvys2VafBhQwOqaZXbLk/TymixitGhTLD+2y/91g+Vp9h+BpOFU4i9
bVdcK6dFESFCLJGxX290W2oyOSQCf6DbHaH7kWnBSQey51mM07BgGvuJ9N4Ad+thlJ74ywuTPcTK
RybAXEQ14inSP7zprP29zDfJU+xlGN/t7AbvbcvghJL5C5LOjK3Q+hVpGWSJYr0H67wUq2hN0jTk
BirdA4XUpZUo0NhTloNcwg6VI9Blgd2h7UsZPtjpJRvQJPsgg0i4AWbgr1MlFk2L54XJXiN9uIyN
dXZ13hKaP+qSIp96zeEecKS36pM+98xba2XXCEnFeV2peeU+xLWGnIKQ8D6IjnQV/dvOodhfm6yu
MbncS0GaAQ4QBj2iDv0N2ydcHaXTOS2jlKse5av7aY5scONKWp3TVMFqGEj/OQ/yf56puSJdAwz9
bf3vLggN1T0X8w+Rv1qh+xAiyhbOza/zHseFgY7OM5pCNNIhHoQzHe8uR5S0nlCiyJE700GIL6dO
1ktyy3Es8QC6W/psbsMJ/mxFQhAxFDw7fwZfGyLevBEsKiJNmgIcgpwnU6Oq7zgRVwQZn79chqkR
U036TL9JjgIf0ytxebr/QyU+1Opk8tSKOpMdfUqdUQz1DwxSkWKQl2m3baepD1WKcDQ+Emp53aQN
eeCewN+HgRzlZXnqtr1NR6jzPhe/9bbPAD/cydjecpxcGtuc+nnHmfOXZc7eIlEkVLpm3e2aewgD
FJUUmeEqMYZPI90o1ZJUuzA8BqecnwSx55TjEB0QR6Q483Fk4ih3TtRXVjwunjM0f0veyYmi1kXX
IhVj19SolTjf9lkZuzgxy2pIxrDHUbBH/FcEZ6CfV0LSTTbBNzUweXCk0LzfsR/OAUf/jaEQfnNY
2ulyA9vTMB02VL0JkjuAGfltgBabT/rlNbJEyJXLKXYsK2WeOwJ4VbHXOxay40JScdrM3TMSAafZ
rRzfD7S15EE9KGoKw+lzMngikDFSPBLKCzEodt6AAcnuaj1pgGrdcOY1jTmuoMUJoHXiMRcQ1InK
5o5r6FxYJVEBvw4qnsIOBKUZojRiWOkPrr5jQAUvY3HMvg9nphOF9LzuHlHgfCDxRwGSoZmAw4Ue
vE67EF3AJCEB6cutq+0hE1YVonoACaZOhr7t6BftToNsQJRKufIebK2NrYQWPlWuK4jkdzRfGVvL
3VErJ9/PEy6Gka01VB9y7Zq14p/33VjVC1Ko86XBJ0IV7H4hRiumgvNp0B80jMFy6fF5IG1HEyx7
f+33RdWq2MeIgePPhSH8itwz84EN4yjo0msSuOGWlxIVmNqewA97zFcdq76lQoHvDIExmSiwbV/2
LyFa5YegvdiC4NhIL9NJ+lMIqJXx2csmQHiB7SrvrXAqXGan3szZrsdGrUsM07A9q4IB4w/tKC1l
yvOWw3a8KmirLYUhRtWEGafjSZGu/GMe8lIDInuwcDspLetaLTXrJaV/6O2az/7eWB9VQbOPaoTs
bOPcANSQ38Yn5RUF7du18itMbQJlUKbh6Q0QfFylNqUZyuGKjUr87VCPgrO8SgjMlfKMdSNebCbu
qjkNULQMb7TWOZkprenHdn/s0nsV6s6fw6AsMb4ZlOCO0mcSD06WdNhJTVoD3srPyUEwP2WvBGF+
GwfdPa+fjS5454S0RcFVzrxiBwR//R5Dp1HkuaOHLGGXUUT6NdpShEUWMKohJK146q1/MVYx6F0j
EP/Raj932x1MiTb0YA8GhpWZwhYcypF0Xdf9wOSBCH/wgjttk0VCmZ5vK4ns/4KnQAKxF2/1m/LE
rFlk59i6qLc2r1oTpxsVmz+2rT2nid641UYnuujBAu35MRzGbhINyecdEP9R8FvpTHWvnhKdTbo7
Nk4uMqu7cG2EmB/xMmFHCopAmxgj7cYsnYa0DbqguNTqOabW5IY/iuoPcxZcCuJI5leF6Ib5KfWa
0X/wEf3TgpomFubg8na37WaQMiYpTKqzBkHFHLbHzZ12RmvOcZevKou1uPJmedQXUJNrdiFERGSD
fD8rTsIZii1e4NsbG+RHd33CtbWxF2yosI5d+4wfG85Q4QudxJ5t7pjNuJIs2+lRH4Ifs2z7e7Bl
7C6jxmhAQyo8jNAR2D5RIDlGmh2Dpq3y140M+j2NGRtcc41ArbexCh7RypISxjIlNQf2akDpAtSL
Iv0+0i7+rOXnpthCGS9bh3hrgp2rsm4AKzhniwOz3bR4YRkx4kUFghy5dNkd72nBrL57fGRb0Zff
BREqFgLD975qeNRy6daSEAQ/lPPx5ZOPlKY8kq0CMDSXglYB1y37sEVYOGlY+r+ou0lhK2CaA4n6
i1Bba61ZfkTqpYqc3phSoVDugrfjYfHLNpuUXZMCBeGBAoqtDGHW09PCkNCJFAMfgm+22+q66zsn
pzzCyj+r80cz9g3BbJID8bwiH0reOFRdhyCuHpbKBAZraiiF4iXcRKR0ooB8Ghz5PsTWUseyXamp
Octna9NUTOfX9aAuJLFvjwkvnAYCl0jGq3/EbU3t7zRqNR56zqKbIPdlrVxapYyUuKTDhS7Xx3aQ
bjIQedjbOcKvCATEFVkqITgG2cag5ptvChVP0pxCtkpe+qrQhr7gbSbhbUymKlxfhbsDEjeYnKwY
J3pgryXjlhGnFJRj03YD9g5H3/k9LOqMTYQxDMNgP9NTYE9yYfYf554qLYmb/+NM+/nAfNPXwMju
gYEbdAu+wAopChQOErRzSa4hgTzmMb6WC7wnjErizZRvtNSBqbR3BveKMo0qv1vEea/oiPSDzDjd
RAnfhgXMDMCc/9GNsw2BRVPA/5m1mbAxfdsfzELAQu42Y7NTzZ4AjkU9tqOJhjOWdprGQi8C/xqO
L8YvnpLLbGRlDtywKIShro+c1RZ7w0lWc65lbAvujCP+OH29ltTOR/+Hz9Gjt5wRXYXBfkVDgw3h
E2c8XHI9skwb81UQ3qUUt6jFf8Me9CHTtpEPL1DkosIGsHA5C75FB7dGgrEwlnb0tVucTZQBNTH5
9Yfq7qigJFNELDCWBZNxMkdzfHUBfAMUaaBEYdWk6E7qRvLMozahTR6rSunRv1OCiANGIdU5MvXJ
/RHWLR2MTJOUOT4rtJZShzccuxPF6sLG8Jw671UVMw2Hqt96meuO99QM58jMHJS1LTG5HpRXxEnV
6AahWBraO2A/uIUZj763rH+FfGxKNMhTfjMpy9af+17TWTs9VZFI7wnlaXhgyl9Z9NVDv99FCFv7
JM8obk1CY9ou+pFgQ3LZ1AHCNTNXDo1etOTDwerxXclWDcUk9biA+hl6o3GOlm55P93j2MOHpUBs
ujlyAHhLNErr8K9TV9WJMZIXgNcrM+y/0yhoKssaPSvy22C8aFTnLlYGwN1+x6SKVUKlIdrrYqJS
x2z0UBRKWYF2ezb4WjjOvFmL1ELfT1oediowj/jCQ4RqLmyAjh0zyQWXuhcy7qKv5WSCNeFYBwoB
G9hXl+8AxJ3z0orQoIjlenNh9txGck/WaTli5HJ5S+nz6U+E0AR8AC47AdTgNbD4lBgazp3klfMB
FCiXe98nSRx42AUmSQeVi+wGcHeDyE7+CK/LMPDmj9lPyfKNYoVWjSWIYxboxu2szvee54ELGs2L
9+gXrLHoEG0mF89hezPR07PjrSI2ZzqDuTq2CyPVHJNJ8m7Nt3qQLMuP6+k5Gsk5wrZhmDBBQrOT
Zvp/bk4AyUMQlbyTsXNTQcbYKQe37DdPma82lcVP43PoandmslpORwY2JFJ4uSkZ1PJsD6LBKns0
LIbnaNXNw0EQx3X4GkJh0o/bkxqi47O8l2Q0mx/n9B7ZW7ShQNOmx8irRTCfecwBsj2Xzs3xWht/
0kpqDK1+X/qodcfJfmUmlblq0VU1rF5hSA6lMtpiyy882S/7nFaJGsH5pVd3YwOxKzglGCgdzmA0
+zhde/wNaL2i5OX61qiIJLL+ruq+Jg37ivxSR0QZiuiOsXQOEReEPjbfCq2jDtV+OJmkoXa5exHJ
nRZjiKEHSdWTr4lWTlFQ/HLfGFCwebpEfBOtbpWIMzBK6QkcmCUFPctcVxJ3sJl+lz4mxejCps2M
m0vfiEmFQn9cdG/H4+778DrSHzhabTZlIlelhpDKbTVtIY7hSWgxjIuYxnIzuNktXcHu4BjT149u
kMXJsfxgiUMu07WLOw87wCgKgkL1cL85nJAMLnR77xJKkapowACmedW11M49E/MdVV7fqH81OCU1
af/jKlZPoLT77YWjLbChnT4Pw/r0/vxLaErTvfmNADJeo+umhAIg/ytVQkQtt0vQCf9EAglKfyGR
gOIEaEe03JlIrFOLSBl4heLJZDeOv5zIWCGL+neN5Vsxtfq8mBFeZM50mooBs0aZW8Hf8Mh3ZZ3O
Zrp3l3elvQ2LEate8V9QDq75d1nzNP73IdOU/j/eN8zMKKpUeLXlWpQglJ19gIXONhZBmoe6vYx6
TGUP+GYH+RZozeCgipYqbrXS5kxuX4ZX7W6NTi09cJnG2AB9ZdGufRz6EQI1ERfBUPw4MSimi7D/
ybyIoPahR13gjcjX8OmUgQfWFwmBiTxGt5WD8y1oSIQZjccSK8gayUEFSQ7LnBLdXzC3bAsvacPn
9paeLkZII9Ye+zP/sKTzO1DppY8Cm/Wi6F1/vf4fxDtOtDA7C6M+i8+RvZOsRAfxJX3JbJ5yn8Y5
gHAKeWeVPMLd5R5AMQDVQrVGZg25hdRSyWNSon9GIl6w5/ZCz2JrPH4j3HfyhXWYxSMtSggqLqZH
Sp7xWAigTpLwwHGgWVOqC6uOeJRXDUffu2qOL8l9AZmZHbV8fag0VefrNKkIUVB3AvmiFAVYAryX
JKyg4LNz1brAfBGqoFda89eKwWlgk7r8i4VH1BehZKTEs0RLH95a6cFqNxjpuZXjh0f0xYWvClCz
pIL6e3H9Pn03YIwzTuRsC39JV0aZR45tJ5oh+WiKsUAx2k+cNG634G7NNAIYSC3B5WSziGgKR03v
eTihFhxrRCGmoUcr/N9iDumRct4A1eOK/xNkv+A0driHolfpluXTc5/CsbfQ7swn+LrTIzwXmttz
Lfy3Tg8VbrUDHg1jjRKE8QSsjVihgRjZigQdwSJ/9JhvcqJd0cF2NFRuNjMT4V/6/n4tcuO27duS
vHcoI1js+hZbQGI26x3DwDkqC39YDblZ6rggNG52DAHuQxfNY4flnFGreRhBqEQWDDoLqchZAOsk
Psst+WCRo0OQqc6JmGAE0PT4MfSBR89BaQ2AlciB3pLJkA0MpQsqFORbAzlziXv8YZFraVIaK3K8
0rLObkdx9MVjTytfkeLclViGILP1b6vC+VNQsOljuoV9O8sSrKLHkfP5beVdQlAAGw2sgG1RI6Sj
a/mfML3cSDfic2mnkazNd8MqRYPOxNWPe4tCAze0gepNBheo2ehab4zwJgj7MLDie+zcSea5aqle
kdKYiICGVb84+YcY5+/ARE97+GpUwr4+/Inyd+lA05HdKZjoPQepudX4vSElYe0dG0Df/lBbAMFD
wHPsBMpjEL4YYJVyrOjxQvlBonrkJlj5/+RN8xOHyMVdyEZjzCaWTUuTDEfh3IgLC7o1XqzjaMvR
owJPeaYfVaMYj2XLptiPSh+byYhWZ6ZXeGKDQEqbUquqNdne4ystcmOJzJfD2N6c4CkUNYx5FKht
1rBnftBcLIJe+gbJrtPi2sQHDSlxPgVYL2zR1mtjOtJTtDkSxp9N9pJZTLNv4C1+b5Bq48ZL5MVK
KLwwWnSLAlBvGv+NI/M9UmmT7FAbANdRveVORhFJCLTEelNuRB0EL3FkicW2pHtAOAshOPSaS8on
vH7uhssEc5dopavBZzHBBbDHwUEkx1smG37bpEfr7WmYcpxvBm6xJS1dSugliq0TiuUdfIFIJoWB
dXbi/DqxaQotBUM9CIC8DWW/ygqwdNve/B8JRPvRwm4s+i5vehiBNvvS/ZlTDeSx2kBRuUOhXxej
LAk8FQcnIQmzTt4mrF1ALsLgu+pSkrNbwfyXpyoq80HAS3oplc5spLAwxUXg4YNOZcvAONMTiTfZ
Qd7UKbbdl/rOLVdBf/BDjFuIiNLElqZP7qqx+nBHCa+/LoxCdi44e/tZ0Puu/EFk/wFIp0CgBuXS
Dx8i3C+117q1nYv4CWE5QF0kxc7v1/OX7RqonmjCWcimDWvgUMHpUj+LxY+kqU5uwdMxePUBf9GR
mGoJ1KJfUNt9t3q+j6aK78zn1ZKkL3I70LOs2qtXRLpwvjIHlervaQ/Idr2oEvM179VMZJgSelE5
Y9W2gxhar6rdowr3X9VDs9qyRL6bucrvtxTbJX7obQuti7oOdYvj0I+xLFRZ3Nme9HHIFu9+lDgi
6x6mLumua+bUivXV9dfgg6Fpe5cS17UUgo7ZzDhVlSQpVkQSt5e7CMd5X3khGAXUMmVqnyff5c83
zCJOS7dtWw/7/Hggm5YJTHWs9T+VfSWq9RLdaAc6BUhmn9gQiri1ETh3hsX5Iqux+F1Z1hYe2VAj
EtCNToHJphjX0CIwA280SPnRkmA9AfqCet+QhZZl/xZNDcqDgm1iWoDgjjdHTJ7FXluZHusJC+Ty
dXUL+zoMSTvmx6OhYIVSUYFu9+JGONuMZblYu+Vy48vErD6eJz+rj+L2+GZnJP6vzAutz6UlHlGz
qYEKAB7Ku0ZdbxkERf75x8dIv+4oe+GbgEgDCJMhh5yT8Q+e2BXD7QorL/J7po8VbaeuUQaUurFe
XmfcwO1XvImqP03F3fNIeeYpu1G25v4VdCtuEdTOjrIBiImBnt4daJGdUaDugZgnGMBGKePE8rJv
B0v+sTNwIkqv1ZBwqj0FES048ug3ERrr1hGdCf8ylZB8XIrtMsz1qlizdIzFRNK1geFBrxiObWac
KL2DQyMG3DyNgVPs8NtAcmZbEKvZ3FBv7kYo70zWlDSmKJMe7A/OboaNF4zuTmHgeFZYG6XCcYRj
3dHRaYk3R8ddnwUNV0XBMgVWs72dNHXJMSMTLCR5QlvQM7cTYnOphVQhcKYYCG4My8RqZpZJs/Fg
O102ZiHikPHX87avgq3BnEXJaAs+zDJPljr5t5mQa6uQbz4fcdop+nYvrihxEeIJTK7OSyr53VV/
8XQOf6YSNJEqZKEkCy+IKyn7UjLIGs7WwFxZAlsECnCdTcI0EXVimJYglFOHnEheA0PNcB4QWoDS
EwSxgg7bYRVDE6UkbeVHSJh5kCAh3GB+yCPmpWFngqRndes3HboV9tAdoc48EDZrjE2Hx8u6AGS5
VpG/OjIom0axWqOZBx/4L0eLscDQrKnfLtovZ3JSuHKfz2L3aL3ZIDILCLxuO3yJ6+ONdliKzbD6
TVBq0Wo/NkKsetlQ2dUNbrN/8tDBev850yzwD2h8XsRB3jHfvU3KNMGtS8IIlVkzjbm3T1pkBEB5
jSHhD2VnMRbAvHiCgRauuoVjzLltPEL//R0ZiC6Cx8k13i3ee+TPNWQj06W6diZooz2sm/dfaLUG
Mwj8dsnwr1UcDe1g+djzG8P7O/yvF+0IHrBZ4wtwCzHpzh1crUtM0382g5CTEkIRN1JQJiJgxbeA
XJ9xgq24Baash/uug1h34IAunK1jTvqiKluQ43ILQt0GOe6oz6wLN/sMjj3tFfZb3zUgTcqAh01s
NJp3LjUSKSntNlGVXWS2eKKy4et1DIzIOv2eI7ObaFzylM0lZ1ZaeMAOTEqbNZyZRLW3zW8kylj5
PTOX7pSyghPeHBKF/L2aDa2CbV+neyIVf3wHmflnxxC2PtUOikm7y/V7EADXI4IT/gXZtevOUB0w
jlSirobbNVmJLeHgoLgR+8EUH7jhUNq4dqKmGlUE6+Y6XvCt804CUogx//leWKqBdy1XX+Xotunv
j4tYSUC2ZFqZjZmdsJihZ90s//P6utfduqTvCBCFZscF8mzHUPUroo34GfhtIqdYdNOSQNIH/GLW
9fNfWdV7d+jrqm/PhRO+xCS+3XqeMabjNmmquEIMNYGG3/2eoLXVPihfMecJESE++PBdBjjQFlkZ
mTXg/awCEnmta9qPOZLG4jnZhz2UioDa5V1XsowFHAEFOb+8Dp0E/lpxGJCrSaVJbLljgnEW86EO
9vs3TL3fygoGR4NciO5K4PIAfxqlqeHINTA+Kn4MIL/h0PwOJmzTWtaKIDX/mVxO70aJyX1ui4/A
3zaLY5kYcO68vh5ypTuDcMp0PsX3aikfstTNqd0GBq2NrCbH1l9tKWm98VrgKMayPlo63wNI4HQu
jzoStiQM15L0hluQ/v4+PSz8S+2ljtoEVy7KU3PAvTzKd7RKnISNGhERBs4f9vimnBEKCe6j7rIS
6ROgWM5cEZIbHg76KuFmzyp0eHOJPcYwzOUMonnL1d8K7hGzZiVsp3egxnS9j/vDolOuj0k51PKj
uYLNwCJQqOM2dxcXxiA1Emh1iiMsDNXzkCX0ylQggo9wafia/wfIKHgcnio1vqN9QVLTj+0Eg8V5
1knBITv5ajKNGZjuOCuGfzcHeNx9YVJsFAkF3p06uPm/ypElxOzRflN/K6Af2dclMgQDFEiFluYJ
gu2ATaXYti3Tp3Rhv/6zJx5g3ytn4uCsdoogbgEwautGEpi+P9naLkdoZMqdd14xB4YY/IIFhSVy
AU7bD4tsNxck29pjFFoJsPYZpo0zuZIgx6STSns9rjdkmQq6q4aj++WNXU8m1yrsPZBBS9lFN/WU
RgvufBA9b2PSsdHbZotISqONbe8xlQtGSlD1RPI2rAYv5QfYearUNv9zk9EKV0/NquLO4zHaKxAp
nhrKep85QkcS8eJwHeOD/zxwEHMl5wNgXHipUukm5IZU0MAE4BsQww6/yn7XZt+fuzWVnkkeTIo0
zegqlCW1RQPGv3Ddloyx0eXIwF6Iqs1O4uULd2ge7yGu1CskDELDdFrucYiafNV71oiFcfiDOT0W
gtsqdevhpJeamRiY6sUQe2qk4oi1miDreaMqOOw6vT3hE8cIyQEDnVo/zfYlGgorMOQ9IVDhG+A2
1TkA7fhJB8TL6HJj8uXWef/9c7/aCRESOnCOlQT+AXltoMIzeuTtm1h/pTgEGlb6mOhB3oKQCumQ
1tdXhtGJdoFgtI7SkCPPjpu/84EAefiK9OqHOvYobUNSfDOyELt5u6d9yDlyBVbQJbgOT+PYiXSj
OvlPTWce0iaiOUY2zXUdXlNq/1/f0hOOPreAULIPGKsLRgId0j4BFgTZrzOnaBvBUIj4Uh6V4orC
34TsP7Q1e7gVrAomBvPXhelnUs1JYmABR2RCG9p/GTZMvqYdRiNBtzpH+AhWo1MQ5AOuyfyaE6uq
Aq0NqwVJgS7WhPkl7Moa92WkGL0sxU9ZP50RRXhTIb5VmDcgi2qFWLl1ga4NDTn8e4ZDi0tmSY8o
QiLu1hF8Ex9NCEh5aGMvEXPr6Y3UMgTNeIrJqx5qoYkSw9FEgQLINDCwOuvvwdnm+Nu8UuEWW11a
LzGZmX5Jcn39P4zPG5eZM/jWrJNEbi4HrBSXIXa9pr4Qes/QDu1/KoYfIbTQMx/m49SWNusqghhm
Gmg6p+BoON980gMYAcSQpQgmOhdDI2XRoj/sMG5XvJk95/SWfdnycPR356KVLRfPDbVXwnNRJ4GA
oP4mafhtQ6qIuTwd3fxDkpEFqs5Sp9lJ0LKZu/SgqB+XCytGekahZy3LWbiK9QtkqeUBD2uCKc3x
tXuNYr6e+M2uNklBBQqf9quBxyGJ4PNLq+gnltGMobSfGt3ihMHEB3a9dgWSDyPbHmfmPulGDCGy
LVy9mYtWNyu9mnSY0aB5I6iTyegRYw3bGIJNfRCq1V8mEY0AEN9cc3Xc6GWBbDhJfWeiqVqRvIQF
1PIS42D7VUbrl1Yp3MElK/ucnt0fgXVwzSjB/OcMaXBOSC5bPxn4WR/faK1UnK1BNjtoLUQg/A3E
yRkFiNEeOa4ffrr935BbJSyRD4ZySm3PjsZ6/tVWrCaC4SK5YaSV0F/bDA/SLAik8gDeuyYibMM7
PJUQGSfbQbNLYut+Hkb7v3fheXS+UlMgv2QupFfSfM0u+zFJ/DNKDPaPVbdLF9f/oujLSZB0oorM
WgxN5gd8TVOorbC1hxIn88ZAgXlZiAwVgwpVbrY/PGbVWheuFJU9bxnMS9v/+nUpSGaOXr1XkkQl
+7qpxZUi9sBVh+g5CBK3xvM5+z4b4k4FoZs4evTdI4IK7vLugscZPX/+y0o4N/NDRyySjyzzq5xW
IsH+tqQxGOi1GwmBM6VCNtsXk2nSDRitkEmPQfTdrDQobqol1WgFDwp936guAq/siCo7Wue3PXt9
qEjg/4UpYBT32n+6nVh0UHbrYyY/zkndYkvJchXpAtCZpxl4gW/AzV3yeFQnkeoysbGWT9aG14sJ
h8Af9OqPROUIZTH8rbzfqILyGP1ZR/XcPI/Fs2MCt8lvjZEirBYptAJQyGHMa95YROlOz+4NisFp
mtkK9hXFs38Zo6Vl1JqL+XVdsGU5WqYF4Qao5a25Pspqo7Ap9Zi2qf/enxsNb39dgL8qXvbNbD2h
Pncu0ZVbKE3XjhkCgegj5LYeHX+P8LUDH5B0FfOkOAYn9LCzfA37cV6PxP1ksVV60gTURTuRAtZT
VTtWYBxe0b4JFSKI7yff9TntlB4a+ANb03KgvOJ/m0aV1VQQUflXiQZG13m9BK/BAbaGp5RZnCYm
DlsDXeGZxXoJDWHp5xPXvm+pCwZaBU0Dd8cMCUoatT0hflWDq6raG+/qAUNi30gpfzTS8mJzu4SD
5lj9dvimQRsVeMgU4CvBp+F04WDIcmRqqulIs2nXNX3L5qtWkXyaZB+AHK+6N3Uzia7aLXwGF3Qw
o8OCMSZfMg0E3HHdt2aLfc5kEVG+8427vdGyMQgHlzeefRZNFc4y4Q6GIWQ4Ktm/jD49F+E9KKXN
cwi3U9lTsS0G52qeZlSyqjrVy4VFyFtM0wsfFlEB9sxLCILophOSZdwWlwTcgIGUnmzswoIClNBl
XqsNud8OttLCl2xNjGRsucPm8GG3HsmBZcJXCSUiPuNuw3hsxlVVgUC9PXL+Zroqv5M8J06FitAr
uPaqA+HObFeM4JtTHFxKj+vKVAxjSQ+VowKqFVzaJD8uTzibfSEuHXxETLAznUKf11xbtREsLN+b
0hnpUMRnQPSIM286D5dUZkM5coL0psUQCK/SatKyuTmtRaBgNx3qUnz3tmajkS7JI7n7KF+u1Oie
0Ui/kJh/mZjWRt4J8hKsBfqv1cjHCQOM8IxNSRTNVFEWAeQtkUb6oPgurwUsUCuCbxRJe8w0/dAz
nAU6fFg8KMGiOrgEYmypTpNF98DhR3J/LSzTWJ8Y0WJqTa5yUfw1oGZkh69TG4qYwkESG22b3UbW
EfiLLgDcG24BNYyR6Z+ZBhQCEH59CkTmYQj42CzglU+lCeS5KSKq1E40JiCsFxD2H+mh3R9Mu/8U
NZ+hxhKdvho9kM9ewPnz7gJMDan8lh4PNq8yjPBh+99f2nwaoY3I9eor311LFUiX1XhQRlfPOyFB
hVXHoI1kyrunrW6Zg8CyH39YhtwmjjzLZ+10PlY6CJHBRHQw31WktH4fZu6NFCWLx7CYqeP827tN
suXVCZRIESSd951Vjp+0+e4E+3X2pi448wvuLOjX3xDwnXsHmK6cPP3ZJ7d+knXcNB5g2PbijmOC
Blsgg4qii8P8gQLNOBjcf0RusdJaRqh2wmQinkSH9CkEzPe5BHdVQRvoP6GH20HxCAVvuXsxZhIU
1dxlds88qPiY7wG+ILvv7NhicU5V3+6U9gQ/HYcpxrfZq85/Q49H8GuDoPWl8MhycorPPJBea+k8
MtgD5zEKWIB7p9c2W3mK2ZtSL6KKNtKQZq0YtSbP9yz7lry/Ck/6x1yPFu1ZUqjiV7wsNCOXToup
td8PxY5Rg4waXqArqH/gqFoGKgLqUH1hwb8WM1JdXGUaXsn8ks8B/BN31nwPNb99pxRxpwhini9N
4+V4D8KS6oAeFEXEl6J1COIXupgy9YMG8J28+6ur/Nl85/SO9APmof3Uh4EJszrLg7Xo9D9XOjdC
x6F2/c9ftCzwuiU/Hes9DKeTHBYonwSvCcSUD0ncPmPRoNclyDVXpB1FOPaPwlgSEYVTp3yHhlSE
nbLOLBgNMRbQF/mdwVNKIeXkwgTMdqbHGXQRG2KHMTo/Jgtv9P81VNCnSxDNGg20wlEnh8Qz/vky
S374xc9bbRLJOeFx6rMiTPFiScTqjemnsQIAkcQgYINBqxEEwNo6N0tcN1joEUUMfehmSbZ7mEyq
pQJt8lb6kB2PvS7bR9Sh4WsL8dpptLDmq6EZu5oRQvVmuimWLhlZuIE/LIRUUAJ6gSoafXLGqDOh
7Hidkx1rAr+PNEANsJMRKPuqY5IsCx3JjmflCdbn+8cCzw1+uJ6G+U/5ISoI8clq6lCyAHWwuxXb
tW6smVNsoZP8jCMtgf1iLPMpZ8TpmbKK4CfnTo5O6a0KcB36ixdogeRqXhLjE54yIZoXnLMGcnvX
x/7TJ0KuWO+DD4pWXLqhCod1QHIK0XI3hYHKWSHtdR859Oa9bkGgJAiYi8m5lE/RLzyO0WKDKFQl
EzvY4kkYPGJYgVJdlaCrXa6crMK6qzZuAJqXNdFqzMMhUL1i6G6d1iTWDgcrux2cL+M/zTpGVAUX
jgoRjTdpyqGtfLu8bQz9N19YP+fxT5gX0+YfwRYISXHoeuupbqwgYD1PuS7trw6MuLq427osOmhV
mV9hc2Nv0aC1ZhxQqw3NcW4ReQD4J/LIvV6l582LErDxWfPw5RaWbGr3npaZNW9hQWVWFDOvZ4bH
SqnETU6hsAhrsQrr4s9TR63hUOwEOwYEQLd2hCbX8/cXYIcc+wR/tBxdPPKaa0gdYsMK0OS5ddMx
UH10odyXQw40XvPHKO8NzvXLkA6/xF5k1kOf0JAQ1zalsbcHgLOSK7k8K7FqMbsPQDpo3Da7/So7
7mVPr6XAQD8scADFqk85LNMv33BdgMaroM1CyAlY77O0CguPAzPF+KzgX4OsxFFjoTW22Sm6mYej
4V+s34/CtfVMGspOgbKM15q136ufWe7aA9xWfM9I3Qz1BNbf5EwzelZv8qYLK8sVmMsnitTbUogC
F+H4fcSu/3R9a6iQehW1rz7nuYD8YLYEM2XI1vRMeSqZZYmUI8HBSm7nXF/cYkF5Gi0gySk5kCqB
M568nYJgoz5WQ8kzipRcIoLqQsOYTR6fFYTozjcWN3L13cmkkdZ1z0Nzx1VESi40c1VstuH/LJuM
kslUUXExj6RPAqc6bC2/LpCQrQQLNJRw4FZH5MwgCjNLrz59fCeiKvAp59fMXV3l305qEb60tLvi
tdJCa2xhWucPsnwJ9VLnV94LZjuz+FDAHdR5O9gyJGQuh9EKUawJYlmyBV/2s6SJk/zAxvFQ37Op
oC3ILw6WJAHGVA904Fgk4pYalEYrLMHAhe+ddBbj4u9XibzcTKeh8UJx8jGFuWt6VgCAotPZMm7X
sp1iIL9K4SIKuM9lytTZtFIhtkn3C2GCvL3yl+0sL0ETo8CEcdhTvbtvyGGhKv3WlZND14Jq4SKo
I1Nb20MZUk3/keYhnzeUXTtcOywp2Qaxmi5fNXXws1o59SNaka7n0kL4ehe7sKHpAjkehHy52K6D
+ACdn/yFYj7yECqoC7rOzl3Fk/y/6agORn4D88TWUHXHzylxRYAJgw1ulisedElIFO7hx/4VuCFb
fy8HyXSKKriD8CE/UVR28vdkicpkpH4pd85d6jk5eTZK5VV/ANnigpqhChABreCINqW0m7pIsufp
y9aPFCSZUTGQBZ8eSibFB6HLFQobnqd60ah1aONiHPjwNquB24seXthpNy1yljr3r5CuaRqBL1k6
54PaPp5yynXTT3OINPJ2pDKFtORE11ez/8anNx5+Is/a9TT8Bus+TUMXFEa9CsarWstuLM6XPQGo
HK+GPkeCTot15GKHEPgZaMWRzzdEKGR4IhOEpZqXaLPqO4Q8mhaywm+7Ptgr2/9vJGhNaSkkRsjC
I6JlgS9ANBMo5HCDOTThLfemkk8fg07k/Hipzbn7xciJBPJIyt6QjD8GNT4OTK7iSuG/i2hG/MM3
z+iWyaajZqwMWeNkVG7kEKp+WbFIxCINl471xCmN8kogDNe58UUIA8rC0GcPKAxj/U2SP49W/qqr
C6Atf5v5IOgwYVSHoT5RKlfzRkuTVAdqaecW7TWhSto43lIHZdItV2RtdT377HoA/rxPWOa8SG0N
RKADzaRHfDffPSZj6g9t4xVWJfV7QPY7I3VO8HHS/q9xzgK/QHE8esR7Wv/N/0f0SugXyr5ZveBb
c8+mC5rPeoMV28xjbl4kcRPdp5q+6lrjqZxbYSdAXPI/h2gzeETlvJyvsI58KxYOjMYWmrN6P1nw
ZYvdTM6A2RpN8RuqOk5F8hr3+wXQcU+5DiWNfet6RKEISYPNnMrBgG7hHcnR76wcVWDW+iPcGf7B
r1Yf3FjqbDTIKQedQ3GrNcGUsOu/rEVUN3ofG+Cl0xzyfEnpRaCjGdCefmF0n/IKE7Y6puMhdUSj
i7ZaCcEBDyB/c7k1nK/Q5sDHkehJDtTsRJCXmjOIHU4WmT39TgX8ayg2gTxaBFw+eBt09ZrtK+ou
kSGKzQkZowKMl98kNu0MnZOqxtQf+RbPf00SvxpiZikXDO08ddKdXzNlL8dN6Z1vp6p0loE15Qiz
KAOzoj7XqtLh3uoHizFMLrO0k6BY4CPwwf6Ou7fSa7EluTcPAY5d4mxwIac2PbaenGdabjb8m0A3
SZmNKMPrJ2viKmlq5Zj3ymVm7W36I/XLNOX18P2gOwAFZDkphB8q041NI9klM+vF+ZyXlMyohnSx
8f4SIfM3C6z8OvVob76zILJPscs8XgIhTt5WIWXjjSRnaLHzW+aQJ4Fo4cs2757cZIOhjEgVJyiS
tJb33N834kkmetWjvwP2ydrDzhjVBCtuwX5u+73kXo7QZFa+UQ4ThSjCoCdyEYBOfy+qAOlfIFjk
vrccU7gIU/61RTqoZlbe9QiNy6PhMbgikS3X/aYaY0bnY0kb1WDJz3+PyOKAiXGu+E3FfOuDYNGk
isQc53FHRMYFoH0wVN1RK+GbDyi44qtEvsXFSBiMdHTy2Am6MZy9B0Wj87vz4dmHxMWb/+jpJ6sN
Y8IT/d5g+swnorA+i1a9Jz3BGE4scT93VnsOr2O32lYBNs7xqz37juY7nHYYiuheN1HaWkcr+UHh
WsnVQKaaQhV2fxGl3p3oHzM/wF5zAl4xNx9Qr3e1biOuP5N2a4/puFgE/0Hml1f2htbZwTx7R4EI
MNUnTbho5g6HcGp+xz0bGrER6ZW/bPPLzbSVPm/CF/Bh926aFhB6R+vKY5PbWAfYLImBVuKhZvWZ
fgzI2tE4j17qqWTz047I4vOz7Cf459DLS/OZP+8oS3SxucAw5qYaCjcn4W7d2kD2V09N6Xwnhdxs
ty1jYnuRIR6JWPTzLqhv2r55QTvMiiaL8N4cwvk8rNxxxdBvUQ2dE2EkeLrqvSF+32NeYGBaXVqk
BXhtB9Z3Qo2kZgUDO5hNUtgW1z8zhHe3RkAJmhVvxH+/DiPXXUF8IBoARA9RC+SEhQyzShx3P7eI
gvF1CdlJElm0kfSuwFoEnzr/IOQP64fRSZcZz4qaS7ZJpE5IDl8zav7y/hkL6nO3NsUk6WrDBuWg
UCEdE7H6wz0eD50UXln/uprlrVE9gVj2wuBh8Lj5KSHcz8X2FqZNZ355gCu+KSbPI33aD/L+RqOK
uqXogXecdo1i6SumXLEDXJsl62Hb3y6ixkR/HPd1wYT0ebSU+Mydxq0Ysy23N5jFHoq0LlFKYNuH
YtGb7niC58I4p6qi2HYRQkCdjONG6Aa2OoCJEtrelhcff39CMkNs8o7rN7JLCqtevIy0Q0gLrWsw
xOzbXTTYSMWTzMEbhrMT2ZAVOtwwIR+17l/hEzzVEeikriZ6b0H7nzW18zaFRC5ms3xE1IU3YGSj
hxja6jKVq1XdPdyMN1E7gX/6XEVTUjqMyBajZRrYP7jxHxdALwzoiOdYqj+KHUn+S++1Q5b3AGcu
fCJejux17bB00UYzWTszsEJj7hzsMUGfYHAniKdLHdlMKT0FMux/FiHTRJ6A1l8FbTHT+6sJEvsJ
/qII6maWueMfCJvsumtpzDpp1M2cXV98zID/pieZ3mreHP49jG/8p1izkBLhlohbhKtNQc6ysqP+
sJiWVWwtB2s0QHMsHHL77D8z9XSk4hjMyaxvo2dKmgpsCdVCiv8rXZlpeJEvQOLEmvrKq9VIVjAj
2MOOMcFIz+dq8pLjiDz5S7dWvftbWXq8G+zVdaquH+OhAXWhEqW4tQJWmiluJ2+HoYC5/yyl+5bn
ksFnqwKiv+RLzyjL751lpI7MSh1U2dLOZDF2B8qXNDr17ilCtrJFYhIL6aKWPL6BfW+2P1nxtm42
ADiVEW01dGlJl7CM2dT7Uc/3uH/Oqu1lJ192DcVL/c0uBaUb+WI6SBSg0kiO077F+F8e9IE2YHTf
26CpfR9SnPPEpysJKHuTgmSoUS0HzjIEe6mN1nuBU8UCo3k/5Enjqj7W573rpIut765hMMSI+H5P
Dm6D2zfeW6oKvthu1Q5Qm7c37XjASoxOkkefdYT6wbr3ndM6KcG0akxTQUHHsfDmxOay/odK5nDH
DnLV7CVDedBCwGuAzx7j3g3JEiEC+UcRE9dIn35tDh3/86ZTV/gNFwVRt5sLG9NdqS4JFzG9USGJ
EmtEToWMebRhygrby7Ri0wjaKTso/vt0HqD2GTrZoBloCvoo3xZ4X25DBi9RK7wtzu4BPZQLvGb2
bRgqWPhmk9HMTifFfMp8xZUQwAXuxek0TWvjODq3Xnc/1BhelEBsOwxn5l97+V/F6lRsChaDNvzG
GqIvhjiHgl4mflhD9WAcS/30B4Oeb6lFwGpVofbyjk9QYLJhqe54AIROLw6Yj2F2uzvolonObq0Z
sQKC2r9atLU55o9T/1eMsgTkQsDR16yW0jYjbC8ZZ/j8cGw4VizAV80kgjaWuOW6hM1YzpK7eAFF
aLQvoRtfPUslhiTOTGkE6pklFf9j7G8UWD4zsIx1j+1ok3xru1VLaCOCz7TsptZRcLnZiGNKPZ+L
LPfPPC2mRhJaBkbBB9uaQqMFLA8cCj26GPBB/32+PEm5UtF0WgofuY1NER6GJ4NRzq4hm9zO9tdt
Z2NT2QeiH3Y3+omL63nGWaHYNdB9m9x5i1K7t2x7GPGsr+4gZUM/rWC7ypUaBMjDvCdvHxB/LKM8
bNqp2fZHN7TMPSMRYoEaBSL6lJp1nZWROwVp0nRU0OFe+00TKKVl2zc2JuS81/1PVQVdP+gqe5kG
zXLG0rnXU7yKMGzRmt2rNQq98xie5UfP4SF3rsaMtzDGlBGYHk+KVES/1slp6AeUgedZb7zDkm6i
M1Ox2y3F0YM1C2QVkEYebJyAR03bmgbHYBv/MhpDgGUiiRFfLA9ursaJiBdS4uEZ1jU7/hF1clvi
fLJXXsrBJa/NMxuqmeIWVdxxQO4SdJI6nfndnPdE9Z+lpLsYJaZF6Kq0VpDplHWX8ngzn0f5Oh25
UR9lQUCh6qntU/b6j6XGNk0H3G5eDk50Zu/xRLWakWKSfMd9Q+Qu2aAdiyYyRqaoViRCURnHagbU
vCqFIuNEJ42IQNReuEGaDoCqPLPAFRZqx5A+1zuGmgb2Z82Y7o+kltCD8MJEgYXyA+gopkZC/LMm
IY0Iu1XNTk6eQ4RAbGZk4fP6mGYAfHwzDtJbpVNTGE7mbfxSeKE31+x336z0jn8eH//+gW7mNG7Z
SyMU4OpFZxqwH39Z8urbeHabwBVUi58Jm9dNBQxUC10TNeH5HuVVhDIcqass5JUbo7ZTtsroxxk4
/R/RAC1ml1b0UjqOhl3Hro13+1cB6pCgF1oM6qvDpW41fgMrOJV4KnhOKO+5fiIHiu5C846j8XVS
6lFgNWzv7kasY+btpICrnwLDk2d4T6580BSXWiuZDi2BFaDPuaRU499hUWFOl6QPEMr1O+v+6M5z
eudIqRx+ih5X8BGT2fZAISLqu/W59oDoX7ybzjfJkcNOuW90AmS53qsCoGlIjUILVrcywi6wjDCU
siFUCogxMFI0rwV9nyHNeup4fUkz6+sm2ztvLpNyWBWvuQQdm/08CcKS3i5aWkOp0s/RFfT5eDZi
b8UdSHkj4ws/ObptUqZn/hbAP2KoNzOG3xLI1yT17fCfFSwNz8WlRT92YYRiRp7lUbqsBOWu1bDH
Q530rejvZp7g3gsYnPq4GvG95mdtQtsJoXJSc/daV6SGw/kOlRknBNPwXqcyIBsVpfgOH+jcwrDh
m4HdEn0fh7c+VPaHP6SkbVCQ/EOnTtaEy/i0rkvPaMf3SaR8gPyVxz0Up2VseMa0rwHePInq0OW9
cO4/XE0qEpeTBLkF0n/1/zNrx41r7Zi56Umt6zMtds4Slavxn1TtM+omjUCRPseF+nIwhGyyBZTt
mtfSEUyKjoInvM49FWkZRoZenxVd4TdiJQ3b8KaqAABRNYkYFsNB9JVJU9UV3kX12t5z/ZDkVag+
1eN9RESulaPaoGvCgyn1eHRwYwNfU3WyvFDq4j2SDLvATUmIp7f2CaRLDxTuyp39A7VjHv09FPSv
gQWSGxNMewC40fdv3u03pKlmk8+iZRvdIbi3i9d/lWP17/PyZDBIGQ7KMwNvIZIyqeSYqUuMcqk/
q/QAGI09us1KnPb7FY6JjCX0rOmuC+SWUb4wEei+Or9In2xxm+DqYX3WkfLA55xzDICfUxFGXIaS
byp9ezvaAoOPBua4ARu5MPgXwFvjWYGekTM+qcmm1QaAaGUyVFCL0kipl3yvsBrdv0Pb0umQOKdo
M2ojU5RScM+Wn165hl5DY7anssFCixUpTBd5QNEJdBrKTkPzHr5evMrj7HGwCqotIrbvy8FgOpkN
frONNBozwT2/obdqIDToNPung/FJ2PAn6abrb6yfgD9GxgN0jSaSo6qK9hNavpdqX29cJoYUvy3S
sTMluDO0N+od9rxzEUA4Hb0Sr9Kh43f12HAKzA9vxtXLhzfM8aKloVZ6dWsNJNpBDJmcVZiRrttS
g04LJJ+eco3MIxCNEO8zOU0HzjNgkPeuPPuRmgPYI0YS+02tlLbTpZMfI58zyuT9PUm+LedVrTmw
ovflo5Xs++qe6yzukeyxObc5/Di7a6J7QRDJFlz0T0wLpBsX0OZqY0fWU3g2TB/VUvO8nggCaOSP
sdvZVqvSmDRQw1V8YJTfi/w0hNNHccZafpT91j/GAeWrQmd5DoM8ElPLFwevXW8GI4cM39+HyTsj
iYwPIaGGL/mMemG13D9HhOwzyx7+UrQ6JxZqXSfJs5V6303szqJLGW03JYA7C7esj39fo0a85X/s
3xyLFCaF4hf8A+VHqKkHwRD2fv/8KyZsu3n5d2D0d/zzWosEKHtTSLoIl8+OISdZMZeKDdsSvU9I
AEAiM8JHqt6ZTVWSmQhych3uQ57vGSYLBkszvwYlqYHkTDD03GTAnIEKsL79bXjx7nNviz7OYVG1
6ZmY8I15Hy6YZgn6uQQYEZ517lsqLgzc5n1tOmWTL/UW6RYt33raBAHZKuzIPipUchVYNviSThDF
UKqBJq5tsdSMIlWf7yzhBFDN+RVpNgxMsKXlTNzSM3lIkyi096UsUneMRkjSgzfL5/v8kA/ivBw1
5qm7iWNy8rotyS3iKvMlXwlaheBPNMt3YnYhpQCT0ZEm1b2JOMwHsgdTGVsvznY5zFAMvXSJ41Sz
4tBrd5RbUNR7FlxvHc9yhV2St2Zj5IfDXdxVYSHIdjH27hvbb13jXmByPkT0Obg+xtscIij+PnE5
qlXhfdK1brysv2uZtJjBvjpqbh1yZ2ZjsBQgZaLu/8nsdF9+QWOAqgN+EMiibVD/GGRFMXmfVTNl
VD3tEKitnWj9TpEWGZTSNPY5FMjKDiRfQE7k6fx11UjTfBfJwkqByn0W3BtCK9VNbTuLKOehip5p
xfurUGBEvips1jf3sjPVVjQGcEeHNnQeElniBeycrHvj2sm3Yuuqzq2yPEr312lHmas6yxmpstBv
6jE813Aagr9fJQJOhT+KG04ZHJ/E7AUs2sW/+zJT1+PHUBsNYzp27k6y3toQ9/QNtIbLicXPRvIb
XCwYaWd/KHSAL7asvb4ImcFmCL/vnXRJiRbUkfWb+P7HBMbqQfGBUIM5GVEl7VZIFeJmdsN6Zxki
B18M43jULKw9J4JNA01e6zeSjdVp82xnlYiy2EnfoDjeDo1BU2P/IUv9CCvk6YIAsTVUx8mayB8h
JkcXPF/gZqR2zBEpDmML+VddOz23Zw0ZNPsytqYfEGo9bD++U3ED8CsQIAj4HPtKDHd15kY/WtU5
2er9Yq5gg+XY+QcZHTKYZveY0G1UXiQrVUVD/3350j2PysmemyCO8bdfi4nKtfaTry2LxUKOEJ6i
kLZmzzqJ9T1GVPSPMvzmUxQG+jZVERT3o4GYsLwbranuSuyfOwZuEbZJSUvzf2/qAYcJv2QT57+Z
7JHuugwah38fDs9K0LI/dOY2WL2MFbc97OW67PtKhM35VNBIWsphvqZit1yRVBMQhXQRJVNUCX+Y
cZVy+96mHRHkDyhSFsrW2O3eXrkjUxT2UrN1Gs+1UWEnROzds2pVVoltHZ/dTm2CF2NBTLQDJP9t
v0HhLsImU+kqKvPbQJBQLNz0QS8PUDAyL9K8RbCiYWGzoUYKswN8BA4XFaIGsLlZjQBnLITPCEMr
YqgfBHUv/1nfkllzb/J5Dg+9J7a63UE7r9STrmdC+heu2vq/RY87nfvCrxytYkGSAWGb/iaV26Gi
vcEPfDGB256TOTducNpM4lrE7UCtsV8fpXZmUc0C8xYO9cT80c5M6B/ygLa80uhdbrB2/uxYgtha
7QvWXkpVUiNhz1PKc0b2rqU0FswLbNo4YJnOOnYCe+exgAe8bRFoOD87UovPlPjzRfxecPGooszf
jZRNGub/j04VVjK9guOfktwtZFJkt/KJfVGTCqFsKLbsYluGJhEM85bY/LgI9bn5JjeCsd0QV2Ct
VF2xmRNgLB+kaLVm9pFdgmKZ/ghRSG38WdnZaF0bWf815ri8rl6lvLftPEo56th5AiQw0dflTxSo
ZOWdbxBmTISshSwmK1uN39nqxIkeYmK0aEPJnBBI4xe0sI1I8B4rMs1Fte4nvUMufreWKgFlg1+n
Z4h/1JmuD1HoLkywXg4/c/LxV9hGW+AzkiH8/orwGqsAn9HxO2XXrDtr1LIo8mlg1ZUG9EKbewF7
lt430m01jSsQFyqV1MweVD63+T5pXQlb8FoVJkXvq1y39uGxSZ9Lv7evTHPlW+PnwyhMOcCu6RSp
DZG5StsoQMSArMgQbfSasDrxcgr7xkzWCbWO9MuOvwnLhq0LigcowRfO+mRQw4A49qvUWFjVYCZ1
WgO0BSWIKAn0bOx1qML7zOJGSSrmW8IK73tAAwGis5TthArOljrtSOer0R/v2EdLiqQI3z4WUy+t
2k54i9ZaUOtsT3uEU/Y4OAyzNJFjJH28ncYQYf3WpevDzwH0/wfs77J1m62iclI19j01RGKntssU
GgzcXN0UC9hbWAnTLjHBD9AiGDdf8VZ/1f5/kkvs2zRev3aHUXC0K64MNbGyUz8xFCY8u3S34cE+
S5R48f+TnSQn7G4TZN82gB16P3/h/n+aRr9lE3VWra5J9neSc+oDL+fvgtWhZ+xYlU5/Kngt8qyF
+DFYMsxDKCVlObGdRdszG7eMxLP9Dwm3EXsl204DHpEwIZ7Ht2Akf/hdj2+os4gATLGbD/sWnlrN
zFgn6tBxcobHfGtAKDJg5O7st5nbpSkQuxckANVkCmgIeMU3CawaLaWY1paqqcoOeZDZV/ywLBun
hl4zfGPRm1XmBOROZMr0bNpdm0sJZF9JA7LnhO6J6Vs7Kv6LUadXEHg890xIlgF4ciNFlyMX6fUV
zclSdNM8Ih1FrzMhg1GKhQb9nrcHV1DRYkj+xuPMgBcdevrjQ387dnwgQA/ddfOCZnR8h4xj78Or
Utq3LxHF0lq6JFbpvLyBentksMugLSoUIwlTYDB2Qh6CS/gU+O3YlfUBrLPu5Ct+ByGpUzwmz3sK
CLP47f81ht64hLN/M3cWj+oA8svDCWfi2PkY/hzcR4Trd2YYe2pQKy3SeEWEi9JC6+DSStjw4ijl
0tb6AeOo2S/k9xQo8GPlDqPIThUCD1sLjDhvhxwazDSC7NeHlCAOdQ4RKmQ3Is6flvZauAqCxX+X
UKo3nP5ADGisJMWpzs+oXn3y/Kpl1UttGFuyrNYeiAbLKCZc+VnrK67iOQ2ZX08HsA+dTW3Mmv5n
e6UuIoJiDPupNa1JQPN9NGT3dU9Wr2S8C51I5JT0WKSNujG1lfE4pG23YP02RrYRiXu0tHPAlvjJ
7WpnusXJW4GGI1jccx0Q/Ukc6iFAWYhV2l9cA4OrFoGWnkjgisf22iCJdDTG4ScvsyNQ23QhFbRt
A1+qAN7EqH82yRowfPLVzMHntQrBWYmWGfjAuO4V/+eFv9HYW8EepGOGdx+j8Dsn/aqO0SwkMoJb
L1RYmW9Wu6OKKEyUPXQuSL20nmNOaMPinNKvxUMtTLFABtArTu6ReN0h/H9SDi9hjz8pJOyw2qwX
2cmw/pQ9XuHV6VkRxPr5BgagHG2VMqkRuINgiHpiFdcGU9cdxwOkl9U3/YM5xH1xuGFETxoKC3vk
IIlhf4dQRGsIeouGUaxDAv7nhaAiXFMkXuSvdB6VxQOV5rMacLPzeGxtJAKBP69zHclgkJijIfPD
8W36y/VzBpmsbFuVJmA/g3hoT5Av8tSWNlckGUa7loLsrTn54/zYmu1Z6t6pVR9KpJmrcRQnCdx8
xubSla/VNXySPS3RC/9reZCbUc/PxqPxaPLY8KbdYSjXoHunKM3wFbvDFgR5ofJqL5lpvvHsnjst
tsVgWGlup+AeY188zl7DQ8LJQRg35Mk3bCJyMyhmRkFzbOuFQyd/lxV+YUVZ1pnyUzffhNg8+ZQD
U14lndUK1xwE/QvCc2UjqjJSvCBKDzDLZRBaDX6MXqbRSjSb5UdpWOxcc+I/X2vWoZqSSDEOZTek
TSUqXyXaDhBvN5YzFojXHNkBz/w5k9iSWzkTLlZ7DY3JBpyIOxSVbm8lcAYaoHA6XdmEI/VvZ8m5
AQRraL2bGpHssvuJ5+5x0I07yiivFX/EaJ8BZShQfWc2WmEXYNgiYycTq3/DYa55WAdCdFOPijQH
ouNlVdwjvFRDjzcLadzF1DeKbUoiwSSvYQxGd3kMpOjYLmNMclZ8nU18WUGVnHXuRxHQmFlScPsv
4+qUCMro4m2UUh4J8UhmUYIom5vPKrzchVDKVRdEO33dFfk5/wzEwQzi3YbKGEDzESxpIjA1T0Tu
Lwh9PHAnSig28ibdlUgffOlgOQ9uPUyjhJny09/I1TIXMamBw7eAr1zaSxOnSzzuLfAreGtzClyP
376jnQIoT4lu+TFcDhLlY1b6jEO990fvXp8JoMdeQrbmk+BlsFxyC+VwZhSXdBm+FCsAuDcN2Tom
Y9KqquGzUP8NsB4m3qGuTHENlddb53oM95BVqf1u1Rlu+Q+pG2brUT/T38cw38SFHCbiO8n6QILT
Cg/9ydzkeNoYEkNvX41XCAyoJGwu+BrDbXWFwUdk1B1/7eurKBz/bhfrtZDc1Z6wkVKu5QnQjiH3
S4T3vPa66aBnSL0w2IBaz09ITErDpm2t4q0on7yzTjHeLiZAg2NKpT9JQ5YP2hSQvgNXfZvfbB15
B9I4uUu6q0JYslMNPZqs7VFrhVrzTJX0FOdTouJb6QaVjgsb6aMDJncXr8E3nFlHVcJD6w6WxcZs
Hh5MdTV7u6VBpMvIX9Sd8/Xry/rMJpFEuckgetZEkzD2vOYpGos7duM4/3ZOx2H/mr0kwDiESYq7
4B9LJjjPlMner+rjmhE2ecQCzM1QLXn8xirySyJS546cRDqkNqElJuGDmZ10QAlQ/yQn/Y7eV1Fm
/J63Wdsp/KlZQ5OHmF1ZfSh2TUFPXV9usXylsMpFCvG2VCwZPoGx2T/U7rcV9QT3slteOPACsYeO
OFjmrBSyS9YBRuwowq8nWrbRGRvqSXBwXi1eQoHUpDATH1IOc9kjy2i8MbVwqUHWPVb4wR4aBAHS
OJDUzUvWJuLWDKOQ9QgvCBKyjgz6Pm7o9gx0W7GgjNqOfwBzIoizdnZ5UnQuBKfPfPfn4XNXMRgG
KUlk9NxMadvAIVFYHjyOe3QocoJ0aON0uAABnsfC2wjykljbnwlyjC5smojX2WFHtZUqE850p/ye
OUeZbfV9Bl1OsNoDLY5JR4Jr3BVs5F+yf0X9uBm48kOeJCLiJgir+L80Fw4mm9OmadhEQAeKw4oY
HPxz0dd40pf9Stku8noMfCmns5d1XvovQnkULh6Wk8/Xy1wgU7QeKk/OcmqIKLFCqnOEsRLdbPBi
xLGwt05a15BQwH0gbqMSkqmN0LCWCcMEWXxsCp8kFXkDb2x2rLrcxvD96R2fmXqEoPpfmxrbkUVo
5NUtal3wdsCgrefTzRdg+kRrqzvEzaLX7txcnWlPD2qyJNH2qtcqZLMUDBUZDXyG1AH9hkVu+mqd
CkmI/wqIeMVh+vQSnrVcaR1qVCppPICbWRrsjSU/745J+ToqJr0tfpJ2w2uS59ySPrWtxDCqIMxc
chlNNfqHzJHuCjScm84WDwcwxPC4hBqVaI3Nf7x7JjG4Sma3jyPxH/i3fkqWm0Vm68KqvcGsdfCn
LtVPHSTihD0xoEmLAxAugXXjxPe3RM1panSMpCHpV7/KEgY93sYW5uCneuYYGpXhK/rG/aPiN4BZ
WeJTR6yJGlOq4fcyLmaeDXCHTZsquXgyU/XAGUN/hdCJrbN+EycyoimuoGPvji6poa9aali5Lz/d
+OHT8MPJ2M8FBVMDCXC3kBn6yzmsbW7FswiqC1UANED9BR+7EZ189CN+OdkawYZ8KVEIWooGg4VS
OoqKdt+HYWOGhvzu1jeWkarPCxJEb6Num39q2+JXbtlRN5lQM6S1Qan19W2SzAJzWt8+zQsYWgc2
8D1IRSHLoTsiXrN/W2RtfDai/ZQj37vvuf+Y8INaoxbZoKTkBS8q4Qy6jTnT9Z+CIh35Hw5iObp3
YGAJP7sNdQdiXwrLbY9PPPrBk9lyZsgWHJrG7HQU8TGqBx5aqKOqJPwaSx5bfp3t8AHJVnllzgkZ
nT9hHw5VEQgZslSmCo8ZP1eG2gUeewxHWwqfmzZyhyuV3SQjdDa4iqvopHJRo8QpcuE7RgcVgblV
4iAJjdzbOWOTObyS6ppDvumVRtDWeRornO6oXIkhyHPWfKM/aaBEWgQX+OS12tmoGvTTVCkZlc6d
uqPMPsxEFg51hs3uWu/kIik51UQCDv1x1P4oCLGDgu+XUknl/wuWNn6q03/i1hFyZ1WozDPXij3s
rXuha8VwwYwCN1r8hEx7CTD3L94j3MAWX42mGFJGOb/JFOikRsFMdDadr7jdTNzfgNLFBw9ny5BS
c+Q3Mti8zpws+herCq4Q2PHsSBkuONKUDP05DbtPM13zU+OW+y9Mx7QFufwYXpo3DZR9v0tTg0pB
eAnSNme3uTGCtNPeB55oOrPQ4cwjiMZJh1GK/+w+xdh9znEo2xyRnXtgfVFNNmaxwFa0RMyAa6nC
Hn/H9T4nCQX6f4YXDQt4CJijrxgNY73rJrvOtBNGA+O2xsM4xcaGyh6s2wC9nPcAlXbJrjWiaBZm
Qb5O/l/fmtXLlO6jNIv91u6evP0QIrjFwbjzq5WGdmGRUi3eBCOie1ywYcZkEyyzi+umnU1OJ1DM
7daknhx2Nq4b17akcDpJXHV8N6sE5D9PkFI9/uzd/A+EichDoZiFswmCOC6F2pkY+1PmmhCjmdeT
W2zlPaLZDMS3HkZgkWRTR2Dqo7zicm8MV7BZ/9sBcnGt74fUgT6SjU4pNLe1QyDRcQ2GTIwmaMlD
b1vziACGETlRiSRwFvOe+yTvKkuroBfqFWoR7IC3WCcqdFUvZC6K/3oJcWyxCHBKm7aBEow90W79
PRv2jKxzLnKIpcC77A5B840cqComtclitV8sftxxjVkKqA76a39kBnpIDjrpKwJ6UEHezUiMgOZN
3KSN+XeGyQQRiLAEUYqgfij0vHN4OLa+LemM8GWkgnDBO5pavxziR7AqrNLAxQomUXCGndIa2W4Z
C6OyuVz0Drc6Hlt425tgEYR6jNWa8lCHgbx5o5ZRJc+Gt6WQrgu3BnpMgk0pSPLCAnkLXfwpoIRw
D8VzetiiDKkuvuxAo8+yzITf4P7YPbBX+TR5YFKKfC/oeXa2XWhMtIDp/u4BlZ1/GWFzfVpun3Ok
1Eluwq1Rqo0npRQWtYu/5sQf7GQ0kzToueoGU4+ZfBqtelh0LdPhFFyLhYAO5aOVbZIg4AYVj/IW
ikMiK0qvW3RFTENxsLwtuuZPzJPQbaZbU9cXVCsuOPv0fKFVr9Fk55GyERJAAs/bGSWn0m0sUEHj
XjLOStkvr2vcBfm9Jm+A+o8F9scCjsJENDirxUAWyY+1JtAjnY62oXT/QZuL1oo/HTJctwQ2FxhB
BlfSvNVHU17V/hv4D+49wx7vZve1oz3LCHAj161qM7VJzSA8k9FOn/Ck0qBM7YYI9nev2MBjx/ws
SjBfbVojrDwyS1l35rLblQy4BmYRiSHETQrQFHngFtikZzsNsCNAEB46FwR3w/nnq+EmHDqWUEL4
qJsgDDRs1jpDS6Ow+jkNtWedTH8BNSx8a4Y4W0dAWrJ03eFNuo38+Ter66vLAOjRMb/1rGL+mVdt
87KiVBvLvR1nKgaaaeEm9BBf8gcvnIOkikynQ2a/9v7z2DqVQpoHDArfpKfx1HbOH6OJXfTTMveP
DR6B7rVg97qQj9wlcp8jGbW9VCFMRJYf2qXJU51pSQckVKanlT0X4c2nMqS1tReAvhsy+ubiXt1z
9h3mfLjwElITR0nF/auhQ8IKFDYePV/MG2wxemZbRKBi4/ywzXBUVLQ5/aY2cYFQDLu5qgqdofY1
3Tr4tImmDP4C3VKU3G8BNwvYe+gzSvaPk94Wz3opVKfyjZeM9JrFFhN3gpKq9WFM4tKR2pIH5RG5
n1RLmL//RcqVpmQVOrip/l6T7EG8KGu5w/yN0yzh+DASMiaP9tyUlPk0gYaastldmtAWgbuMAXSX
aqV1Omm4yRjER27sKAB3FOLMz2iCw7odCAEyJotxt/wGYF7/sJpwcBfqP0pGv9sT7mwFLy4ixOZS
2JmYCCUfT/KkNGHpJ15Ym23fejk+KkBxt6Z2SKMLZ/JHem1hbsxpXFk5t0G7skA+h1dItkJJTQsz
cE33ycAK7go3TwQAs7oEQvteo9xeVJfi6a5HLGyqp2yhEynNkC9EDwUSEAjCk0juV1Y58waM/pE5
RdOEFJDsTtc7Fnvp1BwCoLpd1odGCrXiKTVYkstZCafyXD9hDNGBsawFJX2JovOhZSL/XRqRiGfG
ksE1rSkEIii5nSRYKM1M4Z46hAMDBWyaY+5YIYzor440bUIC0Fb84694EU1S/AxoCe1itWHA3BLB
4g0wCBZBuTK8B/+fyugMYUlLIkqMo67b+nyQzpuBOSszYDib6imm/HXdnlC87r1i/jHbGttF+gFK
mb/G7DolscWBwA5e0B8ecIxlQTOv5WMuv7S+phXMsP7MOQqoAlU7kpEaBc5AYnyHKwaAsbJjFlpe
7NMeABz94D6CbHd1TLmt0xkpwafUBWmHazTcpHzquizZk1jdRAxzGyKs27st8e3a6Zk3Kp7fbrZu
YdDM6B5VahjK/WvuUqk7buEB8DhUai0Tas7lpdB8Gxh7PMjDJePqdsEyf/NicdjHVwea8R0EgpiA
nzm/AnHT2oDSfpQAppM5HOvyIZgKtWb8Zv33AYk1aTxCIWL1aOGs2Y4e6Bm8nWsjHsUApZCTm8aH
TFbK0U1csHPJ2aCYa+1FEFUgIcaQevIwegPNnf4aOdaDfsLErB5buMOjk2XJxa6LWQ9N8IH+aEBQ
6VGfLOA4xxi76maW2THYS+hupDLWw97uj2dVrMzYic+4uB0G39EvUoxhRTrwBw+4+p/VK46ZFBS4
SIddADm1JXd/UNp/5Lg2jnBpvGZcah+GhnELxwbDHuesZ1bmnXIckTLkQRCFWHkwlVeoxWGPWU4B
NDmOzQTDZH7S9e0bY6/5mxgsbn0Wr8uydw7F64pcLbYu/4guXFKQpGbde7kVmSaOOjexTyCuoEYU
CS9y0O1/mdJk9ZM5BoiXYxKcB70wrvblwnXuzR+KjYt773NBrlLmDa5pyvXqhLThJ0Qx5axRvu6d
mLFe+Kz8EtimCw79Rt1tffFQeGsjSrLKRTzlSdfnpjEHw1ZFDwo8xfCdSwbdq+Iq591kufw3uH/8
uMDxfAJteGfTXFv3UqBP/v51e0Ck6+AOw7tUG/WdPN8tHhl6CxhFEK8eBluNK6zJk3a724oat7go
ehjlN0Xq6uTcqq4oS50nH9JcfkdRiajSMey5FBKCCR9oEFAnK9iopZgTyJxSSNeVCBLuczfEg6k/
CgFKea8NFqWyPPaVRdbGJtg1+ygVggnLoFwf66V37v6sf9zgoYWp3pOjEV5XwcITv+uVpLvkIDc5
nMu7yoGRLxNTfZoP7KMB2q0kTmgkTBLvbBuubM05sstR+VDaVljLk4upbLsrYR3FQD+W3oJyrZPh
1cTEhcsGntcbRtUYKSo0WdrAvba652Ax61duDELGxvLDyjvPkeX3quYmDCwA0wdUexasip63R4EV
hybgjrtyci6NlPePExUM4u52fqDaRU4Xfqm1vR+uXvBOnjqYylNp7Q9vd4GdouyPlpYuPMUHOU68
T3ypisOP86HlD9prowCbvUjsRLCMP6b/vMooEouHXk21APDgz4d1FqxOW1JYpxDxVsJ6j3e2Wwbb
h2uV9Ua6tXWABn4cPWv3rF8mcBnyhKhG8UQVpRupzXJZycCWrPz5BZQ+Dpahb27CIcs7pWpDqp5w
Grg/N2vj2UHp0AMNeNEHeArR8/n2AiUe1NI0FDppQzLEtgWA3oeaM70BEBHygvDq3ZG391YyHJAj
AiZEumdEE4qmK1BxueblLZfRtT0acpfkngi5do1N2b0EtO8+Lty2kBbccDdz/aBFB2YUwSQ88AXv
cjvtYwvyaR5ZadJ5f/uxt8uu2GhWNM33f0GPWkhpw0qUexI7rz9HBEB/jVUnQayviUI9FIglrICY
64Xs+bS90etXc3KEbjklWH/pwsZ/nfzM7MnxJtitK3850fol3R/xBzo7+71zTm124UVhamastckF
YB/JmoR7LbZGSueayWeyyVyVa+TQJSz1o+Ik/pAZAyy8pK1YxZLCex67MxNRrRGDsZnPjEFcEfPW
VZ7HgoGkZ+hvhjzkrDv+ecBDXcqd1xo8+nyA4MLPqR8hqSEqR5ssFxgFbC4UvWmPynMvbmriB+dr
2cgiY583bwDO+EJGb1lYod7aXp2D9G2vnSQ8rEZBHnAeO4vQyfOraMJGwgvWpFIznVY/Hh3RR/zU
RxP7Jzye5zXnMF0JtYov+5jLS849Wi8jN2XUgJ96J7n/uYBQCOjoQqhncX7MocRgRrTqc/dX2TBx
4AO0uYnu0X28yVyvm9WCHv1qYUuznBKpVFgb/xvXc3DNvx+ARD2vZvT/gnQnykpKKPcYSxcLV8FQ
WItOIV7D91s3dMtJc1LUQAgzg6w0HQLF5fX0XK4MA/578w5Zi3yA2S5jRxS+PLcF4Z6X3D5Hmrt8
3Y6dsDU0O1RNu59wDfztnTTgQU6ZVI7wuZ+anB3fN3h9aa2qqR2sanjTvvCzl1LYeLTtaOqoJPFo
kh3IsBkVgV2JaWFHyKL5/eC8nqWGpiWcKEuVXZ5HjZMpyJaWuQSOZiAKQI7iHcAeeOezufdnLP6O
hW0fdKArhoULuvt/hCwJikH7GHUzcOFTZ3pb4bRSz1/LWIuwM8/g9hgldgJjo4H1ixy20BDp3ZSD
77KV2c62TNtBGuB4dSmK/qz6iDQhAzIeYtFhFswB9q75NtKDPsV5H7abU67tAzOsLmjS2K4YZbUr
Y7r3o/uLg0+CjQqr97VhyqsE22+QI5OhQPf7GP7Vmea8gufGt40T462wBiwZEP9+n3hgL1jCQKzO
SyXd3jTMihLfWb4Rf045bzfQhQwMAd9Vn2vwJ2hbFDx+RJaH8qHFBscawlUIXHeR9RwJ2FaI8iix
whDkyD6wwaZv3jSwuSMmCcA8NJ/JQV/VJ0op6C1bchEmsAef1J9lu6fI+u56X/XtN8fbYi99C1bk
NYAb3E5ytHNuLy055mPrxblsfhfYPtHJRj0SsOfxXEVYTYSUNluTbeNj3hknvFQpFXJHtGoA8mR1
JRBm6uvJ1V2nYr+g3MJ9vSZOuG15qoG3isIkowHSvUZk1ia3Ulnbvlo3hhAy0BQDFOObmGC+L8dV
hV+S4x2Y7ZXGbi5f2LGVBmMAD6Dvr2Hb34q9jNLWwAX5YfEYlibr88p3yvJE2bMq1kHlo6Ca+FHg
R+3t5YtxJXwW+xgF5p26g2TJ9eyZ+YziR9Y4niP+HmerU2D+g6DbeC7I35kb8HcG0OHOLtRDQrUC
gGXOHxypi19D2T+3gWzXJWmLi6oO71ofphpBxgAGGPt6HcxUKk4lRGLmIAEXizbSaKUd6p1vqS6S
RbMwiRzzh70n9BaImSOpmEB0pBp5IuUVOkHi+H5ueq1B5jspAsxMtI9joanrWdbaM7/rw7/CwnLQ
8WOCm+WPQDbVzzRCnnihndnhG2v2jPQPBmfB/oW9JNWQxrOiNk4l/TQ1qa3eP5V++zJ9zek8nhNs
qN0WEYMgaWOuSdhXZNvy355AU1yG8u41omj2cddLaq1NzdPOtS/lIjqWhCrWaCQIL3E8KSVTQdtV
rQuaROzTLQP9fK0pdfzspYITpBia84ZpTlwoqENQ37iIcw4i3/5pZ0gdjzYE5K60KuzOQIjx3E8Y
MV2+rC8BoTh30BzulCwBatHTzmAt1WDsONoxvThaxER+XD1E44XqQttkwPg6gLjRcTAp9qhasAEK
9DfWQbqOvhl/wvgWCG43sW2lCLpCX8MhiUPnx2SVX4I58g+Qzi838wZO2b66Fy1Ime5zS34Ah9TY
rXwHVoj7Pv8DDY9w0zwb+90zo0F3fu+QyK9vBn/fw4VwbFsBCZbT3BxULSu7dqAVBxwIieLnMgTM
7zkH6prBIFvEwrvbBCgSpSvrM8O8M4Es71ovyMj/waSKqGt9HSOArkWY+JL7zuXC5b49gfFBSGMk
10cc/j2UfRREtbk22R+8LLwykONZrAGg6B0BoESrzG8rQQ524S0mZWQ0aptAgYSkUIccytXxYlkr
8+r0Is+wmQBLsBXRKuWUtNNrRPpvjy8MjWgJvbmpbjTJNPaTsX8wB/iVAkogicdvtp17bkTttlVb
C573BtHz/nAJ6qkWtYPNqU4KmdiLs7hHrDw/8utmVRBZyM4jpsuyAbsfQTSEZtYnMZP7rVaZkaJF
11RZhgMjQdk0rGYpYDZX8Aoygiu5p2HC5tRbbrVBKKc8ZuTboxTfkOiTxTiQj0KskBz3EyjyPknX
IAb2wtjKJF5dB6K02lqrUZITuAyOGIFK6Q0ZQMxPIUOtpaJ7DYKKJsVdIjG01e7EYIICMW6Xwxsj
OJu/WhCA5HJ5zrPAfgL/nXyWv3Z9wCgz1YBWpzKmo3SiUOIWC8HBWwgONU+vn/+DcV/atzPzdX/G
ibue89VkRLUfMDhLAvhuWU0J1Y8y7BbgEVPqZgiY1iOcTcd2G/8AoD3B0Jkd+pYMqRG46SLc3YwN
al6DBkOcXtqQLltuLP/Jm5jjdoTv1H2aS5TCPkqBBV46jX6m+SOrUgwuLc9e3KPthNvi0rQNzUlx
3suFE5qPgyGZDmp5hwu0dEcu7LPez/m1nJKmr7KJmF1VfPDfUM55TXM/ItKkmFemdXmUpXLf1YFy
sTYhNtCxahcSAFt8ebppLW43XpWt5F/t7oqjkg9B1GKAMEgjwnc32lw9Jq2I9up0oI3yegvUMoDG
QlqO3c/FBXwF/AsqB1iKI9YmBdUDc4KdszYLYNH4W9VIf3XKGd5fKb5+9lI06FEpYsduZrY0CLDG
6YiuAn/qXgB9TTZ33pGONLbctEXJ/tpU+WBm6Gwp4ollA3LSvA8Rm0jKhcP+IY5HX4LNH0qBZzDS
9O8Ga+maxI6D82nZG3D7RkMA3WcHJ5Nrb9YX7JzIvYpQarCxuXpYZjnSqiDDzlvHgwm+2fvW6ufQ
ddWhb97DCIlPMsmV//WiXUgQDZ8Bx027ElOHArKBnuxBeVGhbuYFzAsSTVG3upW2OO3VgsGoGx03
slRMAleCvn1849kNCnLP5QdEzWiCtetQqfBeFAymvSrtFvGimkDf58XPj/7GwHjY2oNje7c9OlPo
kV/E6gQeiGMcYttDnHHNwzCFKnLVH/5Hp/5dixTyy7KjyN/Jg1DFHik/6a0NMW7BRXz1fj9CIEAI
zg1wXhJCDZtrAHXqPfiYCcAv7sKVBvCmDJ9JN4j5F1Kw2yWzi09G9HOmlcf5nZl6jryAQekMZORK
iSFeamOjALBwlc2Lam7EGWySW+ReqreCScQUpXTVkDDCaAUdAH6vFcjJqEghZHoO6KcTvOuaIYJs
vQn8rqbRbOSZfe/rH94UNvZlyxP+r8A1jnJscBcB4o+3XJi89hcw8ATKxWpZ4EvC4InHfqYzZxE7
j6bNpfpGr4Pzs43bREdK+0IEuww3/W8zuGvNSasmarhEg/QM6fKUEGu75JGZsNLQ+cZp7LeDiI0S
SONAnN7HiDClnMolvWVccZKdaullGxYxTh3s+Zdn2ClatMWiFJTD8MtW8f6w1HueDkMG6ZTP8bFR
sLXtyL9zMC/z/nhShTfwhTXEAVIW9x0EGIzaJf3jsk7nBV8U0VNBvH/c7tBB96qi2mEADfeX0ytd
B3YjtcFaU25fMl167nZ1RrIjvgL0DfFUvHfMMihEy/oiYOppH1ekqoJ4ZFjf4QCWX3lkHGzteBJ8
8AXhDOYZnd+hEfaA1Did/ANjEePqrE4f5v5v7v2qw5JMgkhK94vhYTkP557MlRG5PPSvMNPl5Ivc
IREHgRWwCsiBrOBq5nkhxncgcwRS9Sa6VNTtssN3VKcacHNoriOBczj+KkWuAI9uRpqt3UWG/HUo
j5oVPAgeVc9HQrPkEtkoYIpaL7SOKnwYEUl0nfdX9QfOFmtrXN6rxTyuKoBuJrZeZrXnPSw1EjJC
xFVU535pSnvgFqvD+Rs+q36UTzVIA6pJWEmIRhlwuhV88zVd/8UsAlvdBD5SUAQWnVAJO4AbP9vg
GUVqyIbxZtGXU5bH/AuSwmBv18UfrXVic6DN2+J8CGqomkIsc/84cAUkNM98HyK6bRn1MB0eC6Oa
rx0MTg4cuG1gEInUupU/mB4d1EQb6JB5xGVWWVfV+QdMtxiF4drnijxR2WAL9q9OOpMcvWYYodGw
WhsimGflSmWDZD3nB6ttg8KmHNa0ut14XWwHZ1dW1m3iPxrq2IIZPkQNqUJaDEosP2I5AZ6GOxvG
ZYOM1hR8soqDpC23qgkdcmyFdu9aUklfq1EwYeti1z8EDq6ec/dRMEghR5bRtKGVYn9x7cUNbb3+
Ripeck8k8dvazBpvtXTlCatDDBdqZbGT0jgTo4LdO42U5PAOa59p77ci8RJZnRYoaBjauTrm9wr6
UMVNrEGV+0NQz+9T+6z5hs2vJUV+fVA+nOkRFVKxTKufAxiqe91ru1U5PshDy3J1b+nKv8INeUJ5
6pgOW4lh4sRqLXl/p4zAuI477oFJFUWJtbft4AqQCTeoqWNcuwG5z5o4Qa83EI8pUDxDeUVUDOHx
zdhW64UHIA8jxIkINYj7cAygL9pFrh+a96B9nverbhhQtBY8ACqE8mCNTp4IiI92ec1K3lvmlRU3
dynmYE+ygRMa3qntUjQInWRsCbsjrRepDKXnXzujOyrB+7PspZ1CijqycVp67RmXQFEPrzB024i+
OHABZEAHu/UzFROJarnNU6xKnyZ58rVROCsiHxIkVC87O8PjWwsw/gnjONB0YqYvwTrm1adLSsRh
oQA0bN8GXLI70Lp77UhWqRQ2psc+wEmJh8a17wHfzMhrxKuquISSb5FyLzgAm2SDxovvITCeGu+P
offtAy0JtA+SRTMBchvCwvb1d5GOKReZClLCN1iwT7Dbk8+j3gNdwl9JqLDAYK397W5gbaL5iPB6
xRb8VBWiE0G9ZQBDQuovXudAeDrmCy6AScvSK7UU2ujnGsvYu8QYZHU3hXFpdAjQwhB8NHjHjHcE
0Gg2yUUTLgwcHsCaURSMx/DR4d51xNdivgqZuN/8iBkXnEShwh6a2XbwDCMIjmPSjh88pCbUr09Z
btvU7pwtVMiipWRAjuOgdCEiDAVZQYyrzBVkFwdGkN7Ir5ZCScIQte9qjICIUwDmtoBe8TwyeeWo
TsblzJ4gm6iYOwFJXU41oDYLICAR9fPkkHUHBpYEG9iRS8ZRcaTcLDy2E3Dd+o1RLYuMTYQY6RZr
Us0X4iAmNRZ7YqLnZvqs4ayacldiDs20dI74lYQgzAi7QeeVCZYwgH40RjP3nI9n5cN3CXbBZdcs
+54p6CSF3EYNpsCW0uQqyjwacVy5aXeHQKV52zaGJOhHdi+A6eRSwvSYvpoTOd8uhC4G1XRFyqbG
SSfvgwRFb9hrU96t+NjWDTgo1U9mvdfsBFFTdpijCDey/Do5Q6K7WIkmPEbT9tP8m+bSP5VUyu9g
EhQ9Zgyqysx2DWubWT+J8YOr9ROhOluGm2ebWkIECOY0kfuP1VsKN4dc/dCISGv9vB+wrlWI1Ug0
Pc6MXtW8UAznZy5LNydXeTUXdJ4IId/nKLOD4ZQEmP1JOJp/l9K1hmlkzm4WNz5fp3I4LyjA2qkl
A9icxSKUG3fymmxzHwaa7qL+ux5oeZW4zATkmu3Oe/6x1+mFF6tlLzbC1TMd5FOGOAB8uMUikfY2
MhasqwzUcJqYuT7wNk+7RnIrZImPOcCItN4rIbCMtnNXK4zr7YcSAPEwpMY9KXfOHscyS3mQhl9k
0JMGf8RvO235MuAJLWK/bjeU7eVxLJ5Z/jPq4mN5iRQiEImr11GhQ90uvwRu26I9dWFCU1cLu25S
ZCowifBAHKGzSohuupXbgLCeTCVDHPUz8LojxzqNEKRH0LV22y70+f2+xf0B3913KzpsSBtp1cHg
vMbB2xqfC2HfH7wRC/q5GR5xp07UQjZfkD36M7OoeUycARxQqfIuoo6Gjxm+ruOGG8ZuWdvrysYL
OyBwTWSUK4JS9TLVicT1yw7o2Kz8pfyGDg1tm68/LGQ/+dFq8EaqHVrBRdODki+/5PxVUKv/npAx
P7SZqmZOmzbYxGXwqmsrkQdRqcMMmPcHSGidFQEvLOQ15yj+R9mAUd8NtbuwG+vug4h+99L+sONU
Q1Crei2zw1iGIq/bb55Ey+o5s5e4EE0xTT6MjBH8PNSbDWIURk5cYWa7WclOAKOkdbVejQe56KTd
U7cniNwViKoiBo6aAaHbULnU4/y5Ly/l59WuwbfVinyCSoLSaHP4njmUmgO9ZlAdy/PDy0BKk9xO
BI5eCLc0p6D6TxVM048E0bz7x3EScz/vHyPCFEbmuVpAkq0qLinYtnhVLJaXl3Bkbx8isnzFONy/
PPXqT8rabUVx4h9MzJ17Yg94wTRkaeWrkp59vW7NmbEa1QgYlhOi/Fg38PN7Qkiv6V//mCXZJawj
6AZIb3f3v0eah8eJnyNbh/djwNN8QfYxRhuGD10+nrwbsoO//5quHU2xO+KWf+6q0ssyn2oeF4Hn
zzNwr/9NlY64NWm1c5R5nYT0G1d3I17mghf+79KtuyXcTbNFb69roh9ZBy36NSI+cp8//Aetw0id
/8aCmALa/VGD15lSpVKVOiEqoB94p168HA6oZWSrersFi1BVSB0/uhuen9UpaiErrYsXsRI30G9Z
Kn2X7m2Eca45TDr49mSgvhjaJyi/9OoMYhvCy02GjsnuPyFb4Gt9AC3tCAjtXwD1SIADS99B1SoO
7kaqsVJnwaglmreP922Hjvl1KW9YF2jwOegZTcFBH+93/HVV3bxl92Ii79Kk724lA92QouTc4OcU
3iZY6zXsSMVXPDz9gmREO5yY8Po2NicuI5E8Ktwvfci74FB15zp9/J1rLk28Q4BBmAGK8pgUky3B
NCgkqryByGVkgYjhyHM0Sa5IdQUTfMlzsJmdh7pchyaaicU5cINLcQLkSWNGMyQbx77o6ZC1f3Vg
w0UlUCWZ8VqgJarCYi7+gW0pMGXd7qNZxgXGK2sH5MAyDUooBl7tXqSDa+a9ei1ZlcN77LS4vhEW
wmTlrQIPFBef33WNRVSY/39/xUcHMEWqR9hp9k4xFGWBh+ifDyxB7eaTv5a344lKIn8W3JN4mCtX
wEK2+BNuoFokCRNyrRvY/k0DS/ZC26tcm5mExBbIsELzOAIbeb7uKwcWU6lfwK9OVLCk0026ilwA
JxdOBUK9lQ7nKUJm9btEcjRwctYEcjhcwfznHn0fk1tPESp/mP+rgflmWsKQcp4O0HtFuVwsrS1U
KCbEQhRneqAGp1TQs9ONTrXnMvUC/57zbjQ644Qqi72/CpHX/Aa7H0CV9BUVJfqnnysQ326XyNLn
lC0LfzIKpIpncNaaY+24zkuMe+h3wOSdfiozwSZrP09deOL8CBaANC83bMGpSk6bAuIPDuBtIWeW
zHsJbU7pje62nPmYWmpnoDRvIGotCCATBQPq5iBP+yvpiRNVt3+zQR0NPYB41gAJMrgA/isaJ44p
h2pzjzixVPbdKlf2PtCDfhRpBtb3w7KcslPlVfjoKGl+YzsKV94AWzwHGXq8UM2+fROS4sR7SbqU
nyAmi+Hfn9V4NeunIp6JBQX+O3GlYXqcFZD72dQwBDG/dseHXed5CP1I3oTc8D2LI/itFUOe/yo+
JYvDxh7GIHyXZc5RXojaoRXvNYDS+Nc1fQu508MwGpyVJAB5+NsnFJ7h3E8N3czH1pwljHnzjxCC
6XB9WLWfeg3wu99eV4vRgmgyt71mzoffF/jisAUY4adARHPlqbydPmMEtzDs9uXQpETt5LAFikIh
9WHpig56A9UbQeZbjKUx2RuvknZGlafKoajJlaRSIANvyBumM68mjXXC6mk5Ls931S+lOJum1HYV
NiDJAZT5ceEJ9WjmmZ8Ubu4RReznbwHHEx9e/KU3TU9We8QLuVufxccO+DePZo5zSnxl3HekU6jK
yqxoNg3XPvYqzyaAkU/pZQDtMEDUr1yRJNFU9fcwr15IL8yLD6W8Q8NIyB+8nUSe/uuMqJJ6K2qh
ZhsGTa5wywNPCH+/bmkmZuAhL6qixLfemhPfzaI1fjwr6u9R40ukL9vT9NnLwBSJD0xhd/LWYgHk
yLW4H0Ws2aKmi49WUuRaSgua2jll07CRryePpIRVw4YfwA+F9FUpwt574LRinaK4nJG/My91UZmr
aWAOe97HHSMt6TzKpc6tb93QqbsYdB+a+SfKDmGTnlHHEoAUUA3VYBm0nc45aFdXaGsN+vrxC81d
bKmH9Azma8kNvUJm6rPG+9QFAFkgrbJd82hw8VdWfny9eZYCqoKI3+adNNzeMWn12n/kBTwHmrvM
S6zKtU77T+ZBiAmXnWwQRkEFJFNFGNKcaHG6DMadr22H/29uGFmqtrw+Mcc8IUshLev2GNpaBrnw
PXdSkT+SUnZcq5KpDZa0hzAr7oQw04vOdwdp1wJtkhskmfdFG3l4fBoui3H4Qds+0sx7cNi5XN2K
gc58jWCN80A6iAEzk2X3ls6FF2MFLGqM/Pg8zFCTc9YkFucbv8u+2Z4kun9ylZTL+tKK18bCOxww
BgQHfex41P6/I3aaCfxgSUewb8Z+HsnT6F8Fv0BFOG4ZvY2bjhfYVc0z4x2n2eI7md5qLnwBr7RE
qKz3Ze7DcS5Z66UmmPVbrjUGV2MwUUiEjzkHko9qPp42/t4pvJkJTSpf/+QXmVNrbbykOnKS4WHA
rFzBoiLpvL9314sJ7F8vHxbF80wersHjzaKQwva/uycxN6HELrcPeZLS/RmBuJqT4uR5DQd9169E
99bBVx/TVKLaXWHvS/5corMIWPN2/e77seXeZ046h3X08lsT2qUekAUdUu3N8JSN0NzMaFbamxg8
8KowZNhebRb1aTsbOK1C71JHx8mQmXGr2/3kVZjdi+smS4dUySi0E6c3zyENA+UQcloUL1h7L+XW
7kNZDdn4aucFlyQZaQArih8PKhJ2HqPqcNVJq4TkosdKcqA7W3KqdxJ4Hgv/EF6EcvJc/IEabGNY
F9AttHM5uflIbjiwJobCoJWofeMuNj35ge4ppqHlOgXJwBxDPgNNQ2xd66q9gSPrv8ySfdybzeDs
FMrIM9ZWv6ucBrYKkrpcsi6L7fKi0j7mPJPoHyuCu63PVcSokVMCjPyYoVWPIG1/ZSJEMXUUtGUm
CUWtjSuj1qiW9pyIwTfNe51E46g8TbmmFnLTtbd6XQV2ae6pWDx9JblEv1Dq+8RHGy2LXFfLowFe
pKepBDYSW4p61jKOn9GEeJOBGG5E9ievLrq/+sEmGVETjr9jQhJVClQ0TN+QaC18c9phjHIQtzAR
8zzbl9Ub+1lYxZMWznTHAgAlBYMTaDkHShhOTuD+ijCs7uoM9husreOo1LhI12SX4VZc+4Cm5UqU
2u11sjYlLPwuuoj4SAUWxdo87ZDrjvpQDxRvYQjL2KxHrde26sUFzUjF7mUc00LAnXCYK/Mj2lf2
uBThw/DU50b8dCJbrHUwseZe2i0F1YIEQ3fBknIAmLGSWwDca78s0FgSmqepR+vOjEu0f2S4p+Vh
/UvD6m438UbtkqQCbLD5xTFrSS1QeW/V+KqljICAKW8MGB1kbRyhvu8ATLxF1LLOqPwr6e4VarXT
+rm3QzQs2s1DZThlhzT2p1o37lbzUzh96iogOSuYM47AWmYzyDfq8Fflf/ICAAIXK9bktos8XZSU
kiSoWVEnzM+ykBA4GrBytwUgaQQQvOkIBhXmp1YI2CMqj+amQJcMOySm+lau7pJuNZMvm83vtOWo
DBW3wFlWL7Kkp3ovMYHjIQjGuyxTfTwjbKuuMT3vp4SvHSQ6JZSA37w1xynggsfe2VMSvUyL9Zyu
RO1rKNVT1LPMNdn+iE0YL8e2qOTHcTzGR+2BMPufhZNji1b6BS7pX3URGez//gDOWvNn8IOJrbyo
FUfpvdtiTf3RywEwDY+ETeBmqvGQH3HoLWFhvp+rg+ulA5yVZpIMKsKlmW8ysuQKOU9MZBg22ssv
lbUdLkGee0QbqDHEeOHwTBdQwCj2tHi15viYl1//O07QZxTmmyxgYMCg61LmQNXX8fId0A0gdGX5
yX+H9nEdoc1ZxtgTVG+1ZKkz3DJBpoOHEmkfwrL8Sd341OZKxcEMuPw35Ap1AwWo2x14JxK3AaRF
DJIgjdPljeugtPHJWLclorulBpsRnUF/eP2lioSLlcy+Ce5NUIFbq00NUu2/LlocC9uYsX/b54dN
P42v7sX/0YO6CledgkudHxFoSNAA5luTCHtLRvKYmsdLImQqXNV5tOipGHOH+jeCMYLBv6D8nfIE
YHvthNybetdJD859AGdtVXy2ZU/ysOA8Fx82mLd2ruMCI5PCfBOt0BbqzW4XKe0I0Ez2HEMkXCzW
wHRfDIcWdaWLxeIY+pYCBDMosZm+QemfLYaIH2nze/3ThoisnK0HLvPCoSXQqDkBv9LycL5vQEAg
IxaGCw0NtzMfPwPM7uzxWtCqZC04ImX+XIbzFEzprDGXG88+2dCroeJOwpxli6PrYIGOC1vK1M4a
5KHUg5+Ym+KXeurSuYxOZwZyTz9VVXfOo79zraTlOv3Ym6kaOLhld6NVsgEmO+VDWk+4zHqRVI2s
4VhXfsgao1dp4B50OdH3TLzul2TYfP/1Cg6p+aLyXlpj3I6dw8u4W/7kfEYo7fUgs4K/lbG1iJ6R
2CFCf5spdhbkET1k2Z/rfjhQ1erWyI3RAGJSzr3hQS02TJdsKnXHoluzv34BefGjMfjocTPzjWRZ
92yOEOrDUfRLXFlZnKqKO32OdcribfFihzqGNEaBRplMNsxGvZf+TtTooXmso3hs9KkTUKMGSeJj
EQ7u6JXUM2/9dp3jGGZCGlnJtPUf2pCpxLc40zUV20YXuLZhrZQS89X+tF+ZvRj8db6cqDerE56O
xsFcIFQ1XNu6kzSTIeDgNMYiadpOYzBL/qb1x6Z2mFqa2E24gmI0/HLnbFRF9sqsSa4dH8t8lZWt
/SAqwcC000RXaSK6/P83LhKLTaqf0sGOM0ppestm6jAEcG5NH9mAl6VVIC8DxDX8R6z2GHKFK4sG
yJ99oKymDa5MRwDzkhTRtZdgIsY9bCv7ljAupzV6YLQ/IDFnL94ohsIOJYDCzjv49Mskxu7xMPZa
DPesxoC924B8OwWJXLQnBwSSVwWhqW6zy9pWAjQpEnW9kBLqcgdDRKMc6XTw7Fys9YFPsQYjNfBi
/GCD7BLLLRz5AgqdROvwByHeQzkjoMhysiFqAiK6jKnr34p7NZXtBaLMn2G2aTeVZunFJFzf8070
QHoY7T+1warXeguoujwtKilhjtWqZYuvvJjNpH2f4A8fkRD49QM9xNNABO8oRZdU2+v3mDfrE4+8
39Sy5QNfbPrFdkp0SQA6jv6fqeOBQNsxmluPFpklj/PpW4+R26wbr+3aW0ykH5s4tzabI5Q6VtBD
RKI8zhLHnvf1lPPCY3Zs6VpPvy1qM+N+M6FsLCoz3jBkwRYP+hvAspPe2sya3IG63eooeix/0dU/
iNIWIR/+RQuACRecw6Xk/CkiNRB8mQLQNsBGlrPN0pAHOj9zWjBol9fJTZA4EiWGbAJHBhkCuFIX
ZwNWN9V0RxqguGRZFfcrK9hzsRqJhqMIzN93IaPTAIiYdZQ0SyXyFWH0hLGHPVqZjXppJ6ENf5jS
kz+A1u40eweBovjh9ysJjBTswDAMWufP5dgM0HIBRFOV+LoWUxVQ6nlLunN32ddSHFwJWNF+uQnG
Nhs1be5Wt6RUrBtjnCghGmXiAT8tGAHso6uLyPY2ivLLcLFWxuX/R/xlbvzTtz+4CpXPVpPTuKUS
yqWHLeI4CrV8NRWxwLT8oUrjpVc5z4mtZVq5JSILOl2iRmPf03idw3mubJ8pEnPFsrU/8uYkJJzw
w2haNFL9JrQBMwcwygZk37dHj4xvwSXLxOxTMnTV1PrHkumT/p4z/tZT3XmtX+NARQz1vriQ380S
F7O/Cui4lGyLouXaaBKZ3B3/V4ZqHMY2RZlFWYxuS9zuJQ4gxzgZO2kXgVnH0EBKULy+KvSvuBoZ
1wWJKQjLi25whWMYLGe4Qz0nOoEKJX7VwyXKfmbuPi9VRpSvDSKV3vdL2CHU24E+X/ryIg8ZquX3
IagaQAP1C3uavUx203rDDsprzcr0ZgEtSy+11Qdv6YSt7REMTAsReG1AR9fx+rdcZfjQn/NJEPQp
+QkLM2qgC4fZGHYlcXXuEhnBMhflQOjCNwGmye2BbOV+VDnvSilWzl61eU2Js6bOlx+mtbdoZ7UA
ypivJ48VqOdD2YUD8fgksjklWsADQJPl+zvDKL/vZJV4hJ4gNZe9ByVQYhukrZAd7pAnrdcyUNbk
vEHXVXiB7p8uSZ7pQDv3C6o3104LM41+rBpBJz8eGHfP+bJIwbWjClO+eOi961DdgLEhKHuCyUSA
N3zfCxmum60sP1bpnwYEnOpyvyjIVAuhtazJBGE+5UOANLoud/ixUrf3WHMC9sEsrph+FOsqoOMq
iS1D2IyvwS0jyKkUImgq4jh+7h1ndQZHtcmr7NmcU2XWKgb9YySSOyh4jeQ61mLJCkG18XYD8ujp
6Pbrzfc1ZSvWSXkKB3EdOC5ErLoXJ+6H0TdVNNZJImbmKKTFHfPMZcgTUBLux2nwoH81CyNvJFcp
vy8tvMkMi5oV799g4HzmOMszSqcvVtJ07FLBCrARmbYx9Wa+7M+HrY4eUbvk2wGDMERkQENY9iHk
RNUeM4jK/K53Knk/RpO1ny0kQv1EokKvziChK7gohMG4PBZMUHmj5+4XbMQV3JGAcFRln2REtxCj
AeX+smej7X4HIuwSVeygkNz/1h3YeZWCRS59gej75Qts7eCmW9OajFTIGohUqWnkQ1wbZbodVWz8
CLBPYZglz2elKVnbB/0ymPtPfl0dNoiPdMgstOrv0NWnq7IeYZ6QNbNYIycAYKqNMilyyMPlPMOq
s7+ow8PwA9A5Q9D5cyhZO/3zWdO4ZbdTVPUWb7J/j87o5f3+ePlFTT5c9G3M3YkPHzgM4TmAYJiV
9/geR0Zuf4p3c3vrejiYdqOXHPYL8HV+yhVB0jBU6Xv09H8tbKOL4So6dym18i7BHgHssxGwOah8
4TDvDKVt3+M7RW+uwExqDCWiCQe2rtSrMxFi2XvcyXKELVpJBbBIYyyZQfZH6KLq2le+ZiPPeC1s
t8dfBIvgGqZh5/atS+l5cT0qZS9UAq/ryKIp3rBDJvp5N+qoZk2PRS27fMNKkvmtjkX2TXiGcPfk
toqbF0wnAAxiQDEc46YchSJoUCP3w+4YbH26hf3k3ymST7Ryors52T5zAfYLT80SyLXZ4u8qQXk9
H3wG5zq21TOqxYIwh0mV08Qi0UfBrYqlFcZrAfTQuY0qZNBYWDDzpUvSLlhIYJsWfjP5Ph/pdBVp
RevIlbA44GVLDUJG6AfSADnyWgTkf5OdTYMPs4RiOOPgV1xiMZ8Q6J7xcPfYEKhBrKbUCBWly3Uy
C6VmxcTnmzLsvCWTdtONK6v4iYfZIc2yx/kphaun8inoq3ecIvo3wl0aH+d8itOP8qxvQfaKE5aT
8ytfFYZMa1VVzOMXQL3+JabgsJpKu00X44ixVde9n+iIXm74BBhiOXoLm7xCrNQN92Yzx3fqo57x
2v4/n/+WueaXZieF6l3k62e8PsdnwioJrELSuqn2MI8Zmcg88QuVrqH+huXFNdMum3tYMpsfoqnU
f7iGn/bYMoW3zz8g3fm8YBM0vsCTxLPhXAnURftynmni2GrjE95gz5cI5JEI2lnqqa9/pmboS7Wv
ijVdQFa2oRK2NGEjdjF33r0tO8LYtobza262uFempeWzAgx2AS/RbJ9VUIkyWsa4zi1wDtHikGmY
LWS2S11Op6oL5iRlcbAi0hhaZuVtNWPQjc0CZWqvewLBP9tNG7+2YZ/egmxdN9s5xXlIJ3LSyR1w
5EPc0Y07bQf9r5eGqQpdgaug5RoiBVFcuEemnZJIajpi20R2cIdSrzdfyZFBMCh3Pnobx2K7alMg
K8RfLCMsoTrj/amtxysZxTBI3fpHQp5gJVosx9qH0kT47B8AZk8/6jlsscEQGVc41yw9RChSYsjk
sHKZm7UWHCkg83BeYB62njPQX/usNphUNxEYHS4yQmOR6FAwsxZfpNjLDD7JKbm6PnqCuzfHQFIj
NlrDF8jP7lslZM05ocJMAMaB22Ma4wjaARTww9w9v1UfDhDo9Ul3Q/yS0GnD1lRwMv8AY3rf+pwc
pe2mA68tvawQEKZCnb9kwB68BZYGM1s5jJ5gIp71We/+vINaUAida8cCuhRgrrdyJ7psWd5Zuqsl
bdlibsF4J2du/pEQlkTsxZrpFR0ZQEn1T1g3k3Frcy4EkOXn2c5dITnH4V70sgH1icZve9yDASTb
yxNS/Zts1jmvBx8L5g5fSzOIxDzU5BN1sP3xkC6jajD02Eu2ynR9B+AgV7Ojzvz6his++jr+F5zE
MZwPH5QQpQ/n8Jf208V6N0Fk8bnqudm+nTxRT/RCP0V2WeiYVtdpdnqOQA9lh/a7b9LXg0eu50Pc
Sm34FBUNN2b/xZz+m9oVpsOY/AdMwXV+3Iy1IRq7sMfU+JOj/oRxEPR7anSLD4Nx9xAztqj7qfvZ
OVhdaCv0nugygODkZ0DM0WQfIZsTg0rw5xyeveoY5+Hx1jYTjJJV/eg5aetbKYIdfaTlrt6T6Zdo
8968ZfLjEj7zWTnJX9FlSnYid8warZuNiC+0wDCNLM4gD9/bQZknGCsERwMOy1z6FfLHNV18VnSq
ywiXfCa/gKfGWOHOtsKm35lbobBAPnM64kuvaP6nuBRvZUDJtpwiSyEM2PFAFJUAjbh2oxEfuJEQ
s0KSpM1MXbEH49TkZR/BMAmHe5jc0nqJbfLBPfyAFZNQrBL4nNFjHTcPhQIVfO6V1ZwOJpieezx9
nAv97geN2CIp+EwrrzJZoOgHRV/qKKOCo3/XN8U0EKpUCYX9pbAM0fU+LJxrWaqU3vc3PwQl+Y3j
nYHXrrrOS3WFRs/VQxcMqXEcC+OzlhzFNImbxzEJfkQ4SR2gNIi50qX0Doijkv4e6o3YSRyZtioA
sHHdWwLFIu2+4OnMRt2ft3s/npGkYBaMucmFTVT0Plq594zNGYxCl29tAaBpas8itrvU45uSP87w
XMYvnhhrc2QSUj7QOASSzhW0gDgg9ushnQCF6sr0Kg4VJyj3P0avJ0ZdJNeatNxwKcVsBYU1Wq83
xjiVe5aNz//zYdrv0XX68KjEYFlFtupXf4ZhhKyS58NyPbpNi7SJJO1r8wWjk5b5Lu8WiLxn292n
NYHSo0oGsZhZTtwg6eCKE74+OgJUF0edFvL0Y67oTBi6z3Ya/v07LPOixPoo2s6nifBQAFrz4pH8
jQDbrQhYHGL8UEvKIxhjicXk5JZJK4/QS04KiSTKNZhbezC3QnL0HofdSW0ZGbKGD6vePJemgDS1
4vkXw4yjwnAGYIKOYoMT8eyDo3jdD4NSASaPXHWduiOaHLZPZfGDvtptnQM6onblbvbAjO3p7yaT
ed19eRd6l6v6fvDom+qyDXW4oBTQfDN0tukxWRzFnhsONPMVv34us43KoGjwZHKCj79iDIzU7GJi
G4PeIIhs1hjPbwP0rQ1c3JTIvwiiAl9pz3BXguVRdwFObUtkXs6sjErcxz/gIXn+3/TpWIKpTuL2
OO/uMgxA4UlI6jfJCEJ3NbkrNYBzb+KRSsIHs+apG2vcrPp0h2SKMsvNGjH9D9QAR4l8yu5AxxPm
ZzqKLYXM0wYs5xWCvBJtdLODIvIT8mfo9MextZIn6rie2v4i3VTVMHkaRFwSPGzDGKtjFapZWY9K
SXg1OFQkCHS0omb7InnufvcI0VnHavtqsuPbrSbr5tN+Z46y4FWFrs/GN2blonpG4op4HlGdvhFS
9oGY+bcCDGjSND8CBdZPhpZxh+1Up+HAvDu96Tmh0lnKzZLvPNzkFEc6kT9pbz6/mwgcf/ZfUDuV
TRibKESMUDl8iSyLXe1nJSav8wgJyVFPXlrax6VVJwxNIXwESYfBbR8+3T4dNQmAVTvKowMDiWot
6tnK1HSBJyNll5PA8EDFa2GxQ8b7fq3esInygPMOuMfnAv4Feb4+milksl6Kje5QJvIUb6edbwuz
kZDbNglR8XdIkY7GrYZ/rIgoP0sK/NqxNeSLuxMCdTJFoTh9rXwok8pX6S7ZyZzaAmP6q/YRNTGX
IUnH+EP6Lr8XPAEx9kAzYxV2syoVOvLwbSSMD84u4pRn9I31uyWTs3Scspw+wbGx+2nYX9EhGurt
DoSSVD1jFrvrxZi0H9ZdyahnNSHvOJtmwmzgV8NztSyhX3v2ul2R1OnCrzkuiON9VKD4AWZ/Fvrw
lwt12njvkxSHF4C90dVzHXU2s+KxFBnE9o6M2Y2YlYdzgH58Nst4cZedQbJu51cXVPPnZCcdzr9T
0K71hPy3Ykwi6rvNpx7/hL4vMPnU7TpNiskiv5In582RVdA4My2+yRX/cOE61bzJ/j80dxV1LXfG
y6HB7Uu25spKtTDYbv10c545IGz4fFBOQYAxuE59HOpmyAlPSPD+KjpH2I1BOBHZUzoepl0WoK1g
8HkNXcrFSkTQX7ePgI57XtYPmf6UCkM7xNSc14eR6qaFk0YakuoHekr0vNmOk6GlZeqCcIhqOppq
0dR9LP8iJZIzGA0ieJnvdsBMJnV+Zj7DOA5QvbYzzggsB+3+KenGfZYPnQufm0ZVLzVIXhhIhB3S
XOn4US7T50x4cnJ6PTmchWaIesORTA/6ey+RweN7du8yUeTw+9TSSJUqnx2oxyyhY9/P4GcsJqVr
ZQs5X0fFcOyR95GCcCeO05K40QzBAV4Ld7P3Jp5/DekEcd/UMSicviFRcpqel4rt0O/UHDbNDVgr
3i0A9uzzBzxbsbQuJQCg61mtAbG8h3/Ta9VsDodToDdorYYDS0wnXRvMEDsv3Da4BGjrxnLT8EBW
rjdo1RsWeULdQsPKGAPx+CXyP06GPfUpSqQsiVhcyQQV8SGzbXkQHeeAM6JcFWxadzXlgpbegzLI
ClEzkHD/5Fnvvnqgv0nSmoLNwIvl0bf/zNHuW5cV7kpxmYgylux6FKC2dovQ8NbS2DbGJZlWQ17g
S5upClZ6uHF8gR6sA0NLs+40bFC8YwKSDyqQV3Xo+Ikpk6lbwpq3vog+u4AO64hPWAlz4smDVqYR
izQuyZ2mUEJEE9XpTGKPcZnonVwsTNmuDfpvVDuCgXTMMaa1AgLSC0xXQZ/0bnQC/xxUTd+NY1wN
VbOg/VbEY0c6j3FBs3r4gnhXj+P28F70XxMRbyo6CByzi0VRRxGhytctvsAt9AftdkS64rSMGle+
rYzKYQ3RVgBstsUNmlMoVf6JnhOCBUzNo298HGxfSUhXWKqrdRjUDxCnm6VEzMu+ASSZUT1t87NG
DfdTW0lcywv8NhF9Ai99c9K2a6VTims58d9q2A9n/1mQr8kvALiimlLi5gX3c5wi/1S2p+GTgn//
mfkBJtI1nxb/vP92fwQzvgUaeXMSxSqN+JtSjOym1s58UBbXOW+7APGC8JHQtEnnO/FT9sLgWZ5f
3bLAtsDxk0RCCsMsQSBZD0aUFYoLcT76tNLl9VGY62xnEkfOf/6DzmQk8Do76w4cev1pnyX1NPs/
JEedwrZh4zN08zG4Re3s3kEuBofjjJDQ66KaMT/c3IBzAZLYk3h4FcT26kkOhhDwlmyf32ztUWmR
R/egtPQUekOfgyd0lZGKeFbIHdoIkbbVDHGYTNw3tFbT7Up7t/s5WN7XdmQT3E0CM/N8tSyu720v
e0uOeUnzplNo2ar6R7a/WwigXS7UaYocQQIv6wiFO2ylAgYH5W1lQIM73sa6zz+zNgXR3TQ3y0eB
qn93UZ1EpY9o0jYU5MfSvrVG/em0J0COiVb4klDb+xTd9pQqZ5WkVuyBjF7DjEGM1LtGTot72ZFH
CNYY4yHjB6BqImAjf2VYrFj3qvsDwXWZlbs8HnNBd/vaERyGt6jd18h7DxVtpRmSCVSA9/9MiLnC
p9eCT8SxjbpFBi1CX9RWYvIXTTReWACn6zJf5RcOK40dc9UrIn4v0CGR4a8QLsS0JnkrUDcNRtq3
ZgDMVKwtAdvAwd6/APqYVPKYjqzk+A438n8jZcVI+fjEbzFgzMNzZOA86Cx3v4aRYGdSYfFdnSEi
DnVFPU21bDshvad8oj8AYxkS9s3fH5P98LSZ850iJbGMxguDL/xPOG4rUvtar1Q6RA5Rluo6fjBg
WqR7AucDchKM018MW7FX30Xu5v5seiojRgoOFv0KOE2ujmFcuwTvoQ7onSJl0ZDtM9v4UltG0d6X
xVPo5LTnx+TlvSvGu5mczjAb5Na9Y5XOiN/lfEtIO++4+e33NsFG
`protect end_protected
