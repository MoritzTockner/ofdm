-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lwBefBLgW9J+ikSin7pH3zw9Xn6VQXDIKAojF55mYXalGWhQ6aniVsC9e+sEeDWbWGtgW77cjub7
+dWvsFebdBitdJfYKZjuvZDhZ/pQ9ma/3UIJkNMLEBKGo56279sXWGks7I/vi1zKTh8wgXwYxdnS
f8isgQh3uTHLF+0pTdqOmIyMFMv28YOxhttkHhpBLAI1j9vXa/0Szsa5x9I5xvip6cPPIMUDHXq7
JJqL3dDCcOW1TBboGQ7GQBlBmSjE8oQbmGaE3eo3w5zhkpfud6L7Mv4IoKiwQil9aCNw9sUeeF7Q
+C1oS3UIQSyJ1AtRKRNYGGboN75sWpUoJUVnAw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
FAAmsUGf1zqvgqD6rAxfvZugWWRejSzTpUiG8HVaUKvTcz/hJvzjkHvOv5wS7Pksr/hGxQBp6P+K
7Oimo1lTq5WuxrpPqEx1nnxLDkTdSLWfjIqf5qNKAOM5evHscIQaMfKi1zAQ9GqTmFiomEudZJrV
0H9PLn77sDxqFqoxX5ybTuZlaqOcVmIS0Ac7S1d+bjHPnrzOLgNF0p6rlm2aCoMWrosu+aa28W3f
Oihb6iJWUIYsOEN5DXctBcu7ED6R1VUxNqOf+l7igVPs34ozSvGepjfj9WrECHa8m1ua9xcil9Ue
8XXJ42bNIUFJNpW+6HzMXQPLPQQhsobECKtmZdu2LMWxuzZbLPaTH3t+Vntx0S/jQIgMaQR1iGrS
jBERs1JY3GKNRDstd3bSiNbdGouwlH6WhXrhCoXlEcpPfcF7gzytkXkpvBOUiJvvLwtDXp1PHp1n
MZn54pRBnQcjHBYdzvMgnOwAcdTUAdYeca9FebwyUrvgVStDxgGmZarBAvFyrNc5MM0YbStBq4fA
tZhYqqg64UBoEWkytWyVYJcFYSseJFdxOEYdRQftNbT1wCxijXkyV7vW/iL139NL1AThOuRGa7+O
cvdd3u+WjWcF0MlBkpcX50MOLjM3JJcOU5ULxGpoNv1SOP2N+9rMDXp8eB5cR6iKzygmGG1LY8Bb
IUPG6V464n4AOh/zKQu1IFVI87gLds6KP1npkm7OLCttU4dvUahUUPTXYtE7JLHzQXIVkW9m1oUi
WwYyZ+5/aKq03Trjc1UzFbWbTc9zZuAYE+okb6ruUbBDzR8BdHM+RYWi7sT0KRmtYPsmulQ3x/d/
vLDiDF/uryi2f85HILD0ClunKYZADvlb5cQBwXPXk/EBi2eso26E70Emuu2l+e1Dpxmncw98y6OV
6uZ3G5Kdn2na9UM8xBZeVCF+F6TsDWaA/tThMYI/y4PUHoToi7VQ8u3s7yHrb8F+bK48JPsz6xgl
ZWfwtcC0GrFwv87bIKfMyGLHJ+O90bL0D7l55TQ0D/D1rTqb82rFE7GxgphV8Xtn3x0gcH3EwNfP
9x1gDa0491SbztJ5XYuNs5bnZLXhcH6rjjZDiVI7kxTXhe8Qnmwke945E1hZuxiKaxSdfvG5YHnL
VZi/E3o6YwX4Sl+1w7ID745jRDUnvMAICBHHooZP1Jf7iCdeCAvctvYpCQw+uBiVufnMsoIjL4vN
hX4TNAG2u0isR5D3EU74JPirY4NSNbRylOjlqheDSNrNpKZZE074OSbCBbBiJSV5PD8xPcZb/dhG
XTXS/eNJF6vWMMziEmO48Uc3ViBiLNscPd+cQ5nGdX34LmDW9+DsxtZViiZaIXUoujc7hUfiEVdq
Gq9y9wuN4LWNaMYJmqPDO8buM93IxpHm2x34/XpNlVI4FNjzULzfkTx3ZnCs1Roce20TW04oRXeF
GTQcFZNgAPnL+KKJN+ayAkC9/J46uZdlLauzYmc4QwIJp0+G7sSLoN5r5uEhBQabgwHE9Mco+V9r
dYoyXsM5vUHLGxs/53N+z6OjL0UyKM7mc4+wGaLdajKzqO0+aQ+56lTGaL1V4IR6t+a0gSFUKW1H
LnPp4gsydTRXOcjCiJPBA9b349HyR/Qv7t6KeRqMtGxXI3UAqvDCrrzMwoShy9kJv0giT3zGan5v
gFvbq5Huvl+JZayALcASHzgMrpoQ3DEoPtcp1J+309645c7Kp9l6fb+QOsVy5Trleoto1uFyCT8n
JvpslYWXZbmKN1tQptMpW01JgLfeDEx88SXa49SgqpEmauVqpnhQv3lpHS/ecjNOwzG4il02kor2
j7ap97c47BP/qH3iPs/deb0HX00KPydFSvvQj1b7Tff35O6unvOg/HeXnMabdyLh29aE4LKbvtir
BpYjmh8dZVros3bcOCrfhQzmkaSmKB5VjrcyUY7K9pt2nFL4tiBBSEwPFR3CNyUtiGA0dD3W0KTu
oCZyjWr2BGrmmfdQiBxq/o8gr3NQB5Fk7yin4GPDRaRpW1zpctcCVSkN2z2bTlKrTgc4IjTaUs3E
nlaKaCNwWXTb8i6XLYb5R1P6aWQ6J6TKwRltHiFrAB0q20ipgtLilk3uEAaKieuD9m/gZcVqQNsY
Z1roMTLLh/dHRtumrQ+94NELIq91j8s4mbW9PrvPE9+vOXmdDJ936/nsHPXi72nNNU+/S4h/jdcl
ttWA8KDvmtKboWkBAphQMqfmpvGUTbFLPB+1/RgUMDGr1Bq6vNYCLLgKH6PXJtuY2fipNpPrmVTF
RonxifS5in/QUHCUAmJvIBDqdWWiDmem98buscjwGPzrUtPYwY0mRB/WH/vmeECUHEBwv67ArkG8
hmD17D4T0FNEh0dMusyOBZpj8aKbd3LfmibLwfIGwLRAw7TAbWmMSoPyuLUEoTpR1xugLX8Kf5OU
o3ZeqyS6NIsW9X0eQJnXuxJh3uttQuWSoKFUj4F22wlxTKghNm/N2g/kJTvcOiQ9BvwEkiQ3PjN0
XIXw5f9PIHZFvqn2oVj58BnBibRB0oWtn0hmJwLbxHYaXa0YoCl4Aa1Or1GzmS53iQd9xDSUU8ZI
9rNol/uBqMz372s2FbQvVicikY0FKg9rYbP9DhHx85nCSFrob2DWfxYd96h532uMT7agiivRlyxE
cQeTLZRvRKWJO+EjFPfAN+1441GohYZBNhCzOj7KZmYCRt6oTAvAe22CnKx57KlVFp/m36AF61WI
BQk338YXMT0tKc1aFX15U6b4O9ZhtE5JhfL9ZxYtrOI1zTd8Bqi7aNbiZCbERJU/m542mj807l3d
wtAkafSJi9Ht//nt9no+EUKyyF/XeLEi3OaZbUIvvQ8nMV2wpFWJbiPLrecmWpQ+idnadM/WJ6rk
LJcLb/pEBVhCm0y0qcmmBokEUsp9dTCyzjHqWjnafZ/q87PH9Llk+gqoxRRkr/Ff0eXnaHzHwxPI
Nk/rfNmBN0QSZILFHLBNSp2FVfNRMzHHmUnzEyhPUKLGC95goD8uaK3x7a4SM/2ijDw7RlGV0PVF
QRGcSpHRSzLJiy874YrLS6mzNWlszUTlxeqMBiOP5Fo6TQEpNWH7Uj2fGI0CKkcfSflUuQPCRpWi
raHe81mJj5F0M63ynS67k6bD84W1QPh0oSYlblDpMdo7t+1hkiJcVc+iRuqTmAUbgdWbS2E1lKzv
T9qNfkyCjXXxVFoAm30n0Mkxz7Rzau0T9/Er35KDdN6VnPu6XEFRn7ZhVsSqU65jhEic5R2JSFdw
r35bLxU3Gx1My7qaXir89uOA3z2Yc7zSfFN25Y2dzA13OxiRO0Y8iDu+Bbs2QPQKiLfei7Tm0hfs
frNqO7honRGXX+CgufvQegw8i5FemBSszs19jbMiO0cBqfIOltSzcm/bGWHmBN/u6O4fk0kA4GtP
hEPZuDUHcLVVZ7531h4MZFaqLSReOlCYSRwiSi/EYY1kqcBGO/6vEHBssmAtFnxfGEoGT0oeur6X
Q/l+oJXHVw8GAjU4aUZq+F5bN1HJqfOyY1qZ+e33xSRFIGvQjAtGSeDGYh37tVVvj0KFsD+d/duz
Di3OCQO1CZzy7g8Qx4ErP7nPP8ntUx8dPcw8PbT+8BuAVJdX8kmLXMzOtqvH4xI6e1HQHaWkppm8
qw8oVIeE45Baz5s/maASUtlr7BvZgpT9CjLbgk+0lDwIKHOV+DY/c5TbdcwvNT8nG82nTof6NuYN
usQWecX12DPyuvwe4SQ5KlJcaiEMMEX5h0M3Wpi5dd9vdqzV3mTQtiP3hgXVcNM+YT3rXc0Y4aMW
AUuVnT1ljBATLHwocG6h3hL7+SxrEEfg7aRN3CE/hFJYcqff8erH+L0nL2C1afA5D11rjFB8VDNN
wMExusaAbvsIZaTTgS2DwW1CArh6W+e1qdzlAITvkiApgYD7U5lcqVQdFZ0YFiyLKe/IeC+IFtvN
cTgTv0kS6f97FXVr3koHwAZzL/5t4z0XpY6rcVXBb1dInSveIQPOOHSjBj0us1vSYzdAxlJgRIEf
YppqJ+cegbj8EwnZAo7g+o7xKK94eEopcABcPhICSjZef7LsJxp1dioFo3JmVAdG+Ddz6hC3vdA0
AmwSpbp4LvCAGdiY28YoboQLAeIAaA7KLB49UDylrrypCGozjgeH/lP2tRwwE6IlzVzJv8v7UFcD
oZVHzRUmbcGToQ2c7zjV15q7RHwfSN6RseS9hQvtF3anNeIXegW+R+f8BKuLKzmbRbeKECD6xb3j
pSEFvcjc7CNcmS1u4cOxYx+Gynej9UJRW3XE2Sa5/Nad79U04LqW5uBEDwwEka+VDzJtiza+5aL8
aqSvv+UrY/vSxooT5Hvem3vQEbI6Id1r1k5tGQSE5FrSwKr+7mSzvxfFLYLP+k7X2iiPisrei8lV
aEwKip4/CfQhml5fOKfEh4tGGd3jicCAPeod/fAaDx04MgrbLEcaQatCYqXhdkGi4wK/6be0mqNT
d97jgh5CTNioJzXE2JrAnIXf7jgAP9ZBehh40vYnasX1fTervRpuq+uE2v+kQU22P+GX23C3XQrU
xQPlYuIAUKhk7vJMm+qFNfvoc644fz0QGXjq2Z86Ql8gEdlXwaH/ldouQztLG8VH/k4vehP1o/1M
aI/hhc2kuYrq4jdF2l0j7DLP0dlZHi4zz8xynWmM/YHqmXTwL0G3hTWo9hOyrs46ewe/EEvu1hNK
QkKvo+eQIwJBFeS96M5I1TzQAbvIXRuyQEcdtwKxZ9UpEKX237Z/1ahvrgWcWJG7awLh17g2AFkI
s+oUcDGjJT4nra4bsPuxmqiKAJ0oD37h9Co2U0585H/S+f6bBfxNbok0EVBLmBsOdpV3ai8IZCFm
crheTF0OOQA4rY8i07iPZihovrEVxyupcj3jhpCOWQ9QyCOniZkhNaxGyz9D/EkgPoyIK96fseys
cRW4GMsrfYsPgLK3x+YBKT5NKGczxjNaY20RbJRn09z+IIB8Y/bIZSVm2m9AP+DYRwJs3dlHE4xy
pp6jzj8obrKPanmeIiI4B0tWpZwda/XFie4tj2Wv0VapRgc/jP1ea7SjpsS536WNAXquT843bNoZ
j6XJ6d68DiMkjoq9Zc4jfBMncUGvukG+QKfCspA7PGyuXhnsMgMAwvc/5eswYnEKWdqV7lHRNv5T
NH53A0JoU/taGtYV2wI9Gmc3x9l8z1us65vbnDpMOveFE/T4Eg44uS1ZdSN38aAe1r1k3Bk8c7OL
UCXpP200Ltxoy4PZn+1xcye44yj4Wu4asN0TUJjLz5XqNYHeWmp7hF0gsqpr3xANlwpi8pVRuA5Q
rvUFUWA3hLlpDhbSFFDgU/P0BhRn6b/hL+KRq4+W0MxqPpXtpy57xaqFeOLZQgc1/ZN7ZUL3ufvJ
3s/ZuR2oXJK43lfoHHZphoaHvvTA55PRXtgLVPpA532f82zkioDU1kd5nT3B0vUVy74TDmpzEpS6
dwK91m9ThTqOgmBnEg7O64jYnKLHBhF9zZ+FKgr0Pa74kt8nopzipb4x8EHhsnmLDJtOngtYLi9R
hmblxz6m5Dg5fwetwG43F4yHJ+rFS+gJ6acaZM/OXRvblasTOwT/YrvbXufqh8bAUU8/SN2mXRN/
e2gzpAQiY6nvxahpt+ilmAvT7lDEAwR5ehaL2C6+KrzLc7IxHL8KixA+jqPa6HX1biOaV/8vqKiT
z28mhxDwX0T79MvKPCu4jIzGU1aTxGfQB5Fxh1815rSqhyYMaji9rmxYCJClYYBz+4nM4jZiiPkQ
Q7w5+LCVqza0Ot0UzRWprC060ObTnNb7CFnlpcnCAF04hstqcFhluCopIp3zO3Q2o0hxFHhqE7bo
AguGf8WUsauzOIVT5x0D7o6vEgmadja5bqqqTcImtB6ORyHtkx8bLk0xSlJQog3mKG/4zebSfhx1
dyxCc+WzIt5c24kKiuwDOLqdKAl5+K/I7aurOumewqmAKG5rrbdlMuGqhY2LYNsK5SMMnRVVwLc9
uXDuIVhiRIcdw7Gbdz9iqFB28pQ1PIJezd+kebe4x82hVOKZwd0yFCK6OpSoCEV19PBF5RH/ZreE
j952nM6XvFhhVYBxPhiQS/D7pUqNsVnaNPd1kEqBe06GTsAbU0U7gwEW2eLHQ9o3BI2KiSf2f6Z9
c6o1QVk2PvE8MwWYimNdMECn47wf02YMVP4gQQWQ9BjFUPT5ChpWN92MTbBrqNOXiDXNdS3Bailx
EPOzWpoueP6Rf+vm7C8HwJVyTnij6oLDK2LT8ufr7vGrbkv+OAfal1j+tBtaq6nGTLXZMtIciH9C
pIewF2H+UddjdNWXrQ1IsgaqZj1F7kmvlZmOB4zuHemv8EGxA8Sl8C3NuOc0+OPoJ5wMedlw1o36
CLbo/kTjTTBzBhsm/c49nxPnk1OBv3pU24B+n0QAMy4VLKa06KntrcDpYcOdfUFx6eWt1JP+sXT4
GjdfkzvYuCwyPz9+cEP7prL1PXYtRYr7Q1vQgXJJ8S04OMN351FZkyylwS5HMFtk1yiQjlzPzo3l
eBnIS7i6H4aoxlnGP52GADDH2ehET8t1aWCn8EqxiBZ2oPzv2EZidwEwNspoJ7UWCyQJFog79Dpe
rmvQLo+nAip7rpyP8dyNO0IOunJ4n4k8PNDshrp7uNt3TmpDMFKq2FTAixb19eyQvTmep03nLz/L
JIM6XSQOG3EI5Tl0OJxQr7sxCePF/w3ALJO6Y2bPcJMA0Yg3Ym/5xljgAZslIdRgc7I9h1fMb/FO
22GmTZBc+VGCcIyycbcSSAYc88qh+svn5hHp3Cn1y3FNn9ru1KYsfUBr53rBbxFcoc9f0aYD92TU
G4Mt/fcEf5/+qagR2pOVctCNjQE0x003MD1ysT6IDd76/RwldPGrNyGBA7OyFg+83INdyVvIlwL7
a7pBAQWVihkVXPgsH1OGtzeWL/uWM/iDob/O1rZIdcEHZpGHqh7Kh09LAcNbMZWMega/iZM2kRsE
Zx0d1MVha09q1GQo/NiwQYHY/OCUf/T/eTyDxnRCw0FG64SSOrgLmGVXYH8gF0DulbQwFv2DhE5C
VPzlennsuy10qTw/sAvBbr/YoT9Kflu51c8vHXVpH6yRQnpECOQExigodTJjXyJLx+5Hu2hLlBly
S2b8AcIaidSVAkdmmJds8JtVtxM15wfu2tmSRm4ywDCtdpc3Jsb+PjVUhQy/PeoiAwzaPvL/ShCk
h+vfaKLhlQuZvvMjv3JLJ1hD9uagv36TEUfBKuxvER75hz0mkZI0Uz8MmjHyIeaaJD+1xkE2Afuq
CcnqXSe1b9wpGLzm4vkKXD64GOwaNq9Yw0lIpplsWvNA07TdiCOS00rEhYxNCJATVKSptiaBhALu
VYNAYgIO9duxx8ARNB7bUGh6nKim5hv3VEzbdePEgudfHKVFKHjbCa2NAKhYiXshQIzlYieGElKx
aYTufnfjKB+8x0nGYvcRpa84Zs8jmuw4XHjZtKhm7ukKeopNkXZlHS+RtsHVNS3K04Fm+wLq8AtT
8VteodRnp5Slv2URrojOYkXh7FOqebwzCtNW9zPlvla1zpGyyi5W13fJ+AGdBN/QMsn1E8KqYJwn
Y2WNid1t678v6K26ROo0b+SHuly9Aajd12kxZOyytRg6QA7S2bwK4lau08BwBwm2jfeGCILTibWo
jdOjO6z6rXaxL9qu9Wtax1+vLLYoQV3IEjgByHlIQuZ/S4NS/PxuvsEr2N3EahANfzYJx85BoXEZ
7i//A2e9tZrZlU6C3Gg1r5z2Lm85jIrEa0Yta3lMGXxEoFs8XHXhwWOElKwsv4iEwpC0ySwHjVVC
caLqVyaOEnNySX/VTCZZOON2uuAnMcwvOHy+fqYELWUplzCu1FqacoRv8nm/EV8KU6D4MpsPRJRk
+Ldd5OxNLq5Vvlsy/HXmSj8aTzg+F995P8R7QxzOgfnQqE3NiVJ2tTFcMIsmM87Hx4AYgF7Sw39y
MVqBQGYL211ZJjyYWba4sGo8Qr3yFDbDG+erzvOfPnha1uFaO60wJ0tLZnPH9uOy9BDzuH7jOHVs
krnefnZQszuTjslZlBGUqhg60ibGIWfpKZptHuLaee6EpLGupavNq0gMW3HH79T0YvqmLh6Meom8
AIO692vfte5xlczjBOHptxrsXa4WO8702ihokbpKs282SNFpp0OF1pocZaf91y1kgg6Xugv/y3h2
PHpLrLeDxWhK40wFebGNNh97anuX1XH5dpZUDRI7TZGqGmjNQGgw6HTRpzDaGVbmAMfcrgdTIA3H
1l/q5ZykaQfYAJd83w7BcXosE+nUn7L1RiHOpPbOlC5TYioe3VAedcE4xMdGXMp8McpsjbIOJJCv
y/QqVo8ExV/6eX8TjBEjs0vUbOrvnahovnI15dSo6N5htxZeEV5Zr4NR9pBEaYmEDyzzuIiOB2Cv
6Rn2Nxq8a8S9Jm9K0oo7HQEixVWlAB9JVHH5NWZzDVuVr0sXkv4b/FJB2N4gEuvNwzg0gnBL0xFo
2e8+yziVM30SHSp4g8Pt5cq6q71OXffmPUWRM2aSX4oEWBJsb3hpOUEwZ2sdiCYyhzJg3YPDVPdJ
WOGen20Ex4/GYMOu+k5Oz9/uhWSVca1fIkJRy3hZjgULP+B76DcOn1iFfFWBL+fzhvGnh0uFzf8Q
h3iJNyvP+Cgj65aGcs/XKgGmuOPscvGT5Lsf90BnwVsVN2bmH/eQ5aF541ftMftD5of6wuolP9EB
/YxHhuLWY7gpLLE17o5qguuumr67Yn0tonjzTihd11NIt6Rtp05vqS4s1VeNdZU+WVkhvHxaY1HE
nDgWtIq+FSEoGNX6dLT8KP7FQHmqwu8XYtG6raI+J2cbuA2hZsyb4XFpj2kO9IqPbono01TeCbwm
vjxZQgxnPZt+KXz61SyswotLrWWKhws/WdoGfdWhk/p7HIZu7dzOFmMw3Ypnc4TlOucCYswjZIyn
afKSGELxaDBSFlBh8gIIW8DI2P5Vom0bobsmgmjsaZM0QCWI3nZwMJ126rDnwiA2dIWBKS9pwVVp
MeHmIKSxrvA8MrKCgCCVfy8Y3dWJTi8gShlLfiFHcwTSQDtKOuIiTHjbPzNMf8MxMX1G7/0Fasds
aXxkQ1iiDqh8W0Xp00b+AxQvTz0OihtYkqDVrNd4XlyuHejY1WTB56B7U3LKMH8fAYrOXoJfaTBL
qp6prmE47XDqgkxk6EW1aY607jjyqUJ0e1jh1+EucM2gNfsZOFG6u3kmvwaTXH0LoEC0QJLXkHKg
sRcha18q5ESt5ygug5HRK3qTEccIqbcjloeVReIKtA+k/xR0IhF8g7dzxvokPKcx3krbrX90laqn
JWd+E3EbEBFA1oRhC7M/1E/uEBpiqjawlVfyVqs/DxdSHq1tRv/7T4uJCsB4uGtA0JiN+owwpUb0
+RKMftQFKevyAwdFKaQzyMdR1UcfS1rHZRQpLHrjruDS+8Cgi0aib+X8G+0O4UPcmfWvqNHh6GOd
Q+H1vbN/p71OYkOHZV5gpPOASXlID9OiQknCQIjyuLNVBrcyhxMpwbqGwpnK2+v6pCQY/Ko9Ol+2
XLbjDbLUGfUVK0zYWOIFcdIHnNx9sJrU1Cym2VuVPdvkrx337wuxCCgWHeYBmEljlZAuy8UlQ3ux
A9FN1XqJS3NwmTVco2mIl0sDk5vnrcwYECvwWeknw8zhICnIROHD/aSd1sKGvEFSXQjZ/o7dAT5l
Kf02ST084EwvWmLeP/O7JbgnilItt/n8SQ4ofgq9rEf/69HHhksTLX3WDUiC3YaKnGzipYnbGAsB
wr0aWMlFI9nc5KsbHCQEl7dew454pUwtS/lIsfT0KLRbZIWIkI+48dZrDHE01ztvo6VO3jjZdJVH
aMXHBrlGG4jHGAeIrVTYKCBY/fxrGRvSIUx49Wnd7BUNLVdoDu5c3LtoKCtV2hObEmut9cyrdiOI
4jFQRWhR/Y1pFutGJ1RFSeD3ueWQbttMgr002fXRKPC8C00sC4S2HzDQ2X96PKW4WGfINp4J8HTd
Rqgnclr51B54AtJQPrbO01ATGQywdkQa/PWkRXbbLIbAIplRNxdqPCWmOFc93GYfESjus+XREo9u
E5PIYnh5/FXQFeOJeP6bEhvIcLYlWT/dcqw+aE05o03tUNNTNATM/S6f2GryA/ZexDYDkE+ZVFG7
elZFngIyrdibJpbw/oUd8h0OhnQeZOlXMlypeS4jdiKUvxF+vH3eNx3JgNRI3a37LaoaHKUXeC+R
EKdHCY3I3iTjEyTdQ5oQvFsVh1Rb6cx0u0j3Ak1u2C69lBC5GknTTQltfk+izsaboJWPkQw6PRz0
m2ldQKW+BhP8cqo12fTov016uZLObP4bBQCQAQiXKVoqsEZjKYMxqfrqk6qs/x+kjofY0xhII1rt
SJAYLqh9lgbz327G34RG3zDIwk2MGw9yKepWf9c5ZMBTcIvFK65QabRLyz1/+EivdAs88sd6QlWk
KiwXpNsIRsf2EbEjK73ln5KNDIIJd545Vfv9PvA15y5I7dQayGquJjrVRU/cbRQGvyMNMfXyBZGJ
HH72ho4lGutXdbhZMAyCcX20eNbh5wvd+5IDN7aNpECulRF45sxXut75jgrbNIfPQmf9rY0csr9x
Q+geNwWfrg1zyN5Gybkw9MAVjCcNLrd0crxRCPOBLtXGb9MmyMT36jjhwgXP1X+8UyZhIkwBmxin
31rd4pfIxC60gGt5Qk+4DLfD60gvyZ9pM1NuIYkNzCz7MUSXFCEJWdvrS7s8zaCofJ6aMb2c2a+H
OMsuS81NZ3jBVYzGneEY3YYvwQWkZ6EHsbxhFWtQ1FeuIKgxeEXkIeaMdR/EkNiNd7f1jZ2yAl9U
pcqJ+MfbAVVp6scywtsrb2aHVWGQYlpTmLP5l00KyyqvMh39nBZW+dEL3Hsv/FgXPAvZSWdd16ym
6Z93A+ED5TEfIHlYXePHZHBA1galyAiSdC+Wnp9+FK6EVR98NdpfkLQ361lwAdlXGIn+TwhVg1mr
6P36OPzXrJJJNQg9q0CGhzCIwh+Jax1kit3hkUK8xnurmlNVA7+LVB1wK9OfOAFANDKyZ3f1JBkG
VdDxkFFfnRVrzQMKZGCt04DcIHE3MrL1p8a1kTBdX1/XxMAj6fHejEG9/UGAu/BhQj+yqr7dtpFx
cEU3EVzRyPWHhA3gJz5JFXgMS28gnMUgefCmi5D0+esu7tKGG1NkxOWnugrQ1cVx/s7Sd2qSX8II
HOQdYqQcXfGJlSG0xLlGJsyDiRY1PneXEKbgzjFLiGUqz+IpZZ+fB1peaN1bLMarNoZ3XEHUQ83g
AYusf1vzgDT6rJjZnE8PfY+r68gkgJcLo/S6Y2dOCfofDX8YnRFmPkHpZQolEb8vn+JuQVaFbkRd
YrUY1K3+N6ijEvTvSAjWwXnUNpctsjZXazB7bPQex+7TAk3Y2Bx3tQE3B+6DPKpjl4enBJX3kbL+
IolIvDMX5OMY42cYk0KpKVNiB0LXDdeJ2qT0Fu1qcNu3pGm+KBNeCdWusl/q5eyClcJFBFc/MQit
m1Wx8Ovh21d8MHNAKo2oz6t9TrEURDgwzTfWE9vKoJ+NJXeHCwRBPHkJg5h6EDXJB7CtYBRzht+F
RO30dUQbgFgIrVxazWOBpKgHfjHyu/NMuAc43t20jKBNcHYuunBPPAv8RrmYHxLEBTxMO2lews2z
R6dniXg+OetQfh02lVyKEO2p5V4ct8fvpMsZ+ZDkBzgjz1djjLmYaoPDjqU7K95n3J7Vk9kKgjpF
hBQRvnTuvuGeI8/pRcOmwO1k5mS8OofsQMk09rwyI/gOUpbuChZY5KASTgqnG+bcp3wW0RxKdNP1
8jOvNi7g61HzIdU8QILjwJaemXiMamgw/RKRYnKn3SeatlZvSxPY4s4yotW6TNt0epbqlqMk83yo
Vsaa5f10tIHnQh4783bF+rCtBbBabe4QvUuYXknLRKZBTVyE43xo/nxVZrPpmcUiI08zP6wsRP7y
1kuUfSrCHCR08FOah8gAPCcvOjlEDt2Uvj+Mlvrci+J2zawUeChQd6xqglrmadz5ljifWHWzHCt/
d8VRjUhHxzrKUT5Hu0MymaJ8+A5qzVB2F6bdmQG8v1MfTWVeM/RPRMgnuFvb0evYTPqB4SZvmz15
n7O2zsQ2P1gBEjfdOS3YUMPSTD3yQ0hifuTXq4oPwgtu9Yx3sG6Skby8WupzSFLpcc/n9ty4x8ZC
nvmga7QnT4+BAaUEAVeWUf6tLasmx8hZE/R4re98gq20FwqN5ccPr9U9/JSbRSg14W0ciDjpf+90
FXGaQBa7tDedMaEClH+eQ+BIB/d1djll5rzlDXxtlVKZhqoDovzggVx2g2aHZ4LBvlrZS7IksZwl
7V1VCbVKWC4bswPpEDdr51QfLf6X1y3UQpnDfkOu97WwAsSyFs7AKyDAvxUO/bJG6GDGw4t+lfvF
fULE4rVXJA1NA+JBYXCSAbMByBq/sFmMT2RerXtTkNLirs6Sj7uELj1k/kqrGnBWOIGGNh/7oV8S
PFlP1AzjloIuzBq3T1QV2At6lE7EHneU+0KetklgN6wQREA5B2mDUBsq/SmMLjBGeA9e36GiQ8NL
ikM0RIOvrARlP+Ma8NCojrcY2WxKLgQxz7OC84WHij1v9JG2Lf7kepYyWmRhKEalgaq/LNnZXYZs
93WMIxyf/Kj/YezpnNd+akP4ccZyJmO58OYB01KjKd0kHGlXHprYCgR3GiKOELxlPzSNBsXDqsAE
gK7kPmuOoQcoafw2IjMW7q/n5v3XSuOZdrREPafxiWCp8OuFqZqHpLtIes3MYXgmLEM2vrGlCQhK
zOzUdg4i2GtcRM+urM0xmJVZlbYcHwmvYSNNgGpczvH1RT/a5YLWaJ3rfEyhL8Km4YSUNZnNu11H
vUNCee4vXDdcmL//6RSE2Bm/6Pa4VPMHSUXdxprnTkscL9OD49kbpFA/l3lzePRMQyZrXQYd0jt5
DfY+QeIi6nUCpwzLuX/Bhc16hCFHiihq+h2AFO/cOo2kA+R8yWbif145ShBCdnDZe9j/jV7IT3AP
euf0EeMevxw5h3t13pGx81jmwpzB4whunbJlXLs5fKXH4Joa9tioXjVPcpp+Q/UtVm4VcCS4ek11
mUD+GhN4dAqQIXty+yo0Gf/3th2hI99kOoWIqNyT8c3nU0WBZTqezKFrvOPnyYQ1dvppeL0ZWd2f
djBMS/B7SWWHDZoWGGQQxmf3rt1PnkigUcf5r0VHfOksPfC05fT7bY077P9DFHMM6St6tMoW215B
ccLVY4juD0eYJoJScxLZDBnO903LLxQg3qrBszSvNX5i9fpUZMFH7NPkpODlFRP6A/zkS10/w6xP
fqO0HklLijim0VV+N+HlMR0X1laIBcNdX43nvdiDMuwqLbnETKidQYJ+1mQ9xtRP9kt4FjzmKWOJ
0XG1zYKC0tNbmq9Q3nLyPRUPFpUvsuTGxJMBhFODNqO5Klsv4sGXIgl1kUqubXeSB94+QFtbrL5u
si8MSCtTNifrpA7i0FTSMu1UeIAE2PWoqiNov4rxWjxRo4IB3Wa/5Av4JSVdGwuwGjPTwWWDNZc9
gHvrOwbZdzLRBWsnmFohlU6JzdxgAXyJhalGn82cwYqnoV353YoEgNL37mWOlvfaTYKyfyT631yT
OA3KwY/7LeviQ/wBetzjdo1eU6uNgPE2fJGJ7ABdIy1LH5JRSZvzqFEoypjGQbcrOlWD2ArqzmOl
azM45Ok6I+3Ddy+gjUf6QY7yhXftgJeQe7tEVZVLji7Mypg8ry9o4cC8KRQLec9IZzf1ncBOjB5T
Ec5f9uS1W/0BISObugbixGDFswsrYxLb3XMDilnG/MT4q5JFgtdJQcV8a7rfMUKM15Y4G7fAWWWv
P532rqfwNmwKYLvO4l7x5rj9OoZvM2tZiYqXZwFUYrkNHt6NvIi7dJxDZTJ6i+zcamAMVrtwdVcN
MheXqIJ1mdH1GYRLDvNFpinoQ6GitUQ94Z/L55v33XCtRetZL4EU2W/38E1umpiSYu5Pq89Xwdkh
HGWUTzUViRsXqnI/ktFdejRF5X+HM6lD3kUrAfz/7ZS6dmq8HAXrsG8MWSMaAAlvrTQAec62Zftf
LTkgkRbXO2tSp3d8ZY4ju2KWKCYbmTfcaT3Ksu5bo/Abot7glgu34QY0gXZSfK2bfiAw/lloIles
ERpxyr8aUrq2FNjXoBt10c3hJw8Nd2cR3P8zJX88Iqa7ulqcK+SZcCM6xuE4lVw/cOY2AgjqSNcO
iEswcT0c4Z2N58f9xpdPsxtlaFQftFQrGlH6Vv9QsJtg0oTPdbjM5EcH2EwBPH/hYzUwZ12PrEL4
ukGsNtkRwbt4vJCQzQaC1oXcaxI6InPzndkVyKpUaOjmnsYn4b4Di/OLjH/n+M3IxYaqP0nALUc9
j9RBSNVULzkiJ6tiRD+EBO/WLal4uv1IZ0eDT5kxxNHLaFLJjW0h7Vi8pAiZrsxl/Ie0pek6WsOU
yJi/6Q3uGY691HLoatRaXsSJ5q+eowX3iAghHlqDqYcnNpUD2YvyEGVeBraUVd0TTnyvmbdwgtSn
kBLcUP7MNy3gBv4rAwyzOzlh8YhXJd4fKmWnVmQwbtvkeMvMfsffbxmIZW6GdIT9L6ChU94W4j8Q
wI9Y+YsHzJtPPPEaXsmjbtIgtY49pi7w/P4vYHUw2o9qP33hjNfRTOfMsqgOc8GvZPTZzpsSt89H
cpqAKjyjlKTLtq3LctR/VDTodE09nZKfYX3KkjwB5JY7xWaiwFDkUs/h4FLIvokQozqsi3Pt1VYr
hXYvM/4/uRmK3IYwWvUzU4fNh7Q8LnD6Z+fo2fdfhywhO27EPPD8+tepzWdz7tDoZlMYSrCzz4dI
PtBIV56SRs6nkFdy9N2hGsTRNStOMP5f4MbpCY+AbQ8c+FQa9eV3K+iVsEY4Y3JvTYUM/hI06p/z
Mgo+CK5zVs3nNXfAUQc+xlM5lK5ZzV5hmTcThhUAT2F+/t7suN/vV8wNQ+uS0tpbLMeE7B1v4PUa
mJxGI8C6PwYFMvc8Stuez4pDygJn392fZcx2sjrGf/0KGG7jGw8z/Ts7RIArKnvLTiF+42ny6hiz
DRHdk5AHCakLQm/ZuHc+5/QA9CTBWPseA5Bi9QR4qz0cf8+LkJgQo2dEOdWIsBTdVQyfpRQer9XA
nE8HxRlejJmEGRPnAzVz4uVbNxS8ULSbYE4H8UPoNjS+0Wx181CwXJFvqbCwpC8wEppqfnc2C+tb
cB/atnYPZVkfGYFlL21zM6HZrLsWQ1RCnApnsFBadbgsA1xu8fCxMesHKtk5a3KVeD1RgUZSU11K
lAzFRCQD4he/uHnjjh89Cw1y+psRfXisipcVmWv+LCDORVKtMGDbejNdxAHdHhHI1pWPYfm2mAYx
hhv1+uvsNijb3yRXiUTYKuTkPAmABuPyYdLIJsGEZaDynXOIvFaeCcwLYQUD72GXbXE5EpBgrugR
RetQy6HKQuHUlm0Xpz81GiQI1fwNfyKlg3yqHvr5GJFUsOdLYgucHlF4EU4MhcRWs/uQXkxb0qAb
GEukw0lUHtd5sP+7TW3U4qpGEnt1WnDPo3dWweBOJD2Cc/oIKLSY4z8Pz6NMHorTXerOADCF4lL6
hohgJf48oriLY7iT9tewKp1d6cWg5Yt9sQI3NdP/r+y92+KX1HhIx1F5rrXMNVCv6zJWiUnkQ3pi
p62rTJrCsOTts695aHTgbOIIBPDAxsnOgHaiyFtU/14C48qm3q4In0QQLABlps5z2yPwu7Iv3PYO
LON9316uPQi3b7/xk2apDdGyU5WadhCic2WOlGmchTuFc13vtBPHGk8WjCCpaXEHy2iL7d7c6jfC
lglW+Ehncf9dAxhYMgIQSPaUK6IYH8KwXdX9kMd6CJPHYipnJxLpaKXSF3+nHTo/+Yz57av7FX02
OBG2pYTmb110WEAbV3h/fGcB5hJ8slJeyLya1DeOUFmaSl0+QiexVfByLSF6JXU0qJO71F1P1xAo
fL12qlTSdxnhTfS8Zlp/EINdq2TUHPUUrueVYyA3FRrkLfZGqonCcD69tJHVPVuXGnmPu8LYSvwc
eckUd1HsTrZzQOm0XuC2p5Z6J1JHdEWQBTZpBR/dn/li+q4uotoemzRTalWJr3wzjFrNY4n9XjMK
x+ylWrw/sysYlI2pP6raoWwPdOJdm2nwbvTqxDzfsIZ5lz39aBknjoY6SlJuKn/rkoL4EFqvSCez
SXpJVW3PXW9qXAHU417z+cLlkUnEh7E2671VsZDMlKUKVqRIoHwYpGezqTACpty53NgwwYdFkipi
BL5wSD/k+kM4MUTf2cAfStOplZUdVAKWQiteq6l1rdaCE6tk830kRWrlHQQ5Qocfbdqe0F8mukD7
iAQCS6y0NxfPKDsGzU2jIIATAX9+5lC6pPQBCisesYWKa/P4BPT5RogGpDuBkKk+qbqyw9TMJNX9
Hp/gbX7EZbDVNH6Cxlqz7RaW65qnkEN2f+X2cmcZFmg0D1ZVKKN9rKt7MsFTzWs6HylmW8RHJRm7
+sYlXZ6innwIGxGQ+r/BAPzjqJD1ZvQuhydiZMbLTVViW6HHOXwm/S6ZRJbvoDoI0W1uhJev4UJG
KZqAj4AY9E1vbDmdXwBZhC/YaYvNGvfKnTW5ck+2f5MJINEya9IyCcgFtIEiSUCf4GS3QxgDB2EU
akZqVuFNSLDyB8jX3cC3RyC3jDDFXivwP9G7amj0YamLfQIr8HvtAhSykOXT2aWWLBxgc2fSSxZU
ctvhp6eovapWSYl4rMjqg3oOQrKLejw6MK/qIrKj/Xc0ICzkGaPUDJKyBYOQ05Gl71XBcKiH2jHd
bmlO1prbC5Mf+giSAXdbSXiH61BhAbYjFkpDXhg1CA5QJJmQP2tfIsqVUKW0Q0/C6YvDzyuXydhO
Uxnjq8I9HDLItwu9CZ5txnEHqsPq0/2ZYRzWFuGmNxf0HHXd8DjIeb8pmmd42T1Mh1bMUzB6Sn6+
EjEVBR1dgTYJVGW/9WWlqmqPXseBFrMLeSm45qvJ/khRygmcnLcl5O6JyD2J3hRUDMc22JUa7+qH
lsf6nCUetadb9syTcMbLsYUlObitgG2NiYjPjuLaXWuXe/HbO1CiOBlW48AR73ySvozP9WTNk98Q
X+2YcgtjM+cC3mvFPqUBNtmnkwZWxIHQdmwKmm51aCdaFTkIc+twa96oZiC/T/iXgdLZ/tpk0aBT
taNHjWKY8zwlan2ryz//Oz5OFjxRMH3PsokBB2g9aodXJYe5fA/Bv15ULLrVKLaHbm3tmWmJF1mZ
0zSUKvCV3MGSkGRouo/i1bXFbYIvvQQarIfnq+0Y3lgjuD5c3ngDqpIL1nltXm9CkhcSqxRhIbOY
BW9s1pDed1FTofJVlSHwO96L8SIg50HSd4TJz67MM/DIoGzTZxDBjVmrOz1JjUA7ZLOTrHrKV4T5
I5K4IDi/rccu10a2dSyiguXmxwKPxxnDW0DWr/AVuqrdzPaZhqn8bgLzpLTfr3E2iQMSvWkWtsvg
ZqCetROB6Tfox7XFwxofsDX8yD6rZjwvEz/AkguT3NeNZ5eHfqtwgEjAcsAqoYXDiZKbx7Nv+NHt
p3+vpkqKDu6t4YkGzwcN7Xg+Z44qzQdX46XispCsFOiH+PpOVXwprr1o4COi16dDWhd6URBIYhpQ
lwImK/4mHWKhQ86idRMU5/yzEwxzFG48Cxf1eI8CmnXTP49/E1iEgISqoLBzA4fLTZO5pwiiZBXb
DF5umIdY3d32wy4AHZ+KZO6yEbfRP629diIZTI9MWFHPARCZU/D4j+MxphrcLW4q2ib4H7vDRRj4
quBfxm1gS7dY5eC3gofcbgAtDSOlwhPsi5zO4OPajwD9DMA29SpJgcLTcWYWurBe5IZdw+kwEr4J
XFv1F5oLjx7sOIbjkPN2CZntA/nK9dWlcljv03Ds1iCsk2UKR6cZRolaUL9vXjAbUPFSg1gUmgqB
3TowRJd/4kK7sDi73TH3HZr/rCMilGKMUdeGl71gETyxjPP532um6/BKYmIpYoEq7Rn21CFpGtuZ
PyYkW1GG/XLsZ3aVY5ZgwMdEdrqSP4fFubuJR1M+RQSMWq2JkViq5uSuQamX7VK0/P7kHZ7xsHjo
mT3NUaiVbwEs8bo3goRBiMtIJV07SwzVxY/5TzCyQGo65HWKLmhMFS6XjZHizHgYKr5iP96dsDeB
WN/Q0m+NpSM7tZOUMy3Lwz7rb9mtQfCSWed7SfykRR+H5BsfCTNZlJEr6sNzigseOe+7d0D+H4YI
WwUXOUMSedUPyev1KuOIwLjoCkKG70J0nC4OTBCpV594Le3o3Emt39F+pnFPIE/nVGMhAmJNpVb5
tUEBsmsYokZqi/B+xez7dE5xhcQZvD8wOjz1e8fuOH/vfiMMSZtTBFCZnWFeoWiFAB5rTsq3L7/3
lBOQHZ3VKSlsPUL2dgKIHIbDHF8EP0WyA/67dgHbX1riKdZQS0U9pKo4yDAfpsNRJBKw2sut916m
nmH+PZ74QD3Kc9xPVAL2DIQu3p+93JBdttMA/XmCm68Mt44+Ki+ACsUrXEmGp+y/VrMG3R9PdDjE
1DPWDd7Yq8hmQRHo8+IiUnAgQADSpjtEoler10t6vXME8V2TRlw7xnlx3X5wlHOO8d4cUk/3HHnn
7NsFBF9a7NjGqvfyBbgux15Bzh8AXSTd8/I0P4NHhNsh8GopM9YCtnxR4fF7LJbC4XZClJtSfcdy
9DapmnCiOEVx5qWDhIn2p1jDZ+0m5YRVMmzlakCMemNrb7fpFsIC6O7JSmXMNskb7aTfJi5ZhJV7
9hXj4njM+6JTJXO7e8V12MCM99VU5joyp0JJ8ZyAtoulgisb2qtwSj+EDNTcp5HkTvyO6pQq0zR3
SmENDsdqPwyIk417rhDqZcV4b6IXGopBWj9Mw+W3BJUWlUW+nvLSsT/QydtAM25BzevomW7js4LI
Q3FCjUDneU/0GpYlGX9saYjLslnv0ReuSZAdei/tJslzyAlNxFq+yS1eNx+/kQbuWlsfJNDqQIbL
0nqbNfvZkDXljV67dZ8IkYvMAl0ntSziFH7ngDkT+iaUfvUk1UvcSw2ZZD0sJzXI9iogU2XaxXsa
MlhyI7rP+tNIfxWhO2os7cQyI4FF7ROSKmrDf5PfbwAT41QaTuRtQsnkLxAAcqd128yzP2WpXDmr
SzrUq2dK2qbtoj4ztmuTfNH8Ql5nPolRFQ2a2kD2u2VwDcz+q/TYY0EQISkacCyDmk+Gty2Wu7ne
lKXrE5gtCjwJNU3RKjhtENjOLEff7EEE7tez1aZVdlkvL94t9ST11jGlsxpgna52D0CEz0IXAptu
hk8rteuGTlujJUjBIvb3Y6BGCWoE0fnAiIow165q476YQ06BZsM8ZpkNIoAEdnesKQyjYHIXSD+6
5rlahRUe35tGFuR11BexKrCNhv294d8dVm7cjxjZiDIygHnd3chpSqYthDBz2r3CO/shPA/on1Ye
htDKt14h3uJnlcrM1M0uq0MUxYaWcLkcNqcgXf2v/xYAr49MjoafajrRfK+Xgr8ujO+G9rFtjEwX
3YphRcVzvNPbQSaUClWg13p7wntpaPSZebCh6cX0qaUWPVXcitwsFHM8F/m7rokZy7n03XhvvKuP
QcbTOjDT4jN+yCB43Hb17vsquK7EfsO1nSsBS5ss1mSHyO0Aowqb5ixf8jQCgJjlAFk50/87ujJd
B2mtJ5CWYz8/LsgbeCv09Gg+7pnZb8uq3o3tKcem+W7XZoDoh+5EMCJTC+HG/xfrYcVWGL1iTIZW
8wo02joy1osZSVF6nWx4P2/xcTJ5l9rDLdZJisg27dVY6yolSD3OmYu3cqlx01mZbvIe4COtBGfj
T567t89y379Gta/LmYjYf8SBdYsEWSCH/5zyaDnJRo/c2JY6NTJJlisMl0SsOA7eSnbrZMPwW8VI
XyJrIuCX4tlT194wM1OySpx3Q8UXPRw7Bv5c9G66Jywl0qsVR7PEShCBPyqTAAKT2TCaO6VPtbFb
payxwslqiD7McQiElZKi4jAap0S0LeJwDGctom8PMQMu4v+Y6rmdTfw1MffVr3bORNV2B0d9/ni7
a2ANSgUqH2aZK6CZyrTqkb8CQjTuEey6W+PXumGk45TaGDbSN5+PVMZ2vW6CfivWBxjWmLiQ2NLK
Rt6J3NlLSvSfUkxDtCQ/pUd4XqxpiqOb3g1Qg4JxN6rspuVXnwWYSZJoRZZzs/2RdBwg2LJxIEYc
0qiZqjRxheH3r8GwRz9qt7KGNwKG/irafKdYmtjxnWska+3vqOF2L8Z7jjmVMvA5dFlOE6KWD83m
yejhy5aJVSXyVGYmtDkpI38lOLSb9pMe1bDB8E5vsx7zoYPq2FQmqegkmi3ho0rRgwrTTTfhUpxS
N7jd80zBlGsQqLMTuO+IeTZ30VIiq/ejbwRtFc0SfjIUd7PqX9jnaH1lmWoFkvdrLZiGByMm+Qcy
9XfQJ8mHtk9QB5XAwRNbKcJoP8uOF7WOs8Y5nQap4tFp60aepRQMm9xZQlwen41nS429aaW8xvO0
6L+9F2ZAUVsRucsK5fpgFwNAM7YV7Qsn9aUAtlukcSgMz8m96zWpKeOcVE5ZoJQPz8+tEB8kQs12
9Y6YCjvRZnk94qKK1CTh07pVpkwfnAKLzq15N2jGLgcIRyiuvxXAXW8qH1HgDobyX3Paq3M5lMgk
RSTP3yBviRmdUHZnS9qHFLguNYNImJDUCEa/NoPILdYCoWZ3zViu3tVP9QsOlShTCCFpK2kvRSM1
lgeKoVqwb+5vzIXBQ0mRl3yQnfIaTslR7cip0OcUJvZtr1ZJXd0p/PX/+9XyZgSvl9PDfiluLM75
fg9bNtoM5DHyAT+ehNI7rpe50wUkuQ9YjfanXkewf7m62zMrNxpGz//BRHyGRwyl55ycT5BaaUFg
FPcfEEYhvS4TgZLeKkRsRNwNQpF114AESFQ3oytWA/jZh2wdMaFOyShY/QTEEmDk9m+hFiJ0Z1NV
jjREPRp0pvbHi1iwh5Xo9GFJtvVCHfY5QSi8FrUoqZUr96lv0iX3wWAr7sovdEDHWEJZgHm+zh9m
ZvmxkpE2f1zq68BLRy2Ix5gBjGqKPiPITtum7mW1fmwgkGdafOnQ7Nxe0GMWae28jY9tQMf/zjcB
NXvqeuoe1RVjNiVvYk1oaO5pN+DCGwpWMMlkIM0Gv4G6tRy5l+vOAeBJsCfKd7Zpm5vGhym3hzcx
7p+/qpFSbP8LVZUG7DpfgdXO04Ov8sorGk4wULt9z39HLy9kzqh2Im0+oVTFZEY0CetuIW8JLBfF
AHJBhdmpoMz5IiuZbDvmg7pZUFTBIJmqPgok+jJGu/itQzrj2wxLbmpIq7w+zYf15mub30ChYg9s
gXhEK55OKW0dCnUnHbIhOdWoBHsvuMiu+/aMAIr+o53zhCgjK2w4vJo/0gIM0gviJTKheZMuJ19j
Hr2rwESMn/YlLCGY7MeZM+Iii3LhW02FCqE9bQdOzDDNgtoAk4/5Wisd+HEaQ8EPILTY0RkdREq8
ZjBHb5cWB+vNn6KmZgOsWzY/OoaKRKPp2JVQqkNulkqV5CICKZCgsKkjFAl2tJs9YPqIvKvrkGyM
vZ2JvNLqUREj8DUhztrp1mn8y9LfZPmDAfbh0Tm0zpFSuF/2U967JQWqvBW3H6QiwStDH9SpzUM+
yW+FPEPD/jyIo0iRhxMTeiUfHFKACN7bBZJyYl+hD9lxMY+KhAA5Fr6w9njtpScvURNRUsMN2aWB
JRvc0FwtP0Ki4S2Fj0wtpvso3cVbGcIRZSOEuRZgn0XvgFeXwlugKJG9UQGZGO6CdN1bzhw0ZVrf
J88ittyAZ19fu+s1N0TLXpg3FaL61Tm5Ofs6RtGIMd/0jPm6mSIPbaQu9R7vcZfHk/OvhJ+qtcLl
dEtktfX0bTM7lTcrjtAiez/O4NJ6ixubcGxNT6zfmIOFRrz9i5CZ4NnT0+q47mSntIM/V5LLkhFg
KXx55TpYEEyU2Hb4b2nVW3rpKcmpl1afSeGp7wzDOMTBNeyJ8wUzyzwNsvSRljd0eqqwSMIRNfk0
sovf2Y7rggBsgZ+HF6xUM0/ZXw0ZZ1cEZbB13epSfLs+tsxjOq0xq9ZU3j1onGjHy8p9ijCcJpUk
Ar7wBmq9+sNmy419c/CFe65kR9HEZrUBQzUiWujw6/0SMi5WEep/+fHdfucceailcgQ9zfFcrY7X
VrrRt393vrgvUmPfd+Sbdp/5J8RNiVI716Xz+r6Kg4a2/wmJttyoMDficpizC3vKvJL5eybnEDQF
Vvg/sf/Rdq7MByvHSC3dbutF2PgNCt5wEvhYMQV1BIfApNt5b4jjzAal0Clr/PfKRAVG9zKFIKfv
+tMvuUMUhxe0DNywojz4Is9vy1CI3RFb+kci6cYlpGtbcJ/V2sQCIICRuo/xT07yrDehzocWatha
w1a8KUF72vu/Bf1SBa2a5WLQ+RM4WPWYXY6b8bPUHDGYboQziL6UzCpqvksG6FUO0U9HkbvXGszr
V9dn4Whgni2ASTlO8iyVsqLrBvkRvMLMuTtVpx0ezTNL/TOzGXXEA10q5Ch91iCL2DLHfOp+t/8x
QOLNB78i5q8UTQbn/nSeGLqy5O9aGmyOlPfHGv1GQZ3fcYU9dmf1O/jXqggSJvOeFLo2+f3zexDs
TEkq6nEUyWioIbTO9ThPtfOK3KVx6RhbQxAdHD/6rRICPwxYGkM14Use8ZXyw8QITRJMuNUH9LNk
JPqMFOOaS5FApfwIZ/NU8T1xp5hhVgsa3bbyzG4i3YDcJc7QYKwic11AygNB0QSzcz2OsrPyEMPH
zYu/BQ+sjNItx2Ks3bLG6gLr6u2VbqM10Px00om1tw505n10g9k7Q0kE+//vpWhVpCqj91pua1Lu
NdXooFIIMD80yU6qt/OfzGcrXzRNro12mFSVJMcO70Ii3qm0hCWg0/wCDX1c4o0dHqHEC0+HG1gD
/oDKmmERsD/RLC0ZxFMi28+AIVQwRx+l/+lONIUxYiHe5fMhT/xFs2xOjPbIeLVrZtdeRo5C3r65
5Y2MC5rz4wGMJoZrrSSvZh++wpI/ONymdtObbHOTBCtvazsU6TFe3PdjrC9EH2QAPLQN67upotFL
qRwYaSEhAiWOMhez1XJNPHVv/G20yObXVnHp4FWEr7rEHNbq5mDmafYH319PWrb64EZ1e1GXrf2F
8YMdC6o2DFtLjWtoVCEOxIvEquQ7hKopB2IhDqhPizeo20Rupk8eOwW/wPEn2bjcm8MBX+0qyOh4
rT+b47IkrOGm45SaAYs8CiwimIeKYEO+o0nkuQQ1ZMALz0RnpnpaSZY5mQQFVbi6yEQuqJfyBys/
yDGe49Hja6EmQMCTK3e7wMDgj3Pgyz8UsmWci2vqNWJR24wH+hKZ1Rd8E2AqNYM1PIgH7iiKZVpx
nbmcYIyPHHW7IjEy4xJymCcGB1X84utCQaw7MysgNwkCWpiW2YC7b0hGVR9vZuD15QgRHqqrU8wW
eJmxeHn+lt/66fCLTHWTDdHZBECFiq/ty2SAasMU3rcEuerMFjJy93Sslr+YBTVZebS3O36H4iZ8
2Yf0gCyDDEnkYplSctAS2cJXOl2hR1qahHvTsc2YUtqPnSWqgi7gG09FgeMRYa1IYY9UBE0ZhPq8
2S5m08b35/p6r8VTGwM5J6p2bfTEAlZcNLIBo0QifDosl7SZ42gij+yIDb2huNE9ECokZhmj1rhG
xAZG/Hv7wCYw+xpTGPrIsHYtgpBZakGKZZgYAmmoi0ekWuDkPKBRWneapZOWD+GWpACyP7igEqKD
t/r/3LOtSwcghLDKT6J9R7wNShHdiwBD+kVxo0bKThOPFrS/gcN6IsvlHoExLffdueMqQrIcVpmH
zANSxActlT1ScK+C/4oUyLs3Hcg7laM0vSqMlDquVu/4YHH68bi9iFi1vlSJCszUjY/WVyStcFdm
ir6KEcfWMfh4pD/rDdQZAPjB31OVklqx4UXhO/sR6KHDlkTWA6yER+Pnpc06uI7kHYqoOMfoA1Hw
FrtShO6VVfnZImi3GQ26MJUo00Djf8W3ZE2Na9xeZNHvZcnmc8K+x6AqdFltfK7l9Sp3g1W14gAv
5g2xuBncDoTJZ+d2MMtDsrxjXFRyRVx09fvuAMjsT3eEwMFio9Nss/ucZBeZfF58p+hrvD0B1Vwb
8wIF9IWa70oSyxYDvFR4wpUj4x4mrLxj5ycrTie6pqgeY1fPZInefNw/gx7uxOOMW+OPcbMgvMUn
qSF/qKsKWp21L+lu3Lfz6kLky+417GoJW/aCKpGjEHU5VSHcSf7VPCDuzc3GA/hp1+A5pB/Qq1I8
NP/k1h23X1g1M/YMj+O7tU9ZNCCUCjVs5F2gI107reqRUmczAwxk/g8mA3qUxRKWwmmS2nTeh9oJ
g3hfuemwP320KNABM1b21fiyDlPlM0w3fbUmDmz7aACqDBfqmlG8IsuvFOGx/IkzvnUifaAxQqDG
bb98e2LShkk4TCJr7B/g7D4+GScD9svdvQTvzgrSuNnbUn0wuOVLwZ1ddnsPoMZKUyCGWhfTfukN
FgsIl/VxPJFmeIOyMoCqbfm3SRQMtlmQKEAvHyO0erGrz1iai85H+qwL3K0rBZQKLpHksGgLxHTz
9gQzgMremKO2WwuuGPR1JIG9BiDoqd7upk5P9//6Ci/nuqRwgfHkHXJqSboVMXvr4t7iSsb9J79M
h95vII7XuYImA7sN62mdE6FX7UZx13mvV0O/s8d5b/G4mL7m9tmbC85xpTvFl6kjo3g6ueBxMyq9
HzJLvGDhDAbz0yKgwD/7wV4/pKOP7PFc9ceJZqkWb6COm0bo2wjFKLq17wU3NI9iPLblL5wDPuXt
bcxqM3rpPjwF2SBHJFDZyBNe196POlZUaWLqhCSnJU+mzQNiyP2NcXKiqO5XAcqWLAIGVLdS7ct+
gxT7NN5Viv6pe5OszzwcL4eIzGwxusRKBi85NqqR5h0u28TYJttaef5xX7tyv3glJKXlRE4pc3HD
E4MR9kFGW8wj83BC6FD1S/lEAQRNn6aFzG8D8ZZAFPsrE6fiAUwIuyYgvky0lUoEr6KHVqrjFo7n
7aPM0rPeIQUmayBqsw8uv8ziGs8YZNqFb0UjXpHDZLgq+7PUIf5AlE38c3TjYit0mUkqxR/Nza+h
WSC9rcQao5LQVOvAHP3rssfIgTJ9nwa4IFw/n/1+YLJSigQqLC7mJyDMeRQgfijTwoewzDZKG0lZ
R9xKQqso3Ar8mvK65nOw1yaGTNc4daiT6xscy44cZ8GHro8ripQ+sveF/GdNw1+5qtnxw103ugBn
5OP2Xfi/fsFtzxWRhnz+upTJdKXNdYVnqP2EpWIKahO/CemtPXPereEjH7SRbQRz2UpFi5awl6Xw
9mnUMAyaxQfgh2vTvZulHwFCE5sGsI7Y4/+za7HQPCeeGht0D6qSlbOJEZhU7Fgb3MYBfzzAADj7
ZJizxOJa9luhUpQAlL6Mxh2iP5+IOGlaiLn3AlMGvY5z5bYvBXN/yyzWIxBnZiwSNXb2lhGyyuvY
RtQe/9ZzJK40ygLg05zhXW2ZdRTnoe15I4jQK+DR+/m7e1VPhkGp/u9ITwamf/iEtaN0eSFZfkpF
u2mr9JKHmnRWZzGbCGHitkqbcyRkEQibtOib+rxHVNRieRpvBF65Sl2vmDCXLmNMbqnbjtHTeIVz
p2emn4oI+b8bLG+tMmZSR0oO1EmrTA38wRO3y4UjRxPXuI8B1dJmV3ehADpSWU4nbGpuuTxINzBK
E5g0MLsNx6zcm5BFz3+ZcjKSncmYozXJx1xfrs2imnJ/XwYYXaSkHyy6/6KGQoqLpNHsAJXlggEY
QblRl/8sSzWZyFw5zPX4rftZHsbnBG6uktLKx5gvARvZw5D7UeccQZiEDWX//TSUbfHC+WLW/vBv
hugMBpw6/xplh8sIpqf9p5ZvqKLeA79a7rj2FBP60B3UyXq46b+7p9eBl3hEcJb7qgvWfBtucKQB
AkO5nRi1OjQqTCt/2Fe07vLpGYOjTgfl6sZuOD31SRw+tHJx+B837RWMLSnTHc6w4J0ryEVb5FLz
TKrucycLEDknIU1X/qCiCphI8E7c9hLegGJtEcmnNQgqMEQ/1k1QimAjuJN/6UAYr8grVALA/HNV
VTL4qHHwPtwWPvrcwvppoUpj7kG3Q/SBGp0wJcleuBi4IoMzFSHqFZ5CwiaBdd4LHakHLwN0zWpX
sH3Vp5AWmV9cEnnpaJWrjbujHFkblASw4mSAT6Ap3am3CxyaLLysSTjhfYTqM5e1WTrUrNvx1cjC
pGn6LGszN2ZN6zMLl8XAoigBefEYuzk0z9j8FCyAgBVKHN47U0M9SkrlgDq2fyNCBJ1UruLv9LWA
o4o8kFiRaqGl4i9AnYcKBDa3naQDzL8aR8QcOwMKp0qlu8mLXlNBWy8hG35ZzK9lsvM6FWS5u+Ge
gzcRJTqfY2L4rSes8Hbc95ElvHluKxFCOBNPvvN5dso6MRweyj6oOhiv7g6vAJN9DK7XkoTwqEdz
tNoZ6uJdIGGHxsiw83SS6IboSrv79yOEwKgHti5TxunIKgroE44S2fCXZ//ZIoNhcPUoQs+lbdXJ
8f3B4X4krZWKJmbaDDsd7T/z+zGc1ZMSzXdgRTdxfS/gWekqjYfD0K4/EUNlVyRUcicXqbDKOUtx
iQgxNuIqXM8pJCLtMFPHS1nV7BivXjHAIzjqwty7EYYqGHVbk1ok2OH+IrjWq8rbioCiajbZt/Ls
EPaameREbgl1ueILU4sLmogAB5v5Z5MGNQNPtLCtHzTSaD/9tIICavkJPOM7z/SSkwOZm0ghSpU7
0mt6SDtqOMA2NOJ7lWxovNVwAxwwRK5kngWrvMQjZtipbaejH4KE5CtSgi/Cp8f1FmtJVEvcGJrg
YDUHwBvlE07oD+Qopab03FAPME1W2NaheqcetU0ryRr2qt9/CWs0yonbv8X3vOUfwMWggyv1hsHg
hyjgRR5xDOHNE2GrenTIASjrg3LtyL115XIyL5FoYqUzkfp/BJo1bprCCnQWlFS9v4VywMidFRV7
pj9Ddq+8ZSzbwXfbLx/5o/maZ0ZgZQwkzDMIEP5UEFRPhJhY4o4Sm1f71iWadoBXO/dgisKNT1LX
qzPfNWLHnh6ihk3HaZPhKMn7czN1j63rSLanG8me0yVcXabFD8cVFR/qZ38tf/eVOnvq7m/SpymM
y9dAmNzG5RY2ADwPhSNxlJ+5TqgjWxf1+VoewTfI2blHjCLnTIIIK/EkI/IfWvlJPxST2QarKUIw
Hk4ToPK87lmFa0Rn/LoINMoWIbru/sFRbsgvZhxTUaZTLmjz87k7GrP5yTz2YR+WNl1xSEmty6c5
Wo4BDWaD30LtY2mPUkGz1WLJNzY7G35H2rR6awKfg/D2zxN/5L3Gyw0lXtAsQsOuBdTn8N4KcKf1
4+iDX3jOXa0KqZiMk4DksKVrIx5hOnOskxgMXWxLtRocdBdVlm96JJtI1DfNXqgOc4Ozaabdt1J8
VowHEOZxGAmLhF21C+ldGTV/WGXtayLsj15p3dBE1GXn5ob7ZTODyI6JzOiGGIuRC2WXtkdLJM0U
bK73Y8WMB10WM370L2DCXeEIbDBdRVaeC51KSJNRwwnv28VtalLIp+0y9GC9pc9aZ6iiSBI57frW
i4EV0co05DNvMuPCbgusEPFd9o23CXr0RcV6iFu/Xjr5Fiea8KDoagY7Gls4K3wfRWqp823FwTyg
+9ywpHSisES48ybFbCVXFD39dka+bsF2juBgaWVXtpWY+EH+3stlrUewLtAHnuMG3P4SOuKqIXiI
p8S1KRzzIujLa9eVlrZtNYgO55gEMLYH5XFC4PSJSbqZgRXrOVz+ALYdgvOQka8w7GXGFq6n3lk9
g3ErI0VKWxURTTfFyMHYXLsqUVAhqYu1dMFzhp1TxvYUH1HvGTRqAMD0K3gef6SzEvffx4oe7qnv
BHFx74Gb+/FZ4oYYMPITKqtiqiPkmoPq4sOeU4W8MyBiD7dQa0L3llUk+GP4+bbH6APGACrzxGxD
udUttuvH4ubloUMRwAjELVZzoboExJA9IhippQJFSCdG19WxuTZx/RU2VazCqUsQZ1U2gmmD6sN+
R3z6WrPyJszxwodeTWV8v8XsmJJC3WV53cPmogNHjiBFE+B5+6ekvGemkhPpExyNEqRab40+HZ+r
Py7rqjKuja0UTwnXctgpEHdaanVDDgwMCnxeyerLO+ZhXL8ikJd7KEz2LdvMGFSTCfIxRN0QMstT
Sx6yVoBcjhvmpKyDofMo/uT588ODdi8PU74cLeB9SQBxU7udMdcCdGY6wQmlfUSnSTrZ+Mqjl6aH
nFfOL/U4fDcSZb407M/6Awzw36euK8ovCS5qRQBNHG5lXJI9gD0jyJqcwpNLna/5zf/UrKZ+5l4k
wUN15unRoAbgKgO6KunS2S1cveslspOZNsu11KdVRendcPPXsZXj/IwxPluuUN6EXDbbOK7hzh3F
reS1+tf0BArqMR/3chJs+uWuN7h4e8LHCHZO9CKMOS7Woe4YwC+hZibiKu7+uvAmJlNABCalK70C
qzzOMl9tRVVfm3+74h1lkwRfmd4Rl/wQu0bq0BjkXapgkhZZ55+HSyJtQW7PdWmwZQn4a5QP2PHf
psBntghBgvrOc/jSYz5o25dyhy1OjR96a+Z8h1/8fAPLiffEFsJTKpCGY6fyU1nzkGM8v6luJppO
Ly+2HjiOPbpoRAwdLlZAyugq0IcV81E3ZTGiw5U2cH1ND7sSYOKH3bvUqE3Mqy8xJHn8QgVPYxQz
Ak1DuuOppD2+y+stpRY0GYYV+Ir746UAvWgcueN/+p7hf1b5gn4rHcnI8gGnidU1NFAQUvsyAXYI
thwDqAY0c90SOUaQQj2H55igTJWzxrIBICM6Hbsao6xsv/jVURLvPo1xOUiNfk0r3fOxvaY73WKN
hsRThXvujWD7YaDpn9myR7MUfgzrbCXElFxoAEwhm8ezCJaoVbGI55BW8iTrZMtEMabVXiS5aKYX
3YHPRjB4aZytZ3g1qagKpz/68A4mF7639mrbWlfu+HQsNbu+El7VOiEWMSwJq11Q6sy9YlEMd1mw
gHeBgv2c76+vyjArhO5bC4HhVWYqbWralUfNO5/VcJmoAfmOrQw5qwCdYfXVZ+7Om2lD2+zM39ke
4wF57ZSZk73gIZ7QNIEszyvFtVvhM2nzktdO3jjsicuqYoxHUlNDVKeiOjWtqZBeavCOACNNoBKH
Yqj9GA2w15F/x3ldLrbM78A85UUv/3uEI73DOV7WMia9K/ggpmz+pfihPly6cBvWELWf3iTvq9ci
Mqe2BBZgG0X0WnFvoJZLGZ6tu4Zw3tfb7wFEahVxEC+4gJvNyO+Tz+HVCo+EvBbwKa6dCGdBCLJg
IpvP5S37pNTYxt8w15BAZhir/lnQPJFvzB+1rP8AerN7SqxMBqY4YpC8E3RAPAEIpmqboc+JVhOK
t04l2Me6XiUsy2bpPKkQxzdVhhd5N/9Fdvck1B98eSLQqLtaO9hvwgQt0iot2Lbj0WOMFUs0nQld
KcrEMpPGlx61pM9mhnBrLXkF93eDkUzjV5pe2EmkYeY5PLDxA22eeZZ1lWPKG+9cwG9w/DtidaHh
YtYZaU8Xp1qF4grFGpDI7icPxinFex/+kfPLMo0Ns7JO9n73/ay1TnykIrvnVNXh6kfOrHdYeyoX
Olt2R7O0Iu/mBDpK77Kyc74s6kwSn/h+tg0+bL++t40fh6i/ouU/UlFAL8ub21UOdZLnEW6nWxcB
FdNUCivqYJrZV4G4o/Pm+uyMS/rDgeJ3uqR+YCLnpmRaeESnMei6nKH+T95HgqGq+madll2/qeBz
Fq+AcxCDAZGpGFiZtUNmF5mKDQFFr7YBwCfZfrQ1lWsvbJTEewOQQ6RLejFOYjBRGeNY/tYTJWYj
DU4MrIVC5T/AkW6b44b2GPXNoTBf2zndYLg1qcjwx4GPQJwAgus9xZwqEAMrCB25AmG2CaOxuyg0
JKBVyK/lKOaEcGIcGPUF6E3HneIsDV/eo+9CtDcOMWJ3/Or47x0c+BKsHl8o7IoawOIveXMmgf+P
+YT8UJlZK/6Lr3bMleu7PazFEGtPbd9Vy810k9/Yto+4RZFNM7JpkJeFu8FhziYiXuuY4iFX2Cuj
ZYjJumMWSMfYue7I2euCL9p0QZnmUYUaEc01HslJ4/yldZeMZnm3xTuVX9fXH0vdxfNBLcaNoLgm
zXIWZmFx8z9/Ty+fagoR4piSxYexgJILVvqmsIb9h70jBnN/Ok41YzF51Rc7XJe+ZnGchL0rVk8m
WUVAn49yLUo10AXLYLoZtXke9/3dyCujeh/kjGtOrVbvogb/XMGJ6092oKIKf+qlZ7Y8MFgQg/ap
3J1MFTe+WeyMaZMUbiYTg4x47huRSWt0BWTG3i/QP1HMMj4tRISNLLThiBxuP81zv9PQQezyrTZj
CuTOASgcXy4Y35Wc/jrgCFdwvFMN/aI/kfM704aoKL7dv5nAyAUG76sw50ryVZOCS154fmMSu70+
sqZ8W1REP5ecdWf2Hor2jPgEAYSBAkPG6jqC0xvwkXG406yPZ03LdKe/xBF7Bwbd2u30UTTErnPw
z3su7U7PuYUgalLpYcaLCasyQqc/t9/goj+KFkaMBSA0QOqyhp5Y6kerkjRLBoAoxd4ZrVGksD47
ihFI+ZprYMLMhFycEjiVqNor6JwWnIQ3wjy+Fs/Im4hydITM+kSOuifa6sGx5J1VE58OYo+kr/2v
mvEZpQnpNblfxpkQUqJEys2m/oKjn+1fWkZVC1h6YH5ZLcxHx9TsLM5mCiRoXYMkXr95BB1MDsMb
v6PmnqumE79sPMaHUmviGga/4rjQ9RiISoGQHGQSWvBbaVyK/P2E8zEMuMeHFS9corh4iHdRrhfJ
zHAlVFlYz27+IgBR1xhJPLq0dKvNCeIvOXqKximZxdOFdI615zT1Lx6aq89C7J1b1VR6Vt72Jd9+
LHGOb6i6MMMg4UTEH5nIMUw+W7pv1oUsIVWd8a2MS1kWeWQZT+947tHL5DdOUwLzzLz7CnO/CCMC
/EzGqjQAuZadUhxAMPzrpK4EItkMqw/VklB7pUDCcEOi6G7AAEClZz88Vren1eQRskpy0Y+i8I8y
wl1DSOlvP54o/qTLpv5FRpWBsAO4vm4RNm1jSIFoTHdGbLTFfUb4yl622Ma32p/om3q84MakyNUa
GVNb29E+Wz5uViycvLv3EaOYQHf9Y4md3wTvfY1VhEQJ9WHuQXEipLKPHXq6GM2zFRGtCPI4YFOX
Iz6f1ZgPG6SPWVWxR0MCc6eRBBI7Ch33CuGLzjCFnPvs0rRMt+SZ2horBA74bvstIw4YKxj5zd6B
AoYwNgu74IZmBNOphdRjvhzlCPPbXGe6m9FN0BYm/qPANCSSqwXunEJq86rlAlB0bGeOWXmb9kbw
1mE1AwC0oVjIPlT23gvYjKWWd6zESVBKj0FM7cNCaBIXYNz3i8EkroVYaWbqdvCUIZLD4n6HnDtH
FkE7Mi37FabJEg7orRyIvKyEGKthD388nyZn2BKr6K52dxL17kwIFKxlYmz/2+CQ8S8A44NqVFNu
ZG2rSTOCrjmAhGp10VZhOHg/tmL/ARsxidoZA4Sgh+xDxzEetTR9wXDlXJx7IibnLbZll/kU4C9V
hBZ7i43Xk8gk0wLwMid78o47bs7qAIgYhT/dxeP7o48arg0JHd2nHEiEltmahjGk3XpNJ/bQB3PH
IEIZox/yDt9iXanQf6KgnJn3ZD0zlHsSP18PG7f3mDKlg72LRoqscy8KdJFw8Vjh/nLxPcyVfinh
hobb0ZlTlz8GlpXAdQe7Q7+uf8nNLl91xo/IOKdRrSGy9GnXRazFI6tosZZuGYanXxDUzgdKVm1A
c9mH9KcTq1LdXxRg6LUO1fiZ4G2kOnjdYnBiUSDmt8KZrbWNiHtqm1CvEt85/wRlTXo2bJ0NqC2c
54crrjrYUm4R7Lv8YMR1YjpOnaN0vjTJWBbDR1SB1mh3lNu6JZZVl55adZQU/A+3hXTvBzE8msTv
6YOCGutD5ayKNvhlsp7jwICEjwAYpwxrAmmpOHwyKfiRt4SNBT6sAwZNcMCSK00GRUp7dI60yOKq
eT+JvGowE41Gx6hOuVkjXBbFWKJhIslgnr6F/JFjZ2N4Ggs/pQdUCLBlxyq3hixNwp8sGCKSQCvZ
4veWZykOtReL2HNq+yQ4aouj5IzcxNU4zCcxUw8Vj5b0id2zphyin5i22MSPF1Rhp6751YYEmxmH
pM763xi6eFuSk+lIm0z9dEZLnW4tZDhlMfvkrdNd2I4JLMkZL5KD1WSoXcaJE71rSD9Y2/cbUjZM
lfX54E6Nv8cO7pgs8bkC4V2eIPz0fKZv38pPBIJQuJRAicdvIN6c5V3SeHE7InyvpouEJEUW3tBb
PRjd5/m1wTqbosR1aFR9Ecnkooj+D+2jU9NB74UdzBfPUFv/4PsJj4Rpr9YKpPeoE/r9Ou3+rwb5
Nc7jvBl9bt8ZLlIt+dzqfME4kuyIA0aBpOIARrp9NrNEbmufi9ok971GbrPUl0kKvcQBAK675Pcv
pfb+xM/LwQNZRP9kPU4Ud7WPyS95rPpGiIsnWu/BFGjZEEciiyuH45+KgkZqrD4rO2yAT7nxPmaw
ptzjaHTOImhhCKTWR0c0UcFt7OLI3+QJ7hiyQhg1qAImo6H0PLzcrcx+Qy5JjBniO+OVmVJbZle6
Fu5ATe66GdJhd5iW2Epzd5l/zmno+7jXBdAe5RdcvzH0OpQxZI1zhwLrFeyrQvb+erYpPQlLvQ8T
gCwDyJyraMVEj2+IvUC9kVz6Slh4A3vPG6dyf2zsStJlENcak5lzDgWuDOuifYSDYdOhX7SFUZ11
OT9rsKI7xZhjZCytXUog6Odn9QrX+M1EPJcOpbRPoU1Kd8KNFHycvQWn8JXbxb2kdvkUVtqnr0W6
ss0DTyCgUHxKfztpoTl9uy8aQLBK/cu5ljt16QHvvr3y1fK4DDYAyb4tpljIpOxHsCgWfc5fP95Q
ZcbqBy/SXEPbpnnYNWv34s0DXznCncRk4xS4bsKrz6rKR3LDbgNypg1twMn/VR/vKxGjGNsJylL1
8BB6++kfjpSUEFISdqlsr4GpwsLzEhut7ddchhp3QB2CzI/vYHwhrByaaMwL3oRGQIDnKjCC6n6R
KpMTdcFboGMt6lnDiFZL7kZPY1j5m18+RF5+7UJuw/OUtAXiuGvjqzzBO6ct3maDE3B8LTHqwLit
u791N7u3rl3agn7hf2sR1uiFHiTl5u3pMgmqWE+lJRKFCfy5lt98iP89ziobo7t1aJq+3Z2OLXIx
aIMCZN8pUQT3/PEwdtC9uzHJbH2L5hbbTfpd+jR+UodXTLjmh/EM8orsMKEMJBDHYTP3lf2+vUFX
AiOOuaJuN4SfHsNpRukItYW7WHjtdw7OIEffqyg3LKKxfDlce3YncXLzEoFl9GgNhh3hyaSbDgrQ
bTNCOD+MmKJ2Ek8wuwXrG8Qe6XbZAxqRYHFBDStSuaDSZfbz9/91rL5KXpO5QZLXPwe4YqkkrpK7
PDXuKv2cv76d4d7cXUYNOby3wcY6nxJ8QlzwMpMgbIalVLX2BxptLgCu7Xc2/6O8Gc0EdZd6k5iq
48+iRNQk4OV5tl+HRdw42XFUmzK9N2PCXKl2lobthkufoECOfzGq7Zn+G0x0EVGQpQ5sEs6YvWt3
Iu2Xvn8yXd1HoNlB/voxJg8Rz7O8kpm2+ONTtnh6pP3mPOEn33ISGxxk2i9bMB0vNf28EJAFsBqV
cqEtYxpad6aXIZt01nNMbVuP6uwPANABABnApbcMvZ/jF4zlNPSkCSo3qFVE3kEISEneIxF0kWeQ
Kjw5KalHWjWcibXkY3vEwUrM+fw9JrJyNVKWOz8oC1zGZ2nrwhDNKQYO7B5ar6f91s2RrY53mloz
0FbB7amjMTGjQYienHLW7KAlcZluVeKm57XuCD+Td608BneFVFMNLowimWuKQS/YRCs5r9nYyxx5
fjLzkdnwLeZwmZHaqCMdkrzOMbZxzMSuwP1StoHJzjd+/bXQG6jKaqcGbm/1aJ1kvGBIy5I5dOts
TeYnbXkNjKSLoY7AM9EKfF5LgcUAuzNq08hzRJLhyg5UcSgLVviStQsp9jz2jDKhG/EJWTK1KNM7
mX0xvCTJcC+e1r+1TO1db2oZ6uBqT6sqrPhGzTv4ZAOxL/8VKs7Bfnspdk8jYc/fgvxXEX/FBmb4
A1n+CYhDhSqCF9CGgmJd8LgmNKBmoRvQSYeXSU8AXnihyBwmEyjh29jc/K7qdeIen+yrgSplxH4/
YRYOgmL+8MlOkegAfcdxF+ZzQoxGV3UVQ+znUHudyZaMVf0oHH6CtTNexdsuj29SD8jZkEnEcmX/
WaX0+ZxuuoFzbh/XU/SKmNXFWoG9nmgTVDwxJwS1iBp9HqHMOAgQNJrCuIlXTrQeSrE9KbWUzzXH
tMTr9oNnK7cMhW1Ib8uokiVF6XLUgTOCoePkUCIdq0yS1lMWoJwn1gdlAB5pKMYwcfjvMxdCvhqe
9GLJeetLBn85aP1+yU86R7f52/XzdeS/Sha4EqnoDYFBGyHVl1tLHWb3mqS8BnC+u8ow30WTQmLk
T4xR5Mfwa5r25PWJqswB/maif+M08gqEHpg2//hsZE9Fe5Y6xq6Futo5m758bZ/jCOZr8ynDZGf0
Gi88MVHO5cRpH70lm0qjSUXSaQ99uN6Gj/KFtPcYPhxmFW+7+yksfA+cCdryboYcS66qTU7bmHqz
9OdINeBJpaG00vvA96o2LPhgnGDMhSP1qoRrP0+MeJWDUtzdysMHsnyzoA96DHzUTk9lbgb7seWy
Zo5BMgAQdqb7Fh5Xh3i078u4x5YT0Kjbn2Lt5LGz0oZ/Fn0U0JhEwyqh0nIrNu6g1AekesjALgAE
D8ObqIDZN9fTvlh4V872JtjGUCC58+1s2cBr0muqIUUbGIbaMGSg6HTSqR/Y0GcshhIcDi4AOObG
NomOXdGcK+nFxUbcagrM9fOA1u6Y+DFMpiFw5Lc27NMy6jsqoKxkHhIyEMEERt6xAAFmfjyNLnWT
0mztoh4Bqrn9CBUuaD97sphmb3vigswIDHh0ODZQgbFKt3EBeAmrZB6Rrnfi/Xvqn7Fr/6aslDuA
O2tJQKdv0bPXW7AWVLNf8vUniA/xs4sFADedr6uK4Nq/XfpzislNu1ejRyMLTkkafvIS/Uqm1DV1
LropSj+LK8BMLq5EFrthfqymKrDwk3dIwNPo0ldcEfBirK0Xizjzfm7jT7iOTU+iv+5PfpxztWrZ
v51PKu4wUY9EN0wdI27XPunHBqjnxMv3g2eXQ8nVIQUKPJlB8ZuRObLX6Pc1+5cIVTWVq0xxRrhH
9TR5eV3Nf3dracPq1BPHGzePMEizsYV77xGgkb0qvzuS05qTOm7qHKPW46v+JcDokCcOftpXOoBQ
00uTNlHwQYEeJ52tt32MsrJdTf11QXJFQCwbpiRAgutdfFp/wn8R7cJDRBNqx4F9vk88nAhXvr6A
1Yj3eeFmUHi8r9m/cyn0Jc8YEjNH/r/n8Z3ib3Z9xyRPnEfJoEMjvYMJAOSAZKjHyoqgpJhYwQtK
cfwfvPJh0+7M2rqLGhWZcWfxFURZxhLpQLxSpEG+eA0sXjm+7TSdqYrwPffkaU2YzAEg3hgQmpLx
mZUgtBP6Eig85iwyRdiH24RRPDBV+ynpgmBBVF24fyM5jb4SqYMUvPuOhsuOSitRqPoKN7jgaCQR
BgtTryMN4y4MuY7/FPKsM9JXK0elfXSd7SoWts9N77XxFXx3NTAsWBQi+Bq9KY4iPN6x1XPuYrqK
bZq2MVEb356ukXVGmFWrbvjL/fyKtqU+5K8iYWeJcP0RhtuXZbslvkLOV9WCjRPcSn92fjGSKD1t
iWFQZME6Em/N4x6xJJ2ht7Us+2KuHgM4xup6b51NMGzwUi/NgjfJCpH43r6XlRM7hX4Ee2Nv2+DY
wZrTVDBcOvaf9+1KNHB0MCqf5SdSfIuDq4xzpyCb6ruLQTN1Bv3g+rO/cc2MSswTTahhL89FZPTQ
u+Jt+R1WASTIraMS5TJWtsYPFzOAjNifszTLQja6Ri3at/FLBbHl1buCMD3mGAcaMdT+LOzLj7oq
bn7U7Zdv+CkrkmRzinEBctMM9P6ZdDwqmqEJ9RXGBFN5fByjzGlDWfKAfuR/6IVJmqF+dRhaliDQ
aTLepaIAWB381GJ6OO4NpNhHDsx1hN789xvkbIRQJhQt5QWoia6mhxq1pF4G99aPJbaT9BrxNdGk
6xHPVki95jvOLQIG+8rrO+5638+IR/MTDgnFMkRIpMfrF59oRTYmWbf3vdIz3bMiFsPDkotugewn
sC9HCjhEz0FmTK8EcBePfzc3RT+EQ8VjX/cbYRRzfKqivDis+Dh1Ux0VEeiyN4+HnocAAHFzYHIQ
wgGdYOgIAfPrrLbE9BM9tVcl/ozG6ps10vmfpXBNfLKh1Umf3VF/XZyYpwjU1eZWMQKbBLt104il
r+M/T1YqRmlULhIMqK4+Z9JsDb0eMEd/lrRuGfG0hPPVar9AE+xwndSiO66PnKoyaEr1MBsouCCA
TlniR6seKTwTxSGzClRgpgenyi8X0QbpGYOJCy2IYJUEfXqYV57VdikbUd8/ivigIpBzGoTQYgHA
gbfSK7h+Co1JK4byVKOGUT37Cu+1B0Aq8wog1O+I7YB6dGGA3RT4uAGou5vQAi39ttrvzKb5B9kh
CTEPP/YUSPYtCct/6r/W2OI6HassSeeyPyb66h0Ksa2pO1GrYyB6Y9HWH+WUGjwHIj/+r7FwaPGf
Kni6dZRgOuMnsopdW56jTv2rw3YxzvK6EZ3XobrbR6oh+gTzRbNPsEBA74YgwFmDOVq+m7iW0z54
TYdWlXWQbyylL20O0hCU435zqImrMHGPHjvJZglNX1U9Jn+iOBqdjrGxh3Lj/RMZYFGgfQ0AnqVT
7YA5D5vQmWioC9X6H0L1URLN5/YxGa0nN7Iuk3mY3G6Z1I92F+bhxK/TSdjsqz02rm7jKtmSqjej
2juZA2HjA+c9sAs94z/zqFxOuEZ4Adm5RZuBs87gmt04Iu9ZOM4WwxrsUzQgcZzkSsZSxxaly/s/
3tXKWrt60rXDSQeK1XCgcBgCApiBORDsBr864DW+7xoHtH1biboE9FT/WezLpXskR4QZJrbvIW3O
Aclw5dvNcF0A6KYzgsw1IFg4uoAS5ISmI1+nuRE20ul9e2BsbuHOn8qrP31pE3qUWJNRNEw1JuKs
R531B9oWIfj66TcMqOdtP7TCEigJtev9PrGlha7xRsgk2xO/5hn+V18SROZF2v1/Dclq0Ulq9PE9
rQeJyjVRP80HN2PD9loqE4VpKgo3LLOaST3uwFroOqK/V5+zkc6NiK+nw9q6YuHEmjMNvtlAGqab
968f3t7F6YVaEL0m6eVVLOs0PL3LQVSPPCIzwJZkwS5J2vyC53lxVRGvdL4vY3k8yzT2Cx8advvn
TJm2SYRzY6tjh7QNDRsJG1jQE9Trsr2224F4kkue1kz/Btbnhj+ivrwtGM4rds6E1g5ga4cVADG6
4dd9OLocF4QlPhToNC3zgwPHdUIiMRly4QZviwvrgE6jrTNdQ0bqGHPP4dY+T7DMEHzyGiYeHmn+
t4QqucubRjD21SMrOTzHBSSJVWoJAH6u4yx15fl3XoN+l/4GvpZ1i31fvUvIFqL5q8/vu3jRiviH
r/+XZZt38fc6xQ2LYnaQT9qH0eP9iYw0CeYp2EfhSGY4gSoLqcVdAJZG1niSXQsEgcVCcIuO+l5m
7il08yKPQNEQOl557MdQU3vHsG4OyvmbHPRt6T6abqFbV7OPq2X/Q1UXNLXRqF4AE/mmoF5ELXHa
nrShm6NO/qpdbuqwdYq886jWu7ahv/AAKRmn/hXhcJPBCdXNOMbXDFIKtt5VQ9WdkKuKaGktITIl
L7OtT9Nuh/KO4zFnF0O1TKw1UaFvc69/QSTx0C6CNbWIWlpfjEBugoHlmOBpsba1HZO/lw7lbnWQ
BPNQer8zx43B/OJW1gYRoK/aFtZj6nfBk+AYyZKcoGVdEurjVHxHRXAja7ef0EdlXcU/xYt79ZwL
xinVnqD2DOZ4O+LoBW0iVuh3Q7Tzvt2sXm4izC6g7FXdpuqFzKHh+kr2vTSc6mTHAZDOEMcwbSn6
W0BfIZmzZunUSVs7StmEBSJZLg9bhnXY8LKwTvFCpLm2n2jm9BItPZhrGbmvRi4xT/fiQt1QObdQ
w10dUtRm9AfTCYom7aTqAX8jPzN6/vmL7uRhtK9CmxkI27LwZqf4sLfQDZAGMu83DbBH3P+/6XJA
hJ3OfSCJikcmZdDxwQ9s6kGTCQ2mwLqEimFzVb4mVecZsStGkqGQ4be4R++buNgPOHKAAHhybIlH
8MgOjuJ4BsdeoUo3hHTCBetuxPiFV4qDO7IXUlNncoK2n/+lA9vodOHpdqvwWlZEJvb2gW/6VpZ+
8UHyBCmiy3ht7z3Y5uLGysRJg/rsqCyFIdfzirZI9a1qCFfyekpHvrQG8tci9P63jyJtIARE83A9
oSrAHUyhE97Oyz5j5ZkZzVyo4SBkQJ/z92/wyP9VdPomHbhveBGVIjsvKRJrjFlvZnrsOdDafsmD
h4AISWtqVzUnZrEdc4B56SQvG5aoqKUmkmcc9DhQ/lnyme+LABdWs8zv8uNINL7D96C22qFvX3nr
2QNA53JgpzTaSdIjVVTGWBHqfQV6QRAH+siB1Vu1yKnBwzcoGsLvcU5v0M2NfdjHlgzS6uC1LRoY
hlvRD8wsU1XiU9NY9bGuOlvApcu2U1JQLYEH7gGpjScsq9mNz63MsBKQ7j4m2H3LIvOKejDoeQUZ
7hHTCN9U/KXbFqKMzRNOz/S/I8ao5Vn3WWOC44tfOs3Sk2mxXsADLEA8POGCEr6sKxUN0/i4Yd43
sGEbp6ZwubBObGNQqcLSO0nQdbA4JQSafgYdK6tf1Aysg5F5+FYuu1PoWsbRuqPpjfatsG0Mhpiv
hrK5TCEyE+CZCzNNELWmDx13OdTUdk7lV+9NFH4Zbvu74/gHTjERMymMuhnGEgURx6ONSjaGIptl
YIfqUQKoNuWIMEVndfvl23xYEC2aIG4wC/tCUU4IK4DVnCYmAIA4gINLsLF5IjOQXM8Cev6HtPM+
RwT8+aQ6+rP9IH2SW4fV/Az2NwAGzb9x//lh22esgQmTQcUJ9MSBQJwyjXd+rK8Kf7VKaN3/wAQh
vjklKOWhg1mfEx3lFm68RwwTNlyJ7OvhI+7ArUDWpD3c4CuPP2W5kn81rCfV2YaT+2RqFAB2eMA/
nnkHmIWkiA5ixNIYguI/cRupLiuYfQBOhadUdMMqV2Yc2jhPXhk/VddhyUDfyLLeYJPcxAcPGe1/
rdF2DfWSHYm9c36ESpT6BqRizGLvuAdQd9sqMZmTQ/DsePHpwc/w5D+Q0yW2qwBQu5+MP3ps7vEI
NB59dag/CTkwAuk/72FwrK7VxbsC9crJKzdtl5QhWQonkgVDxol6sIQsmI7nIxdk1s4K9b9LlPaV
JXhQhkt75Togod8NeU0Scrcg9uNjZNtKhqGFnmzvHy+4UYBWWzcSfgVj/oNyoBiYU4GgwiR9CV5n
Rh9YmuL4bQIgwN5Hulc3MpxJ6bNoFy6sS4ip3xhbfaopReiXAEyswrLfIHZ7JTZ/e6W1M1/qojcy
YMEWatKCyXOtN2kBwoVzRH2ee0pFtERm45Y385Mh+4fsiLSO7pLbtJbA4EqMrM0oJrcTaN0M5dW6
xNddmuEdNfVGoLP4LGuSgB+qch6nC9BfidzzlhTtHtFEtaXEEJYX+gIMPKmOAnpoTvJW5VZHyFqu
b3q+OzxqQnjIxiOZqQpAFWK7tqSNXkXLTUK5wDYnSgS9gKqag/cThBZj10u7e/u7PqAua3/eBBfv
rm5q92L2eeXlM2t3gUPF5OOF9KM4dRPxGSi8zbBqM4OI3eSVGNDKJL2G/8AGvT2JCXYAUuVZTo27
Vt729utDRULWsKJwMUnoG7tuJSEJD+AUW9Z3LIRnnlbqV4kHafhtIh5mvDzDaN6EsGIYIRGEx7BG
j+wZBUk7wG5Ef8UeIglsZF51ugKGHkmwmOssbR+dXirJjsw1XOVJnb/gMp3NmxAmtMz4MdHoEPvx
dIgfN+garmohDJiAOmWS5YcPgExQ8nFwzh8LAk+0Jjgn+D47Josx6B9RJBK0z4sBc3OUUIAm4dgK
nFFzvvOEyhTWzJbdzatbu24FxfpL
`protect end_protected
