-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Rqli1T9BUf2PizgPagyUQ5LyWiE6KTlZFXjspKSIvSYGjQ9X6US5+CVIudTCnvTFmXINtkP9qDTJ
54PAoUUktydtWV6zcRDKT8J3iqxAxejHrTaHuBHdFiER95OrQZ2tAJD02+KAg96ZuPrX5dUi0Ais
PKLM75u7Wz6433ulG8WaWj2K8W29H/U4NPJi+ddwBexJA2LWTjKlLcsnvUvOCX0b2f6wjjumtMR2
pYHXqMnFDSBHaxkrzxkfAHuq9VU1epK7ZyjyYccmWFEhg+UPEU0zv3Bg9PWxLmrMOiTswP3sPPJM
RaWOyd4mzkKRv9V39XVjyM0vMU+MitbWrq4pEg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
t1MgSWGGbI2t5M3xlXgcYL1OKLffgVI6YXJxysv2nPP7Ug6Qnb3YzJLjXmTH4CqGMhBgbcI9Jthg
QwvxVqqSJSQumN9wsekNq2tgT+yWznsnSamYYuowiZ3czAmEyOr+f3WXQV3oScy6ILyKfQZiU6TI
uLJrLr/uLrrlGb4ZuR86XFf/nfItNLy3522IIiR4QEWIE+dUwnrmTRJ17FgEhxhUi7NrwM9AjCw0
0/KKoFTPKZI7qcTdhuZcUrmHqIN9QyO4nuS0B6fUZr9l46HPR2Vz12C/kOLvQFHUBz72EClx1AYy
1k26enlhiBxsriGWnR0zfOfF/UM3S5r9XI5KDB/JOpBrNWbU1/Z5j2n2tpUCx91BrjCcBkeoOVX+
WqRbm78XWsV0yx2Y5I7nioWoTL0+DnU5KImxdomizqlKYFmeegNrDR4pL3i0LyHr/v/u8Z+qvOS0
+BOgguPYogMtPJNwYE1O+C0YvSOwQq2eo8YbRV/AkKGOF0P8Q8zs+IKuB+1N0iR/zVWq0TFcakCd
auJ247QxPPmWb6ul8RPTc0MM7zMcBnPkOHqiCN4PSsbREcd+xhKzgq3gXyqXrAOrMrytyzIA96LC
iggh9gee5jbVa11xUgYTM+UHWVRP7+m6fbUKeIl+krGyKst0QNolLYcU9GTzDV6WJ1hGSN4hpxoc
QGDBsG9JOzFBiD6B2U1pM5s4oSEH1+krybBRl9ykJUzKmomfTfBrSJcRi3+BwuraX3r6VKdS+jUX
uynr5vFpTnkhUxIwnmhQhhgOfAZelrxamJ3LgDOcHzFz4U/yhtVUM/1hhr908QiHkV5d8geBKjD+
dKZZ4eAbrKydaAn9HLxYioNrGxNhFugp9cPjs34Q9yc87RpEFjLWJe4iN4x47xEt4c1KKeFNifOK
ghojOUDETJbih0CeXQg+Q+c7oZzo0iRK2LdAiuWQWWB96Oc3QDdn+zl+9FiaiDjhboH3AHtd/W+j
I/ideM0h6gHLQ5LhojifvxFsFIPFrKsEbniakcR0OQnV+p49yHVULLN7rPtjR8UC+i8ZqKUwBwIq
yqBBbx308ecBCdiiPt1ghxPBblyZGnZd7vHur3Jmbi3NQJX6OQi9Ymvc1tsQaHNjtzDNbFTCywf+
L26bE7AqkSik1R0HmD0HXQ95jruGaHqdnWzRQY+hmrQ6qwNDikSlLYpg/Iyxh1MzcfqT+3KMSqod
OiZIx2vVn7kdTWKfKCsARtjRwwIuIQdZox5lIeCY09mSrzyx5dRUiG9UJc/nC7Q9gtrPidPKHeRq
6HEy+6ktoKlP2mgBnJTLhvDc6z14pXZxwt1ZeVnfswHTwOhhNFkVfEZdn07osKL6Y4RLI+M33xEs
FJ842o/r5s6dBPsW8WDZNBfFASlfUurRyL0NEvjTnUhzYEQqRJFKkwgJsTpozOUJDOrQM7p0OH42
D1GMlFT3t+Omsn9mIV7d0skd9BGjPdnE2mnTyppLg2tG3rhCLpqUOLbIGJXL40X3te81jHmSjmy9
QTs6p2K7NoCXFL2hV4J3+RjS5+6Far32GPcncRXW6qjQo5jj9g22NS9l4no4AoiNyzIvoCST2IOY
BJ9HWryQuFox3auogtghhFJJZi1BvNYXeDLU9JxrsT3F8iLi6kO52Sz+UpsijmDjEkPrBevonShM
gIjfei3tDo28XTdIPtPoAqW12+/7FKqB/CiYyMdYOQ62CQzSyT8vkhyXkb81LWL0aJOh0ePoIMy8
kQ9JAAYo2MglW1c+wSocgDBovjEkTrfRge7yWjwG6oA5pWMYmr8U/3O+0IP5v8KmuArnauPMLnfs
Y6CMpDapqGiIuPlAn9AQybFIwjja4coX+8dxuEvhXIxdUOiz5q31w0kMHwUNSrQsFGo9HJ2SwAXl
RKhSVhdW9wYbOYCVQUsr0OnvK1g6hmISEE9MU3D8TWmnlwD0RvMRuc9rDu7At/4GYeZBtP6CfKfy
J0pppPr1cUVY9s5l7r1e/t2V12wO8P77wvm4U4fZN95u8my90RGSRbfbSpCutYlx4DVTU+H20HJu
/0jBvtVKi4vbn+lvB/dszpZ+bfwDGiI2Fw8JjTX4/CUaDPjcUVP+7SXbQmLa79eho1Nu93BZ6LsH
+xiAyNulUDFr85jMDe2Iidg6JHo1fwJRjvhQ8rQhlxUEQMYArwCs8zLetQW4jRdzPHKMD+eTWYn6
kNVOLau9tmNOb8VNL9oyhBK5w+f6Q7kdkrdcQU09s3w1oUWMcsUIq9AIEP5mQj7taYShvox5jOOV
ErJbD7wtets+2cyHJhPnlft4ozFx+my7bRckercuqtfkx7XQdLGcOVUFuvdoafcEmbeEGni1yz63
gCWBIbdBcK/0IthfE8QATaRXFY/CQ9q6PIg/g6H6RoSVmp6HouBm716tDIOEt+eqjUNWoIu2KV2E
yq3GNbCPY3DJ9CakMAg5FNxdb4hQtuo4kuDZdDObvtphbyzLwB3G3AnilsQ+/wDTSvAtkGsKVlyk
UJ0Pq+Um3u+fMY/czHYl5vQokdIm/R1qaF35+Q1LBisBpxYC6weHFTJ4+Ot80Wx4K2lE9mEicbHn
bjmMKdUqTqTBVrJqE6ec5ZpK4Q4FGHSFXGXHFwQpvww9odCqTjRXMt9Id2nvOADyRVmHajtUe3Z3
/MK7BOQGGaTOWr9LPcGRCdmATuiDSiy4WKsb3BoNkQyoDzVreHJWVa2HEOhS+ck36VlqdAkEfyve
dIrhPS6e3dCOsRVOBNEJo9nfMCheeUzJqLylYh1yhTCd7kb2H79a7qHeWdXSdU2fF9lyntK6xwAo
W0y2RpLQxfsOiN7p0tdKeU0zwGVwiBeAbp4AtlxWHZS3YGNN/Q1SmFFSN+VIa6ggfaIs+08BuQid
UauKXWY2COW/YmQnKVOo+7rm9xh85xw+VYAiZg1ksjf4CKiHVWKJxCZYHfBaO+cgckdO9QtdJ4HP
Cuh5dtAC24BNw4Ys1UVtu997vn6dLVDmCbpGC3d3Yusk5qLNdSK+zSo/Wdg4Pb6ryeR0LbPs1PeA
lw50oquDxDMQXlmPosDt368FzgnJXS6bMRQaeSLxE4kURJQa/eneUCKm4OZuJbf+kBBDF72lkqO0
/x3Cvbe/yQtxXZMMt0JhVEeAtkiIgN9uaSZKTwwhwcqExzjKs0EPC9m+N6UkROQ4/v0vD3efpibA
J8k3B/vKl4ylUKYapFjV0zd6EHKJqdiPep1EUvSYuHhVGLrZxWCSklbAmrxp19lfHSZn6L4ZMeGS
JY0e25ftnV89DtiUw3QgVZ2zFLs/gvxctpTrdaDcstsXgaVGgWyxG0359F6m9EYrjFZCi2ndPpZ7
Yku0OC/LPcO4QG2wgez9qeC7/E0KuXxriAB0edIOvMIw1bLBmiRyzJ4FI0cSSimkqq2Y5nw8t8rX
sGh4oZqoA+baW6f1Z3+2l+cqX4KI9acupxImQqo18H8zvSaaMIvI8/4odNftvRw5j55ee7sKrvYy
Eqkwi/fBOGhMSk6o+bLK7URc1rv6lhdMe8eKj5AtY4K87RVi79rCJQRvYuGEE5cWHVwyV/FujpWc
4hnGs9QubC2Tz+cP6EfZDmvYMnKYu1R0+yifUm/Mt2HYxpKrHnXVg4YpbwFYtJ2yvE2RIFlUe/WO
QPbxwEmjwCa2yWtF3iP/gK+nS83XCtoOVCLOwhHtHdBKlVOuz8SSYd8HXLJIc/jsGz+f3L1NReBH
aVIGRL72yWY77GXCwxglBcC20aIZkwxxXw2ShYresRCp+Zw2SJ+4PUqKh8BUcK0iuPfgC8+6r4UQ
0jvSu3yzaCmiodcypWUqAsR+kkoRIMXoNKREH7WazswfaBzJQdGVmYXbYajFhLvrjrk+TlPs8lC3
spkmb/1MXTKs9fT3X1gkdjX1+eYtSNm771x6fGnm94S1NSEQOXsMTI2TIhshVFQdPlz/tk4b7BnT
sasaKkq7jWIuVFUki+AFyo9WH9iZjp1CYNhMzZQ+YiMqHnURQCOrpPdzgyBYjijwedMVeW5bJcJ2
ldkQdskXNNEwr3DbAlNQ8KjhgZL32g6TYTBMSvbC4k8VT3SJfL13WQEBR2EKOYblk2/uvzWXYdLz
88bnriO6cFkC+KuW+NS79qKa5iVktfq1MgQbMWhYup03sfeQXy+6aJdmgBVOVDEnLpD3q/Zfo/fy
Me+TZzBbHpL/5CeKRJhsac/Gd4YTgHaUeRsn9TLsUUIOI6QiiZyjtSWACQVaPGUn0AyVJESJJzX+
A1wfvsd4pTM6rmq/g8wRBFeW0Ea5ObHJSInvMCDYDMtQn3INa4q+EmjYhvUCE9cCx38pnsz0G/6l
HvVX45duQlJurr9Ch8aF1dfx21i2PtXAIR5eJ9bqmhQcWShXX7KgNHwbJo7WSldj/BoW9N9UkT2I
UrGzXACAOX+PmRu5RRdQB2bl9+5bgMnQv32zY+nOwu8vMlfXWjSfbsqizmNYywFUsUq0eCcwfuuJ
cEXQj0ld1O+cL92Y0YL+b4zV/4rpoZhSPN6TjbjSdTruQVXcV8TZe5Kb1VJauzN+Q+VZK60LD+XW
peVlYwahfAXGQ2EVGvJAwtkSpI4eUlOME0lqEFbyXYIdSOWjZ1j6SlVj93DOlaA7k4Rs2FBKcX46
5CPeeX37+Y5svyyHtXnzjhjmGCx8H+hXa/pohTV0gwqib1jCTYB3KG8N9lMud8XodXaGZw9GpUwM
Hswj4T0p9rxP3+y+r2nogHweb5mNvkgOzJ7ostzjMHlzW4tnG31I8OnXn2rLIYnHOchbfx0+L/f7
Rdy8f+RJWJy708BoZwZL3iNkYTqLYV9DNF6zms4vE3nrmKICCjF45nHe1vfROfXpA5dakvPKTcVK
LFX9c+SP8OpG9If2G99vpn57NCZzuWp3pDEoL3YrlHgJ7D/RIaCyuJjQCNUVhYdhM3O3HtBGdSn2
J9Pf8dDYWhgsVoN3rrj4mi97EX70z6NYgZUDtCm7tmrcglCqd5xHDStm80GvyPVDId6YwRNzBhCv
tZF3OZ07SZx4FFjpUlPkeDb545xlVKG9wo56r0lVfS39jwUsX+8pSbukiQ7oO0zpXrnrlWKcJeK1
mfOmntUJiQW2oTAtyK7eun9fFcqTRMcQ3oBYQ2kspp1TXaQ13VGF3c5tJx7DC/aQAzkjDukCHnV5
6Qjw3n6LJKaCdJ2eHfKGruUJ3UFyUhhsvxxIdqVNPkYo8m97QYNO/qbqqS8rNaPj1zx7mhAF48Be
y+lONSX7HIRrz4+YSJnI5vtLAdyWlMfKTZVeg7pAi4E2QKCpAvRU/rS0ZLpUeqHj4Ss/DJiY17gU
jKbmi3koUr5Wdtyjz4w1j1wAFuzMOTIfUbtxrtpO1jflAEOgpUdwkBN7yj8n5fNT/1+bAcukygch
PcZvgFR3VxSHEJ9KzF61qHUQ/kfmLSpkqtWSm5Fz8Q3cgRC5alpMV7UcabPCwXvzy3cyheue/UNJ
cghoqEBAtUbe4seSp5Z8UNgbK13D6joitUxLq9K+5XYtYKq8Zjec5Y8m0sdIxBY/xkbzXnM/SCFq
9Z1uI7MchNVAP3V0J9q1roEqWLPVFmVOClWkWJjZKimgADvXiqtamoY49wjk0GUBMmFDgFlQEjkg
Yae0es+LJuze+kZGqr6a/LwdQzpJEdtxM8/tS0U954dAX3mrp9uIanUG6gMz7BPk7aDN0xoONklp
TVjKx8b7qUGshibY8FT5kdaYSHqylI0p9Yo0qQpxlFesSdwocDitrDNaOmxpQPz1+UcA+9+L0Hh/
9ksvo/21pHSp+jMgW+Yb01cbBGzJ32YYe4e7lexIIy1ggK9VGQVjnHsfnHDRIT2DF1ZFJ8sx6orl
BPstME4L2bTgc58FZtoWEBEzeEuaGOrxaLmyeO48dwkfAgelDsnJUjiaXlgB4CbmpwlnsnnH719y
66JvTSrHqvYkqteAn8dfhqDVF3E4vGoMn0Daz2M0wgtKfKE2HcLw7yRom4FiJJcX5tYFb9reSKwR
fCouhPnmiQAR/e+PKC2/nRJ3AtkXoKoGu6zJ0QxkWE6vk5KYykpvtv2QAFEH49sqNPA91028d68V
5qzLllPS/V/jWd82jUoKboO8oBXOH1kQO9h1zO7Qh/CfL1okRX0eyZOHjGOp7Ic0c6QjYHUaFlCF
imEJn3uvdqw2h5rznZ0q6ek4xIBwSAelsCrAza2pLOeUMtWIYAfXcwra7I8gZSVD3ahLngAVbu64
RHiMnzkDRWvgG3xXRkYCp3fkQJitA7yJ/rBQ3ZDcXjGVrKxQZ1KX6Vguc1ZR5nsPXuywCaR7eKue
NESd+kpxV7g4evvhALM84+CQk+TCHQG/bXcRiQN1zeqetUVqq2bcJ6u2iMwYIyFrTiqBxoD0z7hR
+sGNK6Mj0k6Zy4wzMV57wy+2pZYu/77a3exu/lSZARaPX0GhxlqjHqQtGKClqKyTEeTphVVy9cMj
pQ+dAaGQOb0ZYL3qOePk4xZDYePPh4JcAvoUwNUjBJb/Us75Rh93+JQ15DzcIQeo/vM7GIk99vg4
Hc6E4JW8KWITKWAM8j9xX2Hzlp0p1g9GQ3Yf91l6PxUJ254RcEyxHk2tYNGqpfmu0cLrM7Zyw6ec
qnFJm2nQwt8q5p7N1prxJ8FA4/RABFFaBRHDW+892/A7okGGbN4RtcmorVLOf6YQIXHhtVkHZdvn
Q3yEHKOAe76jixNbFNoqLINpYTrarp6yNDNRZlE4LtWkka8vy5/qA/LwZemkAALt6mUFKC7zfWge
SAvFEGUIkryEuf4yQQRXtOoxGlRhDBm7H3HEYyM+IhW0fsUrwk8fuK2olrcnwa7fWNF2VkJQMOYf
WXgNOBWKBSr50yw1b/wiqiQL8jEnvJEcFCSjCwNPpLYhjRmunBV4bjtpdgSLTRSDcSwi+Vi2nVtL
lAsjc2zPsnfm1lU1NZTKldYlWACNld97bqhi5wscj8V44apwVDKEfvv0p13Gw5QSo8RSQPn/1awp
vU1lGEuPmTc2Hg8R2SjSklm4PFlc/AaiJkUFaj1DvV9rdiaTQK4SLxywaMxzF2CPIBwnAROq51wL
8brzSozh046Bw0KAZ4q1pzyg3ax9YVxAyBnBzULBEUCSAozbAfpsr2XM+t6PmtYxpPqfzteNcw+j
1nW466MVjYgiJURPfeoD1QQCvnjsbTWUTkDCgvbC++IMHy5aCuO8g7w4d4JE6SsISvRSSJhR9eEU
8dVAcQ2TQJXzGnXY+cPtv5LYeVgvcKwvKP8qVgYLSdBT9T/hwHDG2JQiwnQ1BfDToOVX1psde7X7
5rPWzDCy0wnCzO2c+7DzBUkg8Pg5MazpUlAvoi0P5hgDtioOwFr2ej94wgiEmyni+wCYfC+5N4ln
i8XjFnuXDzLYogr0nWntMMFI4ed+qwDV5Y/wNZF2nJG6YP7r3qUIM6yb4GMpxx9BR3RGY10a6cbD
IEKwgkPZeDXp/N9sCps/QCMu/FJXq3YE+su+VeBNq4DbBtHtHIsn93E7D0URXvih0frq8cOoNWjt
ElXBkdlY7hw63dEZ4L2yv+2dSik96R81TXlNr7Cj93g3oj16RWTwuBaNdezPQijJ1CG3ubj35uyX
cq3pG3EwDVPzqClwMCzLQ7GDYJVxTeI6JsQ2eonxtoYrWc/KNgQ1QZZsUw4cugq+25UF7RfJrfSq
0xCOpMsHd18kdJnNhvwOIT0qedoFFekiDLDSwaBXmY8sBxIFfQzphJ2NjxbAQlsSiVFjv9crAtmy
RBS0anHeaMJrOhCW9Lw56PGXTNEdd3M9DQSuH7hWRGAW9MV0R6jq0aTGqyEx/yOxWKvuWr3VK+7s
vn8PXMT2Xp5lXJAbbi6mU1wSEx9eC1y0xk1WuBLGtVeQ/GFNQyNyfCF0pZ7mozcGLpXAB5Wqp/kK
gqaTtKeD3Gs7lFy8sOuNm+DHJtEk5oLvsPs60Z9TmN6YmTq2pvlG3AWco6Ds0U/Y+CeM10pB7Zba
cC5wCh0QsgSckewJnlUFLvFYj1NNPfLWfl0Do2JDsTcDe+pZ58sFwwPK/7Y6mCvYPGWdtmul6/sM
A/vGIhFv709bO5A4ePHKbc+jC/hUrD22loK6+769uIfXQvJi6fC2zZly5OyS7FnY/DzPNumeBGv+
M2PFzIBJdEcc3lKPKNr13nLCG5cnT6ad0YbdWHFUVE4RO8e+24Z0Lqs+NhjWgfvmaMnsCOewGPPH
ejeJzDdEu1Jo5C4dvx/Ncm5k+8I73pJH5aW/fpDPcDwYsg2ySN/aQo9pw/DK3APQ4N7zMf7UFPh7
QQZne8BYN/WmYBLFwfqbPy+WdHU0gLTaEQnpNjtOPUXI4seLYB8zQIpYnEkDVQF+18PrJ5nPm/vW
2wmC8QC3m59X5OldQw4etz8rR0ul8462ARAWON5gf4uXKurLJynXqL1LKGBPB0/NJD+ow9j/I8Kp
hDzz9/ZDVljaqVbUTGDC24Krx8lC8x4gyuvEoglD0ZXu9cZJZFzyotncdYRdownpowbo07aV/Brw
VDhGwgs7V8MP7HGf+USlqQ3jdTwVZKo1fDa1VeDxoc78pDPhjgPBsfmuOLOEqKilHzemtZMrTz5J
tzw3UWWVd80NowJpcnwsoo4azyuQlLpo4WJ6gUOsqqGN+kWoblgj0yRxw+Y3Mn4lqPKsErecFxM8
eEapqeylkeGaTHS2zwl7SrNJPursZOn3Lr7kEp0dif1ZP32HK1qgJWe3AzyOSk66RDUxXnytPAZg
zA2JQeq6X9hMXTFNkc8hO/zRAgClDuKTO6q8qaRqt9Rmmw8gZiPirEOIjCWd8QLTfGdsq6SWlnwU
SbVh8OdwbWWzi1gRkyI+SZgpuQHlftVbbfS4x727i2iSd/QzlMQaCVm0SImUy+7F7E0aYg/z5RZq
wSgFxRCnkXupBOWJ7xcXF28avCsJnhekZefB8VXJgBdQMGdUASOtmNSjsrnKPdPadvscYCDnyhkL
pNMwirHlKezpSpMzXd65RcaB1l4mtxFjSqQUNs9rmPw5pgu58ZKkRw/lvDZ9FV5HoNfgsX7rPXz/
6QKLdB9k9/TS3kM9B8W03JsaYTetkt4/JAXvPs7jwZTJolOPktnbfbNZovrstJ3890swSLMwdszL
T2ltnnXvjIhe6NgqGpCp8pbsH7JrJGh6IF7HHkaBBqvvwM/CwdzbfqZKq+v4bM+tcjNFwmDsmCJW
fJptL6vccyobr0RvAlDL1GguVODLSx3QAKkJXHr3zNcC5qhwMwMT67ajj+648/KcZIO8L05LaH2z
b2rtqIaKQHR34eL3XJPhLKKw7eAfF9mZE4XxSkdhIfOJbmVFeTKA84EKe6mrevcacLyIygAcJ/qn
bQknnHaKXCTwhcaaJWTMQQBBxD4La+Tlg0DElx9KI1fS7HzsGQGqaNfDY3VTUm1FgVznYDmWHpzR
/VCrIcF6OtRDm4R+qk9iqB3CcbBD4O5bU7TGbQz6tzJTsU2a0SWzQ61h/CduQfbA5d3qw78A2VXg
7bGxcbAzLSNqe5pcn2v68aPs7dB9tQlniqC+b8UBysdG3brBcuAf5oUbcJW9Wz5o1GIbUa+O9Lcd
Qo1aqMqsisyGFJZ+9tkizDo27OEq0u9QhtH5BncrxGOuEkzOAylgDjgibYrnmR5AZxSBfuXkxUTV
9QLHqjcxLxUj3ADD5jr61qvZ+swv1bGX7e1zA6hA5GgXSYX4ceP8Pt5hs+/bDkgOt6lTojF2RsnR
/udAFBEQpekzdSeCiBrdx77GSvxPMODgt1aYljmhob0m2bEOjzGSg5sT2gqbLd4xBshv4h6SWTf7
3OwubM/lXGsESmxBTM9SI9cF/UNUmjhAlBr5l1fWFDqZEvCjF+RRMpd09rAEgACi/4PeJv1/m1xH
LBKbgBhkWDQjd5BoF9TaNZv1ea9WuCPE+ATgnlEMgeWIm65H6r3WMwWLhjvwA0dlPnl9yL3ST8gJ
qdMyklCwg8HR3OL4Bt8S9I4WhHz/XSFOOKBZBzgStlKn/goQH5wykXPF37Twb2pX8gZSPhdFP6RX
pbPk/2eIGRwywX1jdhZFWsJcRdwvPLYI7UEdEgMBSM13ZFWMcNDTnTvO+1hBT6q3ZipRyDwbhU2J
irk3iDhEjkddC4eH2FkO54jxQEZtPywXEQDOE6s+XRfSjE8XdKxKwCXg5fGxAlyPDVXuR+VvyPXC
BK34FU+4jUKHL4LIG8nLxdSL8OGwk0RUpKquxshzyn0QRfg+DNfYKsuIrVHSmOfHj9P7tvBQezUx
20aEk+mnNzUW5mW1rZYObLE17c4aN5JDXZp8EkQx7U/fYwJCoAnEJZSmbSkccL6Ip2b5AtyfzvL8
Bm5PMrP0C9iPEYD9si291Q9uUZg2fLfYIBR3ZrWKljYK38DaZA6UD27vHhMUENCz9FZ+l1emIOrr
PUbao4Z0sZO4HGOfdcJj6k9kHuvs250DCAk/TUX7XyMJPBKGXtQUJ34qxwVMrX3bR0d4yrgvBtz/
z2bKfj0P/Y1xD6L1RBIWrBbAwUlrvfyY/paB7sQfOb6uIgKVt95n73xtNPxkQHVnIwCtHHHdHOj3
sqBt+ro3egBsREXQIMxi+q9UMlFSkYYb2XJqPitGeASmTBt+Q4sh38MJ7VMDI/5BLrfYlzte9apn
Qe9j7Of+dBj3Xyb5mAr2CCFqq6ZBegE8pTvmQRZ3RLV0Umi2uRvQjXRvwNjOlo/aZgf+pHoKbxRw
JAndzZbq8jRxlHAsAf9KFGJKHspCL8HDcfy2GwLfkqvRGrEE6x7x8jZV2L965PuheVROLhg+bPX4
zcTgMmbJO2sYhaJjZsLO2/db82B5jR/nJSFemsLdPpZ8FE9Z85Ffrz3vmNAuFUIAr0yk8VbQl+Ts
hsduylZkhR5B50mAFn4pSDalFoNe/Y21bbyhNB1A4Of699E5JIbQ6Ru7oiR5mzGz2swrx9WKim/4
hlhXVOhCWNP8E9LLUmvhn/xRozE7vBU0dVeZ3B1IlGAEFqFkCPJgbeqL6TMl4GespJqHYqTBFPYa
2szd5xjDHzAETs736gz2jl3tLODyo6HwXcVWE5+LzDKQhdyDorxoRBgkT6JkI5qacv0TJ34Vpl2v
AlVig39u7aPGy8Fra1l6oAFKWNjlPb0emBQ2+uQD1RqsyMyF7IAfys2OBeZlE6CCGJwI53QbYy3V
kceuEwHdhyDquX+5YBJJScf+XIInIiQzyfQaYd+OZGXV2rPDgWpiHPkTqdM+VVXaxI4rEeEngxIo
+qV0qnncz70eBcYNM0HVWhUW6Hx8tHOw2JO6OlU1v/khRDln2YkiC4KeWf38AUX0i2UcFQLRKsGy
Alm6sKafkxKHwie+2iRojpaG4vB8Uk9wsFoxy3BQqxWwLxH0bctVQbChh9vNyJnUItuqjBnd5gj+
PMIQwoSWuLaw5ikLAALLFvn+bfNPAslYfWvpvdq3EqoK+FTEfH46+kbRdsayYW/gsbzxlLrnYVO8
DD/xSE4izEp+HIWEmDsShn70n0NUz8DO8AzTzfIzTP25ePnfOlwFhAqGZak4IaQX5rkXU0noHiAz
Pf8EY/w7jccIqbSoXwHIj3Pkmx9mr1EbbzIWNs7B9Nm3daxHg7zE0NtGEmb1wSfHYHn9cYmyIPx0
oK8Z1dJhLut5d/HrIWY1ex88Hm5SlLgp+MhSN42l97+qdE67EeCj+6ynbtU1BvtKRkWVlwcIIfO2
+EJBZ34fJB9DAXGL6uQM8uj/ERX+NGOvECHKjCidpXu/jo6pwbqu0tDQQqBfPqhpsw25WW6tLO5Y
VYiWj6zu5rd7NO5z6FQ0CnV5a98mWBdEQY58XrR5xFUsnLGTET9XRIy3IA2Ys6Yimq4Qk4NcY1TX
hQ9wJa6E2v++uj7omhcCzzFqg771KGFSxfzvGnO4qRm6KQiQHDiR1OU488ruCABUrkvOz07fMRci
hLfwtNGvcn50/qHYy6R2Wt/0Mc4UkIz1gB7b/j5iClf4CVP6iLGKn+lnzdoDEhUDZtufIrNgTSBX
sMIu6lN/7AjkU+SBBnnudM5rqp52GRwyepkNXBVV3M1HID+TnP0gH1L70+kPtQGY4wqaOV+djbGz
nIGQLheio2RA8MKpd/vnKARptt2PRgxkFsAzfISB0bSvpMpymAO+CPI+6kPvWRZWT0f2Kka4/V3M
pr2hzj1iNpPSz+/gMEfcL3V3GK21V4qp/iGK5XNGdwrvXcYeLwRm4RI/RVk6mCXYEJXqNfG3cEEY
7geIw3woEGVcIACw4ILprNqTqWq99NJgg1l3N3urAORmRxSkfJkcl66tRx12gyQEL3FkFoo+aWV2
UwNOizNouT9PkGjitlp8pB3iu1yEWTQQzcy2uEG+1WXXGPoJb9u/u1dumOO9GUiAuT0MqRgahDTR
UrhvnDyS6MOwYsPWoT+MMo2OV8v4bLUt3SXXTNEzo7c6rgYWxubRxTGZFcBtpJH9VxDVLyCvNWIk
zZhvqzKn1IyqQqTD+j/1i1olNSDWMrwU3Y1lYKSuraF3/ezutiSvY5WhgQryTJecnU26oL7VmcMm
lfdNFR4d8b+laXVy5tNMJH2KTywkQYi5Xcy7ilrDBzFUQOfy+xnky9GXphAnU0FFaowx7BG9+Ifp
lC44SdmboTxJ1bclAdtA9G4P3DQGRBEPjFdMzBnWV9t7DcPijq7peG7HYlN+RtO+e1GaecqAhlQt
EHQhd+l3VF/o4ji0DkQwMdt2ynawajtVlBFxmcbpkNykQHc1fCxg05ZtkhM0oeFkc+1cnI77QCkm
p9MYbaYzzEOubkKFVba+B4f2LNZ+A4tOBXcABh8lHOlpNYrJqxHvh9eQb+GczPgkYbv8QHQgNOgu
r+n8OnGq9CD+lAhCK63AvsknGwZAq+NoiEC7nrV86a/NEKhWrWohvL30uQTGKDvwzx2Ugk5PPjsM
1PMFvppN6wYPcKU2wRmUUfDf2A1NJkgug9TZVc3H4FZJuA3FnhSZEZOvvv3Y5J83I1dpCTNdcye+
fIaeXklpxTxgUHfSF4DtQH7HCKJ5mpVNVslICX8Yf2l0ib9JJ3OEhDp0Hzk4SpN0XRjbFotwxeQx
KyBYTQZMBF/b/KKbcLsrix3YkY1cpVsioNYNP4ij39dVb4FeGfNYwX7qhw477tpj0NYkgCsnuOIe
wnF4cCpUgfwAsr2X9STi3HqxeJfqpzxdfGJPGWDNEMD7765mduvUaMfhKXh2T1Nedx5wdcxyp0P8
RAGHzb6IMvyJwKUayDdVBUO2Ai2yoLoQHki0gdE+DPLFfYE0CYjq0DR4UBwZuPagAarJZ3BlI0nX
iO7Bnx6bKLul7k1mHmnrCKX7LlUrNG8YquIYXvVqxA/SuPEoDKLMDhpAn/RhZy/tac0VHb8XAF66
ksKMIYzf5TQDv6KBHuBqdHq+AhF1T2UbH6QpEleBmwJ20Xgc/AHQd8MEweNkIGPe29K976oQqImU
5OFdP+jRrDvI5ywRnIykoeZaTnaVAmTKvb95bk7xi0u7KJxSQcCCRrqM7lT8akX5bgAv8mS0ieAZ
wEkgfKQ/t6DQFlyWZS8kF1xXBbOylbi596ZuJrIwYUMk0gTVUCljX4flFUZbcsYmVqjjNe4vMUsx
uCTpUAx52lT3qVXJyDAoXaQQVXNcvNklf5SefmOOhv3hPmQatxWrdOkNmCLFieOem3JF+zoKDjTV
3836EDlQFdVUDVMDJSFxZOV5iTCjYLTnjdr/6cOtdRdnReQKTnuoVlMxa2+y3rBawxmj2qFqKmzb
OHs+6IIkxWE18T7JOLisL2NQd7Y9aRVMyPl0eMpw1JxgyUexi7tFgKIHF9IRhLIoZqwXkchwmQZD
n1ydBBJds6cjoSCTei0GO39cW0K6UbhShlePsxaf/ffAm20L9hYY2vfVI2if+ahkYL8xJ7fgMF1z
HM2jmwhtH+40h8LwYe/qiRcSAecEPadzozAsAydSOC30pLRtXJh6XfbGwtV9ph78OLXmZ7hHavBP
jkOuBkQzHNwe0M6580k5NSqW+4JV5m3PmO1L0KyQz+2XxEakI0fLtEuvxunrVzWeeAv/wOSysjX+
JetvANFf8W2oZJommwxh9ZnddfuLlV2BcdCSOfh8SUvU5lYGLIb3WplT0+KNKkUTIMhMZkeB/eNx
ZZbYj9zKnem7woiTAKHeBK9I2RTu0iCKQcJ7FbOI3YOo9LhsM5l9K62JqKscSb7sTlzQDwXmaIj+
fRs8MPg+vB9l8ykNlo6nn/zq6ixJsaROQvxyNDUv7kT3UI0pCArUyXPOJtyGe0GwvaGSHtyd4SHW
A/rzVO2SulqPmepnABxow3IgenanyAduEbwTg306j4DfZXgVHZZtYH2FYhWkISl96CfcZwwPJ2Z+
o8roCyDcey7nxAr3cWaxvbzl8UNRHOs9svLbw79ErSzRkRxo8f6hMHAcMYs/07PC8U4n6CHLp+so
8Znns31Ty2zxxa3TGe9/yOlYBLKygAcFtUenNAAx5zXhiE8+4CcKRLLL/Mr2szr0LQfjV0D4WS5u
qUTinejLHXdG9cNU3m5Vj7a9P57CpvJuUaBTOL1iX4u8r6+/6I7GeTMtNslgd9Mz25HxxrZLc/t8
oT0SFcpQ5sALNcpojS9AWimOMbsKXvfMYkDxOqHfGP88+CyYWNTn2MMuDKyveMFwPHcPo6jjx9Ig
RvRsh5S19pkFesk/A2fQkpPDS4Qp6FXAEd/YCCtQWZgOf/NvH5zUYhv2tiKrWuTxfcRTOL2GoS4C
X8waYKopaJCAVd4G7XqlQaWMopm37Xe7aesYx8OWM3jRNoSHx2PXJWn++WtQfAfLxEOJ4KL2WPzy
eLsZkJMTLs78xNalreuCI8ezXyCEo1hnwb+/xT01jmbhZBckxnnK/zQr8SxWAIGhnrm5nE9Om1tL
MxsvLE7nrmCCUBkb+oz9hTg942WXvOqf88tlXZU6IEzer+9Vzb+wwmrISWJCtbRUhiZqktZt/Bmi
xuWpetL4QDdKPIN3jiAjINXvX8XBaZdV79rRCF6i2AajPn2jzFZW7Xy4aWCJoNQOsNfApo0SDU/V
zVWhXW6E5c5yItXEcgMTdJG2qt1ofRQIGsEk/nh5G1t6WN0RpNiwLmmcJnwpGXvO0ICms9UpRNRD
90vck3NeFFp/4+XN3tVQX9ISj4FcHaDtUscVR4OrkgkR4d5PUqx3yXYt9C5zC65XT9ddztpxvaIf
3AULbyI4hfLudECYFcsYxE1ogIFd+tEppNsapNUYQYoqTIlxCcRlnjZZkaO7cXLEUDZjqWXaUNY9
cUkYVgwLJtdfdEUbBDhk46OwbLND7kiJrAXpzXn/LnI2U3DkMXxeX6SBExWOAoGvAdbL33I7/9+t
uUPAzDmxSq3HJ5GUIU4xHdKcHmqeEOQTae+akz5vjm0HcJRo5dPug5HWwOB0nCKS+F34TrfoKk8Y
AYlWluYEzBBHJw1oJjKduXvkLkTK4GsduyI5SlkLVIUKPXV+5GfvUP5Y2CtU9Z3aNN/SrQ43eIOf
ZTI1GpHVyynOUCXdhr9/OuKAaCh8ZQGcEh2ro5V319E/mIguOomIlp1s2rcD8RTQLGfJkOME64US
uPGQfxTGlpbPSN4X20NBowoqkKyuqaviuZ7GyLe4gZLTJaR+hiCq4E8FbvLKJO4WtklPEkzDtmWz
ajPY0TzMK7c+rfMx4lWdX5wemNiykQBsbAOLQJyXi8707TcALhDN2kPZ1zS3TrnjVvXXeNYj6/F9
SecnuHu/QL1YSsP1NbiqAb5d4qN2yUrgGlDMN9z7+aC3k4nYJborI9dwnAbB7vpeTWC/oUnog+9f
ToOhjNj7BI7KeR+5p1qXqhdof4T0T1MHKhnoIYOqzLBV0zDeOh+1jCB7EN9AYaFMaivPErvvOxtI
fcSqcOjVPvmQK01npE4cbK4ICaLOClOElLQh+T8qPDnDOob3toBY6Y+fXK0eIvYHsJ3KHJ8quhMp
LHqIKJvpYduHxi9AgJefaTn5sa9ILRZ/K+l4NeoHjOsmJipLLJ2gzum+zpXxKTMSXS96qGUs3+lv
uFUBT2zkaf3CM6cSNiGO/iz915F53yC0+e7pwpEowwTXvQrWCW1F6mONmQyXi5nQ68zF2ZWmMf1a
d0Zu8Z4uf2jcLSu1eBGOW9GNh3zr1w1HZVx5ugTjzA/ABFEI72sxt0rxKXgyBZzJej8lUDB+86Y7
Ul/56MMmill5xIqrfYTknzXPZzaVFpHj9EMuQRVn4EUvMQz5C2J7KycFG93cYYhyvyQ4+8ViOvL8
NFj2S104DKbCrhQu0s9j6tSazhcBRcckv2XSeK+P9pdv6WR1dt3E0uF9/d81XHd35d81DNmVc/Co
qB9kNeAfh6KCOMRf/7W9sg2DLwy0X2tDmNNI7njnhUsnjE92yqcjlcOuy4TYen1fsWqpigv9iC+f
k/CNga/p/+lKw9Sbih/ikqX/1y+20QTFS8mb3w+EDpKElQ7IYcp7rcQy9s7tm+btA9XgyI6XaVqH
a+u/3PC5k7X5c9xS57sMHPzin1YXMnWNQ1mIe40/P0AqIMH13R1D69Cmdsl4ZpGbC3L0aMPl9fgp
PxZgkgfnZgsJfSmHTznccXnJOYuPg6ZmTK060nRgNcAB9mwgRt82mEH7JdFLP/SdXm0oMzSlBWSv
xFQmhYJn4YwgtIYX5E3J+it46qUWvNqE0/CXwu1zpb/zHTBJDOfyeRqqVG8M6rxHKw/y3CDJrTAr
o4OAwJOW/NrwDpEpgUtXU0/wvZE9+Dhjbbb6X3/o1PWkjyLyFZ6crxJUFdt2rVFNiffaG9DsnUmv
KYtcQmFo9+K5X2hqdqegAwqBQ5jVsecWz9XPsS0l4XMW+iOlL5Mqk87gqO/RTgJae4jvmCqhl33I
3oAG/D4Yg4qIugNrWl+Ohy6EMltq8ToR4otNkONbqfSQTZW6ePtwl76VFWdycvMGJjXngWXMc61K
SYLrf7utH4h4md7wwAVejH01TPAEYyonVQ3UJuuRGa/PncI0e3Bb5zqysWdX59Iyqj+fueWKLg3T
NshpdwKDAG43sFaZrduDokXwOuW8RBijkauR88NN+OqtcGpMzBmhXy0Ar7p/gSaZT2CM26enJ2SU
0upKABCOl+t7UsbqfMHtK6DG4ZN9d9A92RQXZwT8spBRcQXpUuzXTAFUIFkqI6j5PYkz2s5PNWk0
2sCeLvN8nkn5zvweP2+jTKr9cMBxX+cHMr69/qDKvzAxzeIZrf7xzDYnPuRjomxHLOwbmVmHFLyy
7V4pe2OuZmbdk9PpXdcYxdhhf7EuoEGULqh1fNLv2uF+JY53OKL+Z/NzheDyZMG5t6ouk6FR5JPa
liddT7t3ysaXed717hX2YFVjSxVAYFwxuN+IHOP8feTLU9PhrhkW5IM4Lh1vbHfk18q+tzaEx9sc
KpGCfRhlvR9A5D1+DEPoQoUNVbRPYFq3R1IPxfThTLik+bGqRLD8j2Zlz8UhuukeiDzt7t3CnUXb
3LNcjzir52+DDjiWIWxA520ao/U0Tc1fOVBJ05y1Uo4oy1DX+rxCj02GaocSLR2Z4JWPnBto4KXa
Sx1wLdQ+ufreJ3exgwX99MxcztjthVCDCWqUwt33fHOPxSq+pyAusBhvpdKaxJCjvLS720T6Ll3U
v0o0611lFlCOwkuHSsLYrs5oKC6YAf5UnNYuu1opcxlfVKSPaQo9w7hb/OAwanreTZv+t7ARSr5G
5RtKfUysNWFg6yWBtqr3kLK+DhlbXSC1+3TeNGKC6U62Zjk3XHRP4stKtPNzqVo4gP3xkjYXU08o
U6h8cz126SBCXrE+DtlmvqILW3HYNSx9K6/iTYW3KamAe8jmjRrPXE3SpLhkD3juF9jbSHgkZ9nx
pJ2Uq1+ELEfTQiJZdWesFfbPEHg2+YNvZigpzV3+h4C2Md9mWD5/7J7EDB7JGmRqp/2+Kc3urbxw
3nAXmlPVYGhmPU3tQgFSSeCrcWCwszfbvvTZwSW6senV2JjQ2iAkzWgnktYUIa0MszCH9B0SLDaD
UyhiUG3eVR8039yoWNxCtVKnTxkjrmG0QPTiFNDhRGDHviFtwpLXM5dK/PKBXqmRAhO+mjd8Cxa/
wBYrakA+Rva3qWIDAPxyTFaFQMn+HRyUYmxR/wUOBKqMJO8JKdo3MlBCUaVDwAr7/uJUw9bUNl5n
bJ/gPs4zzi+02jNMzEY0tS0sAgfvjD+ODDUTynxEa2UyfFGNvr69MGEmcBE8QHawTWlw4FG7KN7j
ANfFsxQ1ckWxcwLdCrrrBOw/wesk9yAFR2LEvQFSRrJq2GXwqR9HFgmx79Epqv+0cS6l9PLVh3MV
MpJbMbG55ED/I1GfJ4AcV2Y+7qjYGbxLm5NI3TrBTrNfnRJt9secQMXLKwuNBRALYsDu35AB/ueN
TTb8lK0tEaLIbAZmlz0XqBEhq7wWvVQl7HfiNyN6f+fAQWM3st7BLJPnAka4pEQ1BIgsTLcFwza1
RLRtmUAm3t/vsl2NyKveghQhA0LmzKYV/X8dBpmPSNPAh3cl5GKNgIvLZHk6R82+W46JGGPajDBc
Ai4yVUMOOMIJIzHWjTqxs1YIgOwd0EwjXroxNIiYfba7v7jbYE/nfcFL9MXFAHnvih98nBBwH/jQ
Rtk498+sfl0Z2N1GNCxfiz7tOnH3LZuP7LhotngnB0VrPS91zH9R3L61lGLWMiGVuhNJYHvfOOy/
eIRK6mSfdWArKWk4EW3ZGeKUDtr13nFOFz/awZMjuZzcmiNK3/y9iGCbkSYHgyoCvy55/3zE0XeD
wwInbw1G0MM5oQQf4y2yojP81Gvoz2QieMyNMraRWKnrGUS8bImOtP6G3YYGOeqk3UtKcY/uvJp/
Cr9TWlWadOkFycolb8RZzFF52NUDKNah6aIZNtqsmnKTALY964evRznyWSZ1rq7riGkUSC9Cq/Cm
HlX1V1FztAK0v960QNP3XL4b8puJcg00pYkzHQloAdvffABPEX8UOW6gtFQgdveQoyZZ8xpzxRoF
52Q2aUM07NYBjtacv2DX9yk3Sh6024f19UnEhr+Uwf9j9mgqrjclgHgvQr9XmlW8JJ4aDLqYBpic
+qzCbwvxSOT7kg8beFjzcEM3QYGqwtMFmHfEHdXWX7t7cdszD+xpIlGoi7yJLPGIKdOEku0HlvwA
a/tcdjqGnyzz5kQQsaH5SixVdjFAdFoly8d66xNY34V/4suHHCI6hys0cVuyMtiVL2nQSTsubNyl
k77SZix+a7R/P/RBPE0LJVSSC8JsB4wgHOoOwhZV7z7JYXajRWBJ4ksM4tWEcUqiMvOpl10gXb73
Xhr2ZI5Wx3k9kEFt9ivF6iDvwN4JSHk9C1Q9snVahmP6k2bzAxt3of9lXlHORE45Bq9+Su7iTOTQ
wR2GIjtpgUe3IYF7Jb9lccC7EMbRMZadIuWn2BfPw4n2iKTJ81kMS9HxkV1084VsvZJXwRociOz0
D3wO7xXLyUThlP5lx2Hvs6G/PsIBJPnHg8kVzYBmPtZmStk/9lJ8OsXyoLYIsaFoxLtX/Q9ZVIQB
LhJmPq00sI+mxO86nDKvPcqkzFF0Bv9C70LoPQdUlKe0SZzG8VDloooVxNAz5J45PtlR9fVaeHQE
9P5M5duGuBtSowTVxj8NhMchBESwVdZr9KelkrjM+XtWiDGG934QV8wAc+o5P6+rb2VEAAorLSI2
khWAQiq+3zwul26w+w2I1x7cPP0ayEwWbjTRd5MDO8jdlB5ipbvVe8txq+yCFGCh9ycsGgTcFTwg
/gh5hAJZOYAn/qDlIvAnSgpkJgkdiagXmPvpOh1pe/dls5fXBXwJvSOlSU+E8NaqB6l/g1PKTsCQ
P7tCqBSLfqOiDD1KAp+nvAEi8CapsU9+gOnpIRPPFR+hfwEfbF426IeSozoxfPEugw0Be8jJMQVy
ZTJYrywErD4yRq8Aj4Q6r5gM8PIg4cTqHBPVln9pdBCuPMHb8eF3/WDEJJ4dpjTgHG9fpTmH3BwC
v5o+eejEPbxCBLV9+cKyIVLStHc4WYYgDoWpHPGLBrMybsR6odT9F3IKhLGjjpE9TWZOE12KPPJt
Sx/rHIEqmy3vb5g6P79NR/2fUiAX6Kl8d6ACHNHELbzlpyabb/dr1uY3SimUEa7C2MK+VNWQgseN
n44YFuoJOnEnwoHXCtGYb6+9psV7XqnlzNsvi1ENm74mjNTcIm8CYdDw11zQE1oofL25WqsX4iH3
3lsMMPFLpPt+6Xp6HyOOXl7HjZYvAFkh0qxb6pz9T6mxRnochDF2A8+zTW9llxFP1C5GLXHwwoHs
44T3Ls9uLl1JWXLLoLfVnp0QpkaJGMkxJvRSi6TakxEaypRb62ULT8yQLg2+G+6qBQuOH6CuFVS/
/YDAIqYSiZgRBlPAStEgdGGXNVv/by0mcUJDlr/7fBPtBJpDprP8c31TlZSgflrp8w6pfJXVvQfH
rrQ4712SZjMqggenvWSufGSurr7htclA371wnFG4NkXnQhlHydLxeOEW4TR/7fpc/Y3Bs/AUvmFs
dC9PufM0UuHHVyvFbRZRNP1d35DkF1Dyzg8fu4AcfZwbhBLaSAx1SpQqomVOnAcwOiJ8Y8uxVoeV
wWKec02czWk1JtxxaRrDMLUYl4UcPR5QWSNSukZEYTiaSMa5fTZnOVwgQA5/rmLwoYlHoLhrN//Z
/i9IN1lGhClwIqxOnwoGLPAW/JrGfYDWIHlZMFklzljE0dpm42XZq3CFiZdYVY/270oPZsXkS2su
rez6faiRCHca6V+INXtK3L/UZVSknOdsPG6t+6271TWPPZZ276zE4fMJbi6pcN6Msxt3zlmbbyz9
fE8sVt6LExbMpRnjlT4su3PvuyeuD3fNlGcGWK7awVyX8mDzBFyJt1nuntRrcsBvXI9+oXGUFjX+
8HElYpXvp1sZg4vco1CdrErlPsxF8wKjd9JrrYjll6g67XeZISopvQ+KCRcLIcqLAbv8/B7L3aFv
2KKt2i/KOIaNeMt0eDC2pUOF6MejlB5s8t18JB8XZYPmbIkbxNA+dEMfbSFdG5+41dIEe5FWAIpQ
m/HVNZSPKuOH16gn5whm9GSArfJWnbDqYNYCPV3DCy9lKKsLydpEY/bkiChiQ+qhaTddZEqZpMVB
k8EghB3aont/74t3oNwGXCZ2GrTlmhQE6WS0udYprEN8Wii1X8ZJZjhRgmW0wnXK8PDhBYL6qLie
xuLaHSMJcZnjiMyOEh3SjU0990jMAPU7czdhzd5w0c6kWhB/VngB/pbpH8dVsC9mmrCJPBUJJe3J
67KDywrBakp0hMC96++2IgA6g6xROPe02fa0b666m6hjC+2FNSLrl4XUbamb646kDfKnH8SyCaqf
FTLKREVqTWipGQL5wnQDAdgKV6oHCBxqW7lmwEbM4d+Ll2wJyMlwiFYx9MD17dtKwGI+iPbe6fjb
5FecuBlfCJdI+GzTWhXUmMmM0Qg7svdy+6vs24mJoiHw/td78j644ksGfWUkJBzdV0plOdYqT9cS
McnPUbL5vigBSu00UV0ARshgpi1sJ9c7gFyaGSPm+GP+TN8Rry2QheOyqqz2iNzlwfcloZwdkSAi
ClTNJiEuYMZv8W1ME47UHDW+itXiuiQuAfjr4s7QtrkMQNjzVi3oryb9YNO+n5Mnc/pgfp282vsI
vseKEVhMPJYxZwilhch6zSnv+CIQOxv/0gmezRwK0lCL0xff7l5Ny71dPK8P/D65xFRaX1QnXlrs
tKVJ+wX2DgE9bJGiMUuyeVWQxrnEY66jG+WGO8quc7ix4ztAaY6nfP0bfbq2H92LleOuhdsEmYw/
jMASJebBVJS8Y2JVZfwNmD31u4exkeKVwE0U6MQcgY3lmUBgFhW2LM1RXcQsHxcmT6V4OxgPxrG+
j7/FuRPFnPrqPk7JcK4M22RCamcaFOZjCZHBtslympO3J2gzKZCotkVhn0A/RX2m4N4DYkJSENAN
PbVExCastKQ3LNwR2gt1yx5J+aAOWp0tLej91rpFvi948ZxgzRqhoerynx+Z/kT4doUBNEDyTJ3j
eLLFlwr1P+oFQalnEXK7YyWbevEy485Lo/EDb355XDfrfcmVFarZvKwA3oHOSGk+q902W5+Sjv07
SQeKDbhAiEAi02EFXNOmEHGWxbivG2eE7w+mev9Eb/dSAHyg/ZizcTXmTEk/5+aMq/CQMT/d7Cij
0XYFi9jSFhlxZrQkik/PC/KYTIrX/JLQMs/80/VeTUwYYXjZuGUBpLcE8LaL8kNJywW0n2i4bWh/
GC9WfyatOtpgItfAf0r8vuRZ7AkO1/wN/DVgGU0SKcK4D/2qeF+qaVynbZcioq24/uVqVbm7Aqez
YtD6gChRVq35PCYk0aSb9nb8w5v031Sq0Wlx8BPsfNJdWcIpR2S9ZB1+Rxd9oUxV/lWcyNfmPcpr
1ix5G3+V/UXdyHQp7c9VmAeRJWXqzL8UZNSXuiFPpQQPs3xKp0rpC7ir/h+LrDl+wXHIl8QLlkQW
EcSGVCv0FEXhOuXqej8fHKTNoQcF7OmbXh7LWXyq9owpDFCH/67WxxRCyJ3D2eryWC1kepUzOIqd
imCNvXjOuMj+GRjBvgePCtOzPFagiFPlEG5ctLHP2lGAFLFYjDyGPioUUIjZYLm62g1v2FcSnAQ/
oL694TfoTUPACd2Ad+3zwoWeOyq/LqswMbxm74xBKYma8WUOayFf9hGOqJbUPOj5HQF5ujPWk7mO
8HNRpaktgHwuWYS2rAk82OobU5sdogDMlHtfREqzSUTxkkcki+cgGeMUwwQl+sS/NzNzu0ScYr/V
SiB/KQ8tWRTgqvJ3yqOhbr8lWzQdEgkoq2RAJkVoOgI87M14CEb9d2xNDOy8DaIINjXv9xX9XNTT
7TYqor30tVKCf3ycXeUKTX/l8yxhhhNF5Ol+zaDbq50TWrIORbZBFo2XwWPTmMz2a+k1+jFOScMT
mQqaqS2nmV1b7KITpJ3+N8gUIFMRGQVOH0aRgPQJ+laA4mz5UFlHbF2jWeYHezx9fkRnW1j+bX+1
cy43hQTPH5oFy5894XuCF7knDSFXaGVzRplkVCQ0dprQqy1AAuUhsiDNw2rkiT/QSt6r8mLHLLhC
MJ2nj4k12HA7j6i9+6of3b2wcj+ifLX1bftRiWCEjThevc9EvFN7N8ioumLGCGpPFdlawS1evEAZ
1LJmHlF1uCJrUA6HURntbpQTj2hjVsm0eboycMsOWLA6i/zskjTXJ74D15gacRVSdbSRQIpJ9zIo
FgqrU0PIQ+IIv+y/y7FNLSFtyDbM1iqr7PrnHSUVmx1fO+kjuo0UOBykti6ZhwaNZDRik7FunEcz
lpEQM6tdlzWzG46EvgQpTDWLDX6VcNgKOoNL6r+S0kWp938S+FN8ElXMGPy8wOE/Pczbs6EvqKDR
Qy8ODN6N5Z+iyMeBMBU+dvATXzR1Ipp+2DbohL34xK4gHD3gyCcZkVIspEYQgq5/Vg4w5Uhwua6Y
fnI3iCBzeO/QPiTvGxWywGFEC16Oi8OydKL5WKkrWeuhVk67tJT2cGOq8DwxQHX2LuVmEaDjxBsp
oZRXBvwvOhnxpxqXlmaFlhI65lAHRuFwijAHO6K7L23JsZu2KxjYDe/IrQeXA/iyc63tcM7a1RTT
2gfPIOsf23RJI22zM5KzP25vRC75nyMEGp2q/pb0C2KaA8aDBThb8z1lOmFtwqY7ScQ4RDfIPoQE
hpCHKp/URpvGUYYSdxh+X+TEPoyErdG/5zyEufK2cybldQcmn3h8C+c8Y3KhmH3vFK7MPwYVNNai
wwX/7ulkBZ7WZrgcgvxEoaZmUZPp1kU1KDy1HWe0BOWQuHIKBlQYNzTlAe9d+gdf9ZsEVDe8qzYq
BH/4eijYnjI/+/g3cbE2aTsk6wJDPqMCSvo4cCAIzfUrstEQHON2g9VpfyDTbCrlTntQ29FKlnsR
i89GPK5Tl1kbpnUOBrAGTCOUofbXRVJM/g+mKaKWcCuAn+zTaYRoo8e3jtRxwJVlgWUtB5cG3dD6
wVRkceUNOtQ3vUw4SaV8OUZI0UymOSwjaazcYWnEkuWMlLwCY8X73RCXFRERuXT1nZYhn+FdpSgu
yL27EwVE2Pr86EPwSOaBQAMKhlLGgYURPHfDfSXhLGUgLTlghGvv5tJTUlM2hJkUaf2pN7pSH8in
Ap1JdupOpB9YIi8X1HEJJetUig4eD0AQrgUCv2bs29hCarkOQVKykEXREEG4by4R3+WQon03pHVN
BIP8ejmVrEhjirqdaWIJ69ZZ3YIdxUIvJVQU7GJC8elc+Z/k/FcW+/y1TInx+Mn+cDf3aUomoaDY
AHWTJMVcSs86i5/UKHpV4z1dArG030N5EawYldMpjPiEt0hUtbjq0jAv99zXHEiNj1yNsrjnI9np
6BQNKzNMZSSUsn4hM+Vj4Rdy9IauxG11rK2CjnrAS84lFKNLCxApYJCkQUK4Pd3t0W34gkdd/4DU
LEZvmMvDVSP+nnm8oJcq8chWkchu1u77TeKGC5ouGV9tfcOBObhWgYY1FbThvJGJRdDcp3/UKIWt
JIrIHCvxRCsEgXe3o2yGIQIzvj6xUnK8spQ0foiStNf3LZAhy5dOTEHdj67MkVkwU9eD2RFG0w7a
5BOQwINhB3pMmZ+8ODEmj8lhiRHMLbtg3aM2WNQaSFQxe6WmWqk8/Riqq0D1426m/BqVFUsTJETC
40UDNADkch/x2UQuugWo0xRmG4KL6zTP8QBLUlsgUzI1ia0KonJSvSxzlRTyYS/XqZASSLcUI7Vv
3fA8WLfe1nwFbA7LQRUdLZrV7alKqkcPVgBIDgK82aJBrzoPnPxFPQ+VNVN8NdSy6HXQSDYbpB0i
gKhNTFv2GfWveRHzi1ELBFNkA0SqIFWJ9Xp+wwBKzdE/TSmFYRLAHu2lE7biR3BOHUD64q0nYTdu
cFiB/XwmToEWMuA2VVICnnIBUk61Pa8CXsbriRguzCpCvo8OunnfmE/jEV6IaDHYOOhPCHc5dYxb
nW8td7YoEo29/wfoZ2CEROC/y0Nf5uTgDuJ2emVJcbFz0B95tTa6mHo1XDuU335ezfPwyDyfRVI/
v13PUYzTj73OIP0p8Y8njeHGrzh9KW95zrL83HJ6ffi9Ofoy2qV/YOQ4+8K3aq3TZ0+poGHEpHr0
tS7EE+9klQUeSQdYbFGlWRLcswtG1TWwGccweUUv/AY/zh8Tt6Lq/KDgn76Su75Y//DODAbNmP/C
I8zetWzo4FV8wrZ3yzAdGRkYcEfSl4kZ6OW9onkaenbAUbmelWwTrcKiUMZIn/xS4GACIVhZSef1
jAW4Fa1+pBANYGyMkqw75Uv193zlsat0fzNaJJlN3TNKhQXVQvtuoFgs7PtUUoRM7iBAoTtORhlk
IHEa1rsCc07hagJtglNxojQGmCRY8LvnKYJpIYHw5/6nIlijunX66+LDNhNRlZ74v7CnJ3A4ABmv
rYBItSSXpZsAb3DYYDP1G/N/boyea6jaOwfg3X97NCgJuMPinLVaAqlx0nvmWkHNmJdoesqY7Lxy
vYzLtSHKXAbGMrNaf3K9yfrs/dCxok6ri5Ps4y5PfQJvthnM71UslVnez46Wz2tdy30ViuuhMgHO
fYTy6DqfCtxTjjSChQxO0+mqX1V2eOX+a2RCpiEdANj+eNqS4ibuDfIq7S0GA3H+DMLn8zNfI1yG
HqV/jE3Wzc391ca+ipbW0Ne5bRB2ufitoyRXTS7oqySw0WgLYY86C7cD92FfPIpHhIov2V4wmFCu
4XiD8JsMB3TqY7j740dtL0sIagKZITH8xgyDPtBWwIUpTcMhdFZD00XZvUTQRebpKFdMxKqBQIBo
xX5U3r8WAcHzRg8svbKlkHhJQJOULBQl4bHIMIn1WAERNRVEnOdbr1mIUe0E9oIj6TVRd0ji/5iK
Ao8s03djMlfYzVu5UtLYOqOgkMePkKnJk0EAXwYKOYLh5HgQHMBhhCWafgOQU4esvqCDQ/Co54Nk
TUXShqoAver1YuVlQrzUxkDfQ+mm1f5C9urYfWa36+WHitNZcKMe2mt0X8XjhmysoJaqYyK1Gsfk
OmDYBxmUDReaw5UxIxtNf00uxYY83UEbKfRLgx2xu9hGtH1XmNrQ3ZNfpNInhFSE1LvB2Rn8iepd
R8wfZQKZMZ/QCnF9fDPuVIsVrF3QBOhOCtGjo9PmJ2vuCsSk1nLIdaqB5kVnKCZcrA9hn6uPfeAf
emdrOoYpeAZa/AwEFQWbM9NQxot/Ai1ou6Oiv0lSIpTEH6mwZc+w+7iLfcwi0TNHR2V/+YpBLmR7
wObqc9lWndtB9ROe3FPvMA/N/3IDQuhBhuBjCo+lORY/BsUxNYkXFjtBMJC/8C5owUwZwHL4EPtp
xw8ZETaAcKZYvdbktsyuW5U1PUdUW7gf3Dn1iSZp9WybNvAFt5kZ65yPGeURQRSWA7wigImET2N0
UVWXgXL8Z+rEXYizq2ABjLd1iXO+GS2/JJ0kVZJUUB5MYy/RCsxSI+FogP42CvFGBivXEIJ078mL
7L20Htln8PSBs4weXFN+6B1YPTtD9p1NeE1P4XcgsX9bbaDbmBmIkT4l36waIppgHeNF8Ce3aLaF
H0N1TJSbvj67heEbzsY/7BL4T2k552qVtGu3sCC/bGcBY9KMvtU/OPrAnJKzJviZBd85RBDQ0LE2
ck4NgdCI3se61vutp82UXTet8HGO37eVJux2ny+xwbBML+KI/rKizSAtU1GAh2kw58xwpYWQW7Wa
5tygcHiT/kcF0vN8Pzn1IUdN8GXtvGObLZ7Db0pUZoloFR7tFA7Hy4gUBeRY2Ll6XAlHiSjt+rei
A/A3TMtb4KXSCYmGDzXBQgq1Sp1jjqgBw2DLVAS7k7NSHdoGJuxvvvFXPLOXnzUSWE4bCAQfVXSC
VspWnuLtiZ4rUbvA/rMSVBXufcpWV6fVkNQ0P7BtQbX2E6epv5aW2cClETEHiKsCSybrLzQf4zjO
dYtA8SySs1HOZX++1LvQUOUU5YijbcRyDlkSoEvyD+LiTd9VHQUu/MZIWAa1s21lND5oZZ2eDllc
n6CkzuskDakxZwmVq02hLc9m8gOnfKOxOUJuyPoghpFm3o033dTNy2+Mmotbc0wVaak5QKBDbIti
cERWiZi4rYLG5xv2Uis4wlATE/Fr/77dH9BhfZaFm+U/lg9V1+3032X9uV4Z3iCiZmeXjBXb73Bq
9ldM+zHBISSHcyXwuXwqImb4RO7WMdBWnkxHif50uBlUjkt9KLt4NUZmFh7ryQqe9759XqS0JgM4
nl7JfeLuHOOUNt1yrNHRyX/urwHQmXfkkQbKW1EsSed9pD7BFsLeetCLVyFUrMA90sQegtE9veMO
h8i6jvsOtnx8iaonC1qSNGCiRMeeaoRVkCtoisbjSJC789ArH4HQ8P1PsQ5QgwjWf9uYhWFCYKIY
TdBseX2iRjTtVc3RDCZ04DGiScAunQOIJz8HzmCZOnrAi/hYySmn5IcvXWGYO4wX7vPHWAVpGXRw
u0TMD4mCNOSVQyzPT9Xxn2gY5a3GxsdKJymA7PxStdbTPu/FGbWe0JKsfce2Qboz42CVYd4vJ1uy
pEzc7MipotOHYihV6offiblb+x/LY7+eynboXw7RsZCKebrGnMzP4OqsCw9m9k914vxh//m0jrro
G1yQg51cFT2I5+RARNknkOrrdjJRMySKCLHqqeRwCAm3aEHzQc8T66cefkH/WUO2zhE7uQXbiRkR
57VPTVNCW6Ba9w0ou7hbafEPOgLB63sPRDySEnPvv05k7iEekonIk7Oe24/KftbIAmOOphZxULn2
uikrCRmJAxis15sFWaLZtYSMjD5Q9tEnYGB+Y/+OwT7lJVwv0GTddBCtiYBOQQ9IK9pSRsjsB16n
eTSRaoASCPLTxjDteLwG1t20iyWNojgXCAc3HsDD63ofK33zfXgricFYPimiF2FaQu/u3JamMqLE
GlghhJqKS2I5SCm3A7QIYv+jwjdiI530BL6fMXGLZXVIGIhZT6MuhIG6T3nk6hyMztY8iWUhr9eU
OcWAleb/wQZ5gM42jneexytiUR08lllMmvWwfoOHAMQhIS8iEk0kuNlsbxN8o9u5w6QIjfoO+cbb
f37rSVUEGyvquLgco0gX7wTr8rSGnhlGBqLNtgXPkxibj01azgU2BlfJFYj51+OI1HjNlVX1hBXP
jy3lmV1jDoczVXhMJlCatwZZJge4+Bo8n5e08ZR7GsVvjqqbeokuymedw+O4nnbTGhqt6sRb3/gT
Du/YHuymd54bYo2x2A6jjrZPh6u36xv5d/66xaxrzq3E1tuKhNNGRXLJhvNKflOF3y+HqPk1xBsZ
AHi1emb8zv/YnWeONKTeSpBt/l2ZeE+tZ8WwM6L4dGENPuS6KW/WxEjnvFxxeZNl8FphPhEvndfM
MTewdgGgWwEPZTqhL68fIlgDvD0i4agkwdCTlUF9hW7H6NuBsc9N20+yibBj9ziwTJQrSfpGm3/i
lqczsmz28WqQ0qaS++RT62Yl55OLNMSYAAEVKmfmbjAGqiNShDRte3yok+xb9h7PBUKAKSqtKUty
R1sxO7YSGZgKXjM0XyKhKydFtGNhZSPakDQt6vIsYeKDdP8de7aJqy3SZp1H5DAY9uqtuxLU7fli
pl1g2GgyiNE3S4TpXPi4eId08P83UUaXblVr4DL5o8X1H2P2F6TAJqh1S551uK70upyXuff+Dtpm
BcE2drA+bpejHRj7bvD4Y/e1SYIli+8TrttmtKl7/BSj9FTMCOCz5/03gAqd+D4bwwid9gl5CScz
VppYyGEt9o+DA8avPbQLO8DUG/7WmGn28bXN4IRzmquoX2IoavQrLIkaCcpzIj/x5Vs5wZU8upGg
pszB+HFJ/1Fy1xiGF9jNWWhHaw4nik9pdKD/TpvUOmX6oW0C8tmKso8jYbaPSpkw6fkIpOuZh6dF
qLViutVBfHpC0zfuTV6nEQAttJ894EIZwS7pm6YpXLbf0THfTyhKkfTHjfInRQYdgyJi1NHkt9LY
UgBUpdjTxi4XtiTsDayZ2DBxky1yxt1nXREdsgLoWwbZsWr9rQUJsuOEHtX2YMGPpuriEIEnXApM
rhk46p+56zUQfFlPrqygiYL9KMGZjibNpn3I//5xSWziMypuKwZUPSDVjn64TvFK/8gQBFRDGRqE
Hn1E7Pe9YzFnJC/ibktcO/c67bMQxSq5BEpxdWRjAYAsqAUcL7tLaMSUKL+gS14m6EajMDE4+dtW
BCZ7JMFRObPsUyeZtf8fxcELgmf31R7Cw3w4r2bkhBWNPllBLK7l/mQZK77t7OGE3lxergg4QMYP
VDhI5qJ74z9AUqM5m6sb/B9sNLh6cGUt1hMEvhWRyxUWgl1OXRX3c8+WYTx6OhH+Jb6zfXA6XCcS
1HPj51k57q5Slpw09eIn8R1sm9cohE8pkxl/OTyKG9glqmlV8ez8coiJtqSo4C2rRscNcyFAQh4W
P33s5CprvtsdsMjxa75p9LQIXLHElQm1uSvinmkMmqVhnxz3VnRRB4AW3ZPsC8MPImgzFvdafcN1
PxNsnWPxEHNsn7nGdo035akWcZFzCTMxqdGt20sEkrPt1lCFPlq478/jlbDUpEFjAptRpXwMn61P
Ntp9WF/TNsjgoRs5RQ9i/Fvvbetk1z639t1kKNT52lQZcbJ3AMyjCryC5eBC8gPSZR47qzaPPmDO
UCsa9vHZXqkkZiacAZfLGkT2m+Z0V35b+SlxLYO1POoHRnu0/9KYgw/f6NNzpD1wC67ZYG9xUfdS
3QlmETmfUxTUHweTX5pCfXHx/IoAhkfzuCUb9J2/l1etEU55/oNKwZRClzodPsrhjwVOZ4KnCu1y
B45h/GUqiy9l42Mzo0oxm3SeTbYpokLj5bO+EqusnLlYn8/Vh1XOioxTA8g6CQE2WxOf234V7f0x
VNc1yju5wfuEP81NvD/HXYgFsBXpc09nYB9HzR4RzHRyzCzgCWxcU/gy70Ft1u5GlvqO2HZsYP0s
77q1fQimKxlRJHdmoxv7ojUi8DQzWZR5bjqb131T19Q0dGNdJK+Hxv8R15CvTjClnAxqbu7bnCyx
In+bgEiHRH4m2PuAkfgpcGn7Xio9w08PUIm0hb1unxshC/y6/jE8gByvRJOsY6BaGDQeoVN1ZgQR
WyBefO8M5gLZEbkKxz7bKKXiQNvjzcTEJ6ObV0G0TBgu7ao1+N1zTXdxXErRk/y4M7XD1nBoy0w5
PgdbMD9Ho0gw+Ugb2oFagzV47MwKGmDQV5HU+lCbVOSSPz2bE6sMPCXh8TW6yhfQH3zxALOnthz/
T4bWCFuUMFhS5lam748I/SwoRLCJc5RKaBJssnzc73ajyBR3fSRK+NbP5lYukkjcRYaOMfvCmHM9
TbxIIVodM5Zao7bRGREpifbe0RlGzE8+GEVRA21+/WoF/OzqkbHrJRfqoRNSM2B+kZ04OGKtV4T+
C4+fHyn9W/X2usFvJXtS05ZjgBgSvUK7VMs/AnZN0PNYofA4YxKJr4RgWNz/VopZxtaG4sB3KoxA
KRjWXSIAO+UAYOeNr/1Hv7AWFX42w4ykaCJ5TGgeDsRsnn23TN5lEsiYGoXo2abzGLvXkpZHQCcX
nhf7HUXylmF+eoicqmqKhQV8Ff78TMgJ51MccZ3aVNVi5UoMj76VCYWLSUX1BCTbNFV5fPoAjRze
XsZX0Vazck9YYV2yGlobzMANbTLlK0t4qhSu1OYDGkCCEIgWQFR03wMKVISG1Ec88RUPZVgjgGcn
6yIrKDvUQzAWB4UHvty2ywzu2tLfTRZYnbF40UvqCse7cE3klPIdzlgpLE5GZEQDRgpSYI+c9Sj5
wSwIF05/dZgg39d0Bgc9gxvd8Q2PSiy0IcV2BXile//EP9qH5FNS/RXmj4pgso90EFBZKEsgf7tE
80xO4oaUqaA5wDI6Yk2Y8ZdNXy2dUB6PmlmiVLrtoz9eSaU6/JHtMe6LfA0rB+B7xTVy0/jnU6gv
FtbhEBb72Z99OJynN3BuLy2+hCUlQ7te6+a+XH2I/IJSVt+9XL2lgWKMaCYdztjEp7M9C2VkkcqO
WLYHXezxqUGkbyAaqDO3zmA/yujznOhmug0uT6o6joOAgTpWUUmo75Lvj36wj+g/5dDepM8zYkZf
EuKaVfjRherKUol8K5XpqDakgRL7srMEu5azWSWH5O6nLUXy9ifib73u4yu8jGsvOgiUIPI90sLR
FIt+J+NxGmnzQMAtqY0c+DPcc5wGN1lhLXo//cbCXurU3AdS2JOH+Yfh+jF0fzCDuvpFVt5aPF9N
9DEnxbzLyWgH9VMXqFJhspaRVNl73bSnittMQxAqdfVOy0n9aFjC63woSVSJNSNMQn/+QIzl+ARR
9k4vLg6NHd4lKeQOFvHHQ5D+m3Aa3ce6FDIx1K5au1584d+EWPDEaenmZgQzKNiwT3OWWdViarvb
ik9ytMXfjOksnTMWaMBPpEvgbSyJUl0D9opnKWP4pJkRU7FExeK3MkCCICcuGetY0z6JhdFMB0M9
we/Fl+xjV678pTHZNFnYReducQBHkzyPktvqZoiTDgJsrk/AoeNDRYdSbkndpt/9do9vXTJG8YPL
YVbW6lzXj2eoUGGZdTELMS4v1jiJB7Ofy6QSuETqYJDbZimxzjdKb890li6uvoM2U4Vkjgh1b6v6
c/Z+PtrjIXFN/U9kJ2BSlWzynIkRJnTdLm/FJBm8YP8W+Q93CDJXZCsfzyhVdWlw7w5AXFw7qerZ
2jTPx0buF7KnXB+DqTMcQSQTvxpKvFwrvg2nlrCJWf7kTELavBd9kJeTYOuPfsu4iWD4i91NsXpm
/lw23oDmC2qJQn1VS8HGAfpUpiN5iTPNEvYldSRvXFNLT85qwMZR2jJxKx5nDycPEeRzxL0pQyqV
uW/7o715pwlsmg181zNCyODMPBMo28JPvEUX4CGdqvgQqQs7UCBcExm99fg+OzyQUjdyDxBx4e5E
vFgCcTrxr7ML8LuwxyG4fA3AWxppwtDpTpF6OFTL710QlW+6KvUyU0fv3IXUyGM7tpVzYag2q33K
0SM50/yU+Xyl4PgbcqZZDO+pO9mRarLylYiULW54C4uW/1AXnhz5Xct6sloUv8rPVGMwVTy2ggta
i9EnEwe6Ld0hyio5rv2WYTVdoDRP9X1fobmR3sQwq08VDwf+1+NsYasJ7lj5QZs774bC/EkMxr0+
xqE+7Ndv0+2bvdKWVLsKjo4cw7NXQdP9UjpeHaORONxNfij9rWpj1JWK7/4xqAeykqr7BN1Heiny
YHcCF613WfW/O6qLXW3k5W4pN+S7cBxTRFrjGaOs8F2BcOAu5pfUSHHgeFpbmKJVKa1YEyM/qvMQ
L2dZGg14pvlnflsZaAMjLmuO6trBigzRcRgUFAii5yyjQ2ek+nEGWrZxrCIrnwqDew1lvNxWdJu2
O653P2v6WmqVM0o8ddoqa77teanLKJ9XWRN7CwlQmotLrU4VCArI8TJFg3usTzhEv/1bAH8mVY9z
OR4DhnHmZZ5u4U4k1F2U80n6fMyzx58k7QMYjraqFUVAceMWxysDLMq1zXHrS+brSYJMQV1ZOAwV
8fL4WnKFZ31CEi//lXS6lIyR5vq1QoB4PINjoMRrQqKoCIOD/BIJ//KBp7KbslOVNujjuaxNf8SH
ewN3pfO3XprqGdDHKngyu9MKJnxIGa31RGRhhT6nl4tqQExXVApAkMAaP9ActwMpev2dlf1nC0ck
nPIujd1me8jDSZCiDehz+G+dFN4iEUzEJpu8x6rbGwmP5FZBIfT9PStXFV2FeiYI97Djojr6wA8+
RX7d4nq18G7XdTl+7V4SCXUxS1yT4dt4G5jQNu6WRCz2Ug38/g0Q2mLg3PdOHKYgUVRU1X3E8JaK
4ZIxtHR5ixYweNewqM78lfUA6kg6rb6hmy2+on74PFBOk5rbVTNDTZsAuYdptdDJNKxMb/qhRCOz
Gl5gPq7poNa5DF1OF7IjVSt6+2fwZIfGPRCXqXez6RKcDnwYse4/hGKaE+qzwmcVVbtfbK6e2iNw
YHodIEDpIjqikMqAYP4HMMJxuONtRHK0FtHm3V4OsbpC1o5kwRqzdeK34UjMwYNkMKw96Lq+OCnt
O8Hfx+oI77z8NdmQ7rO7lNj30LPtdpBm+ZWec3NR4qBOXcGIirf4IFm3rKznXRUrYlZt2Sq+htHM
HrqhKgVlfqjj84fYua0TDkEszeHaW3oKC5hGceUswXPW/CnZliC4HIr4s+nsJveHs02z/q8kgBmT
RZ8tb9c5/NGDuMKAydlDok0dQCEQnedeuivQLwLiFcSD82WztAx3zwe/NKfCHNsrXdChRsst60iD
eIDTWl+SRAUQR2hpQmg45f03PRlFem0+DWHFbdOrLvUASybND80djKgYG5uSZGu3HjTzdb+ZBrcT
GAaBo4GvT3sAUHTL/N6g75IMbsxj3jEc41S9oYb71I8UFyKmxRDvbelXE7RckAKazm3jRR8rHN8=
`protect end_protected
