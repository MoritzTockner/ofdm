-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PEx4kn1NLW0xFyzOZwr7A5Dwa+szk93MRGoFlx2gRZOXSASeKSVqScYCzOCqWVoOFf+GhacKKJJc
vetERqY5bcETvO0udvENZEQ6BPkusoiZGc9gHRtsV57ezbapdwzCMJejCUDTtstHeims5Q75iny9
KmHoMVlFuu91MLhyYlyiCbxx5/EHafe8s1FMpzWnADlTxKwevgeyad/Sw7x2MdKLmi3TLpM0dJ5z
Be9Lh9B8BwN5LoLpdagtIto9gvhTvdMSMF0fazecc65ZXhBywVJEmndyT3ODOD0YUz3YPXmY4BzG
JUE5Yl4Wj1KsgJcNj7SW2w+Uzd6SsYfW3FGUiA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17008)
`protect data_block
h+OOV511sC9p/eZoa2ncySpkW03bLVb8Qe+7W+N9yZNcVA8VDZr/h3zyXEnMaQdgPvyt54i+Z5+P
YFdgHjpxlFA6J59NCfCHyqGqz8JPid4GY+D3Vj8Id6rfEdtDZhwcH4u0T6rRH3q1foHlZYcGzxbr
gNFugJplh/iIzs9zs2ZLdBGD7A3q1Kx21XOPhQOKPDPRx4Ptx+PHkQ9KgJnie4tBRrzR+RUxVeWw
0BS64kvlYyTdYefRgfGEQbAALZEvzh9fDwyyHNz0Z5MfjLFQt0Z54SjjQa89TsJgn6m8QQ2QXY7M
xw1qaDvgr3cWj3ooept3YwHEWQ1HhNStWq0G1POBZxcg7OfrwWAC8iF+hObtQpmn5fly9LBUJWRK
7Ixnoi8r4sneNBcGi4hWeIOi00aMtYJsy4eHIU5DtIG7Xoyz//+T5t9TduHb9A++RjldG/B/TY56
AFOXHMK3b7Q6eSjbYDtesUY+tO/GwQagKU+3MCxUVWDnBBCF/WiZb5kQzryU+c2RY7WK5x6c+9SV
oOJIjFL0vWi66gOm2X8Xmt3gqUzFbNqmfVaOxEeRKoJj8Oq8Rxy5WLtJBtY52Om79Hqcqn86dOFX
ewtObdQ8/p7rwAZ6A7iQq57+/nMdc8asfGN10CRHdtmDkxGdB+cySR0H0QgWTYxo0XdpuHtaKHkQ
M40AMWeFXtGIZawqBwuX/lNwULRHQbJuCmWxYkZdnRrTwXnMyovOtNrGLaaFBV6TfP4QK8gh63u0
hT2b3UJ+EWmQCqKosifbqxPgcCQQf4xHOzLofd+0g1BWii435RVYlLkg39q96qyOY9HM8YzTYoOV
EIvetZSYpryQ+5Hvj7mXepMT2UcObWtrsvPhpWTaiiAHy2brgwhIKvAsMk3yRuAbFeaYIds5j5nU
UQGeDqHpUAv79NvAjCRvBYZb3j05cKHodNdZxObCs/syKPxcz4B2TFKJ9DHBfLfDkDvC0jhq+P7B
a+KIXvMNjDsTBP6hUpEOxpaFUUWk3Gs3TmLzhJubDOA4HnKWqFBVzoJgZtg+/wn+7Y5HyxjXTPX3
LC0zq5j2dboePlXS5sb825VZyFke5UvtIPkqmDyTfuYWXS84yq5oRRHPfkxojWAVJH/FNw72hU5J
5EOaWK1cIPS8H61Hhp1qXQzpguEMyCu5f7sqR/dXxnpzmVPU8OrcAa++Ya1lpLQ9gZpL+Qr9lkhi
W7uMm7Sclqs9OP3AGMitJcN58of3tvFLcOeEwlpCvNpjr0E2NigyoyyVc1O9nELDJgSwp3xdlnsi
Xq4USoblw7EJfCBJsYipAAgo4j1yT6Sql7iR4EO67piwbdiHJpvJqlX9KfRmNz0IcJmCl0XkR1yZ
88q/aBepnZtWS2SZSMW28MyQDpCR1blORn9pAtGPQnCiAf+q1mvYmhvnXd7SB3tdYC9YwJ5q87Ha
T92wG96VkJa9Wzm3Bzkdt43YqqPi7u0Tw9iD1c56xWbziuxc9QKy5CkO6NEcquN86xV9SGelYeUf
SX4PMVTfGsUkpdTI931OCBQ0JxJEZXXkqkVXoP/swjddXcoojVbX7g4Z140JbG/QZcXfqdlRPeIh
qSCE9vAtQomA2KmgbXbsZ3eOcRQ/bFx2fBB2Bb7meKNatPThxvtNTfbBFBIzT03QS7dC3Av7fBE4
EV5hH8r7GA7UJQ0HOm7pjh3HU3jsu5Z5OVhIxUMtB8SxktSzoECyk8rcbpK2LWDwi+/mkuNvMyyQ
Q3Fn5bLUB99oY6cwNxG27T+0gf0kQX7PZ3G2krUFAVn4ellDXzLf2LTCW87ouZNJYj/tIjlGbDDj
aE2BHn8pjISAI6Zdu8V7YgKf8/i1O4162JnHa6TIvec7DcQcGMcg4J+MrF9SOnHsDp9she0Xl3CF
KzDYsysf7ySo/74NtBV2uld6RhdtCKlo6OQP7jrnS/hrVH15p5D/6/WyuqyH0i6StF72Kb6CsoAT
OA3rc+hIpCmmSt0LLxmB+qQiD/G1+RftXk7jCRo6r0tmDRdmP/2K6l80ivm3TCJRqZvluWaTf2RE
kuG17M5Z/EVyBv35V0cLADVgPwZyNWVhSofRe46J5mRGqjvSkr48yOawplY+98UTkGMrPo7OP/79
Vyx7JxdcyoFtx0J5N/RtGFdUoWhdjKDHnayyudzxjM3W6ZZet6iJrTQv+g3MAA/BVa4Fp4TYdVV3
cdHSdmEoW/WR/knfZb6wF5ojyuWbImDKMEZDWsQo4KxA8dsrV9KPu9xvkupleHSPp9b/Z7M84ghH
FA2FgCu6/tZiagjRbLwNeykaXdksGipqbZL82QgcWfWFSlwgjM3R/QQXm9W+Az19NLSuNUDsY7Pp
kq8ji8dTuRtDe/Vp2FygdBvjp6XG9JH7DXnf5XhzL6i4nuLOPJe1D8bxD/EnEj63ydkUpE6dgy8M
TocSGF5dlmnZrxcbyzs1omclZGhVr/v4gVO7/7G+IZ6afddnixuT0PcGTS4DhBLNY7kAw+Ykg2PG
ky6/it+lhNd/b2HSpAWPifRKMF18OYClh8mzAj2VMGu7lVPSTC+3SXi29JWBINxd8DT2vQTfFPe0
4d9Flkd+yGaHd3B0/t5Y2NZuvRGxRqXsJrUI7jhI1LN16uA5nkwrA/J0Um5B3WCWpCXYeISjH/En
81G9SxuJotFoi22BHO1m01Ic26b38lFt68PITPKWn8AeGH4OS8U9+HrtrHbtyLQBeax2t5xE5jbm
t4MGiI+aHFQaSNLZoyJ9ezAYfpDgx+v8Zb2Tgn7KEagg0l1YLdREh2LhjIqYrTXeETko8Tufu3K6
JjEIuXC7d1N3dpeHDwS3uqdhtCX9jkzSYBgRqJSglPo70lr0yhdEu6W8r648wwJP/1kBsdqkFFly
oSBqEQvRF4f4SVphdR2zztNbIAL6/ooLE6sJ49EkkTv7j71tlPxd9r6KMWlVFGFq+/auHkZXaNLY
i4P83kvAS0S5pEOr+AgBwzLOIHT8qIEqWiuxO4nnneM+EmfkEkthgU+meCYQxYTpOsFyPfdra349
pK/tWDsx6arjm6ylGZKqvBPf5zrhSFGpGmzCNV/k0hW9YN76SX5KJWFTvgF7Vcy6ELnMq9cs7QiC
OKsW5bsmMJuWeauEyEgcRV5RXfsdUvJialvDzlRNQysdPuugBA9d8E6usQbJh7MS7uqMp8obwmhe
u4xug/0/HMCEziYLdJU0SKDsY6fdzQBsIHFOYlPCONy/JJjMOkawIWHP7kUbuUXxviy1E1lc4osi
tQyY6rJ+A3kCdw1Ia3bxxwbZy/temexrAPvDwg2JFkuDAGHCEuG9eOBmtF6Ce87aSo4fKMZxWrr/
rpc4HpLfln90WGlvp7WW9+gb+lnBnTVW67gUyzjjLqqwb0+w7UpoYDONBLovr+7gXNA/abmXfIc1
Zf3Mqg/ziX1Tx4pTKX9fFDLktetmMFskztCu8VV0zUj4o3ITe6rSgMMlgD7U6CGyOyf5vXCmSdjU
HztvzO/81RkvOXVY9vpriaLwXtpSAQceyw8YeCAS3sMVZIT54w4SR8GqhhZRXuDMLeIdzNY7Gq+w
FG9avd4EOm7WeYkkCkemdHlGTZU+jgGm/fUVUJSJXKBwqFv0/BSDOUGh880dAkDmqwoUcV9AgWRG
ii6q9AV+nQQcML/ctuSYMp0BzhB+OY3+O+iob41cuhCgMAOm5dxdpGINqk+LMN3+EfeRXBN6Shto
wP4FbQNO6YA1uLqQsf3ZJz0fIatD2dGHtXqiPDpi6kerrWzlYsdJKFAnxXwQ0Z03ZvRFKAbW5tms
SH8CLrxjNWyqd23tDjQrV1geoTHq7XDpI6ZM4fHHHDhZwj6hrg+b1bkGYY71PLLKm/wVJkwDMDWs
lBh+iCkhRUikYvsFI4tPlofTHT92Dsn2GgZ+FhTVyvIqKPPATcRYpkV57D5IOFSQNrMsySniO4+Q
d6MnBll9hFUBDDkyik6VV8EQU79bONJSQtIdw18GGVryGDRjWWUlU8ewY+E3r2Xa7fisfc1cFU2h
OqKhLVnWMm0GLz/F5ydX0NCWirhc9Ry8+yY6HPvEICgiOxRcZYQqN5tJgqQ2syozMcDx+aTiNtts
4QqxESmFskBXreTqPeYDELOfg0cp1xZf9kGJ/MY6Yk6YX8jLQMwyPvrNLj9NfpQoUCmmKhMBrWTr
EV11H74LJEqe3PWQyB4Iyczg8jaetZQeAiYE+JBzfioJn6xPn6QaxYN6Gj5FlV4Wm5paC2Lt5yfB
Ja83dfBZw6lbmRW8baEbSctJ8ZnN0WeRh5dxz4NG7OP9lX3szLK465wOfwr7kh14COhPedABHUfX
T4hoH8i75QKiNjcr8ynx5L+uB2Vy7bIqA8fhPWQCBALQ+nOohGFVWYQSBDqWnu6DFnTKGFg6F1bP
N4vWdkurFs8nkD+7vqq+XA4TFRQuKtcacLNFSgJKNO0h1ayZVdVkYFREDuKFkd+yTkGrZoG4cxao
mRkyV0rmTdMJxDzL8kywSC17YsFqEzn8tyIN4w2bvuAzKOujdp+FT+u36/nxG8qEiP5xKoXa9Cxv
A9CeAVI9PSfNzT89a6meqLvJLQb/KABqMTVvSy6REvNctjR7ESWVSCd7bLGhBRzV0Oh7G5YiWnvm
OIh+cN2Erpuiw5tJYcxUHjOwYIuRwqEFnUhtU13v8otRSKEbmt+T+wS5CrbgYNlbr7yrkd9a/Mup
6yQzwXYBiFbIfhy7iUeLap36RC0oM4zeMZ6RhNVyvKmeaM46Wvqt8YDXKFgP516Bj3ka+4dz02B4
uedj97zJ2hw9kkDM6pckWkb+9VCc5WiBWlLEGrdLRA85vg15Chkeaw/SILgL4PrUoPhApkvwU+vG
hWF9KCuj/TmUAtGKA3cQktzXb0+JxMv38MSYLw+mLk9VPsOe27m8ASXoOD4Sj+PzbB4ntNo1izDB
bQAgGFfjIIiJAfpcu4AkEVr00o/vYT/g8UJGcIW0NLlaTnmxF/SjQBGEu49t4UgjHWqq+6jG8X6R
96EdVoc7NVQVAExBdbNwYUSsDh8QTXnk+tqKBzKBSGKMH/EsxhrZixKU/9oC06iV+8UFsLe7xprt
rwk6ruNj00RyDxnuc+w0mutemWu84QY8D7jFmlRn4CZiuFCEB+1DbCMUgtaecG2KefhTJKiKpXVe
vhZubbXHyB5SLhFtOd8P7iuOQLzrsieLoa+DWf/4Y5kC1s9N273U7/l99zj+J2q5V6cUa10R24RR
8GUSsrBHOwR/QELln8V51sg71X7jM48x49UA03DAJQe3E9QhSeUDDz0kKZhOyJN+SIlnypC26cyS
honX7+wSRk5+YH0j7BcrpwPaOvqFX8a3DImrezh7fn2FCIqDIOY3DtzjubEU9Y8NsGZS4WbM1Ege
bvn1aT0iPOReUz1azoPj02JQZbMhWNQirwsDSzjD1yPTOhSW3TjeMKxEJ40TLw4FJyRMkLR569es
ad3/Khpp2ulpNvIw96C4A8Sv+Cae+weHdD52FHrvTRJ7wXgdn0vWrYn0GynDC6hXFrCKG0+tmhf1
3W9HFkfy4/MzhEeO+CWozplZrmLbaf2TPP2Q0Vkw9Wq5TzIM7U+FErZnyFppZQ7P1+EGFVDebLpm
yoRmasT8Pu+owX4OPcG5AsIMgqarIeRZI/MyxrDh6TDTUB9iQHVW5CyWDvjqJZ+hQuhMolkbXYVP
yL01vBSNbQ8u14ONb8RiAC+9klQODugbNwIsSu/kRPzIZ1IuJn+sL0FYUhzlYbOETswUoFyGSt2j
zpyfit/GhUCaklKoW7BDkqss/ferdA8vLfSv2xqD+AvAVYAc8OZacAF33YFO6hEru/W7ia2JnUPV
lFJoFChtslAIKX2twXDWgTX73qOZr/6usD1vy4jzZumvOOpWBL0fAR3Q29Ert2eDjvUIzwhT52gy
5oS1OpAAP+rL8cTkmVBHJ+jRlJv/xzQ33WsEeiLPOMBDlrIIcP6GrOPgyDGYw2ATxtfK5vbuN5xC
M5XbBQJcii3IIkW6PA0FQ/nllTcmIZQ3+8TbPRQN7uvzMThCcexEuqr+pCdgGf7eSDYawirhWunj
iFVzv8O5KBqqlmeopKeVEe826OP5FfG8c0pQtxGPU59i/UEufaEhNV05EsJ9oTbshC49kiHXZe3b
miE/xfs8e8mj3j8/M9YYDRubpJwm3fB1NkhRoJVd0nJMnEKSPKIDLH3mzIvUjAdtOIz4hbNugoxf
XGa5b2Q1O1S/tg0tODWlZqjRpe6X2sUhwV8UsDSISkPQinzdQJXr+4EBME1FwbUZ2aqg4xVa2iv/
wO4tWr09wbUApXXELXILAGVuR/W6HpKBxXUJwtVxhRGFWLNNIn6e8+jHTUPOSIIl83PDr0S8aEW2
vDYCW4mect+FzOyAFiZXQhUXvKuLngMQAQQ2eJmmmc1I1gL1cK4YupHVYGqEhV9K/Kcv33oPrVvi
eXyWtAJ8E9DLBWFKw4usVmvVuzfe6AQ2X07VbwhrOYeYG6KjH8Nkp46B+GGwvxN1BfCOitqLVonb
+ktN0YRwurqFH+TvtHmOXQ0vmxCFuhpK16yBTCx1I/gFCuGo15WNdM+tvwLqgvVsapKxZe9E6uvs
s4s9LRfO5pG84Dc50m/3jawdk0kIcMTd2x445s4BGhVauJXjvWCn0nSRqwlD4r2+mRF00ooLOkZw
K0pvxy2rFdHCkhl8jXhc2gYb8Kli4YPdpZGZARyDFcKGvitjLpraxKUkP+jWKSGtRtNXqzOHyfac
vggTlNnJzgAKTsI8DlgVAVxvL/WEjdVcKxqDkLt4xfFYvWfZJKEsApaEbcWeEmy2emmKfGAazx6P
wSqlCbEodj2TApjaokruIKJfunBZX3LkbELqhFeIuKoAXFn9zmv1kE/jqBe48cWK15/gYdcpcR8K
zggA9SJF/IPmDJWTO6Fp7WVaa0ZhJdKtZm7T4Y403nsiYNwMX6UpF2Zx4tqHCHgrhO47cicHLVuJ
wer9nO0W0w/RBs04kzHzq78MWHPZHObkJGCPuon0zWElXUbxrlJn5f0TsYZS8c+aRRyTRg61yJuT
RZ/IbG5gVPtmecFEmxvSpVty7Tegs59r1Z7zO5U3sid4K3Tx242J2SMsiPorOaaJcrfHr3uSipBm
hY/xl4RKPxyrZ2mavaAY248ADuceb9YaaZCirVsYO9sBhQYbHQoXgQEt3B3YwB18ZVknY/x62Txw
lMgNcfm4V9DIJaVLp6jA7H+HnpxYTY3UYpJjCYco9fp91nN/jjeyBeedqm/RTK/3rjaT031cXfAa
R6lUyrIhvmWpoT0U7tXPt28SbUSEkIvbLAGAjh9eM3irgFxT/vKhft9X0KH7Bvrc7RigBeMimziZ
qTrnIMKp6ra+yPNLNjp6QICr36hlNz8zKcUbPWIwJ5vEvE64sVe/2pqOrjfujknwt9c3zRRYOcy0
EbuN7Wo8nLPXfI3OMQlTiUahSwc5KlXHbnc6x1AUk2phuH/zMvdwt4iQFzVkwGJ6Z5dytS7Q0apI
KgEgJavCQixx2GIr7XzyJTJNkp56L+bDdxQaf8Wc3bpVG3PH+u9vRB52Lt2SOBRC7otxPQk60VjR
YFcfbzkYkgCg5YlcAfUfkOyuV6AXHLaJOfNva5aD+EovpwXDLqrL3npwLTJBCnYuL6c6+uavhoSO
aUtQHY06G/86z/cCKr1wUY4VwSVYacNBO9JQ0cub7bc30pAmmetAA7+StRQ+cnWGAkz+LreWWgk2
1tSmqh/Exhqy4yePypHxs7kUMt6vj/v6b4ElxpW3Ow69rtcXfddzX++tECDzYvprmIPTYRbTTBl7
cOdXoGfrHQmYCjg4uQotN+hhkKBzFpoWlkIKFVsRLc8p5WbXSwVQxHpZ3AYl1Dobmcket5bqst0D
1+gcI7OT+YYwS+i2MTg4OgjJqTjovATDUyufYw2ItMdV9pnAVk+YOd45n4mww6q84gox35YjF7GR
lPPhyIxSAb86dl0voEYbEgQupZo3EgEi22/wekeTY64KGdpK9xGE0L1rlez+ftJ53I5aK6mLVqB8
KQN59y8tn/p2u+GPl8l5czBuOXNjlLPChnrPOJ64WmIk/m1BtN5DEk9QO/tNtltDK35496HSeooh
rKs5hKAOWqL85pTwXqvQoQuLahDtTudAJoPf8XA6qQFWT9TOpCITPgiJEtmrL+pNUWts0c+crjiM
xoSkNlAgHypakkPgIQdfDHwkpJPwPsLX8ZWKLn6E1tAeww5vDngeu9nskbXr7IGKJJOB5N9Qys9u
beseGXsp19VLIk3mz6iCnoUFzKq5XVCa3+AoYA2u2+7ttlr67FXWYhdtglG28GFqddYqKa7xS7Jg
vO/Dda0+OPmfzzSzW8+LbzKUJwKPe65F0Bnx4R/8HI0qQc+Nq+wljFATmd4OYzKloXKdLMvHSHj5
KZYfpbHXZE73FMyYu6yGJiSTZGhEHDQNOsnczs6/SIQ7BxDhF49x1XwWnaDYMRRl1PmP243zZ7Z9
kfupAmEkMJbZCCYPJduF/4r3v+AkBX0FSJxvnYpS65htWKvCNe5mUjw9Zc8RuxvtL55Uaw605EPa
rowfbb7D/XofE0PNmp1CCwMa27l03RHSjAjncsQZf9Hofa/bEt6kv5jcsosxJirbfg9jRaYzCtgc
gqOd9vwWdy3w4Bbv8TUaMrp/T7PUqnEYDVzpGT8li1d6i4COXDIO9OYjxnwW9tFm0POjz+OYkQqS
aB3tnjeo417647ELGdyXbxL7jH7YwPmXypHb+c/Erd/V02IGhTae2HfjNh39QITy6p83poFH5LmJ
F2FtL5NU5ds0vOlYiqKrVsrvh0QVYs7V6eetCq71R+d+zKfR7FraVFkW6STTd6EZUzO3IHUjYu8L
Y9Ie0it5n/xKCNyg4Nk3jrhGLKk8EHmQ6omZaYFcNg76xGQKYEAhU4NykquWzQt85WNlIQX+f0hv
a/Qm6cfJcGbvrT6nwC0kvbxxxG0+8ktr5CMPImr3kGptFvol18GyRB0IVr9RiScSrvYS3ytCUgeV
0DJVGAZM6pgnIN+AVSQAXWHAavGoeIkf9pTX62dg4UZ+ZNITnBobWk7U+2qXcOft91wFagLisEYp
mH1srVlRiU2/w2MSzq3OJWjkepB2zhOCGiY9oSRp8Mtbipq53A+66bBDQJb4cEOCjHYDqnH8NwcG
2EH1CGH0vWPbUIWPkfpn/Ktt013UvecAvvmJ4Ns5M3Z7moBZT4N4Fb54MvibTbF9EmkFtc264vQG
R+gf/iWzubD6vC/lmbB7cTlMAS3RJjSRnLOLFJWMXdY8vgRzeqGEL1abUUBmLRyXfrZP6JCQQQE3
PWiydkJg9VwW/pQCCzWWASn9K7F8ryyo/RPBpb4JYALyoAqX8MB2mGHQesPJZ/P7OyWKNDfYhW2z
jUpxwnrSAj8RITRVXQPAPjyILsbmrLtMSv5zfQSiWJh620pfBrSL0F4uvgpvNtfC/F8JOoKkzoDM
+ddBTDRENl9AXR/gIrgLgQyxYKj8qdwBhLPphbT2l0lCwmLj3jD+1xdA103UChPap93IHqYdAojK
b6iPq394axfHwGKxKFxcYIhk82mNO1ph5QArTFwIEIjc3VlkPCEYx8EqjlueZiKTsjEubI//hFon
/DF9HwDOVNkZW/Sn0sKP1P0KL414NbrgWgmYEpkJTXgz2/Sd3a3cDpbfEE5lr5g5yFE+P9AJ8m5/
Mj/21IdNAtQiXEOVDKAzi9oYXZ9iXJwtm88c+Hv+6r80X4hQoUjygT2aD6VQBMBpN4MGvtfGzuDH
aVabNk8xvfyoQLAp2bUCQcDfI9FEF6uIy5OSIIHXzR6zcYEJyqmizywDNrRSoe3WNtglk6z4H9Gc
zhaUdqTqThoptXoW7+naHggFDJBdey3wTY/CVw3nKs34lcsyVHJdmF/EwPft4Ax7bLRD5hTuQpI8
j/Oc3YDzTZogs3ynmZJLAK7WxnrZWAQAhfgSUG+ILVunvfJmNTL2Nutphg/RYJ3Cna4GMs3Wnop4
h+0mNOSDUo621gVbu/y5o9QtvOeG6viwYFKEFzaSi4I8quosB2g2+Em9OMmbkEswLKHwpSN9B0/P
beY8Vysm9vNwT6hsVZAJ3ugdwHSqsT0L/RcwGc/g1OZc8Ez6ehxu4oCFnMvthom6Xvm8ZT6PF50N
c6LDFqTCH/Yetc0iyXtzNigXscOPnRpAmJjypulgdU1D2/6E4ICFYIeNK9eXadDSzvJ+iYzMS/G2
ykKnvtcaKA4ba/miJWJ4zvWkbkfzp0/8aptdR8BRUAyG96agoamm7iU+sk1NR95AOvBuwGDzsHCs
tpNruBxAfkKLZgnar6cUSrdJc+P3WFF+0LZfaEXEZOB0ZgA5ZgNGcRJdH9eVSAWDyQvpLk86T6hy
Yu9VH66AOkOlrfa4Xy2wgmaOH52WL6IrfacmvNTD3P6OevdZEKy1gzp7qRHPVX51xpA1BXnPiX/9
mFcFNrQ9GBqAMzK8k2aapqjqoZVLOcKzMsCEc+CVs4CFDQDmPTQQZYE8PaDrrWmMXF96lD0zkSi/
8tqKsQVMhV3ddZPMmb/+UxVLW6+US1FCLzSTRtDjTwfj5RQXu2jwNE1joFmbQH58irF+VJMYtD39
We276kVsbWTDVLZBdFcwbQcGKL5l8kwzl6m9k4sLCMRzhGwQ0XTJiPL1Oy4nPOmd8PUAgNS2aNDC
I99b0Z/YLH1snSUWtvRUD8SdbxaGyKdWS1uiI7kYuXe0if2oASuONYIm/VrZt54iAu8X8k6hDVdj
58MAKGkV1C3YnfsF+SXpFlntc7XZQZP+fstAVxGum1TEkk2KH5PfoStoWs1lgYHoDY/zY+UW8b17
fyY2395sHFxCQwajCuWDYxS1jIfxlZz/egdH6nq4gmCxSzTRzGrgPkRiOkWdnbxOgsTX0TM+/LNo
jofwVUuq9GZFV+VyzWpy0Ro5rBog5wszoxfyn5ApYVGREduOQvGtHX/LfvsCuRcMI62A+eHVsn5v
HwQFJmrM1deTMwPVY/fNmGD5oGLx10ZfH7IMRL9lENbOlQPbNj49IKGilMJeyrHZU/CXQpB5i3JL
abG0H7kih9pweUgtsn4LrL+wDfa9eQoLGKlhUhCY1q4v8vcJD3XZItUvVkaA2ry+F5Ae40fVbGcc
OOM5Ppv6gDrJaHA4Mvf8sfPogC+AC6Tdf8anmT0nZCmzKj1c8xUnX8dXPQHLSH7j2/Pkgp1ZSvrD
9jdo9dZitUgB0HE5Riz7V9gn2atsUrKz7RPmWU2EmmpDBh7fIJ6htEBmzgbPjGIFICIS03BNnRn6
WdarbpxpVm1CkxcFP106HD8ukKcPEYuR2+WdAxQRtmAVmuEpFeX4/Zlk0ti9c81IUCNHkIeTgxet
X/yHW2JdwkahfcsqkNRps5enPHcmyIOhlxE509TBt/2z9qDV9wd5FhTK8/Wmpb+g/G79ItxULegw
pWUEnfFbbh+i6APo4uavhMIZSeXiIH7PNQQOfpCX3hNuOKv4hRJifuUGbHKACtKdYF70QF4/5kjg
bny5CaPKyAQE6pmLKtR9QRA44+U222K7NtS99a+OSYhISkpVrJkbNgCa7PTLlCOmrU9fMfRTe1rA
WaEsf5sSdVFfiFlpUHWIzVl4dC4cTq1r/kFZ5xtMY5rhLM9QO5PEkfgjy87c7e76v74V9quNxXe0
HQY5BUh02yYrZXJLLW0hwWD8Mkov/QutcTxWcg+zUZTZirYjtfUCC3/daxVDfffQRaYWHJSxFxHa
GOFNLCnIX6fIYtSGYXGXses2d1K7PIK++CJNbj/zpx6azoQfl3TGhaJbzH5CD7NTevaRfEdVIU7J
uTzmES3VjWdEA2eMy0/PTzhl2b60dXvoOFU6rLtsOuplCX6eSeGVc26REwTSuJYUTky1z9rzSyGW
+Cl308AJtqfOmHwZ94MhlRZP4q0YcDpOZQSM/vFNVaDGpDB5Hd1SI7vLcD5tqr0aw+gAttwdCgzx
uKpCLDS05xSpV2za6cc9bM3RN2sRKNRZczh4qk97XBbHuoNFCKin8/FHJxirRAqZZbKXrp2ubw3Q
wRRcFgsdoubD9+Nyi4OlmrdnxBu6uGDxsOS/55lmV/IbR+FWQFIrxXipS098kM9PyAThW/ywOTCg
IxUErMNUDkcDpZIn17F8ycmn5aQVX9Xe/KJqX+RUcxhwe2gMXVFk0rPn2xTpH2/qzdTB58tOOtZL
zRBLyu0hvq/fdQOvmipZgYfDZcDAZm/MOYKAB3IYLMz3fHA3IPg7JiwcdEyekludUtsslCIlgjvN
3MEyQnrJbRjSPzqcccgBIXXQy6RCwWYXA1O9EKqQzvK8tTHjF9UKKcEnGRp6fWqh/lJKKwRTGhLf
OKoqITLoWPSkB/wwBTfeW0lh+L++Sb4pH2RZUDo3xh4vBhNT/18g57Qj8OH4eYcZQ+5PRsuN1CB+
o1gzo7EZXoNjOv47B4aS8GHKQUj4jf8Bq1pdKkGGXsftTa4rmJy29NExPeLJXyOC43odu+T6C2CG
1sjCkUi4V5eBHOpRi7cibx/hd1U6B0jZ9pa0oez5boSQzIJUYnMuoJJnrQhwM7nkZgUJArjbUQ9f
v4hMv1so1m819vmaJKeFmjU7abfQ3R60kwaUhW6jpKRWia4bzcSSZSH7hJLOt1Leh1ZE9tSOCYD3
+GKuvREq6+N0NZMiUGjeaLpMiHN7cl3/+GJWpj+APaRYlOp5KirINMM0MWR3kWG9PlCAD9Mh5KdA
QCGI6FrnqC/tZDY8wCsFaloSwPQhFr8dlXLdUQNU8XJ3aTrpvJRQbjps/3OEvt6TwH3nDoX+7h3B
L1+mJjXbBWiUXaM64T0CrPnz8M1jRdRSA0uJWLCrC5U7LCAKNYZCF+hKG0gEIaS4R2gcKvHIumCj
TqUJhlkeDio6uwwgcMOJ2/z0KRYMPq0fvGjfwM948Y1gdt0ZUwFbqVS316vT2K2+Jo/NY5hGySwD
xt7HeiBisak2fEsBNcVkCKOnEdTD8KZaWQ7jSt5ncz9RhCh6DexBkO+J0VNnCEDa9FG0YYSaLs4L
rmZRFT0y0hQzlC+RBa3h6ud3AyBFx9FYqw5wShC4Ibp1bAAnKtAgLt3JuxbhFnXb7n4SOQo1i46/
/dyfODZuBwVo+Qf+s/JST0Ydf05gbD6Cc6p/pRWICnJy71flJzyOC1E+3sqPQ9cuRm0+ijMBEp2n
w67t+qQ0uaPA/WznOn1WvtncIgHl0U+gLHZJhWC6IEKrw3f3X83lHvPGp26IbhB0pZg1iA8FL5zX
cgwXaCiQzJEmr10ptLOli7M0Et7EYDf1O1IRQHOClFUtf99BqJIQDSP/qCbpNPBzisKC6knhv0dy
npfDlTYCGSZAKDqrDRldOMK6pIslOqUHyaDrmTpz/tTOlwwi2LUPPE1GKC8OfNxPqcU1jwf+3d1R
Ayhd0prvcbqw8pVEVRJukC4p/xMkNUe19GEQAMqgABhx6gp9tLU628ikMEEyNCejDoA4nO20Vdj0
f7xBimn/qZecLN0EAY8EloXJvp3wtG0dLLX3LBfRwqvBHCYo/BV/o5+yBU7S9QOPSz5XXmjC3HFp
yS/2Eui8g4UbQY7McdBu+ExmIASRSCuH+y7q8WUDuASWu5/yEdPLf1Joolt0COHDyYVqBiA8JDUH
GdRnb9X2bvVOSjf04YqdttXhUNg4eQISF+v8yNkeW8JFttlAsTj8c0i4DAB0M4q7NjAygYwpP63A
wKHurBIfmm/ocnIU0VUngiByabw7s1buSjleu0p0LnFtXJCC+CN6cLTyDfKmR95y/OGoH22nItlt
EujzZM0CP/jOKxVVBwS7BWPmuZaMszWyZFj1b5xgwAfyODWnYDrC8odSv/qAq7gIUbcOAny0UC1r
yCz3yWqW77fC/sLhK0wc74+DC6E3yOQ4OfK5HrrGAcYjcjdS8gq6+OG5dnaU6vaWemCp48dYHPzN
FCK5fUVApgAHmjeQIJT0nglSrxG9Hrwx8KutuHvhiE+dZ8zpag2HieMjuhsTKzBqLO/nEpZ0BHul
+zJaCFbrAtKbuk9UnIvwTY9ffb2lI5zgI7ouOVCi53sj8u8uPJaHtnCpFsLKnvUYbIwSyGrE3afY
78Fg9Q5+JSHK1n2Y5NKL8rW8Au4FIRfytNLD6u7t1JrjlvLq+J+RNojPq7Krvcu4sh6S7FgcaQLp
dwiJEBnOZXQgS16+w3PTVlCdDFEZ4uW/p8OAjNyn6GpkYQVXjdHP9z/L523sVOBnAFcnrCsx1zyN
JIPa6T9qNfNH6OSBCOpw23DpvfiIn5b3CD6e/6WAwTHuBewntozMxf2wP+cvwHFYz/tkB4v74JOy
yEXHm7pkq4uPKJHhpjVTzxhVl3bAABWWt17349Df738LeUP8T76mWLKYQxQIt8ldwISKIak1vv1N
zT2Oy7R0Hhcp0z+OiMUx/d5eqc07mtrXJHLuUFQTG3Txc0ILWTNDc4NPKWWPdop2RTFK63n0CVbF
my3P5fFr3A6hIJJb/zA9HjnOsHwHI2DUaYXcKXbF68dzs7gLmKL4bv05eTpRL5f5OusJPJmiy++d
OtQOTA+7iqThIxreNli24/2B6VPseo199JxebVmI4CoKOVDUrhRiXaJadCPhw2ZHs7JGecuJUzpM
UQlipjOMXQKLr9kVUq0P9K4GcfridYq28/fAjfxcnNM3pm630Sb2OC4UoKb92ojGXo2+tPYrxrSr
co3lub5CdTYryLsmwI6n4jt+kn6mF7zjkZ5t8RiPkLq0o4f05SSUrxaK/SmNGim66dl8VzSoN+/z
k1PyMrTrqXto3/jMbdHO1+tQf1MAqHlYAd7mGjUYCnoaotSWEQyeuPqm/xDRbBAO/IkaZV1RvRdI
WdrwolU2OF3VOIgx626fhcRrVPbPb5Iha1UBIYOGOf/K+5cFoSlg5sQIx/xYrgqpOjyyez5m/qXZ
9XKvxmbScI65rsWlk+sauPwbgr9AX1TxI36mZaBoxKFWFKbqULbXJWxpj8O21K6XbrJwcxSoALYR
vZkUAJZYW2SyhqBv45wwxeGIJHMnLTWf0I1o7NMofgOgJXQ1nH0NQaGX1MsX1C2e3x1jMUkyKQxe
fAakChTGboGNmt8AupqirkE+I6YkImcbmsLCS8B56YMNpCJohdB/P4N+Dc/7UNh78jFIVaTyIc3P
BdY/uoVIi+f32v0eh7ohsoSSD7jZrJiKzNIs5tErp+B1NVV6C5ToyrhebM02cgvnNQmKHfulWBsZ
NITrN6UqOD21nhzoh4t3gsx3h5ERobZQEp3ErU7eDG2O4X0wgjWXLr4bXmKd6H8X41vHAoDgL0VW
hA9JJD61YuJIjrOwdBbYBLcth8pjffH9IHOu9TA7sAQgn0/P+13FY+6nkKvuooChcgB1V27rHPTf
QLkaxrslcRj+jMA7Ye35iuYKHguW6gEyx67jvz9AmolhsEIFIDdQQdkF2eTeSiIcIlxRUDUwvDEe
G08qLTheGcP8Gqt//3gTUUe6Mb07MV4AepCcau88ZiP3FCvqwdTSsvxZIoHwmJcNgpVZQ4VOBGOQ
RDm+wlQnSFrzWa/pkheM+nnabCIKUIMoLT+GQcKvtJVKry44WRTBKqSBFip4cF/AnKCuKmGZ675K
lRz49FWXj9TY6JqfTdT6/dze/Vsn/dd0arSMOn7On/lnzl7vSDq8WDoImdYp2CTnyRHEk6PSShKZ
MZqoyriPAIJmIfsjdjdTxbIDzj88ozWRx9R42VfY3Jo4KPuwcIBbQDV9MhrJdXmMyxR7YfXzznf7
Hc9WQYaTsMAhakl8jJaWkSslSbeQO8eV2V5u6zZ+PjhvPr4ySKr9NUlIKikQed6qQ8fEigc6dT2c
61h/ooAo7ldjeKGl/wkxEgIsS9v+zbRsWZpe9V0LVHgI9uOyjBY0+2ALk15KLyT6G3W6l+iBOfcu
EBeDrtC2ImbJ55TQXFRRZZMCIuVYwTnhdmiG1F+icsyezLKWUj/0Oq+E+HvhoAVnqJx0iZ6U3s8E
DMeZUmXy54QBkgCrh9bnB7eBDz0HiOspHwVJDoEzq07Uvi1zBtvSaSTw8Pco1fkeVK1AzzMua0yO
WmWeUqO1SpOL8FZdoBE+6Ph6moILy2v9jqhid1mxGSYHBuCXVcwHw70rWBO2q5pB6X0hWqcbVEZp
YmTXPw5uZJDCXQJOS28SUaesft2MghJH7wvOooUtyafuJ8wa6qlxZ70fQn7id0YHoqkL4hBgJZTK
Q+A9PG2K5IDTd1RoPDOFojmPcx4e/1sm/8kV1qQkoluSNReEZWYSyhimoUS3v20T4ePaCie8qTrn
mOtAehv4m/cQhThob9gIaK4KMYmOBzQeOSQbCaGL61DBUZ1xDOxnYUHp1KIsLVb9VZnzdK03tRZY
fB3xYmNV6Rf4eICt+owYDFECwxWpHdHSAyLK2obbuijAB1NOwOBv0X8hE3GlRZIkcEx4jtRLy4Uf
WLD79/S4kBL5Bj4rTy0h1vii6jCP8FV1gQGnkwDm05FWfqjq5fkzf9uvrVajLCynAu0h0n3GxPMb
oGYDSkQx7cxdG3E56mkux+ZBKV3ARaDWI7EuToyFt0cLmkMNDf5CYT4QHzIaNxKScowre48WKkMR
uBQ0DN6AgMJOrZXA2HbnciIraN13SI0j9nmXnJLA+WwstAWC6agT7wgKQwcslwH1kxU+sZmrZtiT
8sDyvFKsExviGFp2qEHa+levfRicM1rMDkQPgPcffyvBvoqJF4LOyy0+8Rm30euzVyqrrwP1c5Of
Yw3Z+hnOleONkMiWwPVzth3onvx7RzNHMjKZZGH1e+yCmEyQdKfdB970a21nMw5E3obtk+k9e8X1
rHNdomEs7IBnnOoB32l3EJdtTq9BgSFc/aYmKvZFYg8ZawyNmKf4iPlRnPgb4yzPcHm9nDcd9w0M
/36ri2tPOeq1fY1v06a+p/4uq7/w3n7IoqmRQdU1RaAx1oy+V7v8hlg4+ChfCFWYkvW7W2WMYK7L
v9MlTvGLYsoQJ5Chk2wl5wIAnacnIn6e9xcpPzGA21HmTQ6eBE1k1gEMKYbYn08Snkzy93xs6WFZ
0FhMxP0+cC8nS2xGL4VPRiJK0ZDRQJkP5V3h812BJKc7h25FyadhCf478QUVRNSlS08algHSNjgw
EJNVPlUhK4hng9rovpEh459P8255gz15z/ZxigZ7RLlwwC8xeaL1n0HGMxtZ8vqzSYaGFtjqvf8u
jqt6ICadZ2zZsCKLt5exaDVo5Dev2PVP4ZC3TjNJzjJ9GCItQZ7sPe+ZrLBSitph+uiocEo+tXya
9N3iW5uh7hjwd2DAkr/Zq/nfDXawxuAI3U7QBnGordp1lAXekHoW7wlVTr76fSQXvHmsgKgKfvIS
NNO7CotxTj8AjKV1OL2RH6flvUnb6W0uWqXsAuJ6Ntu+GtF6326XmVdKrM/IDBhUQYMzQ1mGupGl
pgTrSAHnvHE05ONVLe3nT0OObO4XdWuIzngsBR2cjRButAgMqVYUHbqFvNu5ZBDb6XLYidhWg5CA
/sJIoOotk+xFdFpwC8xsfV6DQTbOaQkmxA7rU/8Yq9wIYkEw3n3/4OguPVCT92LMRKqghITn+Nc8
EWXkN2wp4pQLw0RFDj8BJSsE80O5gVmp8p03XUfHjPFD/AqSAzohFoetV63L92MgOG2PmIjicGBa
iJsmaIJh89nqhwh9MPlYYcL3QufdDfOhI+pyXnQpp83ulG5UoEDnbzUxtxnX8iXQC2kcfZevG9ME
AKqEpcJLoTNI7IZFXetXrH/uht5mSBXEsbozw7T97QYmJfuZ1L9At370HdV974J9tk4YIimRRpZr
Oq+3m1E6t1rptTYhaFn5fggJ2MQQ+nnTwzWOIgE8BkZYCNqMjvTA3LTHEC+kCy8pTAAJhO5ucuZl
8ExbM7VvY3NEurlfQju1cbOSb7D7cUmB4pGJoSlRXriyP63z6YhIpm+OUDb1q5X5vBmikmuIgdNd
et+HjmaEQUqMJ4u6kuFbj4ZVFk3yepGPYA63MCILVdva35G8LEUK2vVVUITT1igmwFmz8VpTDK/K
e7Y5lpPPMfoW5E98k5VN9i538jDJM0U28bu9fZy3i218/SqYzVI1aTeirjWSOlk+hf9ghSkwCLlg
5IPe/I02MzaVKNBSPHhqBWSMUDpwxBbt7L2b4HiBVr1wsFvw+7KhhVs7r00zB2S7+UJtSRtmSNuO
G1v8DfKMjIaWJ12dOxtkOrVoDwlhkvyGYRX2co5+pnR3v9ctTCZy7QZC/rcw5jBbe1qKa2VXsbH6
g20+CaYEALoaHeTmu34JAEkCtMkW9I8S3oruoyQoVB8hLotPd05vCBTeqXdiGhOAYOoOIaqiKPN8
oIXOjbZp77Zi0JPpFSoPT4RM3p6U5dWqkAqrmeBWV03biKyK+1GiLdpLAA2NIdUY1FCkI3onrVS8
lc34bHCNSRfI5+QI9DA1zQU06TiKL5EE0FUkjFfA3G/PxK3dZtrtTTY0MiXWdx6rPiNzyhWbp4K6
2ehI3vi0Kw3O4Jk+jIMUp9YRuVR74b80z4C3JhNsRt3bveW3wahzL6jdKsNqrJcBcUHeZrAZ31pT
QQ3OxLyhN9gn4/Es7heSomA5lpU6rRGMXzY9gRAd4lwMwogr4IqOrD61Q+F+p5vGhebYhznHnMZ7
FaujZ570NTdvAVS86j6DiBcJY2ltVVLZUXpcXIY8/vWNEQZgrbe3uob5sjtsUB/kfiRY7tNtcjlS
NoeC3qz1J3h2r98yTNTwZjR99C6NPoFU8L05ymB+vUeYR0wozXy2ByBLftrUerNA4Pc7ZJJgoIGQ
GEZGHlnpVaEkWThMd6tDHhD0CVJdlzhWTaSAdcQAhRbrwdocjSYGSpCZ+I4NOiIMS399kMdRNtqt
1npJFChFOoNh21v731vZb+iPci8Y9qYGjYqlplfXwKSHhbpZVf6yReaEpzw3jyLYBqknCKpO2XmZ
RM29FNaJWtOidGOYT2aKF7Gs99yPTp2WqFDOqkmYg33uNR9+M6F/eDp0+72J8RgnlXF/uM91LiKk
2pn0Tz64AVU1WkYL8sqdo4waoAyKYd3ZA07Q0hv5eh49Qyh85inyahH6I+cMkbIWnLr2g1Aw41+r
XsSudPVp9Bcz3quQeYmFGVtvMt6WvNhM3tbprYwmV4BYaUNMR3J/ItTYcVG9J3QT/ZZwvXCC/sGW
ME9mBYRp+gX67Nxah6t3RrKtoofS17og1nZZvp1g0vhnoFeGHzI3L8DlXHTR6436RqzncJcH8g8w
rbY//CHpAHljE65GRj5BCBgJ5Ny5wOKcQGp96RIY+Kh/dEVrwnw/K3UBXjbAxL/YEaGPkiCfCdGU
cQm1cZ8MBVOkS6O+/RQjEPjOSMoGptAe7SYZNmGseL8YPXaG+4XzCmTLQVfV1O4A5He7XE8HxLZC
WivcE9xB5YnMk2JllEu58hy/eFNphCqKVoFT9N1/0wbSZOoJD9karEg/+0GELgHY8FUgVPeUhkv2
sbmDHPGeEesCx1/JT7edY/oeKQUCHsdWlbbFxz5V7oLNir9WD1V3mdlgX0ALqQU5OI8Bhx9iu8nH
RSWYK0o7zjPUOtMeatjHeTPAsaRN5EfELkZ9fxu2TkF9s7lV8SRO6wP8mAjkmaSgrVmtGjsSHTN0
YHrhYtQlyyd1MYGk5jEWa94SSFwhmNsHdePWiJCa01GZDVoZ9cKTcWc5oI3Nk9do+ki5OLSKEjS5
0hj72ZFnS320/GkPP2hrGem+tbw8pEHyOgwWrGHwb9DP1MbzYrKjXkKIUcLCZeuoROvzBryRMzFH
oPrI5vsaNwLTt9l5H0/ngSr8YTblWqc5uFKm7vrYK/HEQMj57Qs69xzxPZ2zTDRwW1/aYwxSI2lP
WuM/p8/qHxGOP9Z5oCt+MQfGuVT7tG3qeWJ80aDotSe6YiAHhJc9g4FAihJkSkNz17sQyet7duTx
vL9Tp6SlBdWJlwvGwpqJZvxKOJJkg+jIIdRELxNNAPhwd13m+H+HdS2ZHY4hKNSojwg3Jx2doswA
oltPyTW1ZoHYT4nmvATj250JjxpepNDamHZ8ZniZ7/DNGHKLot6bCWCTjVKwSBuSUkn5t1KdCFWT
FEOpO4dEuRGRBamBKeg6zPHf/yzUh8m9uyEK7lAG51MAaa4diJ3uIMaJSkiLpEkEMYuukSat3GmD
8cY77RvHVBROGnaF3/4pQhGD8A89KSY9hHAmwEJPqSpjUr90KL0LogYYFKX3scssZuaEHYciWqDm
vLhy+9RKtBXNWWI0VD4fufb7taMzMB+l16sxggCahRCav+BL9BoNAcvTeoekZa3OcdeT8NxD4xyD
tD2VzE6c2PRUsYf1ME+OS9UGRyWbMiIY8KaJ4vu05V+56KmyRCelaxUfhbtrYo4OvgFxzjn77+UZ
3NM2f7qrhsZISQJA9np7KhcZIQ2Q+02dEfWYENhjVCjLJ0TOdfG4jRfd4ENHS0sqoTejxm45wDdO
iOvCX4318d4wp54P6N24CiGHrRGwg9XgLpD/giQFwqW1+kuB1EpukIDdnQV0RYt9rTxDmOKlSpN9
MO/NSxzYxeRWRCgQMOJ/mLzptJgudZkKXAzJhmunZrMCdzLQHkiULv6pPWppNLazzPhCQc4ED4WS
hplIksD2uTzqj6m1ttTxpyrnDyeHcnzbk5goQ9qhqsHX/F3YHtdOdOVTDP9qkVjLxu7YtScxFzxO
iijKI5UsBr0EXBjuzJ5CL6S7wdl5fp1QQR3HFwCPIpvQibhubNO/O8O0E4Ji6G4xatXEbY3VBCBr
mVc6/XQyw4YlwzRmClelvC5eM3ioqm2pWDtIGRh/1/PABkZNXCXJtQu2M2m/bvg2OUfVuksQtzLn
P3X/eDVvZlMYt0bkX4e3NHfCHXkvgNVFk2Oyo9sKxOA8MwijtEc4IwXp6NtclYDGmSb6U6bzRG88
USuSPPgGE48UYLJ1u4IJfxBRfXYc/aMdmnMbV6c+iTI2GnMORdmOgSAzH6oLSZ72TOsh0KFEiSJj
1oCp7CnmpCd+0RNJd6aoed+X0MxXz6z8Ip5dYzHORRu+xLodDEdzA/Sf94Z0nDOklop68wagFERt
Epl/MOS0DA3VthOwJYWQ37z1LZO4phyP9BH2ZBUQ7odLmDOmOc0mO4xx7yTvwRmW3NCOyau91uQ6
IciKFO6tRV20SwzKc7qoRMseDBdDeqyuoQtPux17ZkyMJN7ndOSLn9VqettHBkG8dkwWV/GPTvei
JOgvctknsvPGQbAzmXtMdPxZnwQHmWq0EUAwod+G9xkMQW4qN9lNl8c3sNRzCSC8CIAYTf6JhHtt
MTLZiEibmzQiJ7fcZ0di8U95mQbAwO6CROVOgQEoSh6ZW+PPHYU381xGtk0CyNifOSq9IHDJqieS
TjOLZi716n3aRuJ+RFVhG5dCeKdBwpyDt9Q/k3/9/2+kFB7dJgvhtBSeaxEGCEbnTqzN782KjSYG
l5yWQlFc3XZr1pupOgb34Vd0d7zoYYdaVVJw8XyZ9KpwGmuvy0hOJHdKQXDz5p/GKmYp7mB6Go7U
jyrJ7GzGEcuPjZYClp9DHR0FZwsrv9RncPGk8kNFMDQEDTMYfWs8vRfM1iERpyqex9JsanZN2k34
v3ROrqmVo6jDxdzNr00BvUEWy828n45yn/AncC/bpazOHpMstCRBFnkWj8BKkIfjAiChhsmI3+7x
7ny2jg6YgYeUsOXv0gh4JDMjp69z2EnplW+ntB9+B+IAGDqKmvhgqvNwzgZZoaMgA0cwQigndcHC
4iMJ9anxpxueyvps6jSkdkECB9HdwEwZOWCfL5iXaRPLwF8oqck4WacGAjP1ey+vXmrGmeHJBauK
TKLUbvBBcaFwidbjGlhKTPl71NRJKfItCFUOtFLCM1Lhrsan5a+ZM2vL2kGGBaIDm4MJrn6JcP+1
NCvEdTUfKqWuBlW4BB3c47KJ9kY3Y1bXEJhVP6YBDF19UmPJ82Ud7UZxzPMqq/XUmNH04Xes3Rbk
eEo3saB0/uCy4BZzqKSsj9eY+p3z3PQmFToqFMIes5Fhignr6HoQbxsLpR23dxdVcUtr7gD2XGrx
nZ9ZQYhW2D+Jf/QaSqiggM5MXypM8ileyphJq1MVh4Coyg4NJASW18b6WVEuTxfLQEG7YUGL1m+K
Xr67tJtK91VtdIVRvS3tLtqFK0Pno1IEt3wwTjUdCwOZbGjcL/c6WYWHNxJz0m6nAloSRYVxGsaG
Qixh3S8IIvGSvgFtKXz5pmbrFQaGr5NPXh1A4uGI3RQJNHX5kH/Q/4mvgrXJwPUyhYidntvRjfzJ
ycDIs5fJDXblUqntckw7jxQn0q2zvJ/JHtRjPA4jpy9hD5gun/trMZ+MIhfpjMRE9ZcPJBgucZUt
NHaJA0ObfB+z9WBYER5QpbGkFwZa2XOUxx/hTH+oYtVHraj5uxat5H6hIEgq20kQ+gu9ZZIRf5Tr
eluOZrbRTJHq2wAoRd5Mj/DGVZSzCcljX8hwXyKyxwUEl1asUP6vyug4YgfkoGoN+SBHNO5rfrHN
7Ys0KpToAbkV5C7141TWtg0EgQJhVdej9QEaqGHy65lkL0kxxQjrSKjZiHbpMU9e1mm8HRVs8UdI
A2m2EiKA8g2vLB+F6D14r339HUx5RA==
`protect end_protected
