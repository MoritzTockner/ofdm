-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XNr7kYbPODFJUj3KaEx5iI0ExkcEyiqomHZN4li44kyXwq4OYi8GDcDqDv4R8jdg0IQ0871+J3eh
wg/5S3FcELRzHOcmhQDa5rllRPLAVHrOs33hG3XZO+MFCOIhr4OunFBR4o1bTEW+TdzpbAV1Hz5N
Q9tK6FzEeSOH0AitAGabuJCDkyeQmYLSn3l/+1IuBHsmt9zHE/+MeL+6WpYPByR4DZYauNIICFxy
orGeIt3MbQB0NRS0FjxQumbp5cvVaC1s32ZY/ff03/78NRhwRLvrj8gzY1//o0guyqM/hvGmoJX3
F6QL2L+Tlf8TFLTNunSpJtNyZgvBIwwANGbp2Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
idDLi0SmGSN2cF/goORq+CtY7eEY41DKAV+daFeqYp12OkGr9Pz18kcFBKcs8z6kGiRDmyiLtd/e
ZF0hJLMvpnkZUHU7RS5wSfdCxczV5JfQh84vML5MsB5CXtcuiGHUDzV7PySCqGYD3QMKCA1QE3E/
unNURPGHOuHf70aikn739Pl3l0yISppKTnazB8aEW0YR4bdv2R2ZbHsjVGrjNJBG9MYRQPhUILAE
9PP+It9+OmwzdSdYZ1/uaWhPX+QfxmG7UFKhLx88fNby9SXI/yFHb+ozg4dOxYlBAWjVnfCxKxgk
oKlUIG40HeiBH/YYNG5FzBsUbh1njz8rFrG1cm0lrVsU06ycG5GHgW0q2XNHM9HdwcYfSLEveXHo
pHQunJdyZQSITNZAosu0BZM3s6OfIHE5w2aOGeOTkQystBrvt/jxWcoaD04UyVATstPevku39pud
QTvSJEQkl0o7HqbuBgowuOIPBEBCLc3sJ//mKkLHpWEmFA47k5dnkm5z7j5hSB/F9anlONIcoU2q
Rl43xulE9eoZbUMwRps1P/r3FNJA1KE3cbQt5ozcJTijWSENhokNpSQLY/MBr3tiwNemMExK/6tb
IA1wLJ7nq5KHJrx4BmarE+nDSh/OlZvBh0XwTTH9FOBtrcvmnSBPkMyKtJFcMWgstHTT8kqjt3G7
VdxXq3HKhb+PA2HrI6tt/Eg6vI8zaQxXZnkYkUOQIA8ZQYvB6AqMKlF9HG6rWOOiFJQFyH8pk22X
p1yo5ERwBf4lA55WC3RDJN0BoWw+EVIMW7L1bnt4bwra+EQVki/b+VQ9g5pO8jIgRdea/cPkmEbF
GYrdl28IoqY1Gss0iQslULzIIAH4mNCNJnY7t09YUBdgIt/a6JY2ZXpNbqWna7wCgb2EJ9xWefwD
Zhk6pUxiZJrwpc/5430mvAtDuzow6xLkINw2ZrmtDErLSY7S0wglEhkJcPf55b1GFfOoMnaLw3TS
4We3cj7UYp30J9DSyRZF/u2OnxHVzAPsK7vvVOF6iwvqTIfy3yo1q0X2pKLbQkb+r4Jm2YwZHcNJ
gkbEbq23a3igb/LK8hHw9TsQ5I6bSjU2Koe1XO1nRGQkGmbh2OfekQMXMg3eC7zFV7a0xNSNV8kD
eEqOzgv+hVePLWNAH9nzz8SOlvfOB2ecnCOSU/CENCIbRQnUR07oHTPKzPSvaQCZJWBLYG9btkJX
IglBK6B5tpt9KlNlDVXpBjOpDevi7/RRAfVcXA1Z1C4ASnq1mKKJhByYeS7S+LS2QVsHcxEodqlo
u/4CpDnU+rZjQCtmnS8R0S3BwFo89mRQLS9f+XX2bYqYwNcHQZ0c/v2SK7tW9nlB4ANuAZ9tGlNO
Ql9i35aANB3aLDjSQQyqzn66DoVpQSwjaKMhhrTO7wwSDxfgsQIitDh1iWnhven4hhgZKII/yVN/
5zmGxoxlE1bNLFPvsmTlw+Drz/cwXxaQKdwNsmfH791Lz8MR5viDz0qwjoX1gxmb8dRnQ5s1mtUC
2e0Zh1WsEbL2QaYYqm/WGrg8AW3tdOtFXdvLJqzKySj81wKVkonYUk8uEa3oH57hxbgJK4IOaw3O
SxlgnHFsz5Wl77hfefiZbbAPq2+0ClV2O0zFwF6Gob/0Q03ywOE898Tx7c51A1TjG9kXEyUNOhN+
CaDeuE3T+lqtberPVFtPxIiEBYIej4GV9sxVgNnPN3e5jg+6WR9CWCjEDsTt5P83CCxszZV97UAP
nlijXCxtyu/sHtuNco3JDABzmM4pgjadBosL3YGCEQtA9gOMn32JdHRSvzshlyLc1TvqNmvza3Tr
8Dhc92vNDfTC+O9R4Xsf4S6dJL0duRYUnbe6ahSYHfuI5qffehYRgfigCEjz9Mc8ZY78JvlJzRR8
wjKen/4LssN6C81JeTsF/N60KwMYATdKl/Vdudbw3U3fUFVNel3NC1hMDwSeGAS5s/g0nRjMogMu
s4Edip6Sr5RWosZBmmnatyzQY4DUCbUVB0EL7ZHLF1nyFKb2eecdRCqu5az/dsY4JTP/8ftVtUnr
xrNx3s6vwWywKjbtU94dhYR2aFIfZqYcYXl2cnXb6Yislx6N77sPjPhVyQFHUslVrC+eaWAzt4Pa
XL5RQM0qAfOt9Ku2NrJULUmNu65xK+CCzPq7LkLJ/9D830j2ElwMApYFrzG8gW9+x84OZxdDAUVn
hVKnpFZ18gl6O9M9ZWZO8p3Cwg2mOguubBpeJao4c4zCgHKxtXkeHUyd0U1q0TLDMyqYA6EHoR++
XXEAP2MdndblypAl3c2yORiGJbpMz4eiUFZH6vWIv0cisGea/rIeRCFbDnAl6RyvtG4kW56/WlXy
NMMISJ5qX5lMAumnBOwgrbp8aA645O2ko3lqhosvmFOlDaMQUb0Tc4KYs8EA62rN+r04hQ21XSZA
DXLJQ7mboC7qopA82CR4lQHPzwRL8g6181hfORVqnhTzQAHOd8HH1AIsS9m6jNdRR9xjmDKwt2rH
LDD/UEGwntqRYUh0mk//eZ2JeGmQAxkqD1HEoNv+/6hF5rDns90+N5YRyyhA5zrv8w0wVK0+8SHg
DDeVn1U1EQorCPInqfwdE6wz5wir0cRblkb10v666gsvifRcvBmoWST0ioa9HoNOv8o2y735zI25
BJIW97HxQTMLZkHL1tAJSp6js63uCH3HpE6gXoQOpXO1das1J8w+TOkBBQEGbn7XMy9wTYqqbZYf
0EEDSKzpLP8WBZfsNcnHDXtSjktqJ7Gz9GRgtoTALV5fRg5AFdxwXpnWEn+jCWYvsdIgHwrdY17z
oxZ9mcrqyOrNaNmN4y59uR+KPkPuKi+TO8WO5u+Mk8r4gARl3V3VttQ4aP3ek5ER6fsNbmOKK/Sa
qNuqi4BWJ/O8616vnHUAHueTX/gm/jeDWZXYN1dmnjjHi5SEka82XAJGXPTM5xnVyYaDBo3cMOPM
v6VRNRPf/opy8Yxd9VAoHqL1ohzC/cY0u3cLlu6lNxDBCnsKgI81M/vbUguo77btjZMNU6GXdwQ5
BQc1lkl0IkcHnQmDbRgPrd+u4g1PfbMf8X0TMd7tOZYMh8Wl96jqtsZQDLkPGXUc+6Tfb4obhOfL
AAaFWFJD2j9c+6A+MakmIbxorqrfTRS4lPVaZSbx7e6hiFE2hF9C2IcXDyLBv3/ogRvG1u1lS9yN
z1FPrB/36LBOuCnarhWlQ9V5doYahLF9/NA2AdQbtEQBNaujLEcvn6gQS6I7EgXnbhJdYmmmHwKX
DGZvXzcExpfiZ+Dof26NjpK7NT3TUXwAH19k/cqnOkRwKYIG8r7U6a8yp+2Ry++XcGnLbynKz07B
uAoVrKGlpM+tbf4NoZHOSeJQVAm7vQmhrgPJ7BpmmEvqeG/yNc2wCBazOwCECL+6mukCHXrQpYIY
p60AtKHXkw5D7d2mJRn8xN+SHn9jehY3A/QXQLV+v2TSYTrF4EjbA/uVRhFuTMR+5F7wnLe0WaU4
B1zS21SWqUwEoVGXVWMAgrBkbEcnpS7VLqeCNDi5veSt138KZPVecPWQn9MnF9geJ+2XUEWJyBIn
VVaEngtV2H+/YYBn25kPHyQwEnhxzehwOcqpR0HcyjCSL8N0JjaOUn68B3XLaNQifExcIXtaLuDU
chBJUcFjFB3kVBEXHainp/MDpT7QLLuU80qFxyxE2IVjoPsCuRdQCgjzd1MmduEPFHUjQzMHx5Nj
KQjfB4VAGtadSdtAmFJpHdjRcz+DRBWyme4ZHatkEgYNX70DggoeETdGPiq9WgcWRD314oN/x6M8
rh0h/MCAK6jUJxxFulpbGLGAmuXSA39fr+mDHoYYoZRUlbmbSoh56pfstQNr7wEH+4/txEyicKWZ
iAb+PY9plIN5DLtGEaXe4/L9WaAM5/KoMlnn6b55JltXks53W5hkg4hGQ4mxTfiVX+UgQ1aln6+5
tY05f1flHJSw2JmMasAI6Ry9qV5twXzI0nx2OnuzZslydXvfekj5xY5WbYXH8cLvge2b1Us6QIXh
SRvWgmJiNyXoOdWXoeCUKJFl00BYZ6Ii2bFDbE0vEvhkdVl34nxjTjkq0A/zLmV39LO7S2vpqYpi
lOpPRDhTpSnN2vlgH6o9Uko6WUojVrJjYfpHhXOATy4yY+aypQJPhJ8mYPyHk7babgk28N/RC0yc
WSul6+0kyWbnWVNqG6f5EKM+Ephy9OZdTeMFgJPHpxfDc+rvlnBEWHOzV7bhqrp0jCPiJ9TQtCTH
UGly2e0zM8dhap0eeOA32pXv9Gd469cUfZh/dwdLeiJRxKK0AMgKC7qY56DPZ8DwMhom4TLFie68
JmtOZ03W98FEbg4yBYUY/V9pnNOE570unRIsuOesJZESmMs8oyMxG+4IJUmO0JDW+EqmOTj3xQFG
X2LHcekv22jVH7GNKKypv11wirTKPWfM5FTkBhfGpMx9jMJSazaPP16yum0TK3MBTE/aOeHn+TMt
JFR1XDhs2LnBzD9LhqpCgFvHmdJHV1rM8GN54XqrSB/JfN0H+lJCGOCNe9j4QjCjhD5FU0SVT5AN
bq8aSA2s20WyAznNTezJWxBxrSm3eqwgCyoZLk57bq27Cw/zxt5ia2bE5S0n9Qbc+f5QyIb/pksv
e1USwZX6VIcI72Ll86dMcdY6sq/SAZq1BKD3EhEVk9TUjgAL3LABXTdTg9d+ILcqWsQirYNSYox9
WPcWXKRoiQSHywI9OwWite/CuKI2SAR1h2sN94ytc3fCVgDmlErc5HHK3ccOw1qOrtiNqvB++ACs
1ifF8pqIWOwbs0aagskjSCNUdSQBT9k4JWGK2zCKW8ErWlJ71HRILISA9LbBwwxMVJJhDBGoz+KT
D1+g4i378hgvDLlK/NyGyOwsQ31YFAbZPIWmiHXOCAXqeu2bfhZXjMPKjDHCuhP0NOCiyoLJ6+aW
JPjUYb4fDYfWQItZ//MjupAmfwqNcIezqMQUQr0oVcooVxggxORxQeb5ILiCjhSqgsNMrY4jJ05C
ZPaoEfSN1DepCtCBFjaekkDnGJ09xRajVSgEU5lZIzCTyD+zD5VtkLpT+2g8F2+0pXg2LSN3FzWT
YUE1cgWmjT5VL3AEx15yQ3AF/a3G+fvm2vQTngAa4RVGzrRTeDZjRCegu+nwEvM5K1Cle4I6JQUx
l4yMBVYUD90N9swnV/tlDpemKodzj4230mbiPbvx4RURTQFsyXUgTze+f/HFVg+Fv/zxdsMml4p2
C5Eo677cJhT9zq13DiUTbWpz2mtWTPOSoNu3a0yqW/WW8BX/OPbBd5avyzg6IbS8wJiAAubwS488
aMbthSR+jZqwcxMUFfxOMoCmBWGRMmf21ZQNYrPAg5ZJAynY8VLOKznRNAP82URf3oyZ55Wp4sUT
zTVKpP+VZhbe6L6RpRTEfhfMGQDBbPI9eLIgUrHomgLxwj6KKBAAk1TQbNPhIZ4FByEyLtOgL2Uy
gxspf2KAqFdOjK7lDr1LOzxC/sFx2w/WfXLN0sLxVEl0mhU9P2XkcNz3OV2eg/Z6XiEHSvEZXpuT
8IkNlWCTxlByLs81FYoGEqTj0k0Zv5Pob+Yk8/QQKyfvNBXMoZwX8F3sKL9fv5ibLUAzD5oPPFN/
oHbSHGN60zJdU8L8chWrMua/XTpMdvS17i3YLxM6yDFTtBr0awKJjzmoYHgw2DYgdkjSvVUKhHa5
GdWUZcCbFnwbV8RH4OhR2KdbEWyPhzIdaP/wwCEVAqFigcS4CxM598GEqqlwXgRRqlRxuD5YOnVe
mpcioynnGdxlW7lQ72qftBag3EjAlXTHq2Z85m4p/3a6cvCg8M8yF1tbTtecgpFenRJWs6RQet2w
tz77WEtL4tnzvBRi0XuvBqNWHbc+nc782hl9jJv85b+Wu9d9ySnVE81PCyUDZw+RTxNjK+2DhDkK
AaKFH0ge7RENX+v/BlNxSEYxGzFSVYrO8KOaQGpVi0xTZWpB+axLXe4h3j55omwq0rZAYgUml2tA
n26GaJIZYnoH3LfT2n/NqE0LIh0DwwhpiaqIKNYvWInUfqAainE1ZCWFKd6itHiCOpGM8943zVL4
4O71M+Q/1oUqA4L00skfwlywxeiobENBNGvTclQAQhtqNEstgK0mJsbTf0U7RTGK6R4eOyHjCqZ6
5Hp0VGmRbhf3YWY8MwvjYhzmWP3vX9QBN3HehmTK7AlzYvwhhovngHhnOdi8beIil2G7SN/6Holl
92x2ZKTstQjE7ORQERequ5eyh5yLMofZv1YJNQeTnKe3anMmuI4+WcksAbkn+Y2InP3BegXLYEMh
hF4dC7ARSK776Vfun4cs7rQpuAGhFUhCzWTWszMVHscWKECVBVjUwTHjezL8bphbpAEuBkxWCVwe
xKlYiXCFdwYz5CW7jUpVtRh9qY30ZB4P9XhyKPSgjedCcmzKz6vKOuWhS6BITKuwbJX7HdOT9SW5
bvw2kYDbQsAnwaMkQL9HvpcrdOcXP0rlDf+YiZ2KS2KKu4gLBVKapJo3Rtv48LwoDQ2pDzPtLILp
LFrp+Yfsqr1t4Io8H/oiIHV/aZtlyoiThNntzL82GUOtN8PLfhg6nnMJAh99tceRNp3OxUbVJ293
U13bAdJm6KSGqR8ylif9IYbP6qejGrLN1GYtCDrCvuRiQgKCvcO2OBGqrCmctMn/bD5OcTkXgaul
haqMdCy+T501p4i3Yo0NrCQLAPThylQ+CEpP305dvvvNfSeOoFsC78yy5ihKjRnep03ah8ZL68k8
3cpzF3zpAZZK/W8nHxNSZZK871IE+930HxrFFnSzjyQlxndz3p4DKaOhJ29AYqpyugPPyWhgr9Cm
CxP2IwSiMsOFr8WqSAYL76iyKCv8V8ABL95QQVFlsEIKCk2ew6fADXH/q/z9NTZWs1AaE2O7haYM
pOcCgtqeoTlw03ZP5FGAsJRSFlTn6MHUVCRqiErlYVVgHzFr2MnRpFQXu99kpt2veXdgZGyQ/oLP
d3D40drtlSirh/EOwEXlWeDwgdBYafbyreMg9GFG9UVGHBFKLm8GDFLuGUKYK6hyrddW4OS8jOpO
ylazBzumTROEqzzxXAIkDkLZ8YXRpqqaHWVmJM9r5si6EDnU4OOMbVMN7LOjuVjdDb625yVDSJ/A
8yYsMuzT2UKOszZbYRHyh1RfEnDsiafLdyWMY6ksx7IEL1Gzpj7xAn7vDIjnO7suOFFiiWCYPaii
1LtjQZA5H9+Xyv064wEREYOiPSGKxP30PRlzbB+3q9DwlpADCyfxtqM3neB/Kxt4V9aQMLaD0qWn
2PQ1nE3qf5BKcXhpMUFe547h5xOKtgh7hW2PupvugIYWdNw6J6AMZWxilUMfjF+/F3AYcMsex+bb
rFP15aFKqmURad4g5Eyz2G2QCg1qFJAF3c6j70WEZQ6nNiVzkAY+Gziom/9qKgBjyy7BycpbAx6+
BD7zQiY3WWxVhfFWRPZRUhmxP9xD+rhSF+VLaHy4d9ZUFes+R1kBA6vS9o13tPHIgYBzmUyArKmX
c9vil7MO3yhjyBX9Li3d1Iz+OjYmaQ2Yh51cCQPntbNwph6jSqrSB4bwY9WkyM8Q7uJa+OE6cxu5
cUaytYT44/mhNG6+0ph9Xuo760BeDyG0jXsdWSlJGYjcU+zOYxT/PhdcnG5Gi2R+V596lR3lMGCt
Mo/eJGUZnv7eqrqvq/EF+IyDyZUQYhKoAzYz1XrbMydG9dpSOEMSxp7f+PAsiRfcQ9YzVz/Yblmy
zdYS7hI/wd6WnW5XbB73tTX8cUGNNsyMstZC5OELDlheA68nXz78MoZL89FluwWgQFcaI6oLDmyt
R9BB+WuApyJBh4NqUzB7tBHj0MECf/HSoGXo5Mu2PojAxrKtuMXhwMD9m4zJyQeHK2F25dORk18o
O/zpju1Aocn2ZJEfCRZd4U2U4HPpOfzgZ1/eWZHEnSDfkFe2/+RWGNSHnEJVMRZfaYsdgxiG3hmF
GDR5S/3XVT8oI2Ib+qsocl2HBbDdKKeih5Akft3uQHUVOvqlS7X21WBznYaGiAG4CUzTJfqt/xi6
CsGolRGRhH1t9Cx0aQJiKszL9zL4ex8iu/nxMsHROtnOnNqHVnM3ApOmYWv66VNfoT0Bg6gJkszq
AaHWjDz++3SHc+Vl+ntNtANgb6nEyt40SHzjSjKe70lANHgzG/1NLAs1nJ4Re8e4vgy5RpAh98hr
FML0ANe25VQpa+nAuBK9CSwZuzOclJu9cTPmvqdotpbydw+qXwzKNKlsUeIb2wlloProGuBOjK1b
A0FbaxhZW1in/BNUBPT3OLgZhulNtumRoNPBDLlOcomW1gVMthkHFaC8o7iAemGPaOW3N1+V50YN
x0mMsoEW4/y9pQVwexMxf8HXHiZ52yD/bW41psWzgYGTW/gjOieGClecCzRtXXIa1kTCHvqbfheE
0Qg6rECD8NxuMNAzNSCCBUyiKh5QJKpHGl94V8IptPVcMmr/y/6PDGLgUfD6Mx3oNvKcYZoyUdn1
Zs93k05bnmfm95qIOL8WeMuHWCoJfND4Z6yQ7mcgyPAfl5/NDwBA1/3IZdBs+gPbgaC88XiBMPZa
BSKLHpzZt1eijL7faAkCtFEBpv2EB+TEHukLilB5+3JBer40GQcFO8vy7tYdSs5ivbpBPCZnaAgg
oU+ptH9yG3BQMczrMdnmLlOtU/0PpKXS4A9p4ulqMoBi1PO8WB/0QRY7zcJLKnJopQNHE1/v5xPm
CC9kiFlf8O+FfmSVqj5qxef7pgPGuK/Lc9hBaa4KnqF3YCmegOrhK0YkT+MZq5UuRim8hQgm5gE3
GsAwjCqGdWo3UuDd5K5CnqCc6au4kyffEXmPtrY3U1z4j6HV2KYQgZC0iGfHsslEx0VzGZjBgjFb
iD+ROm70d9/LHqWz/YMMn1MTj4XL+Vt0vg2yQy/lBBHxqAKyKO5uOyOXybq9GK38xFVIq1HcpHPN
GYQ28gxyr88mNgkvhcikuPcKdFqEmkwYytfHd4iMHwmevSvPXh7WoPpIuKYQOVLbUDC5fVfPw6d6
4Hqojd9R+n61S9YSfPihLHu6P42dTxErBctUl5Fqmb6WDq/ndMRJOqfhvXvBmT6CVNDt/WZTaD3E
IBpZ1Rd713+9pt7COS/VtU7kfdXQcaVEOa3rxgoHu66v569TJC6/fbDdJhWC7PAZVP0XlHK62BAA
H0imbplJ4g3ezawfjeZpub471sMfGbEwoVb3DzS0bPH3plvOdSTOPnmc47CFlQa1n7gl1Z+SAxG9
HOVmXY3YlmYiXBwrgLQ5px44yBK0vIWcVgJMeMosKeAhTdVTyRwvrFmhS4TmQioCFBT5J1HZiHow
jui+ebEjoD+Wi465gYD5NnuEAPJxgZPZwctCjGMwQ/Q7dfYr3Q5gK+HCYqI4YoHolcJKMS9A4obB
H7cwwfQ0J/O3VcFISU+TAlap9Aasv8yEI8bHvNuHfXf/tMgbGCRiRaDK/SxBDStxWZeqDBzePdpM
quQHccxBEXehWM9VZcV1P8S6vLMw0BxsLE6VerV1QOcUVZYyC/7eJEOE8FIwQjOcRgp5zVzn3VQ5
3DQwLb4NLvGwLehzGR63luo5btpngtXZ1uEv3SKNyXnuebOQyQe6FrlBnJUSEI17PVHJJ+9J7tjI
yGWgsnhsM4XfUaQniaKsbOO/uxrhm71/wh/y9DfuekP/eSGen13VLw567+tz03+Ada6pGW6H4k7U
eCAmH/pRra+ivx2vb0+7LLJmqOzbyRCbxj9BM0NmvmuvfXIzfLUYE0295Hcbu7X6YBvYw1HOLYDe
+PnzQUfAwfpr2IVL6k5IoGmSrWMpod4vr1HlN7OjKubdTNAcM4ksVpOXW6OmdbmnGjNqq0GZADj0
U7xi3wqrXDqNCD0/1w7AXFJuOjxC0BGAmAIjxYlzU5SfkYa+AhDdmmYMZQyyJjN7fLMTDorS6PWp
iu8cRUJeKIrXCSdgTKJPJLI86LnxPHXtkSCxukU5a0EU0V31Sbw90dsqRDTW1sW/urpbO+D5Nmp2
plLt5cyP7OknkFvKT+sIcmkrS71k0pVL6KM8Hhk3r/A0UQFG+1p8t7WmRgSUgY4xNgpYpdcB3gU3
yz2veu3JDFLGRFxkUgypDdC6QvUGXwTbjifikXLTL+9ga+7hSibzwow1LyZg9OCMhcZM8vSIMrYr
aGIDvgvx7xlAEOTwdG8Eqd/NVv3qYYFiPvvEZEcEP778lTfLxJ7DD2yTH82WVGy8YSx/G72e92wN
RtFcU1S3VlTUXYMwxvphgFc9RAuX3+jLaN98xaciAEDcD7daV5apHamQRkmDcuJVhgtUA9OS+B3o
o9joRm2/GtSqZUyuLkM3D0SD/ivKsH3g2d7/O234ivQxvZdv5ptk8d/ySI9XBwpCTXJsAwEW9lHR
GyeGm4EhdYbl9qPryRWYJa9Exvb84Vfosi8C1AW+eAtqSLhsCDlgJQgMBZlm42bRcXTFdNta+lZK
H7UWUytgJV2SQ49SLnR5EbY1tyZqBznxAa8RIpJoZ3BBcxa6wB51RqjWwvfk5juw4oUXiCzYwRNM
ZgGZB9yFip/VXy9wh+qYq0h+33iwEUq2gOAp8k4MmT8xHSeGMbwiXbzzFPNtUF5+u06vE56bTgmW
6Qcsm1FFs1zth4AgddUX69DYyPwF9qBpxYkdpg/9Y5svm9DFQMLrWdHsaW5xyxsOEMamByMcg5I+
2BCzqOfxnMzX4LPUBohh66sJDCPWMkpyo2ZjciX1QUQuA3BhMNwYLm+cs2ygZodo8DvRmJKUC3rJ
2btDnWgWapTN3XX5OckiCKIG+OBNYihikyoVoUGwzGPozTdjUntQMpfToNUyjTvzQSgAleEsxIMh
OjA8qqW6LeWL5Dc/1YLQISHYS+UFnpjgdr0kv4UaaJMeR1zgvG7nJsaId2VNeDIB8yytjk2kccok
0yIeewxCylStnTG+bVC/D5L9xIvgIrPWm+0hDbsPuFlhuph9xkpXouXbOxBsRD3csGU9ZPvEwtdw
fWXcONmqZMI+ZZgFLdF2PiDYqxfdyI94+m/2Dao9665gt0pCNjdRjvEnSblyvKKX6b5f/X+Lw14g
GbVOzGoosZLLjnWRS2wqLwxaZmB7h2BCJm6aKB5mZzQLgckAvUGM6aXNHUD0zb13aIEPEfIWZuDY
+0pamSLBJZRRf+ORnNESG4Y4HETjv5LEdZNg3rWfQrqGPv03diKQlxfn77d5kO7+vt3uvIx1YRMN
ZkcBwjlv6w2/KGv3bQixFSxriTYD625GAdtmuOry6rVrETwwX9fXdsDd/OAX3HaagOEvzZ7sAG8A
sOo4NGJDTeoKoqggpRWefpdJRC46Ga9JadQvOYf6avjb+uuWdD5g+LBE2/ekkPSU+pb2xAjdtVzI
q2J3BRe9DfMSNbiqFVoR1uCgEOF1y8IOsaHUpHgzjDLHJn3buv/cVuGuLpJ6RVGvgxsBkaAb6Zkh
Oq4QQM2EpfAP7KZvOdFu1QdFRuZwa67a54iMU5fq3CREh3uEjmwR6Ln7noy3BIksKvYrfPUB5aoU
bMAAuK461oltiIAHj8qs4NkUKvGv3SEVRPX4/LXMmkKIz4b8wLiW6v1XXV78faPSRUUB949yvDR4
4L3mGIgVMHi8Ng6jQfURgfob1GJDtr104z8Deg0QvhmtI2a0kSuXFehzkri3wIqpK/21q7/sSNIU
xl/t0lWWfMq9yMxOfaPX1fxrYj48w9kM5sVGNJLxaH5RnOr9wUdXGV1l4GmxXklH0Wml3p7aRf+W
dEVWx/juozQjN1Py0iR2MxnAL14wb1nwr9f1EWmk9HKdle3Aj4qIXpdXhVUXprJSjS2KJT5RnFYm
EYDp6mABYIBHKG+Bdam/m/WogdlDTJFm09QrUsaq0DO8IuYLCL27Jl1aAB3t1nF/T4DyroORkg5S
SBzk+g19THgMAggcduPmFhXD4oE3RKlBCXZinfPyOIbW96e1Pgl6vJ7g3rLBIidMsN6l+E2u8hwg
EHaNxl1C59FLS66N641bZOGLGTGmUUr0rjYx9/jN/128Foo4lKnwuUk0oWUTJZe1/m2JfP7fIq9d
NIqbIKmc9sjs+uRyIOVqi/k6jsEmR+/ajMxVpuNvR1UXlw0Q1Bng2xjPa1RKp15SfDhdm2Ex60En
GWa9gwa5gvHriGEXelcXkC+6cowxRvGRnPofso5TOFUZwo07L1y4Ke0QDuJqQh+tyTPfEDvqS7Di
3K+SvP444v5Lv4zrJEnALyyLIk2J4nluTmvWQ1j5ES2YHtPUbfd8Wu3/el1GElJ3YUz9t51sfSBu
nyxaceHxnJt0adtHziTBlk0B4B67ZXqgyaN/LDKZFN6YrwdUO3Av+xDMfCdHa6AdaewJXoG6IaQ5
ijZI2MbdsBAMq1m/bUbq6ropwB25i26uPGMML8BSyG0nP52tuH1wXnbSZUgWL9moBHid4ksk05Sx
R6CROx6Mz7xVoAiQF0V1AQbyUqt0zRDL9vOLIiFdpSzjEDAkzSGayDeWXVL2Z3v6dp3uyfIZxQhJ
lrOzY50TmNEVXtHlcAp+OiSD79UhVtZ8FCDqLZM1ZXfxH4vsRfxJ+EPxqBh00nLWSoUj7CuBQtVp
VnuwTfVCsQ6U9W1B9eTs3xDqxB9T2f5sUuS5+dgpz25kgtNQQgBX97NNQlYQpQTxQ45+2eW1ZRWG
FqIhM53rdiUQYwDNGpR1ahiyp6RYIiGnBWf0vb+1MjMKd02eLiXi+mK3O0tVjUc3L0rLWxph7WPM
1EXzkELaHAp7ptXCK08Ncoc49QLRXPsrQ19MtC96ta8pIBaa0k4t9kUZN4AxhYaex/75GxTaiAKF
mCv6gyEtTIr/07zJc7hX7xf1VN943cM9Wn/iCz86shG7NNxIg4YyDHPAXibcbUiqeg5V07DBIA8Q
5ODeJTVPFTFuaF1kFexSweXy4D+bC5VF4kTi7luorq3DLGFvT+x6Bu37E9yZjGmjPK81k5Lg+WDI
O22YRXk+dWgIIpyX1pszDIIwtMnFEyZSXsK6GL82A9I/2mCVibD8dC4SyoWEkCtvzvwOnO9cWuAv
nQk/6P30J9hyPS88O7wimvRfXniVBw04bAWGTYnriHBErZ+urcTtPXoC8pDVa38h2V0Vr58nymt5
4XTeI0Ui7ja4v3Ajh5wMeIE0Y76+gu8iKFCAcsYqs/xRPMHibkya78iLEi/aUi8F646NlsQV47ft
cLC/b18WG8bk+qa8j612Koe9pybVaRoTiWzXQpfC0c2jv7QwNehp+TbdUkni8wfnP+fsu59OsYuy
EP2SC3/9PIjo3Z5rB36iFSpX58W3XX9vNStpLUc8IcfI1cagRwjgFEj9YWYY2X6UFa+YxcUA0aKd
dsLFty2BsqH62Zi6PtW9D7mA+yIB2ozWwDKv0Q60tLRzPd7T0AWUO37cM5hA1weNxx/V/fG+BGAd
UCFpzRAIjDCqZZAetQCPanjOm9IC08KGqgdoILSftWKpdgM/Hg8FHZrbAN+ZbyGdEg8c11bzewfZ
uHNwpjcq4QGk8KpMdJ6S8pOldYP+GBeHX0WCTCdKoQSt/7IoTjNpAX+qNlEeMjkesdCP8vToAnKk
C5GVrW95pGioJxdQsddqka45/S7gmwJoeo6xxVTskb1MKvzOSPhMinL2AaZb1WA67XoRlA7Vlh9C
/iP1lk59JHWutRTq9+evb/hrSJEwptVkBcuO1sShLd5+eY5IzuONquq5ZIMJ8I2bRI7PF0lf5IL5
RwkAvWOFWiX3DZjUpzVMsNHqR/HX/z+9XZyTQKlP1ULZkNkJLhqtr6R4054pNZFOB4Hp9S4qPura
G9Xr0hrDU0fFFzXX8DkVfui0TEfJU5fqtVyIHjY4BJ7Dm+QjDoCAhILXnLYh9D6zgaOliLgcIUdE
Dm7AFKyoJxaaaod/BkjZeUmASEHW9sJFTgl/6tT2RaYrsJbqdEYFEMizW8Ruk9FacXVaaEUPBoRd
PjITVHVhNxOaAfTqjNHqepVUgRRryAsaM8Ao/85VTL93BoiRZtVJV4kycpvbFnRK5f8GxzvSFJvl
3UPvwtcY2b8wRVphMXdup+Q9Zrp+89nCM0iB3GrrjfCGku0UWPT85rKyhomVPPLnGqBg2hoVVFXP
RL5rPah/3h5lnTFHp6BQqBIXFtzWYj0VP9nU73CiXW6oThsOui+pdMKh3hXHdnjWcXxRQs1o1Ghy
TzaIkLWTcmBYfQf14kDr9TmWbRBO+wZVcfNc/dFdidIz2KCUTIoqDkbfYD6oGAinkcrzpsCoRHVH
56ENV5vwsgRKcWgEQTU0kQLX/081jaOcoZQkYni3J5ztGyiOkk+O4hiTdbEF2LPskSPjBLeJiRHC
6FBCUOQ3myXfTZ2mmKQNNwEm83Bv7Ltrpn5QDKXFpISekYem6QrWna5zSwSpGmrKEM7mLgzb5Yvn
Ji0fWkidPhGxNQQE1QOYGB9in3Hml+UmL2FY+C+pvR9GSwVT5nu8JawB9oFDSproSHRpuxohtjKu
UqMzyoSqtbxDFH9K9fCYEe6hHQ8gLbNscImLXnwx1u8e0p03PRtYwxyyEM9fRe/xZz5xLn7aa690
NkzzTyz7oqlfX1PNq4NfrXQoK1HVnkjCCjbAq3r6AT1joelBMfJ4hzzAuvsCVQd8TDRBs/Tr1rAF
qLtIh3zNAHaVAsoON7CPl1oQb9XPd7hGw2uhbFHTQRvIBUCHT+KeK8zErAP3oO5vJfIAcKeXPcO6
VyQwYwS4WboANoKd3eCH8R/1/KULvTW/1nodG9NR6Y0yBenlNPdLWPbMzWe1oJpnK7it7o4R8Hwg
OWBVqGAsvBO1SOsIkAIz9tF4wk3/ZRw8ayoko0AnnSC7rVO0VFf6bG5jmmJERNjx+z5z4nbakMtX
BT55KWHldBZvQ9L6wp4PRc5EzIHzpAbfik/eBgnxzCzWWgU5DLP4UTrDTL9O3jEdB3MOQjsjOdWL
yPRipviV8prrOq2TtwId++3LvJWThm82MGM8S6neU7qKtr+4WfPx1p+FL7GgSmQlJQ5SYJDgLVZD
VuhXX0d82LwbsQx+0h5qChoBKkJNRNY5spxo2it/EaVjd6mi+lKn3IRJnyn6wnTJlkELtPfoi63g
2b06jMjopdArsbIkk9eTEi1gf74oPBEUSKv2d1AloeIKBNDNAAqRrOXGza8k/7Y9RaE4ZXLoIB9Q
e0VD8cGLPEjRsJs62n6BlJb/GSCDE4xBGbdKJNO1pm5w5kDVAqcIRXcYaUova1Zr8Xmg7Tga5poX
c5kwzAM3hTVrWjWfPr942L0gRhKYEw/U6NSzNDimWKLeDkCYuzaRHF/EvjB5l02CCWCluHVxQxBl
kV9TmGjAm8bTxIBDCFBlNLlKZMSAY5IuR+5LwDY/vWIgCxHbpSjXMFpqob9DJTWXiHrJpbByt7Xd
xUrc4M2YHZoEhkEHAWFNjwnUCZxnU7v3h5jV2JqLk+Viw2TV/2dZ0ljSdhHygiz3F2DhpQiNCPaa
kIG5/abdhYzNUzMsJM65PJKkSG1K05X6dKU/KDVuXg1EFHIAiojWql7V2PkenmddlrgNHk0oN3aJ
AlDAZVyzoHY8pmPcGYLJUuOMfQm58WMyBDEPT5EBEIOsmaMphDJ2Ca9QZAdg+tMdnLmyqMcaYNzD
TvgnLrU1ZFHSkddfXPtm1GrDBH5NYfjynbM+yEw3VNZWpK+ambcdLfupNzNbxkiv0TZlCwuoxeOM
9VdXAEid1GT7kGps8nmmzx8hJgSLBsIgyqWlH7zDaQOlBrdLm9LPuNdsvQ/8QHjfX9pD2UZOZLLO
VZ98p1lE+LZaAF/+CYRCyVJwilo+SVDAXKU5WgKV8osPqs7CyIcIwR1jCIukT3mesnY9DgRjrNFs
SDaoiXrzy2U3nmOqUJHut3xyPBasoVKyXaj4T/b41KNPR3yc9N3ujG+zZrJFFj1OFdrD2dusxdfK
W+Q+mCY6Pa2c3DhRVxSDiVGDwJm0yvlWIzM3Os8wVpeOX8s8OZzVOTrmN+WGHfNU0VNUpAbKR9Ab
poKsh3l362yKbcu2N3qOWMPFpR41j/kpN/H9a3M8DsEUucnBhB2SuMc08S0V7QemXXm/OjeX4QYo
DpwxvlJ/tO70yKX9P9AXC5j+WnEBMGTwJRT7dZdPU0DDd1aqcKHXee0f6nn6H3JN8CIOgX2jDpCP
gPnSxY04UPs8oUaPOgeMd8h3KJg8EfashDwDO4XOL7LKZhhZLsgwCJPrEv9iLqszxWVG9gzMfYmS
eqvnPFNJqgc4eMMaZJ89m/AksGHi+yj7tUQqIbCGJ0dZay4s2kf+lXE2ZPsBkvtz2ztfLuWWvcHj
sZRcH/srKOa6AtcDwM2WoUQsjBujsvZMtp58BrrdX0ExvplwqMidKUjixUP2kO4ld4U1+1gVH9+R
QcqDOR9IsYDgEkdY3xIYFnFQbvfoi4YKq34xosJ5FNQEbZFpbxcFMNCzu8VoP26jPR77ukFRR8WT
kCawcOL4O3p/JlocSNhCjqisTsUyd/tewFCIhx0UnneSRuKQY6cnejMEaVDqRy3AmaAlQvUEAQJV
gmWBKRStDL7mtURtDNyLpauGgimVj7x5x0nJzVLI2RJS1XTwVsVgbAa5RXdVgis9N/dmvD593nEp
3neLyPoZyhplcYvHFzZuzOXpcsLE2Xr7Dt6gCQZMcc83IAWmNl57xzVPJjtgrJjwIgaC4vAhxkso
AM/FEw5Ntf5DOZYvoV0VQ6OgleMsUrF3FQi5dtJPghnM9aUpzVQ63VNivRko0AWexYcpMkSzw4cT
Ejw5y4pq09aPD/Zapy2a72P1kgeABnV4WwTOR5PnMLNUzySOZTB0tJyWvOXghfU/3utwGk8pMdwL
c0DVaSdZAUm1zNDrjL2hR4LF197XRccjOxM/T0/dbNgoHKmqN+np0GHQ4e6DYkh5EMvjqFTWB6FX
TGFj6J/dBXVLmA+Fk2E41Sg5Tl5qJKfTYlz1nq0tBp0X5ThrQCi/BLdT77rGfowsSWiGHCIr5RMM
r9qCOZdTg0CPC9B+P6YW2Z7ULA3/knMJioGiqBBNRsKdj1nmvzef/cltgtYjWV4iIW06/+jAufaq
ElTbLLyU6fX0/f+1nIBDvGhx0+VyXqA=
`protect end_protected
