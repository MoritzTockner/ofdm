-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VC4ox7RYaasQKXRMgxGibg20fO3mmx+tvUhMcaDXwt+zCllfJmbEJab6wLbvOVDYZjP2RQfBE6vG
XjCLM2CpZ8OueuJvUvef0ZRpcSkzeoKKP66GIOSFb11S8vSDqEEj6eE3jVxDcWXIbWWxDToIXKg6
i7DSZHSsRkZWFORig0rJIo5e/wySUzU/MmB8efRJpgQ49Ul8WIODAK/MVYDk2nFuJ4AaYxNENOrm
bZs4xfPWYcLCcvA1w/0Vs+kqaqN8zWzqzzaqdiQChTm08OH/E2OXGUun532Dna1N9M7VO5rGOfdz
kVV3c8ASrv4vcnQKCMGH5x4IB1psCwwHRSSuPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
hXXsbGaiAV9jpLaXORTUcJDyBFBhs8pjR1IVcowND/VcWtWWdg3FncnE7xUFU1JTmWzXUpqxcGLk
OZc6/WD8ij7jTsTur4iJrJJoTj7BBAEq7Tkh/TBY4Y3vKdZnHq6qJ4bmSjkiBF/i7peHXONADOEu
x/IObc63ol5sMH2QZ+QWYfsaw0gq4GPDXzrysILR1OAOlZsD9+0uo456BhQBVpI5Ilik6pEqTtew
41BDbkuE3GTaisK3Y7MEMoFHhH7ckHInt97m83U8sA8HOVsP0z96dxzAeJGXY5nHZz+0TRbdGXaL
7Fna1jB/70KIclVwkMyjs3qeQvIUzHhTVilFKo+g9PPns2clVl3S4/perY6+N8n1w9LHGuPPqtA0
vjLKhXNkQ/gJ5q8v2KBNIvPsCCPbRWh3TqUN0jwS6CrrkGvJ+G6R0MAz+N4n5pmJQtZrGAW2QPza
okI6KGZ7Sa+QgiIUH0eB5Q8YBq/HoccAEjdp7eqTOdo1YaJjjKtBXerXxHmtiflzi0BvI3gcqAXx
9n+c693SZCI3/IrVeAp4Ek+5kynb/Aya0nDB9lolDBz3LFagSoOVIpHSreheFzpQMsiCe2kPAYOR
a0Mb3VY5Gmndqm/8vUCP4DzYesLbVPqjBcAu4MEtl5pxGdIcPxyoCxYvGoq7WcpnGFvrXCbAXSO2
dMVZJrM56Uf+JEJEkxipQhJ5C+UvoZvObKb6Q4V5LNyWoULMG9u3g+TfjHveqsSghx/G0rHMDlPe
gqn3fVkcmNh8+qu2lW+8UuB5E3ZG3gmHn3w1u7nH2r1sNxoX9jzahBwYlgHHfzeXlmNmoI7fNj+P
0BbzktcEoB+9Bhyab3QfxupZPybEZdb5rc6bN/zYzAQTZlhsqUK7SKpOshm0TfhY/S6Vg0RrLRhG
8Wht0PspGtT9TF/Bp4uzTFWkBl/R+EGUoT7ezi9K8+uyj/okZGQoHVVjCPOIjhaWu+GUGxb43iOl
XI9ukLgXoiUrko3qk3uYlGrp4uZrNGxLVV8s566ORA678TiuCj4tI0DU033at4XfTsV1Fhz4cIGv
yieK/X3VtnlT98ZRaqyKtwHv4lkYez2MUjkGtBdCDRRKDgluLb9dK3U2z/cjApFmAZWs09/8OR34
5kHza4v5FXZaxj7jVhMhJaSbfTWdh8LjOKUTHlwbFr5x1k9yd39K4GovyQiYRqIjXnvf5LaQm+rI
gDIEb9slxgoJ2AojXHwJfCZKYQeXfKFXUu3Lay0BN/nruEHfA6Px65X3Z2PMGVJaA5j0BJgMCzsU
BoDe7SgjY9TDcMFmCVneCF/bFvdlx3ix7mtU2jgxdE9af9xQY8efvX/ZKbIGIYpC6CsHGm/vhMth
X5qoQ13uU/7NHorDZ3huOSjZvwk887Sy+iBGLjnRiDZIAyQ53IYIlajsJeNDHuUQJ2A4aSYYl8ze
HOMtMHNl87d9pequV6fHKnZcAKA6C05jHG2kE5j5N3rrHgnTULqr9ssRnKSyKvkLv4VMYNwgV6mH
bhZbTgb4jLM8eDRhoOPnrnoA0NBqocM4B0LRGQ07E0WOkKHfpEZIeEYpZdSStiAh0cHrA/pwGPLV
ASh/SpJXflbDh6YvFgrR0IrgO5axEpN9yILzsgf5xAAInxeNmgccuKoTSbMk8Lq9lXdc0cHL2CmZ
7+skCx38PoTXYpKbIcBT0yolh0ElgJ/LdeGtIwEAfqz5SlJ0eow4whGxey/wUYS/QxPrGMzM0+iJ
6R/NpglwOXtzwMZB85NaaNhI2dQKiXnPyMWhQVi0HcS5tgWIhBZBNi95FHgsODTXyGuAp9RpDHUh
na4hgQ3wnobM5BFLDcnsaO068DISVyZ4gzDp3B+y4NzSrdNxt9aMEhNoa4llAGA7Ix4xL+ooewvk
MPMVwyYgym/h4F8+YipwdrHIIvnKazIm89nBIWMVz12sZ0kXgWU+ryvJK7Oi7WCOuhe1tyEll52k
Su77bzkoJvYiYI+PaRTxwCUPihM21j9HIOqJcpbJ7FXTqsfZ6qYz7y2v+HnBvLDcEB2yanTdTitP
YiA+h2BX2Q3fGn+Bqs1OB58Dmd1LdqesfRha90VUY2UbmwbV+FJtMI3w+zNWqyL5FPNcD3JMdj2C
JyATBNwWgwlYi+UeQCrcCWYFQo0x4SSbA9ZWqdbFvglqX2GeKnVVyzf94iZgOpjKdm7nlFsJ5ixU
+i+Kko82dq2kzgppFaOGIiTqBJpjUyezxxEw5B534gumTIBPIkIHzYWxT+C07Wxxkhd9YKjYhm/u
Ct4NjVple2ebWEy7LObhav2HI1avH4ygce9uQrN6vs1KnCbYZgglJHbpEM4WHXZJmXLDh/LiwNOQ
HX8W1cmeQ1nNrMT/5zq0SGrG5/Y5BQXouBAGtC1ZK1gQ0FjZBUPd1TtqtEKvtk49XRjvAnWXPAiX
K6uTpMrtx4zpownbDaEwNaLV7x9B107MNfkyxyrQKHLNVxCIYDwWlMlZPeJxPrMTrCECGtPM6ZdT
Svh+bLrRj+5cYVjKKSN+rMiwIQChSpCyPfbUpFbCcj2q7hwJAsZ1yR2v7P+DZ4BT46aESzkBQ/Uy
ieKhw8y9szFWV3jbdhkE5vUwO+/LiYvgTI6j4oXZidmqZeFrnXMDUFs6f5mXcnp5bS/D8Km7FKfQ
s66Z0SS3c877zbDQTf9rS6sXdqNwyTIceNU5v1ipbmjRQWt+UFBlsQfiEhNro9sWVFcs61X60ala
BqwoMfXaEQJ2bSFuKnklBxbAqg96Nmx2G/VnGNdjZiY+LX0aMsBfjxzkHbzfrM/I7PLZjHHEUsm4
46PlwKCekh1ePjX8rO8W8m4thQZeL+eWBdJ/SJc+UCzL2CFWQKF4mbqx3LjEGbiq8s/qfkRNqviX
nvPh4LNZGdzcc37HNfvKYkCfSqClBY5vbVozS3bznkeb02W8mBpFokH4Kt5dtuMggjQf0O2Oj4Bu
EeIQY0dzHCLJmUQAxTSQp44IsLPwq4r74BpXXGv9PbVtI/9gMTafp2u44ushAaM1sFJ8AEVJ7xwP
X2rXtTKusspozb2tcurkhgTOxpm//5Si6NP0ogjWOBNsP/AaZSjy7A8W8XIryyL4B8L/w2AwaT5v
0VUzukG998EAzo2yrTYACmkNbqC63eu3eZ96RjA0feB6eqs8cs3Tqwpi6wctvXi2VUa5GOI9GeOh
tMH8EB9T7upHeNtLgjJb4SQRrgwbtdc4D5e+J4YE7MxxzIxKs95VuAPw46HPoDS9ZBbaxgkOx17e
h2g/+QiealW/54AKtIuf1m2mL2xgRo89/LZ081ujDV+QfZuFUvb23scvIQiraaNBWjqoPL7BJP3z
HrM4vyuRHRLjWeLQ18MwrliQG9YKhbeKFCsHKQ6oDX4Sppt80lIaMoXFExaxmlG901l0oI6Oknts
cCQYc1bFAEJ4RWEQi2nBqxw/u2nmgGZsn87w8x/63Yh0j0pGQh4kwR4q9hlgR0lsw7EN4etJedWa
aWpfUojtQEVYR8GD+JJFfQxktoDZ69wS+ipHBMbcgQJ2Y9Ue6hBUYQzvjnqtGSNOYsLQGhOfnUnF
5y4alaVkx4GLIf6ex3dNbKXmxSoNrWGIrojn41lpK1GEg7N443e7SWrq1QZk5h3EqzyiJRWZvu9r
NdSjL4/LvySIgaxbGOwbztqFbVue5VH8CLs695qMkYxHPGD0hs0Utge8pW4bYmGd1SXCxGjHfrcK
L0iZlKDK2bUzlQFfuzA324RnPDbAXNDrrXVD5FH4qQBM16Ykn7XJVI3AlqmGpugv2vn9lQ2d5jcz
kytV1LV4tzhajTX/Nl+TlhtMq0+H5cCDyWWe0hU5sUKpexfFOW/b0FCxK/pAHuBmw6ioxKfW50HE
LfyfOM1UB/qo2BzCxggQqC7eF3R9YZJ8rVKyyw9ppV9HBGbnY7ha7HK9ucHY87Nv72h0w/9TC/xV
MQjaSdr6SIPW4bMjpUxVKAxYjct+ecWqOcg9d7Aix1KHU+Sdi07PecoBxu/+ecHb8Nf+su8QrQVN
EHnQV8xs0/H6psb6iJxDl2mFtbz6uymUy84XKI6KrRYaVCtYrYPeGIlyouVHcm4Y6V4n0gmkNZeh
RIazClnM64XkIT/Y8bUXyjdDv70g7jAuo4ngrXGhzbTAHRE+MWTQbRHbwLI7Td4CwGIXXgSYgEsD
lZOhhyPZl8alheLupcgYOxyJEr4mhlQc2skl9al1oWzemz9tp63vbNriItyHvuFiPJVOkGZz1iCM
Zl19iCGdM4rJUJ+eCr8Sdicyqmgn5F9Is7+J5MfsNFH9NLaIA+iTsDoiu0rBr1dpXUuxlJGn53yo
RzV3ZeoGD9aBj/j663LXU+4AAXT4siHpftvv6Wadg4txUTw1ZwjV8gjE+RGQcyqjn3LcKWLcqbpv
HdIsfpdLzQ8zgs4pYhUA0kpClIrFermYmtRkCYWhHW/r3Mu6FkRwy77r+fVbUInEymyETKzwEJk0
P3nzp7STsWCswp49bVi5JrePCopnh26l1auLPhs300MkQ7a78En/RzNw7WE4e/dCzZXhBsdlHGnG
UyMvmJUoToWoxkzEr0Fj2CCvmcudLzCJABDrWnobN3gpvA4K/XLwwVH2uWG6hGsbGIvgBKAjKHR3
MGeHILJbi/0f4vTlMbNaoTctKxttHRz2jHIXMSxd2/rUWq9jwhzk/TinInU10FGIzpVPvwz9/1In
wzvmXTPt7QsI30nNcxGpgS6XGBgFn9VL5tgYa2mEg4kbM2gQvEefEmw+Qnqdiqo+kMiM5rX/Irei
CuMNBW4KaR3rZax8Wv/iYvTu6aGFrFuZ4r8tUflbseWUHDT6kvXTYxCGlMC3I0JERLjgUPMzm5AE
KK/shudEab+g6+ENnLbcUapIiCPM2zkiodP+g0PvsTaOkFiyteIbbBcx9SJJr6cX2wSWMq2ISMoF
WDXKvO8+SweOrrmHDgEJnfZTm0sm8DFl2ikBqOXmvuLqU0J/ZmvKovD2/jOs/RClKnLbmguCicO8
7SA+8mWp3C0pRaEIpEU7UoRae6GWRkemUoAUfAAwTFGR7wbNIFNKTJGcG9WkAlAxv3W4d3iEm91h
a9ByFznS6RVg8z9xSNvDxjpzGKW4RIqfEFENJ+76FFNp4eZOY4i7cPjiJzGqjmoIc31Mkhgj8um6
MSzwooz05bQqIoTao6EG4cfvD+PF/z22Mkf4PthbLX4+ct1og9Q0S8ZyUZdzz0NpQoLiJDVBCUqo
ZnknKekCEnBmwbcndLRLaoYlFpVeEQ8HV+hxFy3mYFHCb4W08Hq5SJPCMXcQZV1Q6+cYpFi2Kn4b
2KgKJaMfF2rAz4fhCg3xJOwC3hwjioXFhQ1w+Q9Gc1ocVAHDE9XGkGJ2wYBRneFrHW5ckcAL9uRy
m634yB20E1U4KWN4ZEFPNSkPm3XEiSErs5zW4PuZMNHuqeLcJHvgGQhLT1HAA+ZcSahsdb/xYiDK
F83mpL838lpX3d244xQQr95qy+wr3W5TzTJBjPc66lig1Hx1HiIxS0+8DrkgI/9tuy8KV1NPQcsq
YVCR1/fJS0cADyELn6GvqzACjvotGYk7JL0g2Q+PgwLecZnPswYVe6hN9E94YKU8tZZjHOKmVSGv
h6L05EUb+l+hiQoKD6ws50U/aHxR0Ft6Bwg4yezcZHNE7Yx15GJawsOIR8nK+rA45mqOUgx6VLLx
Fz3tDDGG/Vj+0wg9jZ7Pu3YIc4335HY27cXLKRizGoZ7tM4VljOwtsnUTt2wF1nYlHPV9BiK9EdM
7n+bFUlWILVDuJZQDd2nkQxkUZLvkWuuW4fLkUe8pC10S9b3Fw7Hj9Asekl8jH0vMYQoaw7g35fK
Vxa9V9FcWkbt++Zy7Pz0z0k3IYNNIwmldfcCkQXiDP7KWcadIyaZxuv770n3ZwwZe0DvNs3XUxNd
MvHUGPhoeON/a6e0KNIenYI0q46v+dy/1rBc/bt+IR8d4z9iM1Akqs/Ozad3HlqlKSS0NAxrmB8X
P3maXwMl0Yto+TpufxG9taKzlCZJy/lw9FFDc7m5AVEcqLfoDjPubv/IiBePh1e8c1D4k88sWsHq
JtNb3HbTXSdV4KdNROcloxsy1cA87VKmh3cAqqBG4MuWj6Pk/exD0gafVFEYSZl5Z6CyXbiWfWBL
AkqVzPWTB3/KOfQQUwfSo0qHHztpL+br9cUihQ7XrCu8I/1WZmULoOkf+GMD3JXhG4eDmtHzPIot
tYJMo9KExSmIhebtDHcfuOGd24SIVAxurEgEAWlAb6Q/56ju5zM0T4CM+syqAF1ZA/ZsFigwZAZl
iITLIbTNS5CcdhyJq9hfDgzvqA4ZzBV62FEr0QzxIVBkEv3npIlfv+6xWwomDu3Fk9IHsfunzOyJ
4oH47O7NAC3UttHIKcetr+z9vfpg8a6lPQV4OXCl/PNhEtRJ2Ehd1qHDn15c/7i8mIkbGG2OmKMN
K81G0P0ynt4pWm00qtlQaPud40BeKJhF5XGK843x31Pomgd5ZAMzp8f6rEAYhLEUcxCLUg2EBtC5
MvKLnVe4pMnWR3+JIDl3bUkK7S+tLhI8f7DKuaSNc+J3dWIDNT69jYtNB6x23kOZKctflqMRWxXj
8D7ir44X3QzJB9QeBitRI38oBZdJEP+Q1ABUlnXLkG+6JgC2vmhe4aKBFAs4+7nizykW2Yl5cloh
hayhqPM9fSSOwHpJxeDRXONTWw/C9yevq1u5Yb31rrkpUiqE4JdkGKeTo0KE82tKg/xsi24u8mh3
x5O0ObwQsvoCA3T/89+DJsnoHvoNsa/VLTcd/rgk86QVwubcE/BvdnI6n0wl6acyZy0yyBBr5BzZ
LiOl6zdrziHDsvCfFVgzv+c9v2j7gJZKdMxsN9gWKDl5QF51xNZqdJJPVBKB8DQMx449nv+kB8F7
+EPuaCOsz04Orpa0XoqDcd+gs4ggpnKVwlNtRm/R9a/HNIQpyhKvVcAH6GA14bBicA2cZqk8uRlo
gS+r6Bar4o3ajUjH+uPir66PHwHGuT36WDXkcLWMz+w35tu51lpLCDyY5vTyMZpPPPu6Xj+b7GLB
wai0mPUS0u6Ht/LQzlQMtSDgSgJ++cSh+xJuTj6h9pcZ1lfldqg0a5qHkvAX+pUqTlfDEUmoTFYy
NkW2095qBDJkMQx2+dFOy4N07kdgGw2OicE9fksEWyp4uIsZe+v2SzBzruhZ2yb8gxpx2nwAWp+t
NeZoQgWFAogoc3eTsdTNpZuMUaAJkNlU5BG1D0EU2d3bCFiBJM2POY6304fgx0g/WtQzC87oToSu
3AQol6/rfM68GSEJ5Z+bD7QGz5t88hz5+toN3SoyGP5OOjdCblItqmdWFeCpE9wbB/PiROnMfA3n
2+hv7ih9qAzjUipGneOALGP+veAd2kHb/NU4eQhvWfGt+wChBPq7w1QKzuZJu3QjRM8XeM0txNYg
vSgQ954jJCY+/wQDhuuqqGz6NDgFvQwDbTQOesWO3eRcRY7H6qd3vpW7rXEMi6iLD305opUfVYV6
/CNQ8/zt/k3EJ6i1Je2to+D8xXsN3/lgNP3XaNHBDz8Ef5fxQffA69hPKAYLOZKTGR60CI10Jh4M
sSAvv0VCz+WC7nE3z2gk3H+7C07DzuIWDsEDJH7afpCAg2EXA/0F0AGxEXbm9y1gAkhEGKXwV8uZ
qmPzY0KlwNNHPvJZVmF2VIz+HKTUBFFx/MAfFXVSDpC4JCMh9TxrgsLkiAq/rdedaC05ZuAv3aRt
LxmiwCuO/h2aiYph+TSvOBDfJ7fLXMCz3ZdBhk6H7GlDjwp+Yrmgr1zErm/0a7WNqp06JUrvSJtU
3m90TVsOUa1YbNS1hOw2A3auqRch9bRBoZ+Da4Yb38p+SFbzZ2xlPunwHCQdI4fxeKQDV8X70p6b
l5QFZokfMeD8UxRaYcM9c73TLBy8J8NXRsQZG8I2Ckj91Is1B7/UoEN3v3ANrK0CtgptzRAfGBMA
Yma/5eV3TNbwqCwuXsHXmNHNVDdUDWGXSbY4oNNsmC/I3tyS3G1H4DVhItfZlXD/ZGZ6FqvwOyjA
l/d3hsabUT0JNt1+Dhh6Oetb5ivcpUy0uixJI3qEJJLj8t3Dra/pOJLvZrpT5WzNF4UViAfY2sMG
wSyxVEnLS6WU5MPBvMvTBnIxcY6jlVy0kaBn2GT3vw+73GhagsxtxJ4MoVbyYQ1OG9HVZjaiCz+C
HQGuFcX9JpMp656J0WWI6EQ5fCqHGVj8lIWuwE9J5q9AiYclCckFL+5rwBxlgCHiyxqEsqCEB4a+
PAScNVuGRuSDgqg1SG0J+lmYZBdhc4XHVaK9etUaLwsAQp/v3Vc+TmPjNief8lss3dQfBRlXi9aM
HOUQJtdJYQ+2RurOvVnG4qJol/msk8NsxU6N/9GtvZHspGQkqW9bVy5RYcpsBQSVww0+aHySN1eH
q2CFlQ14Rc3QNQj02+2EdAhsx0A365ag3zHrOd5PanwZoxGELOrKVAuZsM46b+SIvk/T1X2aO3JF
WvpmN8hFOEw6TRAMa2voWPUz2i9kC+R2n0JnyUQYEozr19X1HUb9CR2lorn9ic9aUftecABYazrs
l4m8pt7NmtRAADMNnUg4aWF8NzYV5mZFNxY46oMiM8clgbMoxvvaktwiY9m8jIdDl5XGavAUc7uD
YpZvulttCGpIdYfWCzr7q8eFFPcl2b2r1DAlkrHXIA8c7oV+LAzvXXxINejOvbEtnIcNuHgX4vB+
UX59p19tbwkKKT1IWKi5hGdwLyJ8XM46/L9/1Ah5BeB2RqhqiB8CTKyLJixrEVOet1w3SlL54Clu
lDH/JGv4kH9s1wy1gtBCm5Im61Gld48OHYagN1wZZ7ewb6XiLSF8GIwb/Ei7LhoXGSDhOaMmBYpt
nXPJ1A6sTkqPvWcOckLL+FRVXIN001GEV6m2AKDSs+mfibnOyatksf8FoSAr8ymnDf049V6Ehnpa
1I4iOLx4InsPnT+Kbs9qrGiZOpykH/NBcZ/dWO2ffR/Voy/sBdbAUgFYV+i47sIMFVEBk7zcnhvl
D21SvjeI0HifOSld31ArxCIdTfKc29IP6PuSqRKvE8//A5B2fVNRsbPd0zLlNbC/fmI527o+UFmA
kPc6rGi/QnStZWpxd9kGYf4E2MQlpOIl7yvDw1CxC58aJXJOLCyNvtZrSkVTCHjTkznSRqeEugpw
yJqCeC2FYzZ/YVfKHG4Qv22cXW8XQpW1ZO4KGtdiaq389J8GPxKzebh59eeqBWNg/V++6/fSIfTa
i6noI+b53aW/0RNMJDWF3Ur6dq/Z6GcnSS0qpU0BKr76gU1bDjlvhmAQK9dzKdlJeBRPAlPu33V7
Vyck0n1OuHQXsc6wlfkkVgPPFrcuZWig6yQ2btW6e6aRC2NqlmlPfUxZyxiXNwi+n9Q7M5uwfGRB
sT9xwZ0HbPsDTQEQkrWweRnVl/vjxGJkRWMo6uXblJviFdOxtTswJVeRET7zQ1fu2d5tHra+km4I
OHXuJSoW4zfnRKuJ3vTLENqUafeDNxhZ3FcOD+sIUabTrxfZXWxV21AotIcdgPjmFvVK419OufNW
Ii+nYhSKU513oeY7LXWUHsiTngJ8FvLo/VblbLe6sPR9lF3x8B65INkJEZZbrushB3ua1zu1fg3i
ojAw+j2bhYoP5ugr8Jazy7P7plwYHWOhSt5UPkwW1eZlXr6xMcx/1tmiwI6a7uho4ChOUaM2hnyX
zQkFbByhkyXub5yZYcwNLPDLv0n7xeu0x8jUPWvsDhsv8WklXRa4pDusL4KVW2yOQIoADtw2WhHO
mw+ARlGKH9neRRi4X1GBOPdblEelHH0kWSn2JwBnrpH8lWwyuOqpU4lqQ2G8Na6FDCLT/2BfY3jC
kGTOOvzRpG69aAcRL5D4qIoE2PoRkMKn9/wRrKSApobLjlVyi4V3twCfGi1hQzcoFXlneueuuEZI
tfDw7S6B54NiQ5SXslhpaJ5z3BGsYfP4jLxmO+K5eMyqLvPnsejApbnw7i9c+U1l+nh03A9MIte6
eTWusnRe5nfZIOXdxp8auDrtW4H2XcRbu/USDcpmfJEpOy3uwzrLpwYlgxF8p11WBhs2vA2WUKLd
rvMI0d6+sDF0y5fi57Iez4JfKOqg+jjcXfPqqdKjgkYUcKAi+8b2G7kba1C3Xv0+QS4H8xTkpXdQ
smZs73Q5Pp/Np8eC0ISjbIQTOjY0EXMNvQ5IF7Swtp76vEb6w1bxAslo6Yv3tfprS9o0cbtT6uPb
vBYRxTHIExF/RIRee0EhNSlHKhi3XYgmMAJpFV9Tvw2iOELEbbpMTvAUzDSikbIbff1f4uETx9Kr
9F1uibmKx4SRU2CMdGf/gkHYi4oy4uJRZCo7NgGceJSWyE30doLPoRZSprbcZJm7GKurDzVD/cok
6eEyRiXQc96fXpDbzZtIjI5FrhIfBqMzxkNS4vWdVx3gAvM1eZc3j1w9KAgFnPQaW/yLfokDSZg4
tGp/xIDAL9EuZX2SJ7nbZBmD/odycfpndYrxPbr19htusjqdrlBasFdmXa9718xqSxponG2yurDS
ZReqtS1Lgb3x1rOJL9vI8+O8mjetnu0NQqX/HSvZtCDkyKIvAhIwO7idHf4/3jm0VxK7ZjUDqGMG
mBIXLb5122lyA15lS6BWhqS5jH5TpW41CqK2WdmcDM1lHT2zU7vBisJcKPWyRpI9js5CEwWDfSHs
Cymyb64UC0zohtUN8zp6TVPt6oxJL+XM+6d2njSg7KhReFfTdZDIC1NTwutYajrs9FxyUf9MDSfp
KTa3WdmAB8hCARxQIr2rosOY8WmjV0QomCrUt6osEWaSlmU9blIMMECFAZlDcIGezmKfjKuRwBiK
wT2TXcEtPLLj0wdc9+vtIMmI3dIOcDreuQgHEYCUekuu1081ijXkLroNmZVEOVvm5Zv5iSiRKR/x
c9bFdAe6oBjBIXY5jnSAoPfnC3DqGpiI/sbNfOaVTERTPj9YE6lmW6aQ89UOzFDtmlBHZDTGJnY0
GwSDtm/DNFA6+rVHe+1fpNJcGqeauciXSxkmjF9o+2I4JQEetn1WeAo8cfSxgq75mjMLSBi/Lbof
9CXWGl0HI9aA5JTjpqMXH7swLjH+lb4HEqLJ1nzQlSYFBpHunA0yAbyDIjZ3nMIKB8ibMlroEqA2
JaYTxGLR4MiGpwZrME/pM8mzF2Mb1zZuv5zPhnUIpJ/zB8vcNikFvjRxrwyOVlYH9rqBChoZA3Ro
9fPGbjqjF8CAx1qOBiUzvxDR8eog7oJNGqTlb11xGJrV8s4zIVppXzf67MHSwGPlVothwHfQH7oy
suKi2gb7M1jy+S2+zZAW/zGPbJ5zK1Eatc827r2rJGIPlvlATth2RSdpZ/5CkwLTLSbAIiMVI9T0
QeIqlSRYOLKXcgd+A0spzX4b+AkwZDJ/jCL7vMKzmpKbmY8O83MYa7oLSdzb3/eUGjWwMhn3s/XD
QX1Lno+c4qLrfDZbMFpxyLyLYfFXVbfUrLTDZLyirUh3eOSTEWnZCxOHo+MHskStgwcgHLDkUyA5
DpVjFcMVf8J0Yh+WD6Me9MFt1XucDv/0DaZYT6UTfpDDmuwK/0jYNjUpBepPmWxntMm91vYIMQGY
utq1/OXMSSbHQw7pm6SwnJcGg9ch5EVWrX0+O4liGs6YzcP9VME6gXzVyN48fd+NuAvDPLhrm6kG
Ur0fpbwFgTiH+vJla4cXp6kxnGJDuS33tn2PaJdV72QAdRzbfagYMcS+fhi8y7j9omNAmaa3W6OH
DSyJFogCyUNOoHHOOlwzaeHsFtmNCefffjOKMBUnE1SsZeU24rfuV8v9SvrI/FFh8wGMOuRnKAUw
bFpUZhwH5P+lOjT5eodQe9It7VBpvohOGFjvGwOnjr3d8090t069U3bm8/uWVnqagZrN1+fIyXRu
OfCbKyEHGxKoDjiTEqxc2gS+M2euNh84+zJBRTiZHZripg+Zx+hv5VozIytxSJGOy6IgOVuB7tN0
Ro3ysGRT/WUEYMmP4cmpNQXlWFiWQVLrAybQo4QG9Lh3jn+JH2sYkGu3Y0rb15xmPka6BKCuGaXk
TrmCej2EnXCqu/aDVkWr1yn687jXVrgJGtqxq51IPbnjmRPCwvLC9bBfeTDNn1HXWsD1LvCI9t+Z
LXV/9aaYGt/QGAKW+4q4xeYtWNJ+9qWSA3DawfKPA5CbMmWRVBp641Mavbga5GLrawemDLycFBCf
cobgEYtsQSL4NAIRbwqMd9ZAjb8lXPUSHvKuBjTRBBJpi1xdu1nd61D9HeI0omueuKGBI06tGWfR
EQEdgjNV5h/Z0NA/yaBnOWeJ2p2yk3GEx0wlnBkc56NP2wmKF/UemI9OaSMhoV93s/ppOLalGF84
y93Y5x/ANmHlpH6WjRNLJ2li6JJnvAVb+w0rJ5WzX4nCdU15tZMIUZiQruANEq4hw+7CLGYlcz1j
NzfQVblPICMuSrgi4CGU2/EiZIXt4tt2UbkA2ks1Ew0IGtvrrIkSE8tFUc9rY/ZOryrTQ9ugjQoc
2fA6Hz04v6o6MK3r/w+WXtCV8/CkH3OdaZNQtexwfhRldH9H3z+HmSXSXiCzIl61SNTzQmpUd7CQ
FmmtxomP1xlMtnuB4ZA7DMEO7RARpxfe7A5lkmulBNuqwdfgJkYNlBJdZsmvM1h3IufDElY1Umze
XCBUmLdZSao+z5HGYpalf0SYOrroSqbwQGvSRo+3yl73zl/ECa/8mA7FBjVgg5lMsA4TMTzvCFPx
fQeKL3cQLhZ2ewViiLkEOQBfkgzRof0saCM+HDGT0yqhW9KcyAqXP/51bxXCiLXyzdkMFSJhTFK1
B8LX7Ex0uOZYfl5ahSvrULOIUcBIekvBEOpGGj+iFgPakosprr/O29wdGGz4JuYkSWFsw5Mgbz/j
ZSHly0L9WPo95gkMkd9t0aRRvHncbuzPp1KcZkjpLcHTX6s7Pu/FiPB9gNw9hszIV9hoE59MTDVH
HQmE83plg5TvHjB5kNbUONATfCPFjI25gQC9WO2b19eFF3lUSGTpmjS3djhrNyeLoVSUBVslzHb3
MRQrxKZTonC5M6412Lbr8ze3ziiyj5+vZG8+342LJcXjHtGU5gkY1DjN961A9ABbxUT3sUC0iUhd
mWA+nTiV1PCxLLyG4wMQPt9hSgqPtzX+cq11PiePXjPNqbrfDx//EhbRnLmamsU7kJSNXZIx5mNj
WL8g22/32J4phsh86Hjs9Wl5uBYLNTGwMjjYLgJKwOW+m93b58+y06yl7hYUNhdw3vLDYubLoQFw
KmXOKnRKS/0LwK/p5NzCNeG5JqN5mWbmO+RDWDlZG+9XDxPkwcROj0c3wIMA6rFCjctDHeDlbP1y
9aaqVe8xSTP/YXhnD5ufd3l+SZCaoH+KZWU2Q21xDE/cRsxBcwl0GU+jGWr0syajXSgo9+1NUCr7
2OInBQAMipqUjzcH9Xgv6+ydRvMcLscUrjoLUj+vocUMtgk+uCEEJxc1Rc8NPfudE4eBmZGXTGaW
zOYeAlUsRhqocqc13TPX65cGMKIc/nVVyDWthi6qQJOuy74orwG3TlG6xMlY5yr/f7k5ZQWzATz+
X4IlwJXix+nfvlvqsFcTTMOuvAF15vUhanApyS4Zs2/M+c1QXFSDseup4TrdrMMAR+a49JQ2Palt
FPkm+678CqfZB7LeLDHYAdod9m1+QGxxQ16PctQdWW5+QeA6ToKALQ9SWEudkTanTN9YZjVntL+b
ZvtchTtx2t4Jog6wjvtPkYCSBcxnol7703ZYxUuEaJtQsb9MtbIhqHjtV+xZ/j+buRJP5o71v8pZ
1l9N4cHOwJrqun5/Faqi8uP5ASQO2/aetS7x9Qf+Ox60IGzB49hZznj2daHaqVfGeoWIuq7Ppg5W
RAwDPFHpiUicv9DCL75RJQq0dAMtDcqmP1WD5MKNWdsEo8fyu33c28IbN26GN1gjYq0tvoHzObC9
0NQXYIvOfGOuRySOmcg76jWZ15MgeWL1IMd3GHtrxBlEdyRq0fHsRJj8diqpiKdcFWhWiQYhQhXW
kj/BTXte7QN5XBY2cx5O2usfNxIOW2gerhyvrDwYVtQcUskK/QA36ZDO9kbXTd7B2KJEsi9XST46
5YBy1xTUq+BaGoYkd0dnYmCJ6qQk5VhqyhLfS3vHuOGdjpWcpKLXcF4tbg1L0nzzGGECX2pAcbkq
NlRuiBOrFWaybSFnKs5Qh0e5oHZvwpEIRd2ShKwZxtoOiILeAbsH9bZRWN18uR8VW0yBCT7dnF3E
BvkNgeadH4DKRPnfm/fg+I+WdEUYe70QkTBPsDqvPJ/bkZaqJaHSZTF8w47zShBt7XRFQSYaMEnZ
V04fZ4m1rh9m09lKD9ykFKGekdkIpS/QPs+C5JF6oorb5YqTnLubR8c1RymExj1xU7UscwGNASJh
ywZ+xrHzvAplbV1U2G3fV49C1v9MenAdsCUHEFToZA5Ql6PLpqe65RRVo5pLZ91+okRlfj4DoqK+
EY1jSoPYWGN5qWbtISOFEi9YOosYetD3WQHS9JI1+Mxmx6p3YbfWSboAOhEQ5a7AgxvQLFKwDDT7
0qUJpFbDsxmF2n/K4PipzKOB02K5HxCXpzUz2a5ouXPXga2hcY8VbrKEW8CJZn/1cPqXpmLOhyLk
mi0FiCAdaRJIgSOcjgAvXTQH0MPVfuz/7pX1dN4/9tz/XULCk88FOsDBN+AvLM3LOYPD8ExIkXwE
5NbWXayBR0ioObw4BPxm1uv9uVzAO4bHLJckuhx2DuauhBWNFUQZ19FC9PYrFzh5ZJv0fNfC8k8m
WkBXokrjozxfngrB8p8XbsSdlGPHId9mG+zUEnZ7BzurMKZLed4jRU5CG6eUBXOU3OTjBz0bIb39
xJ83pFqC/ZR0cQ2hKBEbu4mdOaqkMQmqvPNSKzZN9fF6M4tQ1U9BzfSXnN+UwLmmPq48a8J+g7je
1BzVz05WpdSo+sz1uwQ8GWt3U7F+4OHYlHZHtR0eJxgtkpeF1VIbavjvQwaV212F7U6bO3hdXFeT
50Npacd+B+AJarL1Ht8OlmNYYsQSYqkeXj0CJZ4spxW3/ErcPMYVNkGQsdqqP6hOElTnsfKiTD5B
+5xbqWofnqErPs0NXoQaHLqGoNwlxQYZzbtEchBBu8LmjvCQ0s4iynZS8/5KFseTHc5TlwV4dUpZ
H1RVMa8uQSJbOZdVOPKZ9tqL6EJIKWBKMCHEpD7dk2N5MyNHt1YeCINCL9O2wUKvmXw5bg6gJwPZ
PE7eQ9xzXFpPQbatckvQqb0gCVG2rn5iB+CIUqAUFVaS0QumEn8Vt6xTvleKKcS7QifAUU9g0PYK
rlope9jPiABlRraxzuP6KLFCzTBIW7O/SvpspXyi6766qCA+gaR8CbE0QXLPagfzeg+ZhgfYJCnT
bRzeQ3ZDpa5HACTnn0jitQDRRpyMiUO5fw/riiIagXVQtOqlQ6UR8JvIV95akS/Vyturaxe2m1uF
VJCI+x/gMxwlO0CCWW1c9rKk5hVxDDRXvH70atBejgiKb6U8BTtsfaiuSDqIBD4NGLbpoauSmVWD
yHIR6VFdH695vxHVecWlKN/Df7HHEyEmz3M2gd48Di1+ZWUWzv2Gxx1n767wB/oH0tq/vvDegYk4
jbV3FMMuFnN2H/IOKXZumprVyy9k9jkCG9mURzsv3VpirQT9dwq/VKJiEQKc8iZDUlsOE1lG8YJJ
mYxvr4mxdVSsB/Aa4kyCrg/wEz/Fr1WpMo8dnxU+g2yr/iuo/UnmHcKxVoV/JC53PJVMRbZDY0R1
TT3vbu3M91+ulxEafA1whCyfXK2pML88t0slydzMbrcJJY+yekdOVtKHKGdB4xJOxg4qx2IEc6rg
+RgYaJLt4j5OIbqC7XfQYwwwq2GGKEas9ewlgXEjzABkI21d6CyVUwDJETAIHJ86q3BNW19xYSpe
eWsHXfw9mOA8u9qUmMg1FRmmSzJ1bZszvyEAlVSFG0+Wf6k1bJ2TkceF1bxods5tcwt08JUh0ZDk
p249nvbkxrG6SlqxqYYO/epdEQvhahYORynRO+fPWBmTmuTVRbs8s8DxrXZwaU9AcoH6wA2kVXM2
KEdcMMzQ1VrB3iQhHFCTa9TzZKgX/fmhxvAGZ9tThU47klfNNhwCbieIlaXhHiCcvBWFnvm6wPRV
hC1jenCaKZQGFaAhLzyNv/tIgVbwxwfasoedrBHajUUHIdLq2LBmocnTAEE/Xb9vpl68plhzMPdx
yZo4uBk/1h7W7VKCm1xtmETcWAo7CEEVg7gn4rWEPHty2H68wi401UMj6brAz8t2b7bexxa6fkQ5
By3DGqrGGRXh4i8uroW8hb4gPQPwockRFQ6ebJCsF38kNwk1lupMSkjkiZDbnnGcNKZqn/k1fNaV
DYejj6rPGHu03HbONwbr9aMOkv71RVvOcRqB93CbNy50tXteoy+2vbE3u4EQaJqr/gBXzkNA+MgR
zdml0uZYQtOSVZo5PSpbXK8NExtrx52tG7hSV3W2CmtamsgmHbiTJ4++j3MRn2LTWQo1sArK0mHN
7u5Ye0c30eNTPNkpRpz14K9IBKNT5+THGlYUYE36RAg/6cL8O1MqfI8E7yxhJU47CPZhO0npsQRS
lmab/ek5GrUCkrTOv/DJ4JQzAOofl+zwOir9PVDW2ICYAAC6Jrf3RXHwR11LS+VkqfOBjUf4W3mp
ZvnMa2ik7xyQakaOjNDtGs8E3/VGgujFKYcJk+oZMmJuDw7wGbVMPxM4laS9z4T7Z92wJQ0j1BNA
hHbh+SIw5+anFK9fW3a5bHl4b2R46l/xhYMelr038b+xs5l+qerQ+hvel666Um9FVmNM1ygTVfVe
Xw0TyAlkijvhEQKebf7igRlrnZosDXwhL6I4JJHp4GXiBH9OEhnvKeRIYN6SAK2e/Sji1YeaFog5
YQmeAO1Nxx+m2c6rKDgU9orIu6qhsaacUy+cvn/2LXBc9I5HpdDEG6UgvaT7Vy1gDRDFbPzoQayx
/zCChWR0A7aN5VzwW03+/wiCgpAU9jdyM6nGLPenU435Y1Zih1vEerbQvSqbvR9zcM50u4ufCGwX
pqMZ3eedEfG9Kv7rIvqJr0OCeIdiv3E86dvuJCKwNuLxpm4LA+VDvsm4/M9dqoEOuCQn64puQdYC
MvdQl4HtJpLXYgqJsUAJSiriM+hJsWGnSO2+IxEr0vyKpYSz2Vueji+s2+hEXCfFgDfXxOK3tVPR
ZupyAQtvpOMHV4EA5vHeaW5pM7knH8cvs36lVlymr+o42cRIZHXBVa/WxfDnmK5K+Ufv8Idz+DzJ
5ssYEDutyoPdkjPMt/7OsmbnhoOH99kNcQjRlN79fRTMRH/5n5VGdalBpv9eL6LvJ9zKvmIMBEr5
Hdva3h9c3aQfxjaTqjY0qivGxL0cvy5mU3HJb6zMzhy7M/MCnkLusmsSHp+CSSr4gQp96tmGPuSg
wbLWJyVRg5TRl30rJ1Of2SGQ9EexphdfYSB6/GBR0J/yQ4IA3jFm57whvxTQ6H3jtQebP065fPPW
yA74rxQr84/5qxoqzYvBcitlRyygu+MlAgWe9rpIvbYhh5pzkE2kUtRFadi2UA3pguWRzn7U5HY9
AQL9+y4ewYhGeUzZLScSUDP5S6MQFkbNO+IHMR38H16JIC/mTjHylLjNbcJ6NG4qLYjL3JyYZ3jq
7w8PWDJIgjYfWaRj5OBq7O3n+wG8gupCchrL5jDwIORhqqF4IjlRrlVv41ALPBlkSGSv/bx8wc9F
b/t7+fJiLO0k2pO1rL/pKn6r6johKA6DzYD/n4dE86mj0iU+ulPzkAORLumq/tYXYW08C9qYCcqi
9mNoF1YYVFC9/LE7xZFiW8jss6dt1t27YtX+p2DsNIU4ZeiYR64jTz35MatrhUPxcNy627ig6GCQ
617TWn7T/DNnx0J8ZnBAvo8VPvB0VmIseKJZeoouTwU3LA46VsjPlveT7C0cqm0OrrpIEfRtNZQe
xWSNxGVwZ/Yzq2iF2RmPcUPHxVjwbGgt3SjrpWAzb+fns+Vx/cvaVk4qZDjAVK/3PRFevPtKSOoi
+jnnOGvNNtuwruLWCCVBrmvOuWrU7Ab30N9sXWMuXggDzk91mNyHL6KiA2GLB5FOG8u1lEvWioIj
3FI570Ks0U7nPsVCUTMg6/PJIhKIWf3yG/EqlIRN4c2M9ov3tYtn9nPHBmf0V6XejEgj0CztIBzk
jAlVNQCrCGbVkpsnZKxhhNhqG38CJtQAuCyof6qKwTGZ7yWRKZA7m7e7RhZsBzuELAcV60CKgNcC
XgAUfoMj/FLVJV05AMuewf21uI3xcMWxVC5qWb5t78wtmPhEGPscfMJ5yMzCYTCW+gfcO6JX35h4
RjXT8dp2bt/E9PsrZHW4/PjsseugPvrmsKJEIqHW7lCXuxieT0wRTt1qv0+qPkYXktAYC9D15P9v
HKUJ3WPPkEo3lZb0+kwVU9fo1VQYc5FnzB91RM8M5MVdgWcfm92GEtJAY0ISjpIWEcO0B4H4mT/l
0KylLC0991iF2+4ZdhGhoCT4oXHOuBlNsOhWZvvGpcxFBn9atXN+EFfCrn64VUEmkAh8uYMBlult
SOYJSqtKYxs8O4t4wMd1LY8hIjcjzANc3r7ppV1nPSqL5l2iNrfrtiM7iKJyV48LBvs9CbmhfXZh
kt1R2JKd9kOWwXwwN++OseplbRmLybYEn16wY42TMTlBPJXt7B9Pas7AvW4yYwEwbv3DaTXQeljS
SAZoyYJysVwhzQct8rlGuBw5bcheaTjU8EBOtVrkqtZm8T6vNak21jWRt7VrjZ6huUABRNS0n6eg
o5oMZ8RmVUUubq6sjsfUy7V6V+yuarfujfkLMhKm5PpNnEpPjt/eRbHk97aKILEujUkQv3Etf4kK
umC2jtG/8OnErY7F4uilk6evWaAGz968pvQa+eOlQ4Bs5Da6Zg7t58pGSo44OG/2sQDbOig8OGWX
nxM63iUbTQxYK5BQhI+JxfMcWTiccz4xXtcMaetctoZvytZ9BjM6wBMwe8pDJ0+AFI2JmPpZIvXi
oOrngfUffveKaPP7Wld7BcsVwr3r0JIDxqO8NIMPj1pJEhdA6k8Y+y0Khutoleir3gr9yXu8I5qR
e3HdNlHAgAy0YQ0svDtuVsuo2zU2rjyATdxwy0l3TtfPLQN8i5UswHUTNlqs0FD8F5KbGrt+Zk7m
UzWw6a1Q+ThGLB2K3s+ntPOEKp4rAKKkv5hn6+rLwgPoxDURidjYGy3paFBg0pQa6o6q3AVOIgWQ
ftdjpI0Y+hgKWkoCtLGqxiU5g7kZrvH/9VpapYJAiyeZEn6drCrlFY5kQlAdEMeeIJg2h1wTuqJR
K1BjoOKd8jclzSBJ1HOn1wkwUCcYZ2sDdr0guWQcL2aWYRDBOtiHjtH09BMupujo5FoSQW9oyWSC
jSgSVbOT5dVlrrHPI6Gb+yHlzvxr9c0sr5sz8JEg43cjqSHlgX7QPCJMoe/wtiBLRAU9gbH892w3
MNQAi0EdGcF+gZp4y1lgJy6xTg8B0Afk089RBKMj6kcVcIUCbAEGYE22HbxjflMzBxRWUHXwrQZL
2W/XDrV6jNC7aM0C/lAjByB4ukBTdf5HhbhL6fWRgyM/T81GXqSxVfsyIUACXMmMcfhQxzxdkRGD
SDF7MheoH9zaFX7Z1dfLhVt47BwnW7LdA2lNrMyRmaN/qsG8Ikux1Bz8GPNwP4Nyma4c1x0uuff8
dKqtl6cJAo5+/JVYxEEng0tIiPcDZa8mItBJgZnTu0MiOxzsTWkTTttyya1S29LQkli4mRyp6swg
8ULXv3MhH9t2K4+OBBmtZHocSvkH9FZXgEnrmC/lEAyOX2sYDjyQgfRhkBbN1TsqIsJreDdcpeHX
S6gTc0RCa0Y4HAiwdIZHGT4uJrCr8733SyLHliZqqPDdE5tJtmCPGgqEE4dj+nt3FzzZQ5yDf7uu
kdsjC+vz7RbWoRl3lfsJlaWC4/YAZ1wlJcbX+o/PxcJct0WmN9iX52C2q09SJloF2qtimTU51yCq
FaCyQONjx5ogLc40cobUbEp8i7sbVT7KXDB+xGwWG7s0MbrAxyff6ctwwh1yL7d5KVpN8m9l5swN
dht/toRT6BwmwFfbQbyt9g/p1n1pkzrcY5zW+2hj2q45W25SaYCL9LVUrvbeGPd8h42njxR+80J1
oCzLe2lHB/w0NY/Zcl70lT/k8ZIow3dITmKLPfeKFihfbtejSHyvwI6lIn/kh1r0HzhhIj6hUO7Y
qYyihuzmVPCXCW/ronjo1E8ckS/Ddkn9XKyuIIBtuphNB/8WsfN/zv++f7rsXVLremoh4gTjy80c
kHr8kIoUs1lswHV10ni81VFl/fYFPgUbNoE1QZbeDM7/7//j9AlSgy7bUaDc4nCjIMfKBFimQtZL
KWQ/QqMP3wzwpEmM54sybCCgr11kSlVna+av/GgS4j7ZH3xaKTy/R2JV+m1IetSZzW0BMV5lU8id
kxvpxnheASXAYzc/gtpasMyGilQrCiHuawWctNajSStqe/Xl+d46Q8EYm4ITE1WUAOOehTRZieDg
YkY7D8z7UBhlQA6uDRGKhzjWT6I0Gh/p47kEUo0dSkkS3Giiw2wabGRIhO0TPvCrO+54yOQMfwM8
5ydQxSzyUhfm6Xise4/e7//BFV+bnQlkg9peey7eDdeMUC31Ez8TtoqBnqqNudHOK87hSmsTsrMP
CyGOUk42EWwZhDFVkvukRvnJpqLn0e+mOywWa9+wgfy3e6NhpUChTCNcicvVDYwf9WCuztjsyAoG
6A86T76e/CzIhUA3F4Eg9jAZFpdj5Nht/a1Pcxuf0ff+QLDbLdg0zy999A9/EKecXlRBgcOw2T2A
9+keJgrJ02uZGlB9yq8JzI7MY8bo7vqw7+K+FFLZMo2D5Bd2wes1qLnZE7UpfCEJdAG/X7HWc1qd
8dlT3Z/9T8Bg9HxeqJMoisRtUHo7gNIYArGKJm1z/9knI+EXFSIsBISW87VimE3UrxKIuziOY7Vv
wfCbNB1SBlFejqfi6TSiHsDYQhEtHpOtwgmfh04sOuDPYrf/9jztHzE1aNXJX3EKIVmfgINXsP3l
yv3uZ0NXpuveflkA3sFbl6AfHCbA1+B2XdcYNc9T/GbLMZgWMYl4ENR5rT82hXD9k2M+n+SJ+1vp
AMRLZe8RSiSaws9f8+0uqsjXBdqevXcAoXfclyAmzemNeR+Lg+uV3ltrkNjYJdC1TZz0KbouABN9
wy0bs9Ii05xY/fuf6uaQ/VkNeW09LMhCvKkDLE/z2Di54EMKwI52GCaxKp7ykUXN+nsGZOcB9sD7
qlmPyv/E41sQHMB1Ms18/6jFUqn/sDFjyhQnJBerWzHI1iosYoMzRXxnbxmqDL1fG6NL3rWj00nX
6NNrHPt8gURRiy8cfxlPqZllIKo/zj0o8OVabYTTyMUegzml40n92rR2h6wKWdSV84s/g73h7puv
CVCxBDz3TjwNnmgo0FEGTpklnhsONFqMfAI+ZyCneixuhxTLXdjPyOW8qIbLoLGURPgW3K4ElgPI
7FsWMarCBl3gr4cfy1lBoYdLkbHi81TC7TsvOxZP9Qx172Ed8TVHCuKo/EcSuxHRIKg3yWNZB6Mo
eZC3Cz4xnN8LiNwKg/zqiwC67ZvjdhKndwjn5TpldzH0DshF1rmxNRrG63YcCmGDkY52um63j7CP
G2xLCqBIQVwEMxRBqB1nNM4bh+ePdQYsdoK4aLLHGnHrmPzCXAPcsjUxuRBHT8B+DhvrQj0sfC9a
iOJ35yLWdUSQYyZFEecIOfwp0/8fd83nFn/Q8g2kGuWKXdz9bfa3jTa/2v9LU4AvVPfDVFN+KUKp
9CJL0wPJ8l9zS28qFASMMO0NRWxLP5DkIh9tJ4y0/ukbbNb3sw63UDjdl0oojwQkvgTR+Idxf0t1
UsRhM1nnw5c67kRHqcbaVoy5f8dJUYg9mlwPMJXQ9L53Fbg9Lw8ssqpXE2xeSZqTA/xmat8kiqCN
7sY5yFWEd1wrjaGwftwASgAVY8QMutOlxej1uu9Vel/83gtqU4HO2PVOeMmKNo+JqWAOB45FxOTL
lzLzjYSgLCHQPmVtW/mYo2nbf0KJRwPYLWH8cmxBlsyHAuTS6VbVEviNyRbjVDKw2B2qml+AKuXt
zgR7AkOKbYzVu/o0j/5xYp0ylqAdwwU+BPTCXs0K5XzySFjb9LNRCiQlq9pu2ts3ay8FDe0A1Po6
sMWFJbJ5E7f/JgZXEbwM35Jg+bLcz3qplb33IvbdoeyQ5roQOxYYSSW44FmT5/z59koCCu6lJCrC
BgvK7pT6zzUoYTfaNPZNC6KiiQHcym2onQIcsRpol6kdUXPMQaUMJezCtKSO3yVj6twL4n6yvW+v
klsXpjjU5G/7PaBAxwaUQTpNTnYevbmlB3Rg3qoMAfNpQ3h54OwwTsqMQBb3pVaB5qpCJKBIYhbt
4q5VA02nnHntMAmO7HlEwaE7TEcpQAYWibhxqJlvpVeZrtLs3WaInTM1rgxcA5Y3JYdj/vyka/cM
5nzgpoRX/1fCNR91kEmgS4tqiGaL9WmF+8ber/Ok5452oOPOJEU9afsPDWThWg/XrqRsEJ4n8d+0
C8h7y5GKaL8oYrRHztADhCjZQHP9BzGeRe73ZcEmbVYBAUPtS3qh0HxZ+nnPkf1nJe+GzNkBoduW
5uuK7j/YAT3hnKnOsTQ3B3jM6KBLSagGV4ybSWAxVPBeZenvsFi+IBgJD/0Vs8tFDtF+h1SxLtLs
NPWN6ZGmu8MXe2/aQYmEC+y9LnSXyI4DP17sPRU7WZg5rPlMBmwD1N9C94X3VnVIJf9P+0Qi9s/b
9i1uGA3h7IrM5nUZenw/46DeM88/LDU2YcoBlyEHir7wqdTpckBnW7LTXucRybgXYpZ7uJ8xpq3X
KoIpnTOji91BtfuAjpEpk+R/dk+4yTkLCYwnvlrak3T2d9KxQTtOo+S5kNkwDNAFDUzkEO4vecud
eMfrABjbmzmEMAVyOQMn4LZyUw2c8z9W0XclxmcN5sO8l+D80TpWqABbUuiJDSCFwFMFDv9tn0GO
CpjLLcFoGkzH3xJaFHnX2slErKbNaSj2qVvWebj1lI5L2nev8rs44XiRISsAqlmA72bRbv+ExUKc
Kd637PEZIaZBZC6nbbNAiyhQYgYVz7kKkua/Y9AdIguKGfe+lVIxtzVA/7GS7bJrCtjCQB7/c6LO
gWn0aLgO2TK5pqY2ss2I0FWvoJc1AjEUqUkRakxs0r4JnSsLmwgxvBqvIQ9gIRq+obpWFHY2ZTRt
mMc7JeMqzCwkIUBEQE53IFuVJNihcdKCcHaTkrPl4vH2GoJ+Bsb3qmXnv6xoWyHZrg/2NJpSWZP3
8dpfPTupaH17C08zpw2WKpx1TQTHQ42AGOOUlfNEoxDl1RMOVQqStanFoT+NxJYp/mX4xEsIhRBm
w7KwBCr5HwUZdyKrsqUd7UOI9z+rPnCGGL/TCgqZfPAbH1FKTDjgAUhkhRNj5Jakmn6C4oV61UDu
XxyEkxbfzjf6VBKodptZA5xMD13Lrd23QBFQbwnF5YsWZmdpTAZUzdPIkI0uFo16eWuDOC5q49mW
7xFG4GMfMdZ6Q6dmJHanVy2Up29WvRPTu23rSJb1FlK+yF5U/lOsMdBYje339ALLdcfkM3P4u1wQ
hzb61tRFD/Ga3LBVaSzTxlCfpwoVgBGx43U/2rsAbqxh05ZxU8aDa38KfbPfFFnGSAwdGREWEq1Y
l4sylOgfoqNhI0Yjw7d+44MYnuMk8M26SFm+wmz1deqYqs6RsHIVwugsOwB5dJrDBeqnv4rEZ1mf
ZBM9zv5E8qhTg9I/CTm6qL+Dfv9SRRWxzQoSCMRRWcu3VgHcKGmKOMhoCU47RpWjS8gZNuzSAFZe
pie60mQaLOhQhgyVNf7cpVWPY4PSm5Sd9nghr12UuvFqkTIEQtjzMOr46ME+TwL4RwvnpYQGlGdF
N9p6/dYPa4MVlQnfmKwd0bDwdSQ7puOB5t9WHCiiaFf2cT1FYg+SVEVhydTftt5/IB99xonLuCC7
bw3tbpVkZ0WMGyl55nBT96oEt500bUBhNXT0x0D4N/ENyzDPbxP3twV6fJLMCzKhRQOG40GIptmB
6/0Hm3BhSVfKuhV2yqi6Fxjjv/EbDv4AyssgAZ61iOQgPpkIpPaiDa0u74ilPBA7cz0i130U/mgk
1gXZhUZ1nOs1aWfzTz8xTeLaYhNabNrBMhsWnx68qFo6kuTy4xZxC9DPLO6RWeg4CMYDGvpQiK4G
N1/MBRrQUgQEcJfqk8kXJBEj2238z55Lq1kxkSKDNqHN7jtKEmLDgNWSD8UUh9BF+NnsIn/ZgBh3
B15TuYXocg8bZqbTOP2S0Ub85GTxTuhvkLpT/+atMszqeG0p6QLfYcdNMkb0eVSej8PysyGPX4Qc
nSCumUDYwCdz0GM8kA5gBur9SZTY30FDQaTzmE0bH3Gh1upWvnxKGTlDp3YhwF4F4zAUlivYuIfN
d3PQ8Q7d70rzpRusvm3aVqzRiyjE6XkMDQ96nS8efzEVa37WRT4MUn7UZiEJU3v2BfXyFAiUJTia
31fONVUmj8ZPjjXAULDaHiUGIu5ysYOcDRU/6Cyc6IMDu9WnJVQUTq7QHtSIRskUIeI2nDlyTNxE
syhYWnhTpCW3peXE+G+9d8bJ9Sdlkcv3SHDfEEWOvyQYFFogh8XKXU6gSbPXQQUHbHo3z1Y6agO+
41qFJCiS7HzpKiTF3TIDQvv67XGz/xv3x0UXlYI8V/jbtrGyTw/myiYeEkF9P0f/GUWgnN5kJjSe
sJzuI0zgkJiMdsyyH5+wCy1PiMX9GC+i0kTnyhzateKiNZyNiiFawqZwmLFMiMlDU2DEClWrN88y
g4bTNIXxTX5yKcmQzCBam9OHT5Mp5E11z4NGQXLPyq6xMmxiE3iwjPSjjc4KTUO0jp6z2c/gh27E
4/YzlTJJC2G/R+uuFjjjTfmJ2aEbpx1BwkNVkVKUVDWyml0V6qxr+zAlmBUBuCNVX1z2E+QLd51N
pq9rEzbBDFrj0FsvMUDzQLg+UM2U/FVjgO5HxebNNFxpgAWq4UjI3BylOqxpBVaqFDUwn02OEVmS
QNJRSSxIL0K35LsK0CZX0NeNMIIIQQFPQVNErHYUQJL2wytesHlSU2WoBgkdfu0AqVLd/q4l+JQE
gGjRCw+Z+/NhuA+n/fnE4Swp9iTEMQzOq6gZ4pVb+8YZ3RMXNZmv5pgicAJQRZdT3lwS36CnIEav
Qr0aWt69+c5RqPEtCXYpKlzmiV1Q33TjoM+BifYzI6TlE3CvkrgH2p3imlkMo9WXtCpMp4Qcvfnv
5lAnc3755/NaneUsZsmB74RFjekesyIgLNnB+4qnF4gaGzoWzVmIpFwzPcz8XN4J+Ma5NPz5l5b5
k7uaq5G1g1hAbYMgxfybudv01mWkSUAr7t2StEZZso0XIqp0cVozeuNW2Zu3/s6dEhSlY1z2Ho2W
r1WgZZUaVtwHXlwKpGi5yLR4S+xMhnuF46OrrorS93/AcEkT7gBvUs0l9dR/XvjBq3Y6OR3ZG055
g0iuEUjIs1Uuk22GrEZ0kNxJbBVQ4f59mWyBjuoct9zqK7inmW/Ur1osavTkgytOai1SSEYX8Ess
X2QO1ETKNuGzSRWmMXby+G0O/GYZzAouCWJ1qu4GVyKuMIICd8aKMsowWiLHg3nDa4AGXmAjfu2G
5FXwp63VFgTsfmneCt8BYv/vPlA8xEKWcSj5Y9FN3ptiyZ6inQe2llKc82JBokKyR74B2tOXxVfK
lqDU6rCYunlRXIqdR+R+bmz9tstxoMe/Tbg73hE+3NWeumAo8fv4VXar4x5cjnawENPQRQN353MF
K6XljW82yDYSetDDlM3XesdHY31WcHr47+uNFG3pPsZFGc1/xGykEIXVFFGkmjvMDQ9X6ldoo8md
DXxYYxfoJb4J7aR2n84U/E/tOgeUMQcBeXv+8zdw3067jg7vD4qAricdiv4t2Z1f2fgaCE+IPhf3
qK62+LlTJl0klxS5W3Lu8Y6jP+ARkv4692EdVfmAbd8xTKmAgWWwwipt+aXCh3wpRmOyMssMQe6y
mD4buv0wF1/X4NWEijFrRB9aZgUGrxdWH6+u4kFeZx1iyx8aKD3vino0yzZtBlnu0Eh4N2v/hy/1
o9P2NQDPZ7CMrBjMfS32sWzYJjJbRdIIhW2VDfR1Qlr0GflGvyUbi+IvbGco3koZWyShbiGsL16W
yiedGoikSRtRMJ/p8m+kYRgGI/8jKnr9XpoYPU9tf7Fg5Bqi/vuePldPB5Pd4EfXEs8pcaRf69rQ
SwT/VmnQoSv3UMxEUQ2XFfjzEvUjse5HWwb9gSedd4lu/M5wa/xdmxcmD0sroMyKl3HMkBI15G3l
DCeay2agc8LK20XfZnnQHdzxN9zv5KJVDyYHckqceTdmOtvgGJk/A/E7tsSiHcU1zUPhENehTZwp
G++pCdy4HRhlSwFW1M8IUHTL4O1hUdnMxQVNHmQx14JkOa6mFtzqXyEq0OOySoHAcgd6Bwdhyuwk
41KFYOd+sTlJtH7tBUvPvUdKhKwAu3SQFhmTJUWYw1QM5b4vCEJCXjxFs9sqAiDFm3I/0o4szOvr
8qyx5Tl3+N/9Qaw9VHDA44N5wB8whtEurTQ741rkKpShaYS44aTxrCB8UTJ3UW675ZPBpBuSMJq9
N1MEVJ3+HV/FQai1Div4HmKhouRq5J+JTJWseLCadi8ukdebAweHMr4sLBG/t7spBxGtIQC7Dyvf
6CLl8d5TrigLExoJWRMN2Pc3K78fqJW1tbIVDTxycJL+vQ7VvN6Wq7KZshRettCNTPPHlLkrpfVb
Ef0Sa5r0NF2FSguaLjJ87KrEJEcYGnaMdlMoXvwx1KYXyxnHWzHWJrC6daX2NOvyxM5vxsp1tFzd
iCRxFk8RlV5fKiAurXKHS8BiTnPU7W/Q+iNLmNpCanBz8BGmzQp49I6Ir6JYuNbuEwTyNRmtVuYx
j4lsYPzs0FBHVEOyzTdjh5kQtJCkry8YRh7g01SwxhTRAdLaO6UF3bKe2mfAmdtgDeHLSWdQW9AT
PZnNjqLT/UXbyETlk7YStiybfdS0HYGbgXdWgQaaJkdTsBr15jt4QDSo2RTEqar5iUmk3/CHLUU7
wvA7Oo2NwkEjV4glLBHfW3dr2o51bXzhkyvkCfkTgZqmzjJXQ9QUNauPGFop9o0GEfqbFoqOGHDE
F4xwgur9nX0W1tdsQQ4TXrzAPYYHhMkcS1my6ezrMSrBXIvc2Go0O6IlIw4japRZaXgtuREmMNko
PZG2+5+H78GAkH5ZpAD9W8jy6+MW7g/uWYm5mW3/fIaRmHXj8NEn0U0esxr7/Y3/p8IJuuhGN6mg
qS1Od3f96x1Cv9DmszLpSP5n7mAsbBe7MKcIYkQlaRwjZL9ySsaTq2pG2Lx97cXwo4A+aMPqeoIE
f7N/NPkd8IOot6DBHbeqxaBy0036hLBVrUxgovESJTtA1DkgBNFh6stHOHijV2KQgXBH+5z7NVkG
7gMWDYkqxB/jjca8YLVlWvadZoi9WnoWYMw9670nshQGNdMBKotSh8Jshg88q89opxI3wra65wGM
YwYTtAhefxL2w19mWulaynfkRfa+KdybkdWWOIibO2c08+19G3pGSFuY8Ia3yPlgXBvWh+XGpYYa
2xNQGPg9JmAFO1gEkcL6ymK3xtPSYE+AoS0EZXvY7mvfw+RlJ5mP9bsDoTh36RnUqB1qIWSBg2AU
t7rP7ryqQPnoTroTZyrc0wtFpWZLC8BQXDk4QbGOt7eH7GluH1A7jrmZvAHA8L4aaGom9iAVE8jI
NQiq0/5ImMedLIrJBixcnNbMyo7AXCMRY2XVlPqsPwcS6+e+jO/OxLjbJbuRjq5KxbpmANGYkKGZ
5Fc8YNAaUArhu6p7A/VARkzeVDm5tFKwkBL159Ey6L3aB3XvBolfQyjfU+1JH2DUtXqnfxp5q2AV
XJtLd80Ueber1qMpPezVJ7iUWYFv6gYPxBo7wYjeGMDh/nN/DVMwNW5GUZk6xJO35zJs89VFCti9
2EeU8zIN/rcqN32UFlD1jOTNwmjI4YD0f1NFoE1zy8/A06rN1dqLzacD0UsilJMHnhDUPLChjRK3
go8jFDP321/0umvDvuYuakY89TSV
`protect end_protected
