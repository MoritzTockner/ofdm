-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
RnORNWei7IRd0Nq15a5BPJvhId1MZj7wE1Ah/ooO8OXEnVgEDiHZEVNsH2EkH/g7dhBLb74N+/pX
ZAoBWR09KHgI3y6HtNW31Eo27RDRYRkZoitKIYutSWxGZfV4WrZ+GL3rD2fiCKOI2aO1cFBib7+Q
/MSrn9Td5h/tVBT/qj3vBlymAIBTWxhXh830ThXoxa/4cbFz1wAu5bSuOzQdH8wGfVLxSQ9pl1qQ
nU8wW+YTy6EiSSC1/R+nMaXfqUV/jVATWeTAqLjFo1HSHg8vbXkNsa/HbJfYnZ04wMV2KwOEVXQy
sqlfsGGc9EOVd2Z/3q0GkwFwzvreUjLrGavdAw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
VbsZiGTji6n/jlwBVJee/cTiODWCV/f/vKASxpAIPkg1+AR1+n5e7CIOLu6bv0YyUyo7SZeHNLzQ
lARef4bVxCCjiy/58PzIJ3WiAD7P4yjqewbei0rz1i7CjTMAtUqhfvTi/D5/4w00VLxnBskPmNkE
jnQyZlJ7X0Cqpm1u4W0w/KyDO8f5Mj+7JlZJo4Qw8yv0D1K2b7z99w7xQIPgdVuLC2EDjqMw9Pp6
sH9uEuVfFBtYWJC7p+DxWAgHM988+DUzPALP4KKj6PIPbQf4ryGpYeJ70IOAP+bTOwWCEKgwmTfv
dWL1qeZi/FFjlFsuXoSMR4tw9+eMLtETGDiAwHPk9QYqAvXHF3P5TaubIA1JtWVaYXlhlGaKwWPH
w3KOK4yeHAD21vs8R8+sXBvhnUp5Y25cU1OEg9++ne56MQWDJ8YJ08h1co/gk6vc9OlRrgEXtStg
sWKbhjGEpsiVMTGe3bUpBuryo+ID+rTthGusNCaSYMa6xSI3I++xkVe6Unw2wn33iR0rC/1pQ/99
gHtTIo1/COCdOQmwYl+S+KJ51C5FUpC+fze6Sci+6svlV/lbIR0pJGaFm4Pe4nCRo64ugYBNH9EP
rfqjRaPs5p/f6k9AdMFTk0xzNC5q9gGnO0LjQ9n5INse3SkfvIPG0w5811Uxpio3XBAnKHz32+gX
Zif5ykZq7JHnEnR2NlKSYTd4ckIcvFQIVf/Ojbr4EbsDJyzM5IebNupYm/P2vHVPM4g0POGE5nRf
yB9cn24RCQS9IB/oWaUYTkmnEjO2Po9pHXmVPfnCKqZA2HTIEFf4YRKuZwIXJG+Ip3869+hkgCvD
N7Li0Q2vlwt8wEEQuqQKB2SCdpyqaK4RB9+rB+L1stOS+5zEAQ5f/TLa4Qo6qXXNeXziKuXj9wEj
tde2pDlHneXlnlLwXmZLRFSdhwVS0D8MgEpX1xjqgh+Y5miFgDSZfv1PjFzCMnzVFJzWf16o90Q3
om3RSzHVFBDRKPbw6HupFd305tjAr0OjvoHQP+RwLIcu6XVmJPB2QGGWcVLRp6VguFo0cm7k7wWa
q2tAjSQw8gk3mGkTwDXj2Ak5sRYkAcgjV/tyUSGsMSAUoDI/obecHmlmXPhdC91e2KtUvEex3vhJ
evIqp8Vn/IGEnYeRlgsySq9dINohg1nj0/Byj/izZi1/RAn8yGniQ0qDsMRHTg/ygpUsf09maK5e
udNMP8fN0oEhpipqO2Riwbv+NIpD5wtEBQ2Bj3rN7NE1ANMnyAtfh8QW73zNduLZjZ/j+ovnTilY
MVzagFpUkcAFYRnzFoAhB4e4mMeSVhNuLz7Kz6d97j+XJoYY/GUeUz9yREGFDDeRF5M99l/uDpZL
PlxMxYkEEFKXtqgRDryx/+ebbL0HHxK4jCeFnHRScC5Fm+S06CPFjG5ufNFsL8YuPr/6a5bstywz
3OyLvqU/+wAhXKEor8fNgAGp6oxhcQe3FoxYuz5Z/JeJ7T3EcJLb02bZn1dXsyruIokI5SC0Nj+6
ZxqLFpXaHozbDtkZIC5rMh6HnyyC+aqPwRrQbLCXsseJf4TDzLcX8Jg1yl7a/gwziBf+6qxQc2k4
IR/3Js5HrjHKQwct7iK/FhoBsN4MxZ4PcMHVaB9U7jUXzVAWFVFh8MCLKOwsIrCiRh5uqDfduAG1
ZDCm/t6i9omOW9piXnBhRo1UHWfOfXf++1kthin7zS98gXqD754SkNWfHaOygjvoiBgSttG+ytUV
ZcauPgoR8lYPaW9HuI3VeiuRBkBHr1Nn4qqIP+gmYRJz8b8pfeQy9xGEGMmoTVpzGu3+cXShhfs4
9zlhUvDjlN/+UmyCdhV4LrWYIV0SqhyAnLS4uGHoTqz5MGrxyeir/E6Rt4BF/g3T9yD9UZOVbWUk
+wDo2ZnZeMNeQ6sqe+2mE0ms+KCZDip2tDG5MYodtsiHN1VifXk/PIYPaiKPjWp3y5gZlto2CoTp
mseYA65PbUsu293lxVvlTjbyy2UZcMz3YZptQR+hNFLbCRoNJqTt7bozzdNKQF2/7wcRmD+4vXVF
SFLUMth5D77S40ZOddXHn3r1L7b+Kasl18TAD1+qNx4gBUdyQevNIJa+u9fEUZqsEnXuux8dHzsp
zjShzvGiGUx0jcXIs7xOIhs5wPPDToBhmfS+OsJ1yeb82Yo67LWXlYyEvMAVVXp5av3siWoYP38u
/s7mgQWjH3djjvtGWRessd4o8adsO7+YrE6l9bqmR04GU+9JJKb6c/2++MPVaPIJ+9xv+mGvvXyU
Ud/AAgEFtn+XrYmCG4UlJQiPMqKkqNpEX9ch0hbRDt/joQkidnvCXwULxkzNY3nedBiQRjohmyph
q31Dw4SEwV3ULP1it63LJgSHp3OXMkcT3dEq49qaS0kr8yerCQhJgVYrDzgpbjy+u/G+orAvpA+Z
EDOL+VG09wlBGIjb/1/zTJIHPmjUCQenJ6bZcyBHlk/y5k8Rp3UK/VU3ZkHcMY5bjzpyjZ+Mige0
zhtTYWSLJ2eW8UdkB3tiBbACVepLsGMlj9X9zWYydkb+sxecL5LIC4zz0sSWhJFYw59+lGDswMOA
2cYT3Q6JfzZ26Bi2ncWFwR8qqS5bs6x0Hnax1wTUh//ZWACIIMAbQYFwEV140WBk3eG52THhYBwr
88fPspoUuyOK/Rl5gE+SmoUrTJGUJMhIfCuBww83LQezeiA2DfavmzpWQaJpniup3dNLY+iWD25A
mB8vsiNa+ook8v7HVqp295XJIPCHZU0h4C20Z8WESwHWkrDEucl1/f7ziGbGRWGa2ewUNnEbT0Xp
EBhUaiS0I233ZGAU9exFYy05fTK+OgYMPQcg8BIDxFFwm301XIXovhxGygdUAPymuGZvrXkc1typ
Ksv0+DKUvfEuME1L6sRsmbHmf8oGiubc7Zw5bc4QTsLdDCUdqcka/876M5raULZzBA7e43rPU6xQ
y4LReJm6+Asc7I17sOWJRNPyw10Wh1Ri6C4+tgQNZ3Y/+COXO5hiq2FjVARVCbAL3cLSN8iFsclQ
NJqmwbAX8JQ5HaZDjhptCI6kggQeCg3G4Rllymc1t54BLqREelcfEp8EwGJ3rRMnVqsbmXtmB0cY
CP/if5capPgNLFp3LCF2d+P8HHmwAQcRQKqRMKCIk3IWjnULASENDlmKFiClS//bard03hDyDYHM
Bhtc0nHH1mwlv+3QKYcQ0ajk9VMxUoUudiCh3Xp3uA8N+qMsrJXmrOhWAs32rqKGmfGIbnCEJgPa
c+KzoMzZdm6v53rOMNpy+MJSedEzbX6Vbvv5XhPT3T9AoTKV/hjZ7cf5WBzgPUKQTpnxvAwrKGf8
ticgh2YXO1L66h+H8MOURVc8+UBQS78XCJgvFx4094P5OHVH0VmEe1MISEnwdi64Z2bCr6CjhCqf
ux8DB99f/h/PsQpGcOm5SGMmCJH8Ij0meUuSm10R4t0pLBHNhnvwqqVy74dRm+qDor/MKwYL4PgA
OVa1uCrmObwUWImzVl3AWYHFSQdU10aducn0crDxcMC6CFLhXobenYJ4scrt0DWx4Amu880jQ+qT
34f+apl+lv7HtbFBSU7A+L0QWqqOCKZPxSxz+sGUGIkz4oqtSogOalOIyyVV0M+xm1q/Ng2+C7oW
0hOUtErY80nwEA1eRp7dSat6BqL5xnWQBzx0p9+5lbgdzv0kobLvE2nAIoD0IsQo79ls8LoJGAtj
IlUKJdMCYBQ/oRsL4qB2Q29UJ28/B3x4m9EI196749jZRqlA0ka5MsLcL0uUMEquiwIdu9WocmiW
sjbuUWU5HsB/4Ulx7JT/CwXax+DUVT01QJKEzRA/UGUWXSq96BhhNUnae1rsfryX0O+kGAGjTOtB
UzCMOEZimlBWF28GSgCkBjHSoJ8nNpRFqJ8xRyMXCvadhE9Cx81SJwCvIMW2U7FGz0GwRgqIrz0o
8mywtJBs89gprn26a6mIgXu8TL9e6St97yw7BInNsDtVHNw8fC7HSUnX39jN2y/fpHhtP4Cg2WSj
TB7/qvMK2zz20TjqjXFuf17L+IpdQD4FKfhQpIh4UiLkngVUfGBUAiSMUEA71KBS0V4+/VSJ6Gv0
TSadzinschJF6Q3ymJdt8rFncVw+jypgw3mB92++4b04cfV1SqoD6wU1HXLkU9qCEH5GNfxj5z8u
GNKAoyl21v9N1KevlqSEMcotEnFdHNqNn0lStYaAoxmq3Fv8q6R6v0x8d/ou+O1e7laIqReTbKuz
nRONh1kFpf3y7psEsGquP9VZfa3ZL3CK+MgzEbfvt6B2Vpnv9kywMJ9cJY+mnBWGMF/Xf1eacHWi
+Vpwf5x1Oa696YBKbkiSi3vjdS1eLVL17pulEjKOhTfzS/Qo+WBAIEhtBLuNIoVGSqltvpcn/qfu
aY0UliyA+M+49NtKXfFczpzEVzufryp5yD/1qjuCRZRx+WOYzi6hW80UQ+pRHJ2qfJ7rHtsBYTeH
lBmGyI9kb113ScoCnN6qnyM4MjUXuQtmnixoGDq7qGqs41hpj4yzZTiz12cnlhkFKfC8BtyanpQa
PqGQzqweOL97Vo5+Sa7dwpznGbNTUcJs3G8w8G5z6xK5mxcJL8684ISzSMaDXJbVQ+ylS0roc30+
9pZCh+JKxaaiZpblEpZk4HknhRMI9v4ekjuftNBOtxFEP6kfsxW6v9jM7wEQPuqNMfLd7Br/jha/
QS/6Zy/Kz/1St5ISTIqUjJWCTn320GDdljB5ZD19tn085vVJKlaCQxq3JQQTBeQVa4MqDLqH1/kc
RBZy+bsMtc4DZQ7JfuwEMm1g5am92NVa/vJ2IGBkVZev6Tq0LwveKAdAdhooJNO+bXo1ivj3sazG
36heQ+bxO0ezILwBWE2AvZKb/nVvmS5qQpmjtLR9bnAhywwPQtxx+rJA01dSSpvNkXwCJM3ELPuV
YDL+IsxAP4e7ovykvPjSiQI+PirqyIreDaWFkN/TTrhxQL1MK/TDeZI8hjEGNVsZyB8C3lfVr2Km
5XLAIOKVObFVvImBNjTHJiHwhY1EjLqdYr24Mx0Yk1sEHt0a1DT3YK6V1Wb4BloL84eBhSKIcCHk
40zvjnySYbNh+h9YRkZe3zF60TiH+gckySzFflwXV0OxdNicgllW+bGPtHRH6/1yt9WcdyABC4vb
rJCJdPJv2p4ATPv1YT5bU0qOYC0s4InDR7dE3Y92FAgOPnuCr6Mdz9ZxQcd4FRSvs/l6hB3M23tw
1YXlxnAVNKSZgDYHqvqYAIanCHhoP0MYFpMvpNEaDNXSH1w60k5jtGKQhN299T4DMy5qCeRcgejM
sUXf8uGDlzfcwtIeC9N/fKrf2G73GqLabbjQxAfMO2/eCdcAbQ//jH1J+nhiP90Sb5yt/OuOTr0I
yHye2PISv4bphPmk0Oihmd36/OaM1XL/Sd/npIHgeQ9NsQXL3FG9hVOQWlbvPjNOfa5hDG4Oyp90
gBoUjvBo3z/bwanvmsR/+bNYXdLy3ywYD8VFx2xGGhDUu7fxHZMLJ6pgkiTtquED+NQk769W4KxI
FDK1fjUo4WeuVRhntlhrZ5WrTtz7+xMPNj4Z4cm5PmmH/C9MrsSrec02v/3aeYZlXlo6Y2noUU+P
cs2o0J2+Ohb5duSP5TVtJJk/YdUfC5RcClJ1HOBJjvr6UAGV8iPlNp3wmGYkWLb5CLw1DC0UP1pv
rlWcyYw3XHWvMXK+5p3zq4N2YHOUNOfXDac7ofbp/vZwOAC2dRNTk/fB0tMtq/aCMVFtEq2JwkyO
b+TwnDdND15y46NE1wWuMO0sAZEs/7TH5nNRoMx82cSikgLmNlv/1KfT2SbbT6z/IzfJMjD52pr0
q+ZoH9OQznq15mCRocp5uQidqShkAUAdMrtzC1CHPkeURZwu4uBo1PnZ5oWaVTNGFJ2HVtS+wckf
i2LNhr9C4bDxS0cqNCIHwRHI450tgo+bDgZ+jIAGT/AxkD1V3zuj3Q95NmibDpPMNMkdKLsqTObl
KZGa/5mbmmLKE7UkjHVfYLGRrzR+fy4i0s9XPygu6CuOJ//woZg+Qk3XTmB0ZwJSmzYs8r9M9UQ9
/k3E8Wpy9mi0c7xt+QYvDMpgC8k+FzDMWi/q41gifqgTP2FLx51rGoqxqkFhX9TZiD/9T0eFKLTT
aaw7P41xESlbDStzz9IH7mgCnvQdnHWhzQMyCAvzf2DRGNRkPGF/7PIejfaOVO4PbBk9dDf+LcFf
af6pLF+7MRF/9va2PoC74iktRnlZ9it7ihbYYaj9ehK9JACaacJpIrZuOOYIEHqMkeDtufKF8pWB
OHAqUfdR7PkBsVL6ykQcVQz0wCszSNd34zvPKGCz3BAr9HePMPGy2DaI4ILplOnS7p6IEGIKV0Hj
7cGiXCbH6A3aIH3hVSV90huAFzNnbhADvsICRN3yG+6wvmN4npfoqKF18dGImn+iVJ2hLno82ibd
EcXKNWzwwpFq6q6WWcPfjwVuyKRBdwDfV6dkFGhocy+Bui7+Cn2kMTKWXHD4M3lcXxtNwpYFQLuA
SGnSz58YUX9955YlUPcCvTbgcSVNzQRG5uUAnByPtQJBhYdEkhZ3Qvel9GqpljvhnPNPQyVXAKvG
/ZqFjGXh3wjHC7bcsMNG9HPrDBYXjrSF+VoMTCktJkVQ3nq2oG+sCrib6+4RoOJUR+irVSVQ4kIa
uQ3amY3tvAdNGdrVY9Q2DzJJp+XmOZOg6umlC5rE84aj4efkY/0ipItzPLEIUVrqKNPb+Q1XDv4Y
w9GIee1pS4Hgi+VW+2yiDFJ2+iCgbFbkeS5AX5YGbq67pA2mfiXlXKBBgC/i7t1I8nZ7lOzoMJ6z
p1y0jT581T5+xSlMXLWbnjg7lPr9A91yeaZM+VnrdgeFSJudGJDBv3qq5O1hzGJecZrLPIdyb8P0
U6UIcUGcmr3xExs2qxfcW/EA2ZBS1o0Km6R+2PRtYhfmn7wPOjvOQW4jldJmsl+pTXoi6tKgRFm8
VG+YJS6gMs5Q8U4xzNMzdO5V9uLngQyRFk1Pmw5P/9mMbSdFDYJiIFj8Jy+s+q2jLnJ34S6RBXmN
/mpeKOLeUD8JrcgBwZhXIdgLVN34/qbEsQQesyecZDVEVILqNJHB3PXRkBfMAx5mcuQbKPkVrnIg
+7lwQ7SSEjrNh4q1pV5YHfebxABI/clzuHwW8d8DyocjD5509QYTFQoHQKWBOnEDoVO5whhT9Rg6
NXzjJJ1oscJy+VImdM1kvhv7bYA82GoZaKHjoxGr+BOsdkHEdFWTZORVdo28+OxLrP1vXS7q2ht/
GxgIubyItmE73tUYnJcgW8yZmnj989dTqVzIdENuD7W/m8FLpkoA8rHYRenbSHpkSzvwWP3OG2nk
LZE79Ecv5wSPEJMtC0gH2/1+2g195o0KpfwGz7zIxQIOmswe3R0rMNCBz4AKLfmsUac/QZu0Silc
CJEr+3T1406HhzfDpKs3n1kI41UEvJw28D+lVK4RT3AJpSb58IFt35aUGV/9dGD0gvU8yGs94SQv
K+4odYW3N/fijuE8x1PF17wdyPof7Rroy2mu6hbAbdXPofl5W2qCsQjjRG5zToNY23UB4JZSZeHW
37JL8cqHCRsk0mSWglIgwgQWaqvBuvxYa0GECrk9vHGnL6xAyUvJjLjC7itwmFf4llWABcQtA7An
HZ9Gp5jQqbN8bBbNe/ee+mjcsDIVnXnNqs/CmlAZX+5sPkgKbeQnzj9phrWiXZFqa5KGVzHUj2c5
1WHeCAKZZxNjz7WyarR3AWXgcwkQwYk5lanMwpqVoyKatzrZglfvTk8I4jXSEUH4SzmFUnwyWqg8
xE+0ReYO4ZyPBiExnm1K6luGXWad52npBEEnJBZxD9Mqx7k7XldQQGVp1Z44A9IJaY6mMs6Xb1vO
VIRt+5bjPqYEQ12n3EPBcV+5SZzE/FmS5BYmDyS69kX4g50FeqjRWL2S0s8gSdZLWPSt9kTCeV0y
ph3QZWTEgS7wG+3wueBASPwbzTbG/hhe1W8jwDTi6cFnx0srx/DfmcM1qxh+gBBJfaZYvhg5WE/6
Hxa4Bnd5aaVWyh3wmq3+fdCqA4mTLES4EoLDdeYxzvu5vnJktG+0iSG1i0Ll9wONYptDwWq/tZhu
jCM5K6dd/eh9S/ROobwEFTBLk6JEyiwUDPSphKkAwp8sSCjhD6/01mDfdoz0pBN9UpVJChV+PYrb
teR6jOLSycJ0weu/iwKj61XofDQPdtjyl6uJeL3kA9SyGoo1fg4qTl3Vf7r3nbPsaG4KYEFS1F0x
BkkNtVc+Vp7eZpaG1LMWvgUIHuWABAhpM8IR9AxXneAqMv/sx+j5wZr/98GwHf/x0firgft6knNc
qTO16vtEBJsjlTo/ajrt6CwouFu0J3yydmJbXpCLs6s7PFg03vlbAVkIW9VrDlSDVjg/X1VD8ciR
pERnn3HSqEwm4rcN2XmcGONio4nipq2qQ5sKK6qeLGORyNQUEUh2YoLelw+84WDV5mB4eSB4+Kma
oErWZIGpBv5aQLw6szAhlMNpD0m44oAvQk4q8ahFkNYRSlp9tEftGUw/3HeQ5kee0NvDelCzJB+3
Bse1GSR2HDelZ0tboMrGUsEbMY9l1z81XugY8QDdHRm0Z3uVoqotucW89WsVSjMPJLosNuh80aIz
znLCshyd9UBRmXL4GWjgYW1UKy2eH0h08Ehn2AD8YVEHchiUDwOcBYbeCNlQAff4/w+f5wP5PhQU
wMqSdfwEfJU8HIBHQdFPw9B2PEeWjUJ3v9KIDF8f3IY0TnP1eIw5r7N2Q7ZJ6QqAferDZZDgBgmQ
QoGal+YslKrb3l8Q6qsfB31RklIYpOaGjEOsubWP9mxpsS/GlRO6aKZ14j6JlUhe5i0h5UdiNDwi
CqzK66Cb4UmINS0KAkXomeN0DkqXZAugfP0LM6WALiPwSR8mzoCVMkXDPWmpL9ke/+QeogtpHNJG
RQgCQ0K/mDO0z1h8Wd6gH4LyJVSEWuFXXTPLY0DdUVS8in+8T1xSe8FYAC4UIAOnctHJYGmbIPwg
jj+yt/dHj91/56tQkhg9v4/fIE+WWLWSZkDrLHu+2L0Y1C0wrfOLi+5c9oBS0DL90IFPR3kuWUpB
+xpplamEJcVsqPhVcBpoNvHOtWzoWQiD6hCDXwsICImO8Gfml8KJGP5R/sXDY8RsunCJYFGigeTG
wHmM03oMptJqL5t5eM5Vutu6xE0456w56ggNsT5Jt458QCcmSucKT/TJ9udj9EZ4yEEDyhKUItFZ
umOD+USxrkQ3v0lAVJfl0O0pwvds/rwPssLvb+ttYbF+UA40uyB7H7TpZFrjjVMglnkwWmLUlKJI
tr6ytQbgUWuwOB+Snlhl921y3uweHXdnyQ6HvUzYMwYpWFW0vmn7MDUHJENUOmwu7LG0j+Pqbsnv
UNW+NRR/dvJQLk4cUoQ3LmbbmT9xAAfXl01mHHgmvvt80x7QYnZYUVIbxAWLVymBTGulvt50Z0wh
I7JkQqSLPrFI3SX9OB+bXs5dzlA9911larcwHC0k2SfHnwFF6uzBFbKqy2wyhE4DZmevEu+l4ENN
kry/UzIqx4qlgM4R+JTOn6zdpPAgkJk4nVVoOlja9ClaP/HlWo+Zlfbt9K9PoWBHTSXK8tU31x/r
TdQeFIi5tVAOLpdvka9sUEJEa0leiJ7dh7dW3xFPEhsB+/9pJDWvT/wR7UrYh6o4kWC71Y9mjdqk
tQ4BX5RAcwWQ3co4xIqaP+ZrFMFZk/2Z20MsYES9hzk+mBxSIEiQYpy2mvp+OyFI3s9KYXn6+6vF
MtiV85Sjgz8z+krCpFaQsUh/O7ZRSWsalgxQE7HydZdC0hOJD4fAEO1oxQtnCMynE4YWXKWxrCS7
Guh1AZx0pDT4gypfQzHoIbyzOFQCH5ZsTx2tQQVy7ZyWfxWSaCcPrmFM0ulyemfLPuR6V334Qkc6
L5PGi0ApJ1d2MBM4G4MrrGngf7yI7uoL1DyO53en7KxdjvRIYTOpP1YW41oTEHriAgRZXMiXGkTo
wAMui0kmfPunbK5rBUOc1F5nKIVrkDQWwnP69kZrEgEnFVg+Hkk8jsVEYlLVBYQad86Bc1WCP81f
z52HqhYvpl0ubGtVetmdlNVMb6XcEJ0j6pQ5bdZ6B/xXAyzSZ/L3wJrxdI6JqvsWOE1Xr2SmU3K7
SCcu5R1VnC4UJ2ntXtsHYXoFLHi9nfcFGcrz60yPMH6khzJGxPBK8lrPMr/LB+qfcIteCamDAYPe
tMWgxO5WKtW1J/aFVeeWN4YesvzfX0MJ6Zf1SO3cMJYiNOBjukewga5PU8HMnS4jPJ3MKy0NGoak
qhgxv4t2XxYvDOZL0Om2fRRmi2FjVje7ZXKYV4qDb8UNAyHLwugMj4sVYGVvco7PemWoLjxnuM/q
bY28lkmxiNQ008AJSTcNiUjYSom1KfTtinHArwyY2vmnsZMEcK4ukbosK/lQi/25VL6L+kpmszXF
GSCeSSN2d9swgsWozuNBZ1N1NlLopUK2lHeQG6iEwbN2x7m2YW9XHEOuLyRgL1mQ4+JtKtYipokS
9dXf7nUF5kmjtJoTFf5dvr6iy2NZZcPZZBizsWhIk67wBnT1Eyz+jalns6vF52hL4ufmfx0exS1j
LbTO93iUzxWfRz3I29fEEr1rmRVOuSJTgvfh7orDo1ez6v6PqhnOaBQKtTj0S8fnlgxkE2UD5/91
EFR/ltKdK7aJTTd4lQPEKRb0oaJDN+C5qMuVjE3550UxuUTUYK1Utv0R8cXSQ+z+JiP9iCGDBx1w
WUQbOCV/3W7auTpma7rYKedFvFXhLiu3pZa6ME2HkHXSkTinpRf/FMK/lJZcbNCLzJtw+/8Kd4ds
W8FcAk4JpR8Iz2yOdPLjLjrk1kNFS/n1jbbIN3Ds/MbZUevatuZqfpZuZkvfa43XpXiFVlyPA1RJ
A9+x4xPaaNwuOECalDuiTqB7FnVlvdJOBfE7jM2ykLI+Vl9M5FpmcvzMFyR0jpgVvdBhps0nuPxx
F9rT3FUqAL9K/BU5/JMWmaql8UmN+U9jTjmX3iu59/0l1NxEM/bmJONxKN4gSlE9ZwfcPYt+JS/J
4giffHjx5XmfwAhWjfaHPGNL0qxaTuXJhiC2KJn8PK6p/ke+I/VG5Zr+Vb0D4yeUrmkoyeBA/7vT
MHmFRTsjbh2nAEE9vIB3ohGNI+oFPUpLPKqxo36kbKHmFPeH9BvKe+rKQ89Zou6H4hhq7rqRPrPz
U/ADBDwKlO4TrRpRT1JKIGbCXEFE57xPGjJHcQTbN1kVO1TXscTanK8g8twYuKPb+4E0O1ytOv4B
6HDPhxFDBpje+OA2AiqKpA6J8PzOpxFr96PYGAjXCJAz4Ert+FOJWs3lOClCA/NGP0m4yew0BBUW
116m/aAwoN6ldKlarPMz0TEs3RtpYfzUykpr43JSaNwjXiv3iaiB3O0K+5O2LYBr+lwMb3zxc3GH
J2bEzMPPAhsx+2LkBnMAK23zd5btPg4aU4u4YY4GA8Noi3jKftr/RjpsdO2BZaCZiiIa+TfQSYyq
s/qdxndwvrZJj1pBqq56zVZwpvyP4Z+ugrLEXm4iJ1SBaQpsp8p6fVpOszxwUQc+xy4uyy5g+BJd
XOxJdxZnIm0dJvQvnlCrJfLO+RSHHiEwpuFnNWZcTjPgmEThV1E1Xn+hgRrP83AO3Jw4atqDbb0T
NIYse+2aijTbHFjLo26qKKafJ3pymgf/oV5A5RjRLn1EjZ11zy0HjQkbnKMGQ2SKUfQppt6Ym3bD
1h5aJOtEe6FloKReO9eNsil8WGMF3h/7dHEwB1Z5FXu77wCG3kVKTBUvRYigxv1XT6wGyVGv1+fA
pEtvGScSV47zyK82tGGVgxFE6Azv+SLljtbBQFYQkexKHbxZLmmz15spl5SDnZIHUOsrVFYrMtNE
2MxCHcfHMnMitMTWhy2MaANpKT6i7pVxmnJ6N/YPnMYylwCO3FI7utcX2lDQ6M75n5XIKBMwjmlu
TfpQpcZzoOCAptCwqb2mqxBWEFC5li3NGXN2sl4vfRMo2DS5xSizVCpRJv+9dN0/wiMk+t78+/qi
qltrW2XyL5gDBl7Z0x2d4d57MZJQLraWmYNG7iVKxjfj9T54FY/KtKv8vY3Yaq7WroiHMmq0TjOd
+Ikx4LzaGAKOOUSd5codvcD04kaFIGNXYdBc+isln1TlbJeLH24DbkwDykmRrID6znGvct4ffY07
ENBWYVrRuVjIVVaH3+IZZVP/VY84cXu2xgkLEaYqP71mXKhS8ZdgNU9OmGvZiigsp80kUDHpyqUR
0jxDiDclbTQWoVwIiV6zEp9tI0azpKvmGuGyL9y6N9n53yycVgai7y7BFePc9KK0Fhs7RkLJvuBO
i0TAv2F0pca2NFCQIYAMER9AbZ7J+xNUoZI/86DFJXCDH5R3oPa5O7bSpXIPeCO921q+Prula18K
AJ+v1zhsYxkyaykkN+rn0s39PYZwTj0/067IW2joS1eN9sWEnrFF9JANAFDHZgkF7B4Zn0qxFbFP
dxv9/Yy5EkIGkpli9UQfCnoEn8hw+du0tNi7Sc4vzDWpUdSPYa6DnGcXCHYUCb/vT2w74WcnJY3B
gb5sAzy7DUrsKJo+FzAARalxeufCJq8XdWjBWBMvB+kYTh1PegyCImgmLzIETIWP3+3WFYugKgDM
Xyaug7WJEaEY+N1AUN08/S/v298RHQGBfwYtUdzZ0EI6E90VraQBgphKTSZwPjU1JSk9HO6hfaRz
TLs9flwa2rK9o/zS0d9wFC/mZIMan+ATtevG+NSdvvX71ppjMYH7nZYe7MQjcrmfEAi7XAKZU+NC
h3IaZP1PabfOw+ythAQbULZSRXm7s99YWCQAgK+OwTwgcUB40z1SedNNq0ehmtgzBzzJ7lVxDkac
ItDKSGzZ3oYE+GvIJNNiN9jMPvxUzyqAvd07YOntq6lKJ0yh0lV04f/yuPeK0BUk4syUYdGFT0X3
sLipFxY+mvLFtuQ42cTfWc7sodOShvuKqO//PM/9nKwGMWnHskk/n3L/OFFnRaHom2h9ObLq8pLb
BQ4obCA4WWcStcTTTcT6p89IwpjGRKuUEbyqFzbGrJOOMtYuf3koPK/ZLqXrumFLR4LCor7tdFMW
RGp+R85+aU2OvDNn8sygu0xoyM4pIBkgowCWCcb70eksfgAZhDOA1N9mFcIdHxaghURnPzrUOwAb
E/s=
`protect end_protected
