-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
si37f8gY7vKsNBw0fdz6qKuQr0yClUiFR1lfRQb6xAlHA58gmn12VyjT0OzYpi4imJecZiMJprI6
SeEg8iSkFJNrCanG2iVuOuSj/6nVO6BgRTzCtF8eef14jl39HAAjcYuNtA9Z+/HFBGrgv5rspcWr
9JCw0nFkEoCXX0YvFe+G4BMGrvGTd+3G5Q7jx9J+3b5dIJF6NP0g+0Hpq3JVPsDkj68ooJ1ysnBP
sW0CG027uW1I6tks057LTEWTFTG1rGpuWHfbrPIDdOln0zsXRuH9/29x2pwvAyvokPkeQx+BOffy
ABdM8vjigST4u26OHMfpT3Sd9iNVmSTOIO7xvg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
QyqzA7ziDSCue844d7RAW+esQ+G/hfw0eIhD6+7IAjT/CSUirAkVVk23cm0AOI3dTnjvdhd8PQD+
etgotP5gTxGfxy2YWCna18u8zIwvGs5C++Z6tkjRnhnR64ErWDAD68xX5bYFt/vD6jGC03Opeopz
dyiafYhdGE3ayWJ/xszYFsUd+bRmzQD1ZgpDTbtl8Ilqg0Mf/cyvElIxyUCuvimgmbyhsynzIMh9
QMxmP0i6W9vYwDhi57q057rLwjefBL/uTnMQfSQsSWS1QVh9ttXCOr3V6d+MKj0NU/3TwD8wVv7+
5Hz4lIXN8jBaw5i5cqA+qumcmzF29qtx+hwCOkvF+iMA6slVLHciOtp7zk40iEBOVTMpA544LiGD
ixmbkMQesVGDwrxGuocrsVeBBOd4FtxOPGbZJd0G8Q7EvbF6J29HWwp12SmeA9MhnjsA6BmwPdhe
+Vd3AV70ez0Y7nSbPBelnHF11DeTWu4yOtodNABFrG8xddmkkDORxtpE4RldyMY0UKvMI06cuQ4O
36FuhZy7YA1QImJSzxphHkpQGOp5Nr9nkAiIjFIeEsTeRnXnDUvTKlAHFP86E1nw/d6+YItG+loo
dSZdVwj+yxvbeoto65bYTxlXsVkY7m7aH8/JTi5BhZ/8w8ZSjxlhRKE7Hmbq7u7Id9SiThe8pSes
vA1lgl3ghB8xqGNdwdLMhPZuJKM0WGMOBPg07UG20tAuzS/oLk1IP24b0FbEGS6HKePZINFvpz2T
tTjyFwCao+IlCMur2l39FCY6MxTRm72nT1fTxR9DyOaMhkfu0zprwGk0p7DvkzZwzCITq8REA7y6
NiUW6bh/2636iKOjiPhXwCK1Ywf3oXIg5KIwO2EVPDJdgC/E6C0qt9cbEMTdbQMi/oN7fXsgavzr
2gl4tFNe/joLVqa4douSmAgT+fQlN+eqEZ4ZwqKP1HRvBJyAbYS2ugT7SIA8QORIBBDjWcB36+mI
nlaCe4XsNJvDkqxuVvF/e8OITudGrXR08IT+gFdzynlPrCNUCdVsgJAjVBwtRHtA4H3N3rRvDCkJ
CjPovX5zjB+0FKo+6naI0J+QkZ9HGcwWT3Yvk5jPkAh/b1kyppnvkRrFMMTJ378E+FTb9xMR0fCZ
h9tqW98oiRGkqXkNfQLV1eYlqnePFA5pVyY6hFMyoJylxG0DSrUHJDPehzau2WgHYY7q97q9jjIo
XA9FMjiK1JwjkrhlSyR7qZPWnksnMSI9Emy4D/lfJrzDFfoKo2FT5MjLwjoVKo1aNsPznVceNwAH
bkE5pTnximDMxYaHjFPFUKOB0hKGcas6D12jJIxd8rqVMij0xWToStWGck1l6XM459fuz1vRQ90P
+egT/X7LUpRk4cLTzID0V8BL8bZvVLVmBzRTN2IfqK6x//W5PUt3uay9N5+HiE6rSGho9kegiKgC
+oQmbknkqpRYKC5qN99umukS/Q/KWzBhJp0TBRWe+CguSQLZAUUaHcMrqsRQ6VtK21Q5SJjkycbP
VGvOlbro5dcY/zB1F7gheocORiAkaAE9LQJvyQMdMQvm4xjKRg6QXhqxy0ztI6B17sy50WwYTErw
0U61U6Ztqh47Zo8IukQiYRccnB0qowpLzovwDtBBQaWYhnc3YBSuipPHks1F5/d9lWKBNJTXbLsb
GcGWGZdk9s5H1qHE3HRO35qDAuu+BfsOtN8yk4rhunXb6GWw/DzWiN+BKcDyG3k8vRoqhTc72Whe
3ivt7npLG7RHnmX3vYnTWKsX2mxIffhHP0qSFq69R7izQdMIWHdKclYfegmcqhVdKU2mreXL6s2j
TJxE4hKAKrLzIitGsdeGY3P15IxYHBbmiCkA94sjDPlUrsRDATY9MC3Jg18rNM9nIUzwk0o9Cfts
UV/E/UokRylUnViYTUv/KzSgtUmxFmqugD4+4aJGfFkjQ94JFFwy4onpvyjvtMYN9YDOITyUQmcF
1cR99DFIf/xlD1bLynDtyRsbVpy7raPJh4472HXk+0O4F+JnkN0AuZaiUuuWT9XvCvkN0eGolAM9
MbXvFXmPR2upAjizH3Ac9HiAO+yEmUj2uUnB4jvH6JZg1bl1axqXjyT1QEX+xFEvph1JDhbP21o4
2vpTHc6tPuelQrLUMAtdqO3D04QeVUFPPymdMYu+wJq4YVr4K81EmcBug91B6cmtaWdfhHrKCusc
rEgnFcejaZm708lDdCuqQutqgryzhKi/wG/U3hb5YHIi37ls5BqB9S9VWhJQbj779Ug1onj00r3R
NEzjrAQ6Nh8r9CS5Bpt/v5mr8/YLKFKeGHnnR7qCUa340Nlo2iwHi5YoDJPy3vcmgjqwCXsEZd4O
KUohaWw742Q3Ns9JNc79VEEbr/fpGLaxMdaO/WKPXdQCc5ebEVVCGw7VJK1I/ghTj6euYOXpJq8z
4ERo7jTOZWNOZHa5yNrPqR92xBjVXKmob9frDimR2hv52SONu80dpZ40EsgK7MR8O+SBG2NsomFY
Xk41hTpM0KlmhoHQyXlFIdmtW/fBAJctKv9Ebf9hZrWxl9kO2HLb8/FMYe0rOrORZn9jimedYRbl
iyYlS9GcXuiBBIZOpLd3yE/r9wS+X20W1VsmqPm9TgwLYECfqJl9aYzRNqehimJzEdgTTdQJ6yo4
+RLx/oHhP3U63S9UcDOS86n2S5cw9/I+kLIfK1t4rsBNfUA2w3ICij9Nb7sylL9Nk4IurN8rlchT
hS220+4+lUsZ85GMKa9wlSF2UrNPmtdoN/Jr0CWYf8dP5lsBPNOF9QP14jDteWqAZTDhXD1MIi9B
F/p5Zb2vwuPUkbGMjSg3n9X23SuC8ffEzRJGtpNOn2QPaZGV4W/sew1rUJqsic/JQkzugL93lUpr
teDkz9kLrlFc61OP9puQ/+s3zZretJxDEmOoQfSLL3axCjeg1stquMlqAnLAFs9h+vu/qHDvId52
zawO+Halli1uUpYK45BqtIYI4xmYm9R9aeSuJEY5Oc8S15R2BZC9Rz9/X4LQqLML9h+bekWjEuO9
dk4XYzev6DKxZpGbbhcmB9ZUtm+KPtm7axVKFoea4Dj2iWlQrqVg+LF9Xqv/TWsLR/3wXW3WBQAG
SSlEeJlh0RHztcoEBvsD54WDEj3fK7z/s6uYVCf0qJVbRzyxGPB+j92yu60AGYze8g+CaKLUmAYx
odLb2t9Q1LOsXrJslJlwc1VRH86SIddNjZnsKTSi/tpdzxTfLrMuDgCX9xYIJJN8ZOV/ebZ9+PVe
+G+qh8rPnBMJlHoCD1QZf9zU27iHXUvoEYtOT4VDnTVgUIVCH1dKs7f4caXSAVANnXtrb9yzMayE
01+3BxLmVuyhJROwfT1bDWrWVhgOu6o2AoJvg3D0Bzaed3YPQ0T89nDjTxI+xdD90F33abLF3FoV
K6FlLR/uz+xSEDqQfcnLYG+yEiOv0YujCcm0VfnzTzy84/zbYWZezLoRsraW/5wQk0GfPUtrjhZu
hNmzYlM/88Iw+Ejt6EP9LhN5UmDrVWC8ZcBrXuuL+SDQ+ap6j29W7+UMRHWlUS+GzYpWR4/85p7c
4vuMnV9HUcv58t997r4F1o22qlc5vaBrim32iUjfhFVXmh9/1ElHN5TJRW7nklr0aSmDtvMcPeHM
3FMGRtk5Rp8ZaCqUxOFioSnwthEqA6gsaWImZHE656q7gycwvnKnpiyVUhFq2BlkvCv0JQcX9561
DzJLzRfrH8uAvbRyVp/brRGpyaIRYBaD6VWuyR2u57sicBNn77dWo/TKD/81sz75nsJTVeKEzdCJ
QPKt/1fiHB5Yj5437fYG/gNQ3FffVPVMSx+/+G69BrlWF/rZFbcQL3b60dPJukGU1tdKHpzuo4v2
NrAgcPYTl39vykJapnORDZdjlISj3iYCWT4tJc7wRA1+VeQpTR9/aA1jqHMKg8cJpzemmZ1chSTi
64MSEcVoQRwfAhGXv3fhYI9aeMMDS9mPiHHVpA1uCxK7bi9wVP07C6CDZ3FezheOA4hEtQGcszht
WYRW0gDaJ9xL9LCy1w1qCmzUv30Rghs9mwFYj6rT+F+la+szyHW3LPItAU7KHW2xLO72SRfDzGLT
X5wDnclm0L4Jv8egZIGdtpBeONf+TTAayKIymVN0UbKWsHREr2HHLmzn3l9rYQGScqdWZREX9h5J
FCtfIydOFdOdC157vYZ1FnXFqDTfU15FQSx8rhMu3yBUJXCnk6CX0t9LkDcTPgKOjdMCDwaLx3Fp
q6TanrixPOiZWfa2CaiOToHUiwuyE/8z070pJ7UwPenl9mLCNT/RPfxiAq4G+aJQPoqzjLS90w8x
34sDvdXN/jaOA9j8wV2J9XARkKCtaxZmFPQSh99gXS8mLmVq6IYTYAsvBe3/4D+3HjujAaOMISQl
sv1vHj2Ct6UB+O/v2RnnTvC1W7WbvNpcwZReEz4Wyakh/SZZ/zaTGEVX9WUu9QN/FP2FsAZBmjJW
D3fKbDJOY1HC5EdMIIbzLmIOmZLoUri3bX/Uu/Luy5Cb/cpXRXO/KwSq9LDaZClVLRRF1Zrc/6MU
5s6NvIGoKX/O8cNMvxK8+S9ExUeR8eOViOXYBA9pwnDXyrCysWaUcKB5o3DURgCIHYkYmDx33fNG
umzGzV9FSXlGiIKRmBN9L4PzwjDG2dkzZSNEY6VUuQRU2fo3N2GjxdLjJhJL5bcFGvB8b/1ftpTy
WD7I9N4a3hta5pNLBqDbqZE55pw0wx/K4dMSttNsepyhTBCJCetnFO4wSTK9ZvU/BLQBk9sz0hrA
qDGKUuSKgvelUzULqYqZvv4TNaQTLgP1S2PyaxyvKtEsjMV9HHXA7ZsSVlz7xh/IX/iVzOLq8gk3
zZiEqenpVDEf5tICORyOhinVM6g68W4tF8hf+u4wxSxZ66kIAcFZCpWIYhghZaDgVaOOXsLnsuuy
pWRUDApZhDE2fF2vGCXYDHzcBg9OqoCfqP5p+1+ZxtUDW8KORvX2ODc5O6GDdsNUqyYSou8n4Nps
7Gc5gElknhnymsTgJfUlTpqO242Gpityn1IV7e1B5V91vOvrgZ6X5UtkON1g2jjOtt4HxN8iYG3K
tSZenAVI1eYgNdxo0e9KqBpBrvCZKH77QmSm2bbK9x3ovHo2ReqX63BjqDiops/bPDejrSWFYGr9
h67mU489A5xxkdh4vzxcB5RwAT4R8o56pZF0RNJCpBxOfNMIir2nnpBXpwl/rRdLw+KBY0lkpjrz
ulrwsQzJLu+IRElr1RSslvKQC4T0BxpazFDoBZS2gPoFVTHH7zhjSid4uoo1lwQjNV6OdsflxL4H
TWPdOVdHsnBdIXe/+nucOjBQnjUlXNmdPCzKJfYxSXWW2xy6UveyhGdHqBCsMKEGdV04/g1QEypB
RDcS4E5sBq97IEjzZ/UXw7DjDDD7bfxrriE7Fs1fVUecS1EgVFl49QLsmGxp5CRUrp+qOyRYxovA
af/gFEKOFzXHZzDgBy/kAUZAY1Bs2V4cWptqao8IY09CL00z4Hh5KwbUymD5GIlr8OKcKdZ9Cznx
lWCsHPQNSPKftlP5JofuM+keo24je1U+8W1aObi8iP470cqf9SpSbC/ZwdHjkqu/UqBPLW1ptc9c
t0Wchv2agA9mlslPPZQWsJ9jtv/NdHedxLvj0H3guQx9ZRSLyf3B5nBwXOS9mr17svU4joJzYesW
5iQ7ARFLAw1kh4WN7nnXri4oFTKe/6/kKsDhkprWrPidMIExewRx20JycnRty5d70XmJ01EPJn2h
xDWoHOJOTT/byyPicGc8YfR8MmxJBg1vEgFVw4nc3pFODSLGMk3OI7IA2jlo0MgHqJLk/HKDTh0v
8oKAfEat0Y/wJq9nAxJVpgAxDKsyDVBWHPEET4Kzd2RVGYU1972BQxVa2Slu1+Igb9wcl8GTFcIi
oRE3/8ZpI/d/k/AHUc1Sv+HRP350dm+kbC7jOuU7c8PE8bm1kngmg6OB7N1T3OqmavpO9WyExMUA
ucl7oWU4EWgvyfmr3NB8aL8ErUEYV9voEDpl+p3jjZFnQz0ZhNKbwLidU4vnKJ8h0PzogFmpQDHu
t9SzeDRK9MhC4WEiUiVurmrx6TGIZXF7vu4aoUuP/05igOCdChAyA7kzM3JaRKwniJR89LXFQ1X6
ObE+HYr8u7AP0i2DIVmAB58Yf6c3ySsf8YMvALurmTcIibsDkk9ztoS2oyYTMqSlURllmKqFdfg0
gjcMrEdyEW7yNMRqhpy0lh9eY+NpaqMc/RiaZlFJ9kyjQ1tyiGzIisXuxu8HJydtsiM2l74Tk1qm
uezi8AcBM8RAvdkLlhzbTLYzh+gvGlKCa4LP/eIlWLnqTOUPLqiCY2UxyTppeSyr+qbypoAE+4bW
jazwLHAQO2bXSr7YCQ6ESFygD2QqfVOM8z1g6pmGobH7HaXoFSJJGO/37R62or0KYy7K/Im3LWWw
7PotF3U65pMdf5dEH4MU9BzQwglFndA7mLnOUY8iwmw6OWz4HEC/3xy0XVigUR8IOuAJaB91/dLG
M6ZIhQ15yVkGiKKG0MKYAmwvL0l2rANsWuR9Lj8dWaaS9nsVaIgQcwkoHWm+FkSsN68NZ2MMvZrR
i/lTiDODmmn4i0BuPvW08DeX81o1ms1iA1Jt9neMcloUly490QCsjwQUVEIHnZ9UGxlsBLb1nqN+
kzV7rqw8G2gwLUUPPL8WBEatVWYxL4RcZynouvZYKoYG+YLrcyBfPyzbolJDFGPTH/9Dalbr9p+P
deuCuwxhEYGdm4+2RdEVBeG/Ou1BMLyPzp2BDFqMCbi+01tYN2N2+f5XIZO+97G1O/ztqd97+OpH
uaHKL3sa/khkmLXkiAknuAsUHhNihrNzMhYC228RoWB7ifcxQCf/olVDf58wstzpr8rm20Jsi4H+
/YxvWiSLbsMI9vTTDnBHD3xGTXXhU8HWv4S32+JweMg+C5O7NyzsSt0p6QiXANTyMzLEMxKN2Ywe
6nXqstawj3npT2Lb7Gqn+7owgYno4pWdT1trB0fLw0s2jWGrvnygcmxBIjCeD54t51Nib/fw+/dS
2l8Mj0Yp5rKWyk6aXXtiS6+ZHwyC2nXBg2SPnu1pLrD4UBsRVRY59aRsLg81TPKYHaFyB5vXr+mQ
c+I47CXOtG6ztNm29d7ER5txEeulQslSJbaoi0OAS0CrllrnrJYbH3K6+TroGcn0ax/T9XxFtFbU
EPxCAt5jVCofp2CCj2zvjxH9lVbYfJWRHixU4WzIdoX5wdrab4cz9oMoJvX/+Oslin+V9665869Z
yk6PE6GS9ZOGD0MjLQ/bR1kvXzQHQUEK2vy6nS65Pqx4P+f0F8V8U1YNSZ1ttKUR3X2tCIsRVGxX
YHpYNqg52u6esZPOqAUtdrvX3KxYlYJsbwm9KYW8GmDKuBY+eqmjmAUTYX+tkaBPb236lupRBI3y
7Io1anQwuQdCRsLlCV7mRt2JpLJRXfwsj7oREPBaU1ttV1X1trarRp7jKxeGFhzv5yggn6ovl8oV
j4ipYSHqOmvpYcAmGk+K671vyxbyhG7cDhN6nOQPO8g5sjlA06lggEi7qfCQOsuvQwbmH58aUePn
pcFQ/985TrJ8FrYY/GqIR1bFlyXh6o1RXj4r5P4azk5VDJs5ehfykZLvBSn/ZVAr9y77zIYENIig
zy5n+0dYNPGvyQ4u9bcLGS/faMDOhwygszcRmDxMwP8uoTSEwyiUMuMuRFzFAx00o/g+4dR+7GtE
PRMa3jE4xk2V3dzm9ThcVl426+SCsEd7luQotCwiCeF0RPzUj8pR9oca4N2XYJZN+7F8nxqeaLgv
6ZHJjHHtKyuME7ueyhrFNFf7yCuKd4ltWMvZPpQI0CHn1rXKs4eWzfF5QlR4aUkkZeu2fZkVmj46
lziJJYw/MQA0t+wBea8L38t8uvqWzD8AwSd03U/ga27qMb6vAyBQ0vCMPcBo32N9P/yN6WkDN8Bb
Vq+a+pp3+jvbb2Mp4wr4y7Uuv23NJGSkbqbAlfWtc0I/835lZbcbr5R6r7PE9pq5iL/J6xDzkHFh
2Kh5F6rfaD3h2CYvi5OvNgVfJ7atgugfs8ZBtfS5VI0c1P6ktLywwzivKmUfEe5mXpTl0a98QWE+
Zd7obUB9+sVhd1GvOjy9Hi2VBGOW+pqq+KYV8kt+nnzHKGzRt4TzsDhcSA6KmP+kT53xq1AB4RU1
SMKJATvrJa4FDJvzvG/kyh9nYmPIUeqw590Y2uDtimYcRYVEMuZ9V3KD4ffdok3w9toe0vvvuP8q
f0ki4iwOP6SupDIJFNYCukrwXGEK63ggzKvbtKd4Uu0hOmUnk/rUkCfLIxMYw5TEoZFak/ZdcKnK
ozbpoAcwDUdtxfV24J0qnybnz4E4zQQ9RdHHlUZYPMpduAIY7sf5fCkjpIS+mMjs4DZpc6jX86Ms
4Zoyt8sRLHvSgJFpr6fxSb6YHACnGT074v7+qI6dzxamibV7DKo+ZTGaY6MyJkCCSnjmG0/1bvdm
NRBNwvO9X0A+h8HcaEZIUE9mKle2ofkc9i+97LqGMpQm2HxBIfLWSFU4sUf+5JdxKCVhOTtRC+F9
bsiIGwBIRIKOPJTsEvzJsDHeqSuo1+jfGGcgQoJvE3PS4SR+okgN4qiq4eLjfzShXAHTvzR1Wk5k
1f8mZISP9EHGfo7Nm2hhC3HEvbzhA9XV5Svpyl6QPiO+OBIqP+pIJwsKcAbGekQM2Tsafmj9xW0E
hJo1otTl9s1xnEduQYiGqmeQCVdDPTIL0r9pEqrnSalt3ve8qtIhLSgMfE+fYjkpMpSNckquBoY4
512VYh0li5M3LzzLw8vsHJGCMnbzbIkTo9K4PSqix8WhPMhmeE6FHNOLEmLzl9xEoIcLPfjcRc9A
jMqAzAJIIoy5v3XDSwT6WC/vM9R/an9DS4hktC7OKw6dY6fpe0dHEJmx2rX0fWKY5lUySFGQLp6t
KywWkED1N85tehiWNoHU4C0Cu4QdRdvMlxz7+z1PJlUdVgo0djQ1wUW79SbQ/nbY0Skgi1O8tBcM
DLIbW5VGTTYinyU83wwXaLpDKaoBN84Uu/xXTgQmbmGmqn0oqR8fK9et4jNN57w3EFQWnn3NMEpR
vI5sYrUMb6dJ5nPYjMnEyKxddY7j4XEgpkNGqydsowpcbaauHuCYWVPQrhsCOXHOur5Ag7vAXvy/
goAPAweiXXTj7kojq2W4jNZRqwbDyVIMlVTvB0gGsW1oTdd377r77Nn2g+svwgUXb+7si1vty+JS
hEI7G76rFjxHRRB+mGSnKfFgIpqGXJ+5ceX84Qt+XNYJwrBgIF/cw41eE9sp0XeXK0NW4DV3NDWk
EiQfRAnBZf+buQt9LV0JZqAJV+tdmwgKrnMdLCUWFJgdSIQDjfQ7TVLpT/CduOpMPvInRi8fdVUe
zdOC0laVKp4N6pAjT1sP2gDLSybfbPEbI1yvld/945yYpt06mlX/0NHt1Xzp09dJiHDdbWfoiPSt
xj80ph8pSOkPyDFIlZ1oxv0fywzdLnf2y5USItb+onn4H773UXnnFHPr+4ugI6tKFPP/HOpwW0Yy
1vt+EB5IYp2tFVgRQ9VZCi8Rx4Y1uzMCVchktrAvSCCDEcufLmtMbFBaKhhegM4z6aUyXU1wA6qY
1WMl/ePv7mbnOPtfvLaHqWxhks1YjnuvG9z/9JCIZMEQq77I04YpU8VaXoOKPVbNCXoUjwLjMHf6
7UfGF98VAupZ+EMqAJFvGgcnsE5Mdd8ArVaTVmDK2p7GVxP9lDHTBD9U8GNjEFJcVhxAswVYLuwl
99f+L+xcGOPO15azrdtVL1bueJVgVyuKS0//k0xRqVyY8/u9qjl0GP4NPz9/j5z7SZKEsKIlYMXj
RLBwTp178I3WUOnDfLH7QACOkJ7FBorxZPhH9pApaBHLUghz0KUzaWKgpbN1mhre0LTOYj/a0qCh
mGa14W0/S+yVC01avQrSRLNpRGhhaoOEirJEa9bHh8LFbaio/5LoHfUs0w7hFEV4VVuDmuUYQDY2
Q7RkT8czzPO87PVidUif0PjbZJnAbXsuREEf9Ful1MjS+KB79Q7Viy3e459pGweSe+3LlmBcVAsT
qCYM+RaZOiNZdCnmvqN+eLMy1bz2xPBUFgx92d09h1eLMW5xBqVNuLtnF/vmNtpuwe23tFK19d33
fafityfIr6ydD4AiVucR6LXenbDLbNhLeN/YX71xNrfQ1u0rZSRMdSxEO5U7aDRDgtgsSAig0a/v
rHIdLyGth4CEESi70Z9iYv9q+6WwE7gHEFysh6oYSZfNjWPb4njl3FkUwCQhKX/XwEZ+QG4vNl1F
Xx/5H5AcPYhSbOKId/SoWM5+gfnA6FC3LoGqB/FEvu9tnzjYSHVcitRCwxR5wdc/SE8TCPq37A7B
CWRDZQvtH9bG787tSgdYnks9PnXfgOryD5XgpqK+ZGGu5W+k9H+1+4L0dyCHaTXV5mO33q5JfbbS
iWHH6LNOUcfBIlyG4NuZnxDWnJdzWeVc+01FV3hqukveRKCnCFxSq5nFX5F4vH63kR7olnO41bMz
9R/qJsnxU0WP1Wsqv08HsXjon69xobrcvub7MrY5BOtK1OF9bhNyG9saxc/aGQV4+vmpsAvVZdko
ixWq7WtQkBwOqLhtZCReQVz65YQAvlqn/dp2qEylLdn6afyYLXGWI1ANKSeUhHGXawhTtbKwuAYJ
Dx8jT1886GmWYvnsh+Xr27crOwDVP3CwAKioyxBp34JkoJUAhqZE+2328zAKi6Lxkslu95LF2/yE
L/Nvx8fmbx7cWG90YHDtBjD+rPm5uUnQipnbcAFniiqsbmXQ+BEXSh1dRZ0JRv7CHXuPk980LoYw
ttxZp3S47+1ItlFzXxZXh2KLEG3+cxNRb/jirHasv+Da6xUpBp+EwJoYpYWjgyBlpp/N92d360Lx
L5OjsvbKKD5h5ibFyn0vaEplvqjTFkms8kDjGkhPP3BxwKASgWpe6KOstLk1JEkpdDNsjduBFrMA
+KtoS9HUsc46g6hZ+KyWbWGMOuyK0IbB2SotaxbOz89ylHOaGkXXNzKgJ2zuGHw75ZFoW7NlpDjG
WN/PR4JJZdiCpQ7bJl0WYGpqyGI12eRZ2Gb3MSQwICcljBhl2PNHXpZ3ZlxQ5zTQpjFhERtWAAaS
kb74Ed/Y+A8757qTKqXpwAMPfgQnKrXcoigQ8y0rut8GbUluBhLPvRiymyObHPv3KOw9xf8HE+F8
zYt3MaJaDiEG1UYuTADX2MQKVPYNDB0Mv/qwha7P+69OTtIywqr5R0LxgV9RXUTYGTzrV3BlLrXW
OTeTAp3gsU9Xveyo1mzDBnCyAfPqGyhPvZ/YU6LSuyRIh+LI45IfE+UnURu9m3ckDurjWTqcQdeF
Egm4V/cP5ht5niOkzhGgUu5BhoamObgXFrB9HKiPVwyeH6p6MqEvKcHUukVBtNTccbqfN6PmaiUm
mqWuSEIzRsmpXAmXyAgFhB3RS/BWTJrsxrJcNJ2JLWbD0yLGl0iILNLy3R1tPInqaFl1f0MeqrcD
8vIO7UZHpJKCpL7iRZLIacIaWSdtAzNgCu7RmKONsR/9BphBmaljms0lV3hmoxyM9mefIUkfZrWh
WXk4AUkUmF/w6heNW0URmQ9UvZvjFqCZ670z4rgkHfUlz2VSOWSmgLomXL5cGhoCiDYYyIRDJxbT
uODpW/ie/kiHWs4uyMGLiOyQk7ENMywsDeGzq3DurjEWYhZ1Eg9leVQKBrlUt67XxKbZsKFbk9Np
L+ZT2poBJjIqgarGym+ZR4aYJWYkqVjiuhTvoOA2rH0OKdgUFHBcwFKFpygcr39fqFDIxD15FTj/
1MB1CzkTz7zY7EcP2LGUHnakRu8grCeKL55p9e5DN5x7UVJchOVt00lmZRNYMwGQ+fnkuU6OfsIX
AiyVifZhQi2SyBm8yJvo/jMme0oKF8nNRt8nsKDVnuB+ZkJfnfgRDRUTJguGseiasnYuR+Kg6Dc5
/bMAdtHiNDhzz+/ewdPnEhCvoZ5v4wZQCv8NdzoWUUJLnjwj71P2n/KWxKYwKqUGf0zaKzomsKXP
6zrJv73BSe1teKwDdzHLeVuqabfNfR2Anyooj6r/C2v+v4+r/RJD7q4eOejycpoGpIDXpGzpMb4G
W2V6GOnzR4PfhyutV8ix4RXjILnfYaVkdCMDSaUaKqWmkHTuIQT4nppHTGPmZ6QBqhfPyEyG2Kwf
aXa+IQiGOA9yrLTJYpWXJUY5exvKPRG+YAo0EGd898SVASE3/AQjKT8b6IIwTKRCkqsqS6BO0BMC
cIXDxwPnpvBl4/VzKVvVF6J4lK/42ITa5kmDMSy1biMIkG4FEu9WCxEQVUVMI7bgL18bNlQr8GvJ
lew+fP+xJH+YnP4ZCPVedQENPVkpt1gcjbIeuibEZQnSetGnYhA9kiWz0m+z0c+WUiqfFOBZTLPN
JB282/hgdpGzoNXhr4nIMOrZVDeNDt/qWLkZkGU/a7AdKUF1kuuFhGTC6GzrwETDLZ+icMk3v4U1
UZ000Grae4sTXCAXxsA3Dak0hzhO6lWoD0hU1Og1so4CZILdkcUyzfl53aID5sizJZ7sSFrueVYq
ELQUArLAh/ZS+5Pm+YlHekISBFeVa/gTLrpLSlJes01EkSqSP4hKgwTjQALI2WzHownMLp6p8vL/
8fTI3ga9DcAUwzpNJdt7aaXzkR2e+5W3WLrckQ6V7aBYofH2B6XVaA7fY/QAQ2Z5G0YgoG1PnNQ2
2MJUckQIJ0u2EulHdktQQuVGew/97PExDY0n9bVU5zLDdFFj+VfltQgDBNuNTvWDY94MlASD4Kkp
Y76SOYvEQdLdC/XdWL/DRbWUlwDy/osgDxONB6HkvQhC2cQZ8cGQoZ7N1rsjW53Gh+wd3DWopWvb
DEqgE3qi809DGiLQEbOBFLK9fZyvmtcVRk4INmIjkUuUbG3olc4Y1Q7E2wKhRvt4xEux79vmMa0v
MGcfzDeg2zbrgTFLrQDAACKT+cGTpT3hSTzpnjfs/8rcf6E3cNh46aX30lYGGkjaVskog6HqULLS
tlBJj3ovk+hxWp6gRfXkEhBYH0awHT8JxTRXNqGP84KygbEgKD1aFGuKsQmlE1OvCzPHsl/ffQgy
SH8UG0x0mZP6yqIebaEycYve4Pnpk+Ghqhf0PfKjXrysOcD5PpW8v0+JdIWpYQUNRY7hSDvwgJ12
DhOtMOXABLvIfl/Q3tt0n4YhbyWE5xskrlHrglgJuSrAUHF+4gdcVpCQK7P369PWqEVWqLGrEcVI
WPNwb9JVCPDzC01J9rR3KdrsmTnh6eQk/Wd4QdWpChoQ4IK9CSfcjHeb+Okg10AQhaPI99BauRhy
OQDRrlbW9/Spagj7m7kshrUhjYLTTWJiiNO521ZNwW40Owq+3G0CpiRDgqZSUyH66cK3e2UZW3w6
StMn1nCIfsBjyEscpbxaIof1CF0ZIStJ74fwXjxpfI2CY81CkUqnxRz315xi3DVRkrl0BAiOZF3K
C9RAUdFv209mEzT9RUva9pVYd/ToIn5NoxjKrxgatF4M0sGu9kN3ek5Kn5g2Ah25AX4n0i3kojVL
sbYTVeO/lFIGZ21z/LDzVVdxI+ayPVc4bQkPefkEkzS0izjRzbVnKca4s8UIk/C8spSLX0g=
`protect end_protected
