-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qbsN+G9MsHKgYRILpxWyN2PgANlClqhpuUOs9YDktz2F5ouGMIh3mHKMPDm+trfWaJsbYJCfvRCv
J2UBDTuv46X8U7fjJYstxs/1kqHdjT1lFZskJ5JC2uR/2HuVtKzakpGVopGrsrqdlbC079eOysA2
VXC0DVRJsKr0uApmBZOFE/uC5zMGuJ884bqRblLX7M+AcBHcqGtaXEN+VdPvJcrfUkIaxvOgRWxT
cCFb2QqIh3ue8rJ2hurqrpOnFvvbbCVz/iSz9vmH+iGStj9o23TF6fFZWPe1j0Tkzx44RTdkFeyX
bcmt1HVIY1t2VPLaDg/8qSUq9TK6nS/7Tpo8fg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
rSS0kIpZx6QxnIIE7zEvYti9rOumHWTMUhT74Y0N2GDyhWrmDtqK8930klJ1m9sW41Be3lh95aZN
iePTAJmHyi3JS3hFzQBIFCERnhMCYa8vrmV+KNmKpSFtKGLLoXD0gquUK282pb9k160UyIr6zmsd
LNl+pLJHLLVHAJE9k4lDd3ZhdOjhh7Wn381jCgWVwMcBerHZuFU+1kjly1uMT5hLfUq0EidLF7Yj
v+j4IOQkrDs55enX/t7Fxw9Xc97AKpbq+OF3sYSXAHq4qNWTYaT/v1RTj0bZnEL3GODMJaNM8flP
tjvtip9mEdDyfr/Nfg9k4DdRFOc8r61sBsQ4ZWBUFevytZbhj8AU3TVNUGvXzPce6ZNZr9PjXIz/
oz/bBLhYBJ9nQAP+/Eu1nin5Cr8PtMQ5YOUelsQasza4+JhiZrPepSxHlifPE+ot1L580mrM/NIT
rZW71YiJAUYKzHHGbzrlRgYechR8204rRyNIkiNi9rVRMdNaKb6VU6FtFDYajExnEOYmmfZdAlFn
jAaGpqVB6wc0nrW9WNf2Qf7xFTXEK7YXtT9Mf3SMY13eVoXlbAq9bCZCV0c4vZSIRgXTgx3H9/5y
Rt8g2fX9j89mD4YODYLTu/CvJTuGz+Vdg0CFWWaEOr/T8e/glMg6rg6Ws+6zS4HRIGc+R2KaVwsW
OHxnKBK1Sfxd0nseB2l21rR7TevN0EVbY++sFhjEZZtbp7uZXzj+dsG41kMzCOx8Q4eeJld+Anu+
MKE3ZCtUxy34PK5AZjrxANG252L5XTUJvRCddrxw/Zege5q19dhsPgrdD+HPSVlfG+Kb4Tbr0Eil
HDN1keLZez4rChsdowNSjEtTfVcaO6w5XRxbM76hwgAZLHeFNUeKpy09amwyUq0Q7jKI6gcj4F7H
scetg5VCtgRkZpUtXtt6ks/RDO1j6j9hjnTDd3Cx7ma3F0sImDOPR0jKtBySGEByvhMi1oKngRTH
AsWn8PM+qBfxRYf8f9tFyS3rIaPybxe5CVegBiJXNwqIbcVDgPULuNlXvRfVTeoOVZ6e73e2ychc
+VM8r9Q1+zcLLLMJcY2xjTQ+sJvtCSD3VmOVaWHC8V5YA3U32Yr7+JREq7SvzP1bUglS69bkxRuB
fLULNgC+xRp7aJIYsXpWHg1suAyQSvo+JuLqgv39mA5DsicF5xXEc1F1P5pmNAAf4RT5Ypc1mGbM
Cbzr9tPqIURdX1OslI4zMhWElTaL29vQBvoovvIQJhZfav6WxAbRIP36dwojhMRir+5EnaEcpxeQ
dSdW81vH2E56rDDrYxHCT54uhvKowzZ1zothNWfL5AOjHlyL2Zbef+C9J9WXdJQKl2gS7zU3A1uk
/ZWCi8JtgxcA5EJPQPVJwvsfQNaVx0DoAy1ZqM5Ws1vtOLppHCWT1ffmG3XaZ8ai5mejNE7qSLZ2
eQs2qE+QEkgHwMb2vlZWLT+JJYZrYPZDYmoai2tkP6JlubOKDr1rPpo5/iIROeiPJtKjlOdPeIHE
yBXf0ytYfOEslGF8SSSbVDgVkvaXyeGFl1iHXNb5dFmE2n4ytF4AYOToYoKEhHxw0JjZNNHgTPvH
fZyRaV6xhxcLxTaxh85czPv3xaxO+bmv96YtE96FE91xEJj876hxx8FVs1xQaNU81EA7YkDjScCy
pyYD6oiYl5gGJiKvTVRvMhc9jnJSxKhPtZh2Z4rRjxU+bUus98U9DzIYRSSf5/nrx01XAgvbNhM7
f+gIVpEv6/TElm/mNAT0GmMXJIiWYf/gkmajnJ/rreyfelwpO4PSW5H82z2HxB6ZaCj3cIkFnVxc
rCmJ8RTuUybNIHh9LYL/MCbOaQ8gbyY6GXSALCSzsgF3VaUDaJp/T443RVxwD5V7O6pKhgsIuvQq
YV77ys6mATwApw+YLgamVsAYFdjzcIpaiuCCewKdandN1hwMfvUY8FYHGxs3plhRJlejNaAcpK94
vLy+BA3bf0tBYjeRIQq8JAXFbwgGoLdE6se7je0d+7Xrzy9Ut6AR/EkH6TqCa09j6BNxQMKi2mFt
xCjOW9fH44IkVGUc0jRAzax2SwEKkuBGwORitKxsiYBm+UBQ9gX2swOGjW2YPaXSTrDYU1KKfNZL
Ag9m8dT2dcnK/Uvzz2n8NaTP4yMwZVxHht8rlo/P0pwioOB/vDPW+/8J/8jJyMqx9/BdoGRW6uXn
lqBYPWAvwA4rTyz7Ojfc+Rce8HLNyHy9wnyeN5uk2msuCFjcRIaMxBgLcl3WK3jhDaIntXqfRU9J
FSQZxVeyEKowI3wPQo+CXOGVI5Xx2w/6fYws0nMFHSv5SpN92KahwZ4iB7cSncjPDlXcEOFB1ay8
5fM0sK/E+IfY2K9IsvC4UfJZ/KRw7KMb2begVOqh0XVMb4YrOhXeBedymp2pDXk3QbpGMuxs+c2R
DuUz7zhspONF5ePtx4X0DaveGrspd5cI2XCSX+hoCnW5K0zZBuYCljAYhgZPB+/ofr3ZAFD9iXA+
57nYdxYsOaoNDJ11auMcZD8VJWYQW005Y/GRquXsL7nHjXvAYFQJpMds4BlfAYYnpyo1x4M1qnhq
7ltQgZ5iUq1v0M206W7d/LFD3yb33QAGyz0cBLE1Os3VugTg13h6SI92ij+/FdxrjQY8CSUc/iTL
lWYdo06w3JM9FnP0evNir/0XpYFs6wFW/U68vUH0g/pifsdZIMX6re5iWiyrkY8K2cWg5iBprtoW
8C7agFp9zxjcvN4wb9z8K6pBgTpGpCegA1+ZJ/aTpOQH0VFiKS3VRkOVbX/WawNE9AHvm10LqRZH
lPXNPIpkRL/D4iQYATZERTiADl7EjuzHHFw4pZ99W0roh2cWYP3PjAEnm6aB8WwWKP3EkS4LxJgM
Gtc4i7S41LmsEr/Gs6U5KLIPyCs3tsf5UFRlAdTd+bCil0Pe6lgT1aGshfK+9lnoI1rXc+kJQkGv
tZhO5FCXxbWnZjPeB1vrSctw4LXKJP9psfId0xpjoz6cF3ZU4Ewvy8EJnzZnzVhnQHPLWLL7YvzT
GV18GkB4OkFZmo/aFGa7o+IPMUfCg8MJz0mvdz3rZ/Wjg5XQTKnt1byZfMuI2jvAKJcIpuz2CPOf
xmJIiVrpMbZG2zLPZvvrrFSDV7eTl7ONeYMpyF9UsOUxhtsvfliIJhPg9W4aRkkKI58dTG6b0jJZ
+Kyk+QUtZSreIivmu3jAGk9epI8Hr1LSGHQj42OstPqidgUTW8TQHOUaQRswMoMWesWO4KCIdItH
A2gOIqviCjJHasaoy8r9fWFdGWo1Zu7H8Np3kpXcGuaGDwh3pHz2a1TookLNIU4Ha2B4vF0gsD+0
dKIf8KWlzrixSAVMHfH+Z3MjouhLgtQse77VaiJxFWlSENZFv4+qiHRvRzrerDTKbPNxQIvsSbjR
JVNYYt75p6SkZDdaiyqYj9rHMx/uRrhTV7u2JKNjOlV3oNbqSIbddNklTJbBefdLqxr520ZUJ84W
z4tXysiYRoZQsOY3I4w9XfH3NDEGbkpN17z4k5/1YFsKOlly6nvC1SqHjgMbpPOsKiQXm+rVr4wP
0Ocq1b6Ng9yQwnz4yoLFmqOMIln5YTvosf66V87Lh8OPs3sA+1rfZGcQxWohQRWJbvJHciE0q+zU
7mcNMwBypO7eleJYQEsWOL3mN6NJa2k9qrzx5TU9r41n2CNqJ2g0BKYiO3eDCCoAkatiq47bUZzM
e08oD7W5CkzSiThvXkBRLU+nqgMQX72JwCs+B6/vBRxlvb+WDatXAYZGfae1zyG9Z19WuuCg0I+T
L+iO0LIO4m9PToF4FeJyT9osSTlLTTr+JiFEYReAeQZODhgKoTzmWGR3s4XFJxxaC2fmsvj/caPm
r2/RcEN+dJzxjOX9Hr0ZarVybyyNkTfPnmkjMzVJzds7t0N9q1T5lK6UV/2fElQ4stY/7pexwpjS
2Cr0e+Mwbr+ILRHutUUgjDsgeyA/0nFbMR9tzO6SJ/u2zBVOdkDLmJ7ZpBtSOCZ05TINlw9b5eB/
x8jg86F6MM0yJbXqN+2/vH5FBG5iRo3wwxuFnGXtijjsjueufZNyy5V8aXSyWjvGRU6P5tv1MQ8l
dULW4oiorVazvnE1KjUPrtfezeoZ2BIOdKw8E33o4E1ev4hIDd9fxKct4CTsiY0PfCeVlL2Qks39
P3jnA/P9eRwXa0jt01FLybLEoBiSVYp9mMc+Lw0d13IKRVn/1eMdzrMaNeptdUAPD9U1GScMS2AN
+AsV0RG52zyRAyOUK2EuP/v7caYCCV91sy8Kwx9DzZaqX1RlKsGKBFnTtSQBZfLZ8nko6nUl+cKN
3RC5IZJGxwrpN1cjf0TqfIpaBy8hIzu8A1xLdjkjO1f5UXGSOC9cN16IXB+udCt3qMyR8ZyyNV/z
SzOe60uf27w0e8axd8ip5ghqzo9Jf5fQZp1M1Pki0aRvelxXqgMxnfaUWUqq8OYti6rI6x2sallA
Qt3slsenaR3k5ZfTLAhVKx2y6ukE+ExN5NTvZsA1HxiOM13OyZnulYjeINo7t/U/iyZtjp962J8X
3BTw1hRVFAYoprzWMMCQMe7CrFc8wijdg0/6+nbCi0BR6L+aUdAhISHTLJfjUk/J9OXz2V9lE0T3
YcXj+lGNRLZVGSTZLUjGarJFf0rpaK3iufSKJm6RDqbmiifDtOQq9zD2MQjw2MNeXGnUnOeJt4je
CUoTHCk0Y1mqt97gHAloYSf91N4+mJGxdFR9crVxB0FloRQ8lx9OgmNrMfn5uKPKzyrXc8i+EdhN
xRDlFQ/91JkA/qusXXvs6KM2JEvfwdIMyPSzqXGmA89Q2QzOhW54iKvT6V8h8lqPccIKnhZp8cyz
YSTeI0LfIa8u4UksLQ7nIbAfjc3qoqA8BYtc+HMweHJTqAM2r4f4sK/flGlzABI4RxKsu1shLL/v
f7HwFYdW7HZm4ZoAPblHtdxcGuS/37tuzhJqc1EwSM6NewB3OabbiAkJN0r/2LSx9sb7pgAPvLaS
AuGlC3n+ZLfo6XFLZqL9WuiCd+vhE8ul5J977ojNG0TP2kI6j7TI+fTAf7hHj5k0J0r/YV48cMip
lO/EBpzYKEV/A5wxPhIiGKpbEvWJHe+1j6aeHg9HVFRdEuM/GDDm2iSbCLFGXp3jZAMPpCCauwMH
TbS6r09WARb29rheMT2vhqPR6LzPayrUMc6IN3KqCGiwUEK6s1qjWIaBWAMMZSb06il2Z4OvbFoe
dzNoN+9biZHPkLiW8BD0qSBRVmHprl33EnjWnofsX0ClpxBhhGlNj8ZOjeQ3f3TSrZho/akZUNFb
7OxlguG/6eCPEgsrH7hi+BYC2U35UmDiTn/9CTqZoRlv8DEQSV0XxUrHmewFxZpk83qZUE4JnTLL
/qIrvRcTJvKTh4Z6JxZT/nOT06Og1I/X8jVle8C6kNwypOsj+VmfYdxLXIp/ZFg2tH9YaGa8znSN
aDzApXrOTK8ifDVzSuL1CVPytYZ4XO3NCgppqFJId9tTNxpW9pkMP5vTeRdRqS6UBfWMvZcP8LBR
rbpvZxvRED5ylqbxHKWHzteOgxe5m0Wg1ouu1AEvkeGnmq0gAYbmsGtwboQD/XBM28ZvEw8itzOU
VbjPI6hH/hNkFcANLcYUx+00SuW2Jy+15hfqA+IdyemwUBOhrdK3BP+rOHvj9SnDKgNSxUZRgcaP
GAn1g9gfGEdI7wwbUxIQ+lfpNbAxNhrarF9/zejvA8SqXKYUREFbFdp07e8xBBk/+QNDuy72TKwX
65LJAQCsQiC8Y50VmjYDrvia8BCjkKb7XfI89hxs8CEPl0VwEyrJ23vSiSB0WuveRwZ0bpdH48G4
/HGUxv49mFXTJMY+KOvm9+Ymv5SJgUsWRPQL7aAAfJC1X2K+F4c2AjZgr45OmfYK678KubYh724e
DGyxjC1YKMZiScr9QNTE8xqi1Kkihas2h3NpfZznB/tIEx1dN7079WPIKhQW+ZQQzFP5MQ1Iz7EE
OnFId2LJkx3C/CacjW9emUzG639kyJbK2Cd3imUCmZwqJP6LLDnSF0yOMCIMfmAeuif/dPx3SLof
9PVZVfeegAgAMTPGuTEQPdRSpgqre3rRmxdlYxesR856tVpEChIqBYMMLwhV5CPyvx+k7i/Lvd+P
/9lC9YWhTf30tY65LcncpoTF4VKBS4eZBUCcvEzuPk8SQXtTAykiuDIzBC4+jZZjd8F396KQQK6Q
Z10zVJwYDeR7l48KE8uCg4eVbOltG4nZFxbesMqz1fFX0LKWfTVGZaJZ0TMQ0W6icfU7vkSWisc1
djZf+yl8BD4+CT7AFI6ZonNZ5dnKSmZBriH5LJcaXIQFtbB/3WavZuObk67AC5aGYwSEaItNAhEv
eLbB1RUZv8rgUXgUIZq1pKsvA6r+pKEtYPJD68FwZ2U1pvmUJYBLAdKMWy7TeRijEY2NBs8aNN7u
eZHyTKnajF9p30maLndXC05iZmjPCsWQciiSAKXaQz7ZQqb+lUPHYA1fiywR3S2vrjeaufaQB7C5
9YOc1gtBsCQeCnRMv8ZTA2cYIqjJzwD301pSGu2To/JnclfbnWeZICGZwgDbMelAOUeISZxAbj2N
kzYVA9h8HwGxyKNmhicdGJJ6OVVsjU4UthWApgY40GeX6QzkVhFN5YvHC6gCwYwSb0haGa0cHP9R
n/s8gFRDhYfk26W9M8pzdVYk8+S1kNaLoUB5ZYIGo585nhUselrNTpk5p/0mV7O4gsePfx/MT5C8
o83hnjaePfiy2s9uXYGQdKwSyJXd1dFrdXI6XllJoMrqtTt8fdsFS1OLp1W73QW943NHlaS/1Xwy
w9CUtEs4JqNJ9EOV7nVmg7o+lZgj5YsgbcwrRU6f+qKHOcK9OmF505UJ2TPiBJhNsdMd0GI5xtRD
ow3HeBS5KYxVZfw7zo+MWFXexhQYchSYieoej+IVSdFqA6UkFEYdQgAhhQyNjZckg+zFT46tz/Td
w3mqYmNt6AM+I+AUeDmhK9I98fMSZZD2QxNcrp5te7hsVSMG5cTwqR91F0YftbNvXco0KfzDMKSj
BI33DCIwuMifbcf62kewZaN0QYffv1q/M50JhvLzGwhCB8Dwn3FxzWFZ61ejAHqgm5J3gZqcWZ6r
+xU/8jlg5FyZMYaZiZ2DZl8BuzhJIBXHBfvzraTPwS7hoOZlyu92oIP9ff3uK+1dB4xuu0JLOF9u
/2CP49qWSLpYwT7ZsVnqGOY18llN+vVBaqc6X1N3pqi7UAXVE/c/oY9YvnURI/qHG3V+F7fX8J2V
s7XVWU24qmgCFcjpkTUgk+ulpmROqEf/9BP6SnGE2fcvop92INW2IqrQ3QdEV9ZE8fvqa9QMtQlp
LiVsuh94Ysmb8LxlO2uhsKk3BGUzFM5OzQu/KHXkjUg1OlxckA5/92zWwbRaHOhbPOa7JcKt+pkU
t5mjKvVhdUS5FHjEob6E+0ew3/Kw6sjuEObxUzzusOyXfBl2IBvXPzxRv7X5xRYBilg1P3ao02FA
TYN/3J5FQJ7tMATIbfEnIz5eY8QaID4s0OoQvWc4i3c4XbThDO8sajVnbAlV8tfNGAYkhEThXs4M
5jgTPiuAJFcqkz6675edSY8YeEUPpbEj3SNZl80FtvWhO1qxvBgOF/IF7jcVdRCl85oRNO6zSjlX
JAelAqiXIapSNEG6MryB0keaX1r0Wp0v9/aTvbUgiBTyyv8xAZJgvWu3WVG6EYub3VQzUFpmJLPR
n56T3UGfqmLooyQ+RHBq0XZrBmcKE/7R+2D/Xz5LAT3hDUjDiuxeS9MRhNgRCZzJet7qo2JZDZBb
Gbidbzjg+vTVoJFz4WnyTfIVgE0AS4jZIoFjnvdSI74fiOSO+uTDrMHDTlGB/wU33Naxz2Z7zbEC
xvu+eGYCYhdWik7CF6ew+iOj8U2hN1VjY5FXm6uYKzV5VLs/RhxhPn+zjNaLvtnPG8SYM7Ca35DZ
Rmo5+aI0fwCLvx9LrjqM4GhJ8k56DRW2e+P45d74bnsA60ZVp8cZlAB21+oAF/OH3uBOKWvgUxQ5
4FNiTaCtg0p/ud9Bzn4fHCx1jHEUBe0HYjbgw8/lCUyWEl/GOeKMcFwbLHjVsY21cp9fomc2tbKs
TnIPAH1B1PcHDDDPT3Uiizxsjo/ab286WoHvUNpDJibIhbXxNiWERanoUU2Pm6H5uctlXmdM8vU5
f5aMM+et9MavHZUdAZcwxBd2pSXVU7cBXa7bDc5gOijhPbA4W+zClCcIRDK2IhYbG7fs0exZ/GpW
afJa0/cS7zrj2Tj095z60ZW2jCiAJS2CacjKX1fT1bn5ZbiWQCELQXHU1Mq5vRGdG/1TZI2yf3vg
wZpKRxwN2eMWPAzApKSmB4JRg/BeTXhP3dzYwqAEsahmXbgxJX8suB/KBHFHG4WVBWcGhBE72Ncd
hEhtYdTvhu9WYKxjxaxSqfVbd6OvsEBk3bS53JPCSE6eRR6hk1+EPOWIbJoFPOGNfR+OEfm3TIIz
7wBFkWtYDtVHn4BEtrTZQHnFwfjVB8vsu41gCVSXWUSJoI/2Ai5i2139I0vHWPm5T8sINgCFfhnY
Zw5gOr3MGj5GIes9XsIwWtMT6XoKMVXKWksOWvhf2S0EbUkH+GZ8wiFyYJSfI4H2qeoecxKIWbMu
9M4BhrxbkNHf1cgz4l21OwU6p9rZAdi+G3apnZgGmdW5+XzTQt5TPB8e+KWYXVM24Nol5tpk9+WD
trO0maGLSiAgFY/9py06lvjYFDyI2rHEMKZTlLGWpQItJ/yzeX9T5CD8q+ljvd8MvL8s0gqDehbk
NDVhXA0w6nu3uakxVCs6LLF5nTcWrzBAFVDmRJW1rpPK9SAeNZCTFWI+j22NRyZlihwJKCUkc4iC
BAGu4c2sLTng+MG9Qsx2fRKEpOPxk4yGUj9V17WnPtqz2l34cu9pxCoYBI+/HG7wUK5eo7lIKv9A
FN136bf/vo9Hi2x2jPC9c9VLWN66zyS9oJ6xtlb7yEua2sMgsfeGklGxgzDlTPvSRMQP8fUhxx5A
IEMxrsJKrz+cQewgI5icbHwinPTxoqqiANieLXuSb3JFZDu7jiS551UgNGlSVfAH1ICZJJ31JbLE
if3sgy6dzMsBJMj2tCJpumCMOQ03WoTLQ/S13SM9ynZynbATXDYcoZ2kJU6r+t+LAHT3tw6SZROD
qHc2Xr/doC+zDo3o3LCLC4nFoRJPoiWiwKfJKP2PUMyS6sTMOJkwSXtG3FcR8Sx4YNMd4U61aGnH
SpQJmuv6yhnEgJbEZEXgG5Vq9ugt4A54stkz/6veCidk05VJ8QY9MZDwUURZ61ce7fPWuZosnbwH
sYouPTEAOXkxNau/qBr+mwlajLZPHnREqEM1X+NREbCSrvY++BcahTO9reMVtEYKYO9zXC80URCn
IKwBf79G3ddVwxBmCQmfXnVSPqaHiub59S9hdLI/3ytpJT7Gnr/n7JxHMZHck3/Ia2z8u/29rnWc
LCW027q2NdrfeKzrJkNYMd47wcKFFieh7ZMA6z9oHlM3ktgEA8F8mT81GISbMOlhzd63NgJjRgI5
yP5MCUuY9UVuNQWyoHEA+fbyd6uDLWwsCmfSZri2ExSnQtT/LPeYvrCCiEjLvL4oyYf2XoJxtwP6
8BofBpfRK8gM8CrocOhOUUzdsHfkVCBfrC4asuSY7jOHsX18m3o0MtZizkjYfc328Y+dMqkvGhbs
iooWZfO7mXzMmbZOk+Oexah4gfkZcEIdjO76+NvgL6ooxqGWoRim9Kkyk/jLhvoAHu17z5E5RZ73
utpB+aaDcH21AJkhkAxcPDVBbozN7MyjScmci/ZfPmTO6DLvcY3NP+ADP+tdBDkBBpN2VKavsL3d
eesgXJ1KLjljACLmEmLLHYWwhMUR5vVp6wzBOn8ewKjmKFfH3RI7Pq2NtqMjSdujMszT/DMLRxk6
kwk70+fhI7DAljU4bItjjhYC/PTwgEsJ/5/eNDPssx+9acxu6x6+8fL5UeUiqoQV6L4kadB25jRW
KI4Lal9AnfhVHDo8lPTW4MBPmxRxX53vSwZqheco1EaOc9+n/xOpbxTCeZQJN7sCXX63cYgrYTiB
BdY6Jp6lyRBt3RFf9WgiVqQtH6pHS5RwgUPTqgM8Vx2IZgZJeeHX7mrUgn/7wV2zGRx7REwkAFod
g857VmR0tFW8TSwiqw2hNSM2O5eBjZqO0ujefdzOClc286jSfCcxWQhcG1AqhxEiKydFsBLBoskk
akDBNcCFG4okg6TbVox1QWo9NCznOU/JdhDxjyQWPGNcZ6MFF1OhzsQJddbC7esMmbJbt+jIxI8L
qRmxz6yneE3dzDv69c6hUMb01NHHHQhrQ0foHQzrkthTlyN6cGHhy8cMHzfJg6pnW8S2uZoET6HM
v7+nhp5KDmtwIDE1eBBJEFZczm+LDASxnpaJVCwqx2nX1y2LakVDcOF6qY9sjiZ9CnCBduZVfRPp
Wz2BwIBYMxQ0Qt9psG5yCjotDlY8ukeInQIel9NQkutch7bh9457b0+fNSGbQraArV688AKx/1Bd
9ZYAs/N/gIX1E9lfi6+N4uqhpOFM69qpEEypZeZm9hQWLr+UsAlX/3wRzGDEg7EYfZwm12Wcm1TR
pQKcZIBU06odt6esTq0pTlzi+RFdt7p4nYgXYwKfMD9GIuF9wudWRUQx99RKazWxdpXBZM/gJI1u
Hn9R7p9RB5ivtyO3jrPHntyVdN66WEe2A2Ry5QB8aO3Zj7Qi9I3ZOuuMa8FOgCQGPdfI+s6oFTBv
v1KwlVoEE5NHH9hb+2tc6ycpjbfCkpDwHkcO/kasz+dGSf5f6cwBrbmvdd7sDtZouJqo8ZwCZ8n6
w5RJXMFMiqM5hRIonjBLaRM31O+qNlbvvfDEQ1YZ7OfDr2rYuWO65FGofAMpiu6oCwPBcNn2lcpQ
QTpXZJbRu+EXSDlT50eeIYMeUJo+82y5SnY/Bg6GRIpi20YSB3xMzRHrkKhvlZMHHGZjoGCEnteb
Q3OG55Lfc4KXSdMMXlUri0fNPEq3nnxgPV4vtYZzznGg1FPqqretJu4Nqn87UyOOt9q7Ga4eyEe4
zU1RAiNMhY2Rq4OevDIwEqFxvSlm8W2XhYdnT6nffKknO3z5nbGf0jfdoFhxDE1BC4PvKoMpkLYf
/DHqf71bbdNlGWqMB78vLtOP84Dad5D7ikdyv8UsEPjKSCLNWJ2DIXxi7M9JX7+932elyfslfah4
3rEFPjicvwHHmaHYEMlN/DRtwabF+EF5YuysKtf9lFc7B6EAhcE6X8jJ7Upupz2s68W44MpsJMY1
fPELG5A18Y+JzFkKPHAMq8U4jgdY0z147LAeKQAQc3D0kQLQbfSeU2Z1HQdzHqTlyCd08VON7DY8
Ci1QxLDvUyqqgIsWfFCGRFC0onqY4oY2SRiC3yjFCRKWDnBWJ46l/nMxojRCplgjG+nevDGmavVm
B1lrtJ+71ZFQFia8qob+ZHFR/g30XzP+QjYwNuFH/zWZb8HS/+Vl/WNtAPJ4mxzLjZZ2a4MnGxmI
wMChpoF4Ic3Bu004oRizyJVtkWYLlWSUAUoqfvV4oTjRk9CChDnISUWD/oihpTtKvclMWkLsCT0y
if1Po22RP5HhB8/vDptoXoScS0S9dR6lGLFF/XdOslZrcfA8wVLzx2aXJkMd2IvJMGJfsJslEgL4
gtieEaN8AlZm5y8iYOkyS0KLC0R2HTv9fRPaz5lYbft2NPOFKamBBNZu4yLUxe/NJhtgsvodoyGW
KCy1kWHuNKPEbLzuylZtWUz3XtNJMw/5pSy8BsgYvQwYfF+0xegppODn7VOX/yHxDWGIvtuS8OYb
OjPKQuIvVmtUiAkaM0hnuaqxW0OsVeYPczQzT6F3u77v5xe1bLhOUUloXqLDuKjHbhNFvb47RiKC
U8KIpo1DYlaHFzLsTkO+/mJhjugpeHBPwKZZSYLlIsHRQ4PDcTw+5TGAZ4mpJEVVhp96sWsb7IDm
0w8BHt7zVK9Ywk+3cCsQO9hhoqIwcIC50L8tgXsFktcJKWqZmHsiOvtbWxDJ3TeHD/3fqMirE0mN
PqJkDWvtMcmZw4bVEyZtOMJzcsn8Nqsr+WSOFzZh+zoPSP1qahfsTIrU2NCeVVqYkQW6GO6RCTOJ
liqdQCqIZwySVo7/9bA7J6wpNk24RWMsEnX4kbOQzLOTgMN9TePV2QTPJ4KX9lXW2TSxayhA8Gjx
rHda5ArySuWadlCOsjfwrulShxD612hCib8pnmGNLp/bJxqpAeOwgcJ5zjw4YAuq0OhEfVhJZCKM
nxgzwRmqYIM4CMC7BXRJ4Y8m1HRBwpZdCwc0+doGJiJ9xHcsDJHyOoNagYsClvtzb196h/tZVhmO
Q0uJhT9b+pGs23v+780lHSpvNkaX0w5rDTjWsoN7NDjuTfoevyVsj4Wj6ZU/Cd/kB4hRp3IJDlFN
nN0sH/O1eLy2TR8F0VU+JdeIaSVMDEUnzBYDT5sFvvKVzo3s58b5G4gViSJ2n/9OF/hBuihikpeS
B9cHzioJ1ytuQt2DYCVU68DmTQE7uILNSoX2GwLNnSuJ0BCSkxadlRExoESb1oCkLl0ttl4gUmFv
go/qnbKD5s4gY/Oxwh0HXnd3Uyg9jYjp2qqkdJUjCjjpCE+nuia8nlS25qBybw/ZVgwRPCMyPxmU
MUhh8bo/Gnf9HQP7wfCI+4npavQ5C/BapXrZtTZ6IdavVhi45oCE7GoIgq4BoTyfX+Zf92NKb3RR
d7LIwoI1CJY7cMCl4iTxJWrQQ7+3e/yMObb+Sx1rMbxzpfpefxQQeTKVzLNTQ4PBVqgvGEPJFWbS
Seps2KNsaj0pxxgwpHobSM7+qrvZGNfxOj1iH2C96p22RrmHxT755sFOjgIkpdK3AHiQyRN9Pn4m
qObT/NMu4AGW4HUjTcbXtbfw5hj8YX/rPGEsiBsJL3YrPzx9/Vi7eOicloWInce0YmWjV8TDsDQ6
T7pI9eGO3IK0N+0jzxGs/iNuxeWQNrwc/bA0T3hsdf+aYYBpv3GxmgoEDOs4NyvhnokZMTbRdh3A
62KzrtY81OZvMsDdIhCghO+/jWnpIgPAvcH+m5buJHEgJlz7bPRMTdmKXgojArBHRAdncHOOrdFB
3o/N3FKVFA/uSlQjUb7aVJscN/Y7w4CNbcJRhmF/dhvq1Zyd8ge7AbesF2YJjbur710L6xgMdl4n
6fr9takWQ78i4sJ58cbhb/TQ1t95cjZ+tURkU4czER8w7Ygh9hOJ0yC+X5hrgHYX6iyCCzBazCpO
13pq+U8J+aSLn8Hbkg/VJ8tI8Ax5nZPB4RBVWI8AKT5rPsLjZ4P8ZGY5t/HvL2evcvl4tiZMKJqu
KrlFjO7fM2aMknRvjcKBbh3hrDxk+wxKmgiblDmyE0YNEJjq4BxfvO1dG80V4AQ9aCQFg87QyRAR
D3seOkfqudAJZTWn8bBN6IImCEB1uNtw2SfVZIKZBcIpaFQDwTArm6jZL+jZVFICLgPDqUnJRqy7
Q26rxrZzfUCGTz/4eA4qX1VPta6FlzNtlFNVhB2fP/wxoVt4QhPTTCWUITfAJO6cwrznBUQW+1h4
7nAP6GbaowboYITzAbxwZ5L7MSFZntkw17RJp2QmdFL5W4Be8D2Okmm7CPFIF1/h1FTTmrGxV2TL
Nbg51O/l982rocwtcfBHhqyp2FdFd3cOODAn7I+FoMWl1uq6f7w/+UNJXM/Wg7Oz5Q8SC69+pcLP
QXexZL9g8NCG+yRETuvNTBXiOep+Nau3McsdfLuA7KU0B79ZMsYUKB3bDBX7gHXYHqFv+9B2nSqA
+pR87yqIgqLPkU19UXPu3ACfytE0VDr45ox2Qtes76M8jXqlgpUzB2MCSXGDGBZCtaHrOcg287kO
rh1avLYSqIgMJ6M2+t9AbOl+Nlar21yUUaLKQ2dVxEbFkI3yXjKG2LImsR4UFy39499yJPFRl5BV
YApXCD/jOPX2mFKbI5UpZneaoyaZB32CBVPNxcVZrCxr9VPYgAVgu1cVMy7TX+AVqEyq0b4ihhk9
hP+Bc6P1y9dUQbmLm6igInzjX0TUJpN5cXWDr/2c8ER3AYCLWSuXuthWTDHF2CoSLwdE3GcwuZeB
B3u5k3U/HzkBCr4oh2adBtJ3egLjmpLr+0sLVfVdoMpDgQDhLFe3wbqpBdfu92+QQsF9HDDI5JIq
hKQFgHBRCWVPKhZcbYKI4IIr97ZO73+Wh9sJehzmWlI0rmsMy9XWSp0ZBWdIPRyUFgHorifHeZ/w
al4UXT/5oPsU6pWQBXwZS35rBfgllDsG1sHcs420qdU40H3oHzyPUIKph64LHVh5I36LUZaN71vh
0JCXPLPfE/kOj4Vs3ALljdKv7fXpSkatMOEjrkEQ0d9JCroObLJ8QFwM5h1ALHAeBcAsnutRYdrq
tlcc6PtmuDN+EdndQv3MNq/uSni0EutfaH2FdUg595SC94LfyHyvbIYFrFjjBgWnVHThkQ4yb2PG
F9I/hTSTo1SXMlycJ1masDS+KlmZpnaJAv1g6QUhml3C4BUsmlSLEp/9urPFWonK7ifNlmtnhgM6
DjYciJiA9YsKNjwz3diyY4ULuRSHYcw0IAtsIhRAZwlzuA1YQjyJRHzjLBOBS8mUM8pGH8fwBsTH
xskuqhmfLI9lblIkKWK9ijBcPzzRAGfID8ft3ksT6wv8EfWwksF2ZmNBS+v7+UKenGCq8gp1/8kd
4KhlEga4BmmUI0o9hsnw2UAFrU51Q6C17YHVDQoPZWJYWrcDMvGDgIrvzGgN9v4vNhS7l2P33ktX
KrMNvHWBikq/9b0VIRfOcOoqccvOyiMOIGnYYsROCbk1sC0/Ry5Eljr3nlEIl+3rnvVofcebki6N
DbYSP5OFGezlAfXAHESAPY+6HSjpIV/qRfinHqu6436TEvkKWpUwodT/W+xLV3dmRoP89MG8JF/+
rxGt02OhOCpInUj8Y+fcn9S4Tj8nV5D5IdoSjAb2Jg5sqBj/5C3hBsP7ZnWtzyN+BIYcptbp5fXz
bvtSDpknPxWJaqzHQJfyt7FzeiaNe0NIOSP5EYpuCn0BFV2fimhINeqB3qLqlTfrtMEoabR9aw/L
B76cAjMoBJgRj9gGz+ddGs5muHagN1TeRrTeMKYgTPehb1ugg30nvBCr8aBDgrPiqsE0b0nNh/0P
iJnTAfbNTetaye5rCG/1JKzwytL5RI34dtxOrJH2LXB4pTAYMV+pBHyvfYYSz6mxvhajOY8XOL93
P9IpywbxJ4kfW+1TsByDzuBrVGSGV6oB7veH3+79BSMDTkBskuzMSqzMx/wk4FfCrIG6lmz+u8ZZ
WZCx+smsJptVszSkpr3SW8IRCpQRAs9UxW7e8WOpArPGEYqCDLWYhlwOvXPxGIZydM28nB/kGvnB
XF7MWePS3kZSJ8ikZrj12SeyKHgDCddbUoQz/Jkisuc/VqMcT0+3Afir+aM8JaD9BgBjFFGRgofj
00hJ2cZPnKAldKbwiBXMObDclQ055i0P/biHirvynQ7gV2LP+VaCHiK9Elq2P2fhMsms/agF5tFo
JWYtntSvU/ERS+xDQjWtsGNmRDSevbZ+pJjrf7Y2U0/DjRh+V8RSaCEkaCvpa9+rUmWUVjXZhlKZ
GS5Kgwqjg/tPjB2JKNCOVzuG0DW9lphp1j+NWLvuvrHnwETktyERRFTq83t4qSws5iJlMstU8OnN
KffEyOmQYvzqPYI4otg+jPQjm1WXIX9jCCV8mC8sHpv/JzfjVclRi9vE72b9gfAtTMPQHrikFcLA
1sjtvXzg0leV+lBjPpIxDL/owCUWPtogAwypA6KJN65Db0Dq+l50bERF8zWbfLPqvc+vkNkfAVBW
uYSSowChrTAtvAxCkO0njDKgSz8p7Pif1akiGpjz1K09Elotk6Ihwf1x/cQCYIiiaAowir+9+YSk
LwmonFMyf8XYqbJWwdA0mpZO7HRaaUH2R8Gqkv9k05QyMWTtuRSlEh6LE6gl0gg+y6ny6xw1HEVA
OOE0t3ffAKpIa8/KMavZm6uuZh9m3ue+1/e9Hg3wAHoRgfi61FEjnMZtSM3oK2QjaF/BKEmkcew8
gXsITFwvfcYZ82Pt2yFmL/6alwnbNuboHL0W91RRRhrkp5FmTFoyhgsGB2TInH6+xMe+rZieq00o
zkefO+ibdSrhjhssDa5tlsTTshl3TnIy0h2DmcxJvOW3R5M6ncKB4hwFjRhngYzlFcjoa3f4QbU6
n6k80kn+OPjGfCutMJsc5qwRW9gLIkk1SVpTRRfLolA6Fb3+zYidg/lkRANnImC2zPrXF+1G0VdK
LrB6k+fKFsfZRrjCwwyKRzkdQ68LDn6vHW1CPmId0+3YSFSxTplV9yt40xNE8feHZzJgw0IHArgT
NYgIJYzP8BoeKfPtRuuH45sB4/FuJj5C5TLaUmZnA30meBlKX0YilEHpzH+TiZf+ulyZ8/1Gw2Sc
kBlVetE85ionQareg+sfozfCGyuBF0N6cXp9lbsCrRYfyB9NZh7pdY55h47JN4UH355vDTUxc/BF
6EowM3txovLumqEQ/WIYJnGMVlOsSk4jmPcCyW5O9Jk+gTYdnvo50LhuJ4iHrt//05ILM4/bEi8P
c33+omgmzvHRQWHz986c3qgoU7umtMgMl7WiNr/iJnyAev/I84Py72r/KB04h4SLZHTDZTXjarQe
AKSr26/joZlPcS6q/q5ROYiL+d9lz8KyZd/wlU5lYDadPcTt2zjWUR9g8Q6+ek87hxAxbcRV2hK2
kUakbqPq3uX6T7+kpHoAtSAuhIhS2++vR1z4dlS5TshXYCE/FUGN8hTSb/WYUoOUg33xPI7awTFo
9cViiqhG3/HWNOx1K4UUcWSLqcOf7OVIMGqUvdjIO9Pw/h9b1qse96yo32JpUqOLCXd48QtPamp6
7xs3frQJZwChYQFkBK8tkCDWE5wYsHJwWi7btKOIUIBYurqceBp6X7rZknFYzlvT9bjG+wMH6K3m
KIGc8d6ngGjyltju+5CwSjxSnX/pPSk2RAMCakCN241Tc0ruuHZGpUtPITIbN+xoThVSipdH34Z1
QCe4ZSixbxW0/C0zX/xXeezBOwhPZDjfBMSpq1/HV8TrUgDcB15y60fkazwCyqaiM7BCzAHQBR+l
TzhlxXc4RyD39JV1ChMQszs97w3iZOvWcgdlmyV2ZOwX6jhLuQgPJx+uaaP5uPnvRoSlLiSxPRD4
sGN3OhhWnqXGd28HpouWcTLinWbze5R+px9Mzl06vgtZaLFo1PIS/MBDmICRTmoHZ3tyXTiJfggt
OL2RIeON155+y9AX6PbxJ1SqdJIn+ky1uCnHesxVVMYftAU8eWTInWLtD2b1AxiNwyUNhtFEG5RS
h7O1NDZcln41P+HlgQeMtL+g9YiIpGpxMGQKb3sy92iqmcmnYj2sUJIp1/co4fE96iMoSN8kKX4a
ePrQB7QQ4cKwuyoG9IDvhDyR/LtUUgvVbGdIQjiOt+nJFtyK/fMTH0KKb4Og01fj4cllq7wP7bGP
mXVcPjKUEuVYZ27EHyHmkKyA88mJpO8/tsQCftywrizbRz87orVFHLPUagt2Q7Ituug/lhAAazeT
t202bMXmFsUe2Ook7nOBN7WZYK8gGlsBgmL5dGPy6DsoCM1mRUXkN5UsxPqEIZWQ4rDvlOlQxfld
6NYjAglKfhM0rDW+1aVt9uQGvgk5d6+544x+mWzt6P2UNnQ2J9J4IQiENd3iBQNhPg+zigzcypS/
DNjMbLOa+fDR1h81d2wwUkVevDbbPeKV1YU4xF10aCA4Wn58ZjLg6IPYJ1RRR+muY/aIWkNzNP+x
gTcvKCL3zptj6QGqT+9j+a0SWZsQ8szf61A/3oI5PFJNRyTiS6mgsUnwkRl/V7HeA9sCx+T10UTy
y1be1WfNJHYSHQZeTavgzJpi3cpKaSHxjTGKPlaio566l0JmcaAdAUOtAY0Lq0hr1g3o2UP5SGbT
yb85nhtcL/fa9eVWF9tjtfECOUHiTbMriRKVteKme39vTvSRXPR5YAf11mbdc4AjOc6vJ8EMnSV7
92xjF1DhU8slJ2Uh6BV1TJOYFB7JuYq4dPi7V/yQYKW/Wu8Lh5Otm+vXxo1IBF3MzvUYjm2I1eze
sTQiy3Tz3oyRa/p98QfOIxH7v78KXiQeDLpffRLlXcRxP6hsjXEyQPlPGHEvj+PRbSwCcuGg+FSQ
bbjdnh786aaDrBd6tMEfwsxZiJK1gv5wafWKLPEu0o04RfzpmQdE+aXDv0974FpKlDpegJtUXq3j
TFZwEjuynhn0DU76dTUQk2lmoMS7Jd+srEHkKPqSNTsUsseiOUDG5daUXcZCHPbVbFqa6ejTv2cD
ABnicRx0UjaFlbPWuILcWpcEBx71TBP4njFGbb2Q9qEP+wkAVFW6RFOyMccecMD4J5WgU8TWkhub
U5Wuwc+kD/ibR/zWXbSIQizER41fLHwph2sje1EodoKvrdKL4lCD2xAmw7tNDbJjrd47d9wPlOyr
LtxfEYcHnFGWWgCOrWfxd8K61Y+yjJAHEa5i37qk/UrHkN4KrUJeLnp/Q2FRcUgGJGYuJVvP4Y6S
JFTyRoNBSBqcdEZZp+9GXsrMecHfW4uY6DJ+tZaUf6BB1j5/NbPgUqy6JA33mwhCjba21IxkNqS1
vxv/jCgRY305LUWB+RdCKp4BSnOTfCmzhX5dZUzz9/HbU84AA7ZMjc5716/k2Jv3JfkAFCCe7iMr
a3HDW3caITEyYkfte/DnvSCujm+F3Trp+tz2pyJqvOsC05/QPr8pmbCsI+RkpxZlL9XE2ijwzrhL
R9RKcdure0Wqzbd+023nhYxH7CwLeW5jkOEoycSGDtrRvLmgkenDs+iuDQ8pZu1U/4nhjXnUrc1i
dFoqdrJYrkjlx27OMYM7Bxj9E8HR1RxZsmgs9qbj9/WF0ndxSyRDk5/7iy+L6bviHnSUwaQI15dY
glHseiVk/Icnm0TrpMyVDn4O/HuLyxbFE0xkHje6Yi/GCqBV82FhKUM9pfLTeA9tg4rKyOGgCMDV
v7W41budPDN82FFuWUeWKg+Odj9T0JY3JuOG7Izg2e+B6eKZxKkuhRcUwqAg8J6vEy6Xq81Vlw/V
Cp4Zd+3OCSBwDOdoJbwjc+0nknKU/W0kkgbeqzCrZ48r5GvzttrWnyW+TJV+N79zvc09AkgsPKAX
/1pNOdRqdCnWWSMYPGQn7x3P2hahQYQFU+5KU0201/RymL3hgh4SQ8kWsAeKe2fLkJ+svn7RB2Ti
0aREsLfjwOw6F51fy4T0grPBfuYBzUr8ClwOktxCEkNXjngOt/c6STdRDHbB56ZydakWGtmjqPti
/PMBcj1xp1kOeUNg/DMY1KE8CWnwlr4Ia5+Tsqxe+P2RwfuoYseISjJkU0o+e3hKEpU13gQxhhYV
Gl9OBncnMb08t2XbzQSgPwbSmTOfU53ld8PfE5S+sWHT2aBMioYEMN3E3LopEL67oFQxqr4TM7xz
c1snbJSZkQe1laviogOqUZe6wwahXqCcJVwQremzlHiV8I3JYVWI4H4KDUNFaTcfnJvpSW6C/2bJ
8uuINXagiWUZkXhcZtV57ogAtcRBhsfeFljZxbb3uuAvWbnvCjmVXNrNdvwl0Ce3sIdpdotDLBa/
NWGzbtmk6bgvEnbGG0YYz6igJqfOoziW85YjOq8cNkkeiGq/vsuDHG2y+4UEwvpMB5o1OVd+cpaS
/eTsRVrNndkMW/n0eh6svdvSXLI0sYjQ4pkXGWV93SzgZyhCz+OvtTkgXhPkhFX67v2iKaKr09aa
9AZuWK+IzeiTE3h0J/j7mct0MsgwRieKTEV5q895jjZGjusQnLgEGHKIYGv0iniD0rM14ndixPcq
izhAgyAyNt3+iO1nTVUfWdCo/pHchHpZGshSF+z/zT4U9R5sp6owNknoMViFkUyg5xqVcxJCHYQM
+w4UMMco3y4JWgr34GQQn2IKxXYyYvaNuyjZxxJzTEtEn/6hJjgJI4jKL26s2dNBjSVcJmcu9qE3
Rh+iaojzsS/Cxww5cviYdB4LnVkD5th64wGBs7rrW8I0JerM7bSngVPfzD5aeqVOJQ+Ruo++fuH6
6s5RG79DmnSUK8XOGfb/aT69OzmoFkUCopvpM26sFmlZX5n5sI89nQlxHdyZL8KeC2JvHDZhjKQV
FpF1lYySWQs40H8g/XhkRguYOB3z4BOC3EVGGEfSHhNZ8laR6TiEErbGre05PEMdGgTLNxVUUtc1
QeQZKsAPSR2Yd66out0oXrTJBMWk5srE6u5M6tpF70qXhvnwSH1Grm257HGZwsHzR2ffaf9MDwyj
cO7QtYahUaQzdzRAbp/qtQHBnRlZnoBikom0MWTj2KDeJUPgtOP4OMpmmaaeZJrP2QSZ8LJ4FVM+
QbjNU36D8p4bxliKEgGR825PHkU8ZJ1lsY6t0pRB9bT2g4NOSr3COpIshMYjNOZOmGpst53aZaVh
pz68rFN7bjcRG5Zln65ehWAxUq3CF9eFqlniSf24EqhmbAYpisT8zrhFEc57h7kp/m3g7oT4T652
AhZ0sVNj6jwKdCAK/K23hPe4enIE+ebKk3iXq4iMgD+wXuBRUGdPrFwiq3gkeifVB3854ZSfjtW6
qZB5QiM7aCeZVwp0Xq3W/Kr+NJss9i34SOLMUJWDmtdvppvOkxR+BlXCj2Oh1PppdN/3nkhyC7+A
xjjeBJrwxQOg/Wy0uW1Ss1x4wWeZMx+N54BcRsEs2eqSReMmFBW00obzLFv1djZXeBNai8OpqlUZ
cF+tSSpMuWFfAdFcVe/S2SrFXDrEI7iptP4ZJs8t4cW2UTQ3hmGgXhkl8OnFk9akEkzKTtf7I98+
OBlTQduedxGL0obv0zWN+1T8YwkbIFpvLmYYxoK47JG4/td3b24GLWcmi595t+wRmC6RYKTWNMXf
DgQv135rGvM8qyDLJXQKrKSOYeSy7DoDAS4BFDYU7DapZksYBMDoe9CEPtvo7uIC0FERfsfOcdZ9
Ds0pidC9pqDxI/XlhP/8ApLZhwWnpcMkWHRkfL+605/c+uQr1U+ZOxm3TL76/RLyOrILvHFq2qum
wjYEEKreSB+fifqC+AXVMnJJZarf7BK1VnNMF83Y7WzZeiMQtRYahSgvKbINo20sIcFkz/9ilRwZ
V5UoWdayvmDe9mDLYNfzGLW31RqwdM3Ic6CfCCHhuz2Ai9Sui1uJBerWtsBNWObVqjMdrB0IQSfh
mcXV9s9J/NMUwMTKLpIHizFF3vS+SlVgzLta8P9ek4nai/QTCEkEua+jVhUsElsg7qqmEEwKpHhV
d4Or6DdSqYsHNFleq1FtFWKfCGYil/ibE5FZqCIBo1aFm2lD5pojNVbOukFiSdAKImw9FgBgGi5Z
bL7FhkRCmDJPe5PeASXoLrpzT9SsvUYnfZB75o1eVtbyP0H/ZyBFZaApKTo8Pkf+7a79636HlB3n
aVrjj/P30jPL6xpD6Eg79tFrDnVxzG6eh3eFGI7E4Ps6M7Ng27Vusyn40OD4SI4aM+6XUtleqduH
1SOHS91olgz8YrlnCtnQ0XM4pFgPuCF3rlOmNbczTI8Lyu2819G8dTAdqU/9PyF9EPse6Mpysj9Y
BmceC1GiFJdnlxgQ1eP+IgpFf93Mpt/N9PDNrjwDH8Hpfvizrvs34Ex293M7rHySVyuLQZkLfF57
wGoCXaLzc5UMi7cruhMjtk/PZCB1u1zHTRIyU7tmVNN/BZXpHrsvNTh+Irv08FgvQZcPSrVUacmZ
hL0wW35SciOe3o2W46fqpzZOe/S4vzcJtmpNlmJ05yZ7pLNH9pcFo5iqgqLVTDYw6DXR3UHurh58
r99Cvd7dBNWdA3uIwdznzoqxcLpQDcnQkvEPmuUY34zSpR19cbmU8vEzrClWLg2QIojXlFUMpM1M
R6x0zCe+FFOWQLgCmEsU3NExDSa+WKkS6VR2eQ3kp15H3/uXciwubbo3lq5E2kP0dgDFB5hQz8yd
FsAbMA5pUP8woH0PFI0YmC0xcQi3Yj28D/wpkXB9Qx0SReIckviQHLrbEwC4LzBTVTkCaBJ3yo6g
yhPWcY67I63RY04+UKFUQTTZQxhfcahGKQW3QLukgthYZbexfI91x2xNDex4W1P8JTJr1YoBBUSX
uZ1X+6ZoFCbN60Us8L6HX16CpLyHwdbSbfBL0dRyTLTaR2hquDjO6O2JpXSMTaOalMUcGjJzbbjm
3u1//llPxbFmxj7cy/N8NKlDTYDY7nocAD4rZlXkGeMEZLEBC9sJL5rE5RwnTYggvPW2KKLYR0wF
onn3Vsx0yQihbgSJv7/t261S3UlXmpIVP7rtg9Cex+LLo29h5Zaiia9221WX4nV9cBFJq57A/T59
3P4sKdzK9qdfnE+W5zmVlo4NCvAJ7Lz5sFp9DWy8QipPlgAtSQCw/UkNctfZs+gTbPsFlg/xtydA
XZwGpoIKXE69tXNVcJuoI8BzHayVzsSNnK8Xr3Ox5I2qFLiJsm9Zo+4Ht3OIk5B17xbN9KgJTG0J
Gs/VIBEVPRDQJhLZj2G69sNOZDggqNfFCacs7eqQKfhy5FRvcqeg46VCB35AKxOS4+hYX0H1CxJ2
Kht3q5FiLerhxfTod1j4CsfZ1nVtET+pOMH3MOXx6ZmkJMVECOtXP4MDvKZ1CA8tcUKMdQzRGkRf
1EzCWbY6vicezvZ9+QGETMmx2nMI8OYsjqNgg8IR+lBVc0FAtQF6mdG9tK3VgcG4URH9HZd9wZI2
anq9MlSeu8Ib6RAnmBy0Ofe5auUUIAF3ptQlfZA6UiWsSfRjbYEqsE4xz6qeRFTAeH4fYMrwMuC9
Q96oHnD7B/aTe72EiO4wTtdPIzw0oQSylRDZZNtj8XqXGCWYRVQasm7/373V/T72Jz574JCLAIE0
eBiYYRdSQ9yk/r5NRWgR7/bd4RCsjFSrUTe6no8uNe99hxvkpJ4DIiC4JHlfsWdKKdqflXNYH/5w
9mPNdkCLHlxYplztHXRtNYQuC/Kie3jOZzy/J7Ed7rpouACeD36T+DHZnwAohK2p51U3UnoDtMTt
lmCCMp1DHeEiJmDUkd47/4CKd4WZk8tWMnCGX7jEPekU1zdkAFs7qDpbzqrl51DcSTbO3M0jt21F
q2dFXkRt1FyUMsksbVhMSRD76WyutYa/Sx/LfN524TZBIJirHq6iOlhxzJAgbLH4G6q08v3J+UDx
E7kcSaHBvO0t0yWVdb0nf7QazVYODYE8GsBddT+3QNW7JczgBl/qSh5FvvGrJLOVkAab/JoQMoed
pqCfl9z8d5qedfafXtp+KcDVjw9nLF05vYTm5YtdEB/ZTp9KeeiftXMIrNUPCSW/1YuVsuMKKWyT
a6T99dXSgm+RGM/jauNIR40trQAZUAK2kAZNx/t53v0SVUcfP3DEETQPB+KSzGhmmFkQ2bg0D6mO
C1LN1w21YqAbP8qlTJgn3wf2AYOZdTheNEzlBAiDZjJWkqVhVr4884Wu2FSi/Jei3ZROwUov3Lpn
8T4ZU12Xl46mqsSHu+K5o1Ri72Tgcxl3MfF76R2RdJOMuAzdv1ggqwYghwAzNgcbsb0pxBS058Qy
xdhUPwUOkCwDVmgDLHfiHVpNUDC1FOzebtDw03cS7+GqhJCvts0esromrC/2wzvA4Y8+1CUB9t8s
bsG/cvKJeAUy7KzQbp2EMJxF1tnQ05GcxuRjyO8GKvbpo/mD1BsAJIEiMhi76GLXB/G2nHMdBgrq
qXZlz5tyfpm7928k17gz5xx4PCMMlwfsBO3hl16sv7D8YYdRKvC9tkolfhiFLtTI1sQhcmJXt4hq
noqKaDyJK0cGsBtPhl/d+fOSQFYozDckQ4zNnHF69TwcoPIjLKVLyLn1uRr5SAn65WPAt+T1Ut57
Of8V8yOcwG5OyzUFMaubjyiF5Od3rR6Z/L4ADsp0hayuBY7bkzwrXmvQZNqpQJ/wxSp4MX0Kxzoo
atEm8LrrK/dGAv0YBg6gUSF8VgC+WXfD1lAKoEbChUHe4EWYKtP1l6rdkKc51uDEwfZegEtrZCD9
OJ//3clMv0lP3WKFnDjpiyvTs3Y0fVV5hLyqcyjWeF6WzAvjgIUpLdWDRfKIXADtTnpPQBoMKgAT
GQOOV7uSe0NhsAz9QMuzwNPa96dUpJxL/msu44Tfc0CLo3BjC6BN7icp11yozpnCpSA7lmjgHujr
frwD1QheqtZNu30KMzqXRIUEIi6zpaAj+JG0cACWtRdo1Ve268UxfYNXOgwVtF0GpaQ+wu7GffCb
syBUe/ze91vyIe0gSKGwI6cme1CFDHOZAiekFCYy6XZkjan3NeYy5jayu8tnA8sofI1KYFabBX+R
qTStgZXFoWfmyKzQsEKwB1zr858NCRaLvyAmLDf8YZ0FASvurwmMVjF8w53TxzuU9wgNkaLxlLYv
6+ZjSaIZUXWEIi4pCMf5k+v6v183ouB3PaPBYu5SJ8rlpzTkXx5KDOk4Hi5sqi5spJYTUYtDgVw6
C7bWYCKSv2DHzfLMFS3Nvbad6CF4jbTy38eArMUYrUP8xh2/FbZs6n9rVjIvO1mpyXRVzc3iSYTZ
MGrlW4OId9nnHOksFu5qk6qI+by7tLNKli/oqw7/lEii7kY3lvo5BhXawTqNJ1qOT6RW0AKpRIqB
9/Txr4XzudsTUXUzFpTXPD68LqlGb0UQracDMtn/4y2p2fna+luoRHg78+6Hxj+31Hd/W5rz0HvC
vFz1k8oTJrkTDxRwQWMoIyiymAWsMVs3Fg780s+QWZpqvJS8VqVvG4GWWPtDA9kIU8V3oIOTplE7
47iUR5LDQmPE9jHlOISwk0qhEucvksOQqT4g1w0WqyV5ZFlxLMLOS5wraKbyJSBMoz0++VkIZER/
wLftidgSgTd5wLGetd+NwUddQqaxmMgAzG0RkyDSSwlh0yBDBxxzORs693rsLg5/IQ7kDF1TLzqU
4Cf+14+1E9CZe4FJhM5CXSUSvUGuY2t5lPfe0I48f5jJrpXaG2a8jsTHqbUTNa/sXivhJJ3zVcRF
rsOUNfTxJV7Salg+mJZbiaC7hefnYoGnwPPJ/Qaa/1WLWF6C4jqEAB1L4bge++hY63obOqX+jUPY
6eqhNJVJPZAH3qigV+a47uRpXl1U3IYT2LiVJ1konu71NRDjjWnJG7N5orS17hvFKUrFUtUoILuG
8ZUSDLVznZznebcsdnnLy5LU9XeLh+HlBFh04EzwOi3iIgIC6QB+dlx0vfxgRSKOJOASUlOV8UsV
5lp/70Pm0CGPMryvtdg2sFPoAig2SM3JHdWcbuGcFwCpMRKvdhYUPaITLkrsFuaWSGMXztJe2OFC
YGpgatzm8aFBIXrU+3SaoVL8PrrHGZX3GxFsGGsrOE/Yj3gbZxP0O8EZdueft8OAv03IaN0Qqd/e
sgmGaw8A0Vsj2peEh844IAU/Vcc785b79UBhhMSkyX0sbK5sOlnM7c4zyByJismh3a3J10J8NAXU
i7Bruw+elcryolpMixLl6v87wcfd+xaX7520n0q+AtwvbQaMXdszwd6GpW/fotMKM0Fm52ghEQgO
drB9xHN0QFj8ehdBTd3e04+29xl782k5zAWhMjulUViYCDC3U6nUiHYQvCNhtL6gwCmGb9w7MAHw
VECsbYLjW4fXjtiCW+ScGSbLAZqX67jYOCrWwl8NvIpaQDaUH0tCZlSSeqrNaaSyfvDZ1ktx+md/
bnxcwpaCyHsh0E/LdZihO+Ae4AHkzW5rhY/yPH0NjCyF1ck7cI+hJj7sDR3uBkwJD/pNG+4wkr0S
6LphfSh86L6mQmhSDqleZcIzIIWN0PfJDsWnQ6UWOjOUsCPahD1ZdT3+EQMRC5whNz2TgmNgVgiu
zUMkFtGKsZo5un/WMotVWxCaLsLimLuR44sS25oSBSJ3ThASl0xVlcjaqC+lNUTO81eYzY0NDGy8
+dl9DgNEYTr/mACqfxHpQBDYhK6iY/1pONpj4UH8VeQ9xCl/pAFWSJQR/ryx7Uh5dc81TaU3YvAb
RrLf7FNLRJcAjxNRAYv5t8GHX7X/kKX3+YJz611mGF4h/WCawrskY8ZUVM99VUNzmuhy8IqFbw7r
Oi4jvMX7hr+H7MjSOAz3/EQcJpcksYpAmHrPI7BEgnYOTlhFj5mo86xg9zChHuIaV1Ky2yHtJHhc
q2cS2YUNjhnrEzHXHtSfQfBji3CbxCJb5CtxAZz5Q9QVj+gPQmxigJVpHpqPCkW11o1lHcvoQgv9
uNJJ7xaGFN2W7qb7ChOeEqug6OEW4CsNkhgdzHsw7cElpqZZofHrzM6Cv+nSNaHgzMCp6edw7iDx
raRIjuUa5ht0cQPba/JfQLeAAOWtV8gYXrT2pJhvm3+OImV2w3wzQljHFZoJ0hj82cuE+nxe/6uh
4Or2aJcDItd3jpf5ciZ4vS2Cj+y2Ah5zVSKLX/neMGq8CsZNrabj3QJthcPovJchABqs+hW/p3uM
cc1K9jrdfegajjhZ2+sg0tMcbCjr2whG2So8Z9r2DO1eFQQddrbdFzXYtYG9tYk85cR8QNvo9MbH
eAnQ8nOQA5SlmJ6NahbuBrnS433X4yd27IhNQULzobQfreSuHSgAJxxRCb3fvxaIPtgjTVjX8ByZ
qdBTydxHHPNaPwblQxU26x83HgqXmOrBFZtTUozLfj2oqk6ik/qh0SqRZZVar0FVYHySKYxt5qJu
fz9IqpgJ5YT4xwrnxUAjQ3lXiASu7s1hrxsGlm9nYYDcBmHQDQWGoopB4XHOYS4X/R2jxBf25URk
DqhRPbxiCMEFCZGCWBl4TSmHXdGQAIYDyzienfiKIfsrZLNyrOTG913U42bVqxehWRxfce5vsTeP
yhUSlcqrG0NQlq7xkz+K3dwvK3oG3ZoP5yMLr/eoExXrA8wbLwrT4IYjEUoq++K9f7OenMZ6VXCg
M3Jq+bnpltMJ5IF9SieGIgHAbMnNB6BrfUPXyK03ZytdoVTx6iCXJeEox+/JTIdYU5Sr5APjg1Bk
EGWHmn7sjaKANlREQZj5cZNm9OskjxHJ56xTNuqXRHUlg2yj4mUlWinVdClGsT8pQYXZ8IiFY+pj
gEhEe24YVFtes8edkGz0Mxr/MHx0hi9uuppI8XyI6PCf/IdviNz7OoRTCddAOQCnJ7jL3p35XvM8
ZgFyAXw4Wr5IUxxzTB+KUP9ZlyrqhQKhAg7mXSb3fb3jKuqZkn/CYsfrgA2A7U6YGXXJNtftwmFi
RQzTeUA1UN1M8UxVWvIJTsZu4ajYBPp3sJRkaqjpRRbRJFQLBWvsfjvJQb1nlSKyTH3zJBY1Uio5
EZ+GVwCVeAnxRCRoq/mq2o6uPFfte19WblSKZadRkrJ7dzG8PREQH3laEsRrq7r1dfsexSUPcrz5
tH0s92FyJfvlnycHWm7JXF0+U0fhYmTzqZKQGTC4dKvlAsVkfsQ0rx1GKiCRXk2IgiyAdqqKpigP
T88ic3tKzsnm9WWBU0zTouSg96y8rvTR6s7ByvPO2TOD9dYKWtzolzQEuwOTIeocHsAqbMuUVdYG
UYdcGdNcJcWwTJDm4xzTvqEZLfh2V1Yq/8IfQasS7DHmnnohUbzjSnGqtslRuXo+S/HB5uCVzjDM
T42fuS+k9cMs+0kHDwl7XHM3k/jOcLhueUOILyVyzYY2sZ+MZ7m1uffDhPzC1KxRqKIiW2ce4g07
zGwl6hiEmwPzKBjoRbOH6CNWDNyRJ9ehbA20kh+hrYBUsBzQNT21uIaPnNzI5WxQ1Hiu7U3jHRvs
gGI=
`protect end_protected
