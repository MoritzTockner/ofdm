-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HOV/PDlPmyHmhtaA5FsQrkjSUWlTCUTpaDWWEd0TRBgY9AUQllwrYpigk9haEXWEOPFPTwCPYfGE
/aDSCyEPeJlcO5M+CHd4c+SqHl49sAd/N7OGLIztg3X9ezfcIZdcAtqeqNTv7uKqlWYF6lDoWXPl
GWVsvaUtkQeBhJtKCCYyBTMxrNzyk++IiuEA63qGJsj0Zbwl+NuiJ3gJ0abJww3ik3o7bJ+JctnG
0+qjHq5o0UJMIE8yXwZCntVApbWY8B15jZ+WvDqTzFEdaN1ImNpFgMkdfbgMVO36R9JdF+MK9Ml0
v4HkNrWpC8fWtS5EWUbrw1Oqr3s2bKsynM3fxA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
0FZku3hP0gb0ebRIsJ3AwX3CADyZprN+HfAJiJj06rIOhPS9QoOxEVQ0Yetb2+GJjMYfzM202SGm
kGyKfhN57OYtmsYwngG+M42J9PjZgo2GxPPqSW0KFa9zu8LVZTqeAN8dCFmJT9JH4cSJMQt/D2Ot
fhIuPmrScaP7FJ9fjBkyPIhRB8Vp6B3dm0+AlHFlW6A2U4HZou8gaMu5SWGNdcQ0eXoEVv2D/kLv
/XVkZECUtuN4dvsvAwvlRdhHP1hptEfUwWU467uCv8mUz0svAFN3sSYLucKn4cymRs4Eib53X/Ii
Nvu7Yhx8a9ewwEsPsM7wBmk5qC3p/IacSHl9e6SPHu3/IH0z2x+hF/8CfNhtK1eYSoXBadUZDqkC
egxyj4DMFk6JUkr6jZtxJMd4DZRQDyBWaN+u3BcRCgblQyYjtlCCyajjZavtpkwOc8ko/YcIGs7F
iwsd1WpIR/P39RdKDEpmN1pYqDfPolVlREGd6NUPH5pVUbWXuwnsE9JMnB36VVfENFJMpmmVbRLU
GK9O/CiEV7w9Pcc+TPji6DIRviV+ZynqEA9QSkeH6+kG+HnvIOYqrcA69WRlSv8PSS5dgU+ab0eI
0dBFcc2+h/EIrpPk2IPlNXBtnVDcKa0LCxKT7nZIr0FxB2qxrptAPhn5kqy0Xw5Drhtk378lZFi/
uD+n0ba1yrWxnSpR6hZN6Wbrg8yZHo5lsFs0w22nru9rHvfYqwZJYPuykFtHep6JZ4ecfuOMEOcD
/OQlkT9LtVGL+02u1HnMrqLeMO3Zu40b5900TvjTqNGIi7EE9ITfMOR50VE9DSZvQUmmJ/Ue5XbL
/aYBNJrvTeK7Ki6mCkRW93Q2zlG3NBSZbM+TXDLTltgAOTsh5y/cp9nTni/sgOkxCOvRB91Qmi6W
AsmE63g/l9MNPXszj7W2IhxrCFo+1QfS7WOZKa5cxqeXpgU09dAgGurD/tOH9BXo8CsMn99wvlRA
+9CFcIj/12UHVDVJqewwuLv81qYsHL8G6N+C5eXnvTuBe9qX5MyDzRk67ITJbXX5P7XbzPO56CV6
qDjAjgHhux096ziL0vVlKqBDbkww6Q3XyJ3Wu6CqtWriPEcQT1sqelGgS1JrnpEVpT18MTcCbMxV
32TDPk74T+LjGNNl5QAm+K3PrrmqVDGEgCgElVbZJu0uiSyFCOtVSoKnf+IQTRdklFtexgO6CcbL
yyvMA8+gdkkhLO7mMB/6VYacrP++KeEg3vAH3efA8LhW/GJxyiZDDL+9/Y9xyMo7Uw1AsawsWqYk
B3DHtITdctsnO+gHZ2aNo+fU+PrGYDheVAH3HjPXcvxG9i0dXLQf7DOjBfygGg0ZKrZ6oWj5vwGF
1IDURjHlR/MccAOJBChwe7qWoNpBkPCRHzBYIXMPTvzbcWK+svaRpAnC7/33NAeyTHKpFsJzdsHS
XRccjSUzbuS7OQ3MUgD9OSJc6za96YFJe9ejwzrDj4tSZIIWV2Yi+8sdPSpL5jDIGEEDyHRUEJhy
rrEGkANwcOHXYO1Qb5mOnKWfNgvbfbVVci2CrasNHoiDHZOqhbP69c9OY8EtQaMojcxUqofjFioM
XBFRVEkxQHEe+48Uw5unamYC52kXHrXygO4xM4q9CiF5cUcm3lp142PH6szizRmqWrhWhdONuOml
afquPuoHnC/0smvEiYBEJ2Gq1NZfVN4FcQ9l/7TXMeHuDjAAQ8Vg/8zM/W3d0+2RUXTQMGMMVagu
E99KsRnw7Ew9yNyG0etGpxdqtItRv1IgMPlfbIwyED7a8XqbwMz1i+nTXUDonFILDw+0D7c4bsHy
qfvCYFWtuKCztp1Yh/RzT2PSFdfbBROWRUOLUMmsVePlnjPCBnX3c3eywp9smZy0nOOVamULOkr/
/kuaKVXjevGn6xsqJCHP4SOu5UZLwHyqwT4zRntOmeNhX2wylPeQh/tcbLz1OJOlOWU/XBQxuSk0
+Nrkws1DvrZOPUsMccqRbYDO26NE8tNaj++RgPjMzrETgZX5uC9bty4M69s9hBm6Bj8PDTzUaqy5
7xmmDApXamqxTuBVAN8KD1yMFSUoG6+PNdZyloYpqFHVDDzfq6U6vcdhsr3Tykp4N3BXH+Dweh1E
Wtt0uB+j1JlTc8shHgJuaXPhxVhXOpgLyLxmOyJRM280XtuIGpjQiqkG87QRsiIrE/foZnEpLnQ3
6KqbjJgUAFd8HBA9r+9UQ7a97cdPW/GgIto3Lxg5vjVT/KYo0Fmkv5GrZxS6Nc0ruKPolI95fy4g
VQUGWpCnGgSLUhXLfq42KC2t41ofk3X4csjcGSxR/NbSXXaCIl3PgLYaiYoa315nHgD//YUii7Cl
Gdc+hfNZG0pSiNtIl3K5bUk4OUpdNwXwAqvYvIAZJjryZj39pmMqIqmvKMjmMRWN+S0IUHb+/5SZ
UO0YWMA2O9Kqw1kBIovZuKpsXgJyqnnUuMbXFrbGddECP5hMQ66fzBRkKMNnE+EygBDthtguQ7Ag
l13N5L0CGZOf8/bLpUWwQa9oQzUEsvpBVMLvv4CK6UDLSE7Xn8Tup4Ii5z7Q7sfDBXk71Iagxusb
RXhzKtpHADIhH/tF1vkjts+od9/RCAmw41ZgeqWs+dKb3ObaUepig+STiAMj/6jp2kG4U22zvkPb
6ClPF6lvRoaKznjwKDprOfxnPFfvT/r1aXml9xpnPbJxip7cLCZ/doe2OvgSpZ0v3g39+9A9GQoh
KiFG7dU5HFyKYpy3Ba0VNcDgOCq339L2HLugYIMSMqx0FgwqR4ZIztmjDWRmcqF+me1Rhm948gyw
8g4xXObX1Q4DZ1xD34kxep4A7pPBKK2nOSam8zaXWdlxeXcC+BUfVz07RbDoKZc4flvD2JeidIN/
RQ2Hr7Pyx/HiBFn+mfjAyX5cidXi0UX5sBtsIGXjR0TMnqaCnlykSHCtf+W/tA9sXXRvnIaAGeNv
ld+19jt7wX7v2stCLu/j3xA/ISEfQMcI+N0CgoXfwOSuH7kgD2QanBc4zl3DAsDW/Zhg3Jnsex/7
1kCuwE17U4Oa4TZ9yOQPjNOj0liwXUSD2Fd6gXOhBrqt1gUcfC5VXh0uMfusx/yJQexqcxCdAoCX
ca2n6Wr2PjfLJ4iopS84ExgBNtQ+qgo7nR+ji7asv+aVVBqYK2tpfYbPUc7sNRJAGRC+70u/mQwa
wcZRX1WQzcvaMVsUAtcEtfVlgwRl3sRGpC9a5s97ULte8H7Py0KWnvD++YsAlcvhj4EXx9VKwTov
leISo/XIV5jbih140GBAfyFqZt+JjCT2pRAkNhu1dwaEpZkt3Ewq+Of5tu4jf9IZuS/xn5AbgJuA
yqzXwSwYjukpzB5vDiQlYmSolSuHA4wPPzvvxsD9DMvUpvKGA0iKEMCt0jCXWHuBWT75uRGZdbJ+
xHyPSGct9sRCFBephmlNqPw+eSla3qL1z4tBnD4utN1Z33NxGL3DMsXn9luyr4vlUm5kd2nfkhyO
b9UDS8/oZ0/EI1KHtikRxLnlNnfPMqzyMcC3vcBC3/Deosh4Czd9SRce2Fe/Is1jfO3kZORAyBWB
aRpbOL3MLcfqJFPtLvloOzg5dY1jcJ9hjjeR1zkk9HmGNo1a5Piki5I9HZLRZKP/R/JX/Nnz5b89
77te8LJwKP8RV85b3GgRIok2H8MLNRtpVirPO5sf5OsTxhTTYWe/nRL22dtsoL8kMQxDmU1qiAE9
Wk/kkGzXHp7wlM9zMeFwEtlbEca+CkwuVE07bwb8zjtFhacc20ApGWMUz3TsHrX2nF1GVapcyvkx
1rOKT75dhVkrBnY3CrFQKUQUcldiGt1WgQOzrEyeK/jKfYiSjwA8MHXRXQm0+0YA8sm3CyHqx6zm
2LD3GN9JeqxH6qu8TPiXrgjgQWcSi+pEq14YJ5iGqSwdGRuWnpIPfObuYILSl3X/1LP8r554xFZw
FK4q9Bxz0NyoT2QY8eRgoJpyC4WpXyZJLhvFMZnz5zS0TeVgH0UM166erA5UK6nIyUVtl9kjbSns
piPSyVo4kqVUXdgLQLMqkG6N6d5qkg4tJneKx0MjVUHIEcbiO/LP7DqBwuGhnmCSc0SspAD6GDm5
8IwcMsu6lIv3vEI4rOV/NlSySPRiuQeWN20qqutcEDx0ZgBkueUdhbUmtlT3NBPPoTUmIcDBAiCO
tqI/PHxxzncgvbl/dDCs3en0d5VQ2ZsZvXd25frQsvvbrliKQUi4s7DSmytlPQq/u5ZW8l88tugj
IyWr/2kd23qf5gEsH7cUVhB7a0V6UMsVODh5hU6oHWfgGtjF/gV2Tfp3gemQCsnyKLsXbFGH5+1P
QQjw4gETdtMm2bbgg8AvV7Usb8rZhJLirEFUlWB68O77trprYOkjyz+BkHVO/zPEnNwCrd2elitX
RBIE2D8Q8+XM8U4gqlLKJtYHyqnrR5Je7YZng+W3/pQXprCWFg62jRUv+ampGJjijN+FE7BSebRv
m3iH+iV2utDE0D0AylTkqycKafuzy9tHiEWKtk0+NaU55BGDoYayG2Fn3n3+L9gh6u5XFhI2VgAV
qjIESK3LVhc3bA4kfX3Zatsnt6sPzn2YZChJvWvUhkh7kK30dOP804lflO+hXaHjRqGqFe8Q26M3
CRaTSsHBTbwUvY2bkQv3FURjZYlUcKz/nLI4rkNNH57Pj+8yl9zUTzXT85PjACvDRrQVy1CF5D8r
lLfq4rlwZSIMojbA3eafNbaJya5kh2EtJBvFtZ814c6afiCQM5EeZBsNcAo5c5x3AjFRvqcGZntl
gJ8yJx1OwEDBk8I9/OAX0bCAYCyKWJl8Eoc6dVk4wbzGXLRMCo1PBgKg9HfDjYKccf6NZ4JYPmAt
5ctBSlisrnkGkTHYeHIbjM5sW7B20e/TqhFjKHRRfrnEYVZ7h9bwulj359gt1whMcvAFZ8TOrQKn
2MViYWErFZktxEsmbfMVXz6+eJd7Q4O3KKb8ifzFPB8OZhX2UgwzfR3BQWGI/wGijJ1HoBo/IuP/
2XW9kLERxezU1h5+3JVKKeK+QBuGLqUL347OqoU1uZohvtOj6MIGOJu+FsDBthO04oYlnspHimBn
lLswqiNCEAIpFmXHAL/d2JiNpdFcDnsY6AapDDR1Vu4HcyEq7cFJYcVKbPeJd3PFdsyArU2XNWKj
kvoXqGbvYlB95bGL4iWJuu5AFov7Lu6af7UXREFZxv6ZGAKm6McgHxh0V5Yx71fS5Ev3zYBrb4Zk
8tqmvyjBRXm2P4ze1JNNq5tqXUOX07jHLZconVRf9lYgJ1QNhruP/tTjl0IEq/6X1oII1SSsLXS3
KZr/xOPxKzb+hXlz8PRB/6Rg8fHh9XLT/wdbB22FdSdY9QUBw7XvMR5aNyW6sv8rlRRWMobT0kTp
YryyvC55FosCdFSdr2vFfARk6U2kkkko7Lx2aNFoDxNzq4LqL2+IUiHk8duGRhaKfAtGkKUDIefr
EuSyc9UJwc3wtN9ctWFRhbZXnbFgxeq44DavWyvJLVetvt2S2Af65P4HYr5zX1hCv50v4Ddhkq39
SOtjxAalTYv827Bk90/mUVoFDjmSakCfmKbdLJowlZRMOywjvrhAVkj1tRPjXBETxBPYINJohsmx
zFDVjZeUz13hzQMBx21VjzkIJsrs7IXqrSuVeVA6MT9dRpN9v45MdprQ6HgemDNt5BmDoPKjIiuN
ERWjmRjaUoiGjUJYgQVMp0bbdRIK/MPOzpIdwFdMjWUHInIromj6oQ/RDsqe1QW1wFoxCktgX3Hb
qw/fshGTnROrkmArfrCBt0d0AVsreTC7y+ZHNKbgbHoHc9aCcyGEBBUa8U6EzenekyWu2DrvYThx
v1YKHsVkJIXvHo5VV+f8ROW5l+mpaSqwMYl0kstTEOnvNGFQ2G2hy5EQNyhcf+CH2APUlTkmn4cz
NB5/Z+u585yCu2DG4aUaqzqnqWfnpJncarJ6MTzHTOw9t+iHwnwUZrsMQw8LYRNNzdqEin4q6vac
z8Vtx3cJw8ePf4wvSg0dQ7iIOIh6ORQ+hwwttQ206slSQLJ4UNv482LUMTm7VATn0nct+D12GfLE
m7UIfYSw7g0OMY4KGNkcgU+SY6ntrLgYMHL3FA1wqiWR6ADi37wR96p7VPgXnfvwQZ/ydaJbcBHN
pIu/xz7dQwt0uhU2H5P6F0UcXuuviffKgKVuHGLKJ1dcbtCpgLfWfBacJ7PZcAvgvjfIye8xnmtQ
MQ/N1Z+X5Ff1vgoA8bojoombu2CFhOghTxII4CmD8EzBy6yhlUyZCn5r+r1PaFHWq6BUkmBuSgN0
4oWVnIeV0svAJ1ofBAPupFghz4wsy+0BR847qugB6R6ONBLSLKtUPdJ6hUnQs37AXnLXY1mZ88pu
QGCP+iYpdhrwqXA0b5N0RvF5x9QEvyKFwR+AGO5cFq2cBEaI+ODT1kCDenk775hrBkoj4S63LM1j
kfeCDqJwwGu7Y66RaJMH6XoITqiujMtLEsLBzVo8NNqMCKjNyWP3rtY5JUN8EcXuDdPQTidVSIFN
pFr1/1uToEyCNEQK3X+4akOelOm9EVai0IBoYJdxyySr+OVMKEEol5RDKb7uW5j97oBOt/lLZCM3
rEVKlCWlkx8Pu9MFkNailkMwxTuEVDKl2CGgF8szFziw6E8FXZ8wcce76YvFv4jN2/E7Mtk/h18E
dWUliGWz6nnkibZjg0cc/YEfdy0oiPHoWw+Q6ISqNcsO3Pb8I4OVI//1uQ4/c0i5qnaMolEvnOD3
coiLv4llM3J0neIbas+h7yzfmBIpItxBv8W0j3AppQqnMZ3FnrL7iF/299QP3X4GOKvBNrx3BzC0
Kn/9r9q6kqhsM4ZUdX9cAqMtz95LUt1lKzw7B/nxC4QKCKgbyET/bU5uM8+u+nMYMmHvQ/Fh8p+r
uXf5mKmoxvmMZ2xlnpzbHcHbFyDdbLaAMxJ+u+cE6tt0wh50VaRgov+pVJNWtz+CyuX14q6GyLbQ
OYvd1AcofkpsdsPhLKLepPMGOgsUfez9yjV9tRb4L1AylqWk
`protect end_protected
