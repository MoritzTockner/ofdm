-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WObCzryKQnOalt4AFjUjEYM+s72364mezA5wRxOSxtsz+aGgCWGpWHfeHdcDc+yy/6JxZjKzbImF
Z6ddvjMRp4KOcomJ7ZPhHXGLs9WZhswjkmqriRwEh/RaWAbyqZBC6/o8S41e8TH1e/aEGRqvJOBo
B/5ym9rd7rLjsYPF/n+Z+Bp/DAMGPFVdMB9Ffrm0bpyPg4b7MoIf9dc8MdAAagCX8M3HDlRCvacu
v7PvY8gaE7DHkDm5YbJWi1SV8dmXQvXc2cs01JvDRc0QeOUmQn1ltrhWNXQsFf3Zj3fLJoTEStI0
uAFfusomsT5R7Z2S0uyJlFmwUVq5mA4bLETTSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
oY7xKCJwjay3a77Gn97GHvC4CzPqOwK5bob9NAqeLL9Gp5tIU18sm9XPzMhAOsD0aj4IKWDLqteF
tTVC9iHcAtsBY7BiMAbiScM8eN4/uc6FmX189Sof1a4FNfQo6fRZ74u+oPpmBZkbqnCw6tCgDbUg
cVobHyHXNN7rIZdRoAA6l/dNxslnRZGW8VfrA55qK+An44j/WQBypQdh3sm1aAvQ7Wx5WgxwMSpu
uqb6p7RKv/gbILd1F5TshvQU3HWR8oOJNo4rhosEQ71rzL0mXpLobYu8vJrfjQwzEKJsdTN8jpui
UswuWRFRnBOtIacHLO8hyNfZxQbVldSntixm0VLmKKgRrjU8579BPwA1LBbeSRH5sbGSLDgF+NYS
uUHEfbDiIyga3oaIZavvgWTKPrb12G9dCMUvkokqCmRykyN5z8JkfUCQ5E5PcgsZ9TrxkCyRPzGW
Rw5mfyZbq+N4hkTQVDSFmfDyAkiy9vU/C2i7uCqHk8Z1JlC64/xLxFgMYHYKs+hg301CZxtlJ41J
L120OQWqC19E0SUXlCAHyyLpgoE1uYfeL7HQ/hE5cc5ISHSv06MPplj2Vo5W9iR2t1YI8dj2mMBB
ReAF4VDXWtu+juhX48040VHl+Iq0CRr/X/I/yMP7nZAgyoS5Yd8ydJq8U0eH3VAtyerzZBkbdexp
fPN0YYUZgUtltDinu0UTRrK0QEcpbSha+JmAAnBklysXrqFqIQ4DNkxLPVVy/HcvuTSWUzCe/IHL
i0VAsjqUfLEK/fVfpTzATzoDmODZ/ZHh/t+JmdxSSe8Isc1QSRrb/KPoQlncEygv0BsHfb8Le5MF
5cWsXs+GyXrnY+LELhofAQ8yqFE72qtGl6PCdc3UOrpzqY9IId/axd3e5tdMwlLqyYhYSL8ysIT8
91ndIbX16SLE6v2LEMa4sv6GmIEbIEWBHrRs5YIlxj0aAcy4ule0jRtX9HtUdFKWj9pKGtBo7koG
pQsOvhykIIIXIxxvL2OUD3R5cWBZjJXj8Z1DHoVMDnb5lULybvzNBHHyTLtFjHTF3Uu003tJ+Ij0
nKFSoEa1KPwCG8CHB6CcRynenZXmkrAIOZgVFcexQfYAVhqVzhUR2+DIispjX1M1QQAJX1xgrJLS
LJs4RS1gpyK9N5Kg+LxVkOVGMQY7I/aXR/B8ZbYlKCkKd3eOvmixEQhvTXwZGxrm0+K2Cj0qNoW+
ajEwBQEuGSW3XHhj3C627ffbO9EPF6nIOrGNKazT83kkRNZaY1P5GrsSCkz3Ubedog9uLXcYqh+A
2b55iGFjFTMWOkWncHLNVP1o3vrAMXKvecS5itJifRIuQho9tV5xbipddVv4N75f+qeZOeT3iRmO
lNR40p7xL9xES/vrbcvj89gnIyWQ6hWnwQjg48GHQJLgg0GqpsUckDP5mshBDjdvrckR3KkhAjqM
DBk8ROVMY4J+8Qc/HQcW5jDfpQnmiZoKVkCP1PsJw6y5yZtDWDRwOa56kitdWeYd+8tCCqHQ+ZJm
kW51NudVXJn4uT4QJsiubneJ6z4dCwmEUV/Fiiwc6qC80ffbu6wvLVa4K70nw7g2zU66FIkBW10P
UXmRuxP20rf3bvUkxrB6RNQZUPltDv6FjJvfyNu/SblaTF9udLNsy9bbMw2N6k+3jrGx/Izxgk1a
jg6imCDS+uV/ClN+KT7tCVhvUsSdAA7DyHDbA5HFx7oGfhDNm5x0bU0hdVhgagdXmfxENiz2XPtH
6ANlQgC6nEpncqY9USiR9HlYNDPvFL/hNAg0PXMxExcZ64s5CpkHo2tkD+3GNEH/QGsMRsUqKOKd
kLS/8SBspOBwGKY1miCMVgclb6Zgl7sK+cSevFmCevgClQCMC21Bod/vGG0+cLP2sDbtcDQc3Qj6
5yeYi4TJdSoAeGEEZsVEndjfwSQiXlUcL+chRic1UwnCGteFYTVAMazusNyWvzzHtsrxYhQvamda
PdesMH9wfjv6swwueDlYJW8NyVxi6MlyanEAYJPL7jEyJdbwd5iBuT/4hZ5e/v0/mAli6CVrSSnn
akArUcch1mcgxCVcb7Tc8H1NaVkYEQ35nj819N4kv4f/BCQuzgnc1P4ctBKaEEHE7fUD2H/bITaz
4kGjEeVvfF5uSZJCT8r2QTPK/mJJPwYhbsrFhcH+0b62WOWn0XnWJPqLknf8itmtxZG/nXfH9qMP
HBBlFhwbCMSwCwzG8ZVJqRuC8XF867ybBPM8uD5qQ5NKCXw6AVwm31W0H2Uam7H7mrjb2b4HDR8z
gQG9pCNSoDajJ4FAw5N14Jg/4auODXS3vzsUHPVOMjA6yjSpsQLWAuRfJVLg1LEjNegcMCaDSpjJ
L3pOAV5O7skBR/xBrIgFXaGEM0Bz2vaHybzxkEnr1srEGWqY0nyUabvFrOg6larUqywcDflWVQpT
zf84dfqDu8Bjvurv6Z8U6mQk86sWj4V6du5woGeErvDh53/fVOdoQRDpjCwx3WRYR15SFYdQHxnK
C4HkiCAzEjWxgUndOX+ABpl8FRzPf7yFYO3X3B1ttwqT1sijDiKawdIYif4siGZE4DjFfBEiGKWQ
Ic7eYvkza/NGqLF635JjE6znAQFvHZ10fpvwQ6ljTopQKGJRJtLDjUS5wfa2na0JsftgdYEPhOfH
tWsEqEZROl1nQwlBqxPX5uQf5Q5B/uobd1WPvh0LJ3WIwpfu1YzqRrBNXcDEEGSiwDKdKEb0sxzV
8fj5/KXHZzmt7xtHDP5UlC64Ym50oPb58KSK2ic3MJQRwiTh5zmMEp8Z0MDuWa0MKbpcIifmUSAZ
IrDo8Fq3FDRMNQqc6+u2OroH5QFiykzI1Xe1TkGKRySITXvgN8yfSyYsNrgCQh5Vzhh9kL4N3U8j
IamVOaEnXXYCdyFSO66sghuBtWdzIBKuEJdLFgKq+g2QrDojq0mkoyht6iGHcEGSfACE+DwPmT4R
dANGkwO8nmSYf57V9Y5EsuB3Kxbifh8s5vKYKDC5BPHM0sO4u4Ihv8Q19xfYi6qqLlbpozil3Z2Q
wUh+qGePfTq0u5rikPB1vx8BWrESsdHv9AJH/msAbi3xB/JtxFMcgwRZ93iN548p8ld5z7sCITNO
CL1r8vNAXCfpfleIdtLs1PCv1Sb+7x9N2JWUenHY7+7m/R9V9at+zIkBc6sG9ioXSdBDq1vt1URz
Ze0gXKXuF9FXZrdGCSxf+flr0rH3nPv2Kuhb8EALVhLc4Nnian6TElY6jhpUfC05XG85o6B346Oq
N/UGoaf0FruyciqRrvjVTHoNNFRpjF9riWeVWDkIFuu/rt/ZKl/vBkwy9AZO4NwAFtzgqvlKdTWE
6DI3z1GOejeYKnz/NeWhilFzvLXyJe5IUC38WhQ3+HXEpnsX65BrIb6w+BRs/ZwWa9ZUMSoMeZdG
H+VtkIwAUz94jGNs8SpZCOvWwPSL7SYiDeOiA2Gg05N+ytY1nDFIVBq7qYEXpPwqIBOf8pF/THNH
kAeg9zuHXGWF5NaCIZiL5u2nFHmdldTilkvt9LJNcXTqXBw+KbpbG9gNBFlOTd6Hhd9SZDsGOra5
PQy5b9O3b2Ll2XDUei7eHh9apPJ/U6ZsJxzcoCjXKCq/ifcrV/GTqE3QopetQMghhBXvn2HVzqvQ
SAAMuOKPjJi5E8RGjJm3Nk9LwyDTFah8KT+dZNF+qmWeZhVlYV7jiJyFmGLUifyUR77SnsVy5g7A
2LfajPw0dtTWl3lonUUviWGXZoHsgshHdccIVHd1BKBbTFmAvsQM8iEDTDyLGHATWXz/byoqMhrq
PonihxT9PBLyqrELguqGY/6vxaRmO/dagYfpVBhRORgTU9kxryilO0KMcVN6wcMrF6KHdq7uqwOx
xDWIVOxuSedvUGYdjV1Idg/qD/Q2gX+PLmo2ciABwKuPiJy9NXaF9afMTF72NobTHGVuJqmHwM2z
aFKuaNgu49ZrcolbY184zwouohKTg7W6+7rP8M/sG7YSbCeNlzvEUugHFtS7axP99ickBYIWQClq
qsYW8rpzX4t1LoKtVaOysmdWPqaQvfA/3FaSHnKkLK+iFwCF27bRkcDPO1ElkMg0Y2hzOtEUywSX
hPrms7htn6gNnVcZulsuWwB+QGtdPbcNu730VC9AUUZlOYyRAb8srl66y3RFt1N+LDGvrRT3O/sR
AypZ1TxxRv54A30uUtcVFEMooNrI5GUKa8+ZV6OVHPRG2ZC6pB4CpZ188LshTxb8467peTI9jG7n
Rvrn9pWSpiAyBJUraM6CFOOUpD9ymnfuz++j1cO7naLATX+j/IICgEuwIQMGIj/HyqzMSLDfGvNB
esvBoCz4OAPcHednTK1rSLkABW0tEeGQTZfJLpPOQd6BKuGXsJYdb3ybtoMtirOZRGMxynzdjkY4
vjKksbI+0lkVVHT/TnvAMdhdhDGFbdr+BP8Xvfw9MkXML1Wr1qeHZlDTJZ1QMnzoJUm2Ah7KgG2A
C0DcwIC2J/plGaeBAiDS4pQaiVEC/YuyhRcPHVGwxHKuKNk9IgN45EvRBEU+73Wo2hETcPW3FX5e
oO12fIxE8snPSt7pPb2HojqwAOAn3Wry9fWAK6OtPM2PIUxB1aBDGokmXEc8IlJ5Gr4wyyrop02j
XXNmWP0hO79TIVueRlVCtTydSneZIUArrZfm52K7gL7N2zImnfkPHGY7EEtVgjUbsKkk52zS9yG9
B1DLIa8DIlW9B4cE8YQ1lBh9mWxeY9skJiCqUTJEwum/nEyahNtJ7vNfUamhaJjul7f3xf1Jy3bC
swLkWntloaKeYWqrBIdK4x759kGwul1mADZBcn0/pUXK6kcLMDUo64AS1hF0jD+2PbFPnesTACUB
JOq1K6OW9ykYG54CLNsmCHzfxnQUIbjv+uE7i4XrBFzEumLdJH2Zpxd4PDYo+9uAOtObg5mG2TJa
AOMSncyGVKZjVZKxC87RnVxFW6u/5PW5oLY9q+logYAMcl+yk83UqpBMBg2XCj5zcMkqbd8J31T+
8Z6TsORmEPBoXvcMTZnc5E1XftjSvU9xZ539VDOfLZPq0S2fvjqJmGfi5rjp43sXVrlMIBZAGmL5
LBX/hSxaB7pugpcReJlYV4sE9BGsBF9dU+NHDnkUt7lP3TDrLyzG28X3fLTEuT3owXmtNHxamGD9
D820fdcwe0odsiehxcOK6LIA3tW9xt3ATpDwOOKe4B+bC7v1dPZXXcuBoc7hIwByxO2fD/MAbX7a
VDJ4Gc+m+im8KHxzafphEbtXCwLyGPhdGF6qzgRmt2VCKZMkpoFjDrD5MBUllkFFT7wYz5TPkbgn
wGhX97pnW56EQkVNRcle7t4Y7ojCjecXO2xwN61gYkOFkFbmmrmpLa3Rf+HilphB0KV2wegqnFOd
xQ+HYXACVV6DIksi60LBnWBJI85QkQIJM3DZ4XQhx0ip3bNTuTMIP7SwiH0i8vpnyzj+wGKrLOaz
SqeNEBiOF0HvY1JX6Ozhfc2yQiRVLpfdf3wMmJnR0nYfIoXflDduLiJDghE1xdW5WLhsPx7a5LHS
/b2GxFzbig1Vw6Xw8FnutmjfrBw042T+YQiHRqomiQ2oQD3Nj5Hx9y1XaZAIgNylFxXWy2Adp8Hy
m6jlTQ2B4vdeChkiVVT/C/9XdnJvguc+g62hx09C418GhUv8v2ib7oFSWQ+7ul/xCEXsJFwmrczX
VVGqvU+OPoqwcFDWMJXrRx7wZuXfzVCqyAJzMguSpxiabjcw044rUxMtCgt+x89PKkO3IeNIcXZP
XYQCi4IDLhMOhdzWCWwHe83EuJMOYyfe9pnpHx1lEEQQj088kEg1tBYVJPyTiJEKqUgCiRBVmKup
TasqX/9mvGzQcv5de+HFyqVAZVCoRDVcopHRKAiWsZxIyOY1NUELe8peepk6VU1sEq/7Tl8ayg3R
XKN0gdqJchvoT/8AXDLsM4wmUIzk1NvEmoI45ODcac8CTjpDdGnUdOP0DhdJCugcOkR+uZdS8HZl
7sVgp3RuBRmtYONihe6H6znzcHMxjm5OlW7U1jdw8s9iC+eR1nIiBct32f9OTispbR9siPigW5XI
cU2NAjbEYeyhIJqgB2cqGu5rgYx8UKpJqYI9APEAyCMzGU0fWVqKMzixjzVsiXw1t/1hZq4ayTx3
gRk1NI+lQK3HQypjvxsoFc8QL7VKwAIh3ZjG18fTIpT0xFeJPqlnT9l7jgAdt5TgE2ZH4BnnZ5Ea
a4qi/UpZmVHaXSDD7YZk2ZgoUBGbSZBDinzGIBdjWruuzcRYBAng5MdIduOToTuk7rU2A+JTXYEN
QSsUA/BBi0lpqBPanx1zLuwWMvhAW2JgWqBRpzn9i02CrsAjzh1+2uaZbG8ucC4loYUw+xF3XEiL
wRKioFAoQAWWSueRdtRBC3i96ylKWuFCrJLquVGvRSyExRmrX6G171cou+cX36B2z0emyWQ+4nYr
vmynSI/u+x5qSWuSSo9A2/JRmKe0UJJsYpQVjPDFESW6Lsa3bC5JIdEWqoG+FXmN6lhy6qSneXoA
FQH7CmtDCQ7+01J9xpbcjDPxlVhL+T5VSajo0YMElhvvtKTRfEiTRKMzH2LHOKKzKFDb2npMPKYk
gK/se9Rn3A6RxgoObHEJFSpu3+t0Z5R6BW/EBjWOmzXGhEIR0nDiH9W6vjC3F3/e0FTSjSPNinlw
nO9EL3KxShrpIH4EYE83u931sIdUcCXVlaYdyKkjbOH5OeVz+oOn9OySV7aemFNBVdAk07Uj6pKI
7bz/bPNjEWLd2vKDTbAIabbefp7DPVEUhsVE2mu5X4O7g2DEAwG0e6CoqHk164Yb8Ct5L6n1n/2W
60hZ7neTw8isotcRDsEQDQ4nrcM7s14kG/MY3nptawEjYFs3WzIMOJ2aG5w9hxTXCW1WvDuliY20
68BTM0zUT8vATxQa/zMsSkykl4y0VoPo2IZzBVly+URZuMILkWFUu/zqTU/x0w3D3/WvYqax+g69
fdDZSg6B4JawAvMm1cnwdZyx0ZsWN23IjGvQgdBc6pkBh05D61bUqWAE5Mtuy1/FuStJ+VToC7h9
6O1Ilh7maLXzEohlC0ZRztBlHokISg3uMEyd0joisLvXaRpzoOIwIkAUOxiMhzRSnwOfoOF9cHjD
Oit8H//Y3jDLNyH/aTUNhu9oT2+Ry0bXI83MOiY6JhtDr7J6eMz6wUi9J75KvZa2bRu9cX9WaxvY
gzqLyuLp6NtOkAeR4HgbMLAw1oRsJkWh82etFTwNj/MXK0wSKUthTEC1w0rQYxJyvNFr9s5lFJXh
X3xWpoTmJd2xe1n2M29XxUq2tWOUmEI2lIpJT6zelI+9MzoD19LMzd+JpAGzlXh19Q6SEyAfCYzN
FhwGvqxYsqusIcKtqWjEKkBndduS0ek045uWfdtY5fruT7ih9cE9ThEXZ7jjlEapHXlR/EIu8CK+
w/gZ2BOgrQwVoeMc/kRyGMGjo9f6FVzqOZINtPmLwo/G/QEhODuyQuy2UHx6Yj/nk2I0bpOv/ofn
IzeaH/a4FiOo9UqMiZi1lBuB4Kr/Ettnf0SvbkZMiYGoRj9avK6g9ixLmiGRxGGHtUJov7Qqq69j
+f7oV+J6nid0JFVzmMSKtWBuY72mXU76iL2v9GvwXeO9h4eHS6l132en8//GJyiuRXXYQ/YtBhH+
l4pnh72qYU7zvhgrpUtxj3hsSWZkAB5QRnIY4E001ApsWkO7jjg7Zf70ZNIYVZhQELbyWXcbUMlI
Srm0zCLpjlxw6EhDxAxg72LSWKqxeUmxgeXoK1R1a8m5jRSH5DTcau8HUzU2Hf2w+Qw/FeXCNpH1
o/8T/EX3pMCMrt4LKrrpBcW358NnGAVXbBW0TtnH2b5CG4WQsXcO3mVOOLNM7qYxkJ4r4Kh/PYK+
rC9WzcR4OYKSSWtS9Lv2puBrUZDQ5bY6gfr6ixa6dVpl8W5CBpUjvGAaSaf+3qFyGpa0Ub05iJdG
oo/TTmqzeXQmK907QjqZOH5GPvRh5n/MgvRyWolOu1X4pVekJln9TcUY1wokL/K/wFnqIIva/kVM
RapuXrZcWIsJbpT671l9bvlAmRU496enrZtfpecA4IJCPMpsZbPh3h5QEBQiGcniXb7JXqMDT0Wg
cM12LsWCp28Gux8yC/VhSeeBT3qX+KnoM953GQuHAZL5UmOpOPHybR21Xy0K4vX+2UAV4GIegICT
PgR69OCbAeVVpXXiazO2P0n3unw1NlIFMhyrKkzJ9kcIX0aHTpwZuwnw2oum7FBPg7sj2FnhHtz7
1ucE8lb3b+Pip9LBGLNQdQQcxAK+9NSQnhV+r5n4m3IjufWkuQsFrreJltnKQz3A8TIyPT8svFUz
+M3kKRf3byor3KKHEhPj2u7S75lXuPazmrQe7MKM2nzc0exYqxW7NP9MvYPo2BTzQu0a0eLdhhIq
ZgNqIx5RpH1rxFWMMGD1xN9G+nigtyM33bWnutIRqobJtEjbCvrvbxl5Lrno4teUQx7MjYoXKwdP
qkdqTf1LD4G3m5CtTmFn9PV5fKUgsbtelSXVG1JBMgPwpQNhHcJoYsQFKXHzmsG3Joii/m3M5ANc
/ruQX3mTaOjM9M3BF3bwEPkUA2HLwjr1ucS6AI9MEv7TLpIFtCPGW1ySyYCkZ9dqyd0OC8nrSWvT
fbhJpSF9SoKCwLxZ4uvEzxHToavRTCohz5/5k4rNaQlVaxrqOW2Obm5LYz8npYIsYZR7C9zlMS75
+ubQvmULh6MrK+8uhMRn5TwAJzbuNR0pq+uY2omPiD+UqIlsM0gB+eduqqc0iXeJWU/Q1CN3FrSq
6Ol7CnHtfvGWbFgRiP8pl1onSRpJisfansLPMi3LQcwozXYbCSayRhjmgNP3W8xbKAwDkZVdziHN
ydx4Aj1WDu4odFeABIRSUXXhDAtthkAMOTJWk0Rzm22y0q6GD3LhdRaWhmaCnNDL7/+O4yJLwiaz
Yzm6OwqqTZNkEwiQ4J2Huxl1MI3kTvDaG71VoQYxM+vM3ItKkSn8tCK5xg7088hUPHni9mBn1fSd
Jo8rTNseB1rfCgEhJlThu193JydLsuvGaVGAf4HqvBMxSABqHZ5SKez3wKckvFKBrG45OW1qs6BM
62/J2CuhWsF55voFtfvHNLC3Ly/iyHhup0Csh15B+B5HZX6+GEe1hFwcbHnPQehaa2jQlTiWFYNE
Zr0v8TaO5Zp+I0i7f5FLle1JJo2SOOFiOuNgtfiV1GgIT68HeeZ5lJ2ty2ReMqL9h//kVKxiV1YW
w287PKyURZGxv8VIaxIZrQq7EdrYjDSIAGAzqo8iVpxmoLgwEHfB5WVLDh69/IsWDV+EK84JESWj
KTmLXCHaE1rWpctMDFUZT3CG1vYpCNSuTWHlM/TGZIpJVoj+mkuqiXokoNFYJfZxNRbbBbluY6eo
Dj5JYXbIzXveLgF2R2zv3drLjmnfrknZfE2Ujq4BLWSH6chM0P+jYS/96rMGw0iJ2Iv75cdyKIy6
D4yEw0qnrg6kwE6luwEmF2lj2joT8a0QFCq4dwp+GPrR+pFLDs6CEqh9jMdplLNbC8LWjzyEPiZZ
rdiOJqujrHXDMc28WobBZl6rGEVbZ2wm8DYih4tu1deAaCXihho5tJN6EF7dLTEcRKH+0EIbPj1H
Pl71HUDg+BYLhuhqHchd2uQw9QZgoJt1Tk8agjr+1VHIlynCWAbh6pqzAOAApVX2nvn72WGOx2AL
5clakHiII3c8UBJVd/oFZweBcOKyz6j2r3FF5nOmbSOtoxO4hLeV685kFigDy9dS/C1QB5c66Wj4
Gvyqghn4/XGTK840n7zi5PB5r/UpmxiDXF7YPdOW3vor7fC8dbULBd2CmuW0dzsTtDL4uOW8BZWV
2PGdR0GNszbE0O8f3F5mZ+Iqo91Fn1hkBqBDl3bRKD6M3qynYFVuxwEOmQwiN08fXHuodu9fbwEJ
aaoy0eoOOinwzT1aoDxDDjCvBCuKHqXeJN3o77g6GkIwb+wOGoz5fYyhkrXBZ6P8DVUl7K64kOhO
4+15W+4xO5X9SawABUuA8gAw3R6I7txMVGAF17PTNOoO8XOHdY3HQkjMVlQvc7+4y6ar2Q2+/0IX
xF/soFWJwSPYERhzuddPCXRf0L00gihvfjl4aADfenCURQJDO9N4bxFYg7yAsJgAIH3QEZ2D8ZrG
6SatA/A+trNZzOkF4lhtJAzFzCnxHEYKjaJo5ytuvqnFGTf6MOdcmFtnB8DYGT0vnI+SA+ZR4bHW
igz669yZxFw8yNaqXbVmNks+hnt1OVpW7Cq30v3+vGmdJxXaoOlLkSKc1BYWzaNo33jqCvZMzqCO
7y40XFaOSeLcuTPndbXItc+VOyxs1UOKFU582u1wB9UqyZ49SakLcrZ5dTA607b4VgbQP5w2Teew
l6KNNjRpOiHblM2RZY8kKTXMXenxgYN/gLCRkuoff7hHFLauq1eQFx1Zi5QqT08J6e17gHeE6m9k
MMScfTCWlq0pGH76JqGaE4QCRyz7G8nROBCnb7j9SYMoEmbr2IvGyMHjrHudNDYFLuoQSjeJub3a
L3IwvboF6dbNR7madJai8KDRw44ki+RfGZ4hAWTJKW+RDxrolLceFhyJuGKtlQuG5gDoyrG1o+04
Le7Zcpm45stMcc98MtEsZPD9gTQyWsl70NTeh/ZoEM4gRc9h81IrPfSPvEKfo75Pd+4q1sEgPiQb
7ezl/nkyE9lkVSC7YSKhTaLOSxt1lSSFjunCtFifWmTqtOiYZ//OL7CHvhnMSFNe0Qdu8SERD1QE
LmlVVxhMblENk+ybe4NjlYS8BmrOMcYpr8+GAOHRv4M8AuFrDefuo4EwakiBwD2/OCdpdfmmeSVF
gpYi+q9Fl07AW9usIk7EFkkruo2ZzQL8RV7mlBxHVpWaD+sVuhQoTC9nSUrWyI1iKL9lNr3u0nLi
bu0uIsT7V2ce1pQQb75YEWvJGgU8yrgci92oXt9z5S0tS5WnIFLmR/UTSg66PSQTdMQrECjPQpwN
JqfRXv2E1Ujdc/dIfudNuTsgzAb09XO8Y8bMuvIwcY8je83qV3iQ3fqJgNrhrYyp4Gz5+8JgoSDQ
yDB0XLVTMU4uiyxdvLQtfFb7ua1idaTUA8dnEG1TAgTBmL/ey7Nar6B9KLPgxdmwT7h0XgRGDnJz
G3NrACsXkIyaqdYX4r+gSt229dJmqIhWgO0qUFH7ZmHsMy21t/vp257fJH2x9jWJkSzLVFzJFTLS
9JB5p4Vc/ltnMvfX+EYsP9JiH0MdnxxKzHcqKG01uLkgwbVq3N2kHcaEt9PNm5rEBvymbfWyLBdR
1vCfeyyaBbDbIbB8/CtXfuM1cyyQVxzGZqi2LVtvL3Bsoo3YiK7TEwwfg1iOoQIxdF4dPr97eM/6
RNAFxXZuBqYEwOEwA3HKc5vQHRAg5KNLV+FDwmt+Unmal2+zDrmuquNv+LESeBq2TLYVa+96PLtn
ZvOI+nBoARrAahtiLmBpVG7/yRgBvXU5Xon5d/OIU4IFP/Yhiw9z4btQ5IA8arqWhD30W80fRtTp
+aovt1UgtgjxZmKg0GnKcUSjIB6ncLMXapIZhzlyM7gjO95+F0VIX+Cj9rAMWjX+PWvLOL/oJoML
aHXViB4jrYjgifMU0wDW/5NK5Hnzkn+UPRWbF9V50rHupLnNwNgCrQmmWZU4dz3ek1hb6bGu5bf7
EwJE/eC4VFUybpXdO4RDzZ724K71gTDP/mh52CAG0/u4M7Fa986EBoo+B7x92jCMyzxTrm36Ya7Q
qKhhGXYzVq1Is2sF00Cyb42CaCko7WR4YeYB1b7bJQMJS2Q8OO4sgxIVkXRQovCuBAU2nZp/Oe3H
PERw/GJ/I/c0vH8JEYuSbfoLZuoNPgkdA+ouUO+V0eV8J1xbtfiMmRxLpO369oGXQh+9UDCdVOwK
/TBHXyQ7AC1Fwb7DNIRdCWpho3lsSObOe4P+kjbgIOnOna5PsGKNRJingd6f6OtUWudKxY7cSVum
x3SyIs31ffkLMdxRTkf3ioz/PTI0PlDpf8QY9XLDaivOm0XVnZfiN6a5jShnYbYtmz9DZI3vRWYW
arpS1r97MHBw9URb63K8bhT9lzlktRObv21M4mxTaPDnkxyDL91bhvIf4YhgFxt1lAiAcFkfkXK+
WHXWEkOTDwdA2s+MBN4q30Tc+y5dIKwp7zn/D975xPnVIU4AVuAJo5LL96v3jnO/CHQEqjLdJX5s
yp2yVM6qzwzOB1MjA3utLB9v078hHuVdDYczz1lRacdq7YTDf0ABjxO5HKpQg1u/QvVbEz5MSbNP
m8W5J4bgACj0z+xfZGEx9z+AJi+Ql2BRfRM3AvlGEA60+PPSLjQssLBF8LmqKt1f8uUjdY1onIcH
h6fAjtYJt3GIB93aH98SQJ6Bm9X2Szl+qsF41hGyDcGFmKjF2rSDvP3/HooZNu2xE4vCOrLXF8FH
j6dnHBhKRfe6NcaaU0qiBP58uYs7aYb+fKmwaHnRBCA3WuOAdGvEvcl+JctedFpZEXsOLDY6yGHm
+DlEyCZJmEaMgC47emiU2smIEeRX8p7GRFUV30rxQ5Z5wPC9ptmy07r1jVgYWScdU6rXUeIjztBa
GYgpslDx7qUz02kiHbNc7b9Ajhf8UM85DvkgEp92loqgxlO0z/i1q03PyfDktOrcWDpOa6PHPaxC
sNalfdom+oafp9mA/HpKNHHMwiCoHglYklEmBqdAP+wLqEhq4o8oYSiw2EX+e3qBj94GFPKOJiWM
MgPKIoVGbgCvnKqUv9ABPlf9Pvwmf6n2WPnopbky04rYOL3NaORacZA6enlA+EV+1YEntmRrKCqV
o7+QcKdJRW67q14RVdlNf2u3ERDG5ugPmvMr/pK2wA+5+nCGqoHxExHjF4Ze2jtT/fZTO60+gzpj
YhfwnexWaY5zqpPWkIO83xaGe2Q/++Qk3q2HKjgkIr7hJoMfR9Afqs3q9LCYYBrve4Zg+pQZr8LZ
1uh1rxYgRoqeA35LgRa9Y8/qgX5Y0Ay+W8hDnh/3X6ikZteET2X/DbtZg0W4NE0UoXbH7sI7fThR
kZAznwHfOmQaQ042JQVuLKycwacZeA2f9kPTDF2O2AP1cnH4iKDR6UbFE4ZWkBwzo3EEC479ZreF
1EGfJNYuDMijvInbLSIE403SBx98FI5GiUH73/v71fiMTLki+4gZv862FuYTdd8Dp/pRY36kQdYm
0720onNY2SeNxhLnUVU72Pq2DtgFGZXqs/cTUI9IZZiuRupcWOK9aMKbYnq3zuutojtT/yuQNlzc
WpZCcpm45SLs4nXB24SvJ/lfZjiIsOJxbiqfEmyoTFdawKOzpYp+pmtm5SDxf1zr4SYiC3rRC+/P
kRsttB56IR8f6tdSlEOSTna/s6xpTC6dkfKYlO/VjBfna2G3HVdhgbbFfeWZa9V59I5eA3Wp9bhI
DDPfFC1woyi/uKmP1wXnrzJGvITvTUmHRpCbsVOtCNEKBmOGKxlg5luZZoyQhEyekbzbuyJ3bIw9
BRQ1NgDSGhx16yTkmhvE7Pcyrecszsm1Z/Y2JvnZk9gj/a/eKWMi61vcqlEaal9VI6YLcsrskXHh
+5RLfPLVIgSACru9WhPt2j6L83LosKlTyzsKWzD5Lx0BgLyIqWtQ5O+6trOjws3T9Ifvt0HGqj9y
N2igCEAjpcsYu5G97sFGx1jeXrRyYoCbs/PDweZxJPqzLzpXOb9AqBKXDElu7cHCOq6ekHMRCrJP
WhADJUFeBcOQ2banFBcqkMIK+E9p9Jii3PBSQyME5Z22pOi4jaSOu2gtUPOx1IfRhhSKgRfddUcY
Yst9RUbsIqGq21f72PBwPUEx9bgp9aWMlJ4wlo5RqQpp9lV0txFcMGUmBjhyB3aWuXD4FdR3R9UR
kiVgdPE06Xp+m4uixKW3HFGg/nF1Gz28BlV9eRKtB4H51GJUio9MWct0iiIWmzE5hWuA/qFqasdL
FHy39j2JD7Vj9+zhKDzldYd8TuCxAicPps3kKuDxo0bmZBb3xMvCPSq+Dct7XmwtaiQGhpEULi3N
MoLdT/Gr6VQAg6IySSwpoZMfv4AHnr7hoWqmUGpi9Vnq0RDzmzbvtlnDCuo5ubJQzUBphb8s8wRk
M3HLs75LEF9WVq3rDjn1Eps2fcpvf1ICAS9JEvDHkaNM/TBBhy0v/deshtW2htOksiwF6l2gcyJM
KvHNYt5fCYEGehcIUFPLmmNdgvFbbZfECtGG2Uo8HhjUQrrVHUhjQ5VdPHpoqbc8YIbzsqXDJRly
bZYEA9+y1S3WkjuXC8YRIr+vSLKTGBJq94cwhCRBp9fXOm0fSpPZf9/ZORdyXFteAJcyLcaStd7E
8x7TR0bMTQb6CE/S7nMa5aSdWzhcT4MOerOFBsCFu3GPuLOvIVcZZdzObBbiaqzuE1ji/7t5gbI/
olBowdHOtt9g//o36TJbvDozpm2fOm6rwqoWPX4nrzsgDlwAzKb/WIdP08QB6A5rIpeMMhYnHIrP
Py+g+r0WX52rW7iPya8lbhtIgci3B2ha0TnMCqZKcvuUbVHK8ra+1fXtTH5518+CwojuvAluGcdt
ISBWx9nw7XYuW0Amo8WXIwrcSKf1MA4uUuNF90712/HorLL7XzzqP1yPvolYFb1OfjPuuR9iuz7h
u37y0bEPteZq8y155X41zO04sa2y4xLvv4MWrXnoQLTgo7Zl6Ax7/hXWD6/Wp4UbqjqX6q06eYx0
ScxILrb9axJ14/DXat6+FzIqeBM9uCLH6rtkG300T4JyUMdhzxihDMXKgHxmAgbsKGKq/0n+/9Fu
E+rBfFRQLFupfQ4AYTOx8keN3Wv6C6a8ngi3ed6W//PR1BJGiPutVB+BrqczzAIDkA5AsaHYuQg6
u+aUEZIF38KleSDcCpKsFto7CU8PpQV+t9kuiGFv5aA4znU+IwnYRUe4my6zbLofXLHGVCGp/IqW
o0Vr85ub6xoM+aUC43FaNkSL5WS6dadzMFYgeELAGXRoYhvqEzULKM3yoOUppCx61h49dK2Pk/cj
Q/+yligZ4gnA3Mt1qC53LVG6KQPf1jbtlHpjXiwpxKi+sT/0i5lqOQzqOszlfQKVj5zxwEmR8qfO
A7aLyFHlFllItma9L9o5OazbdlQL/1ll2qoze/lk/RUmfRpOWepsyWmivGZOCOF20w7Qsvkjlwwj
b3ZBMzuNoiH3KO1olCW5Anm97nMP2mUJzpD/wW+H5MUIDsc6q+NqOjUe+RtXv/vODWLRVA6sZX73
ciFcJwmfv28i97VDu0HfzBp/9tO571b8tODgjxeKsmg25KPiYG9xHKfuALqhqfaUrjP9dGQgTXBk
enV3SYfuQKcubIOUYLcyafoozD4ZENWp5C2HCJoZ59L8d4caOe5A9019jjpKI1NXkBh5kYIn/Exb
gy9HetECF3bCUqqChjGO6T0KbqzWJC6UtiGbtNV4S6EZ1XN0tUClrQqGNiQ0M23CKUjAZmhySYbK
wGx1QPVWSifBCAum3EXXzgbzVYNBrQEAuiosgj9Md/sGfWxzDYXq4v2LYRigMTyylBn6mUWzOUYh
h6LB4YOIzK66mcdIX6iYGdMBcsoFf/NLDQlI/pRIJtMTpn3t/6TQeOdOBToGA3GVf8x6uk1ptLyo
nS0Ebn5+GFDpo7vkF62dT5vIv6fd+SOp4+++PRXA8I/umIZ1pMG1+dxLivm0wjirJt3AH1xsq4Wm
pHGTVRWFxjYdZ9aCFBLOw2rDhiAJkPIfsGL1YugbilHMKSjOrvEwbY0INZZLkLf6KuPRT2JeZe8c
DnV9uZzrBqLi6tfqhP3FBOptwtA/yuBpY7PgynHmHoDgCDmlbvR4JXhFXmQ3b68OMxbQ/ODsEYQT
UFflXbivBz2ZuHy1nMzQb0q9omXCcLt1f3sBOyjqRaFR/+hsgPMurWHqm6hfhRwbCGc+kcc5mSD9
sByL6HuO1Onav5soMOFY2Ber2z32pXrBMJH855wXQFWzBNLDIi+f3emw9K4YdaNUVOZpo35wmDmi
MAQ7zHkta80mmVDtTYst0iP32F8uubHvRePElzEvp4WmhDlRro6u88VqIAlNvRJ6RGvDQ1pLCISW
cXnlBn02+BcwPwFgbEkV51IEJecof/BcncVV7mFGUQWIhn87f8Cbonn9rKHZ9Bb1ErdkGuxIRWlA
WeEj7yJ7qXe0ZFoib9sMP8haCN30VF8FjWbPZ+kUYdD/Zn0j/zvM2d2Zp5jxhyA1Eg5iJJIzFHAr
qLuU1eFmHsdqeR6UT6s4bTElCslAiJ3T46okIKCJ1Y99hzJVvRUaNYNtOnWq0AjEIbbPw1YBD0+4
U4fTJexeUjT/gN0kzWMRELfTg5TGAfy8fIEhSTNadcq/iKqwNjXFlJ0mdR+ityWzYynsJCfy/ZRy
6MMA2hwxCfAoOlptv9NWDxMKwwCoGJcevo3INc67za9L8yeXegwf4nbjOyZLD0fimasDviXW77AX
AXkogyfoUQVOnCfcejeemMZLwm/gsVVEHic+5Lo21w==
`protect end_protected
