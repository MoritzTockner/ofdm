-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
m5WSyyoiOQugO7rDTde+BhOVpAA8HisaozuhH4vU6vu3fnTWcKAYbYDvxNMfOt0UTKeW/AYFhski
N3IKfUnbSnMGdLYbrH0W+wzNbB7QrS10qBArzaoRYUo62kmNoW46gVMRYYP8bmowHHKQ5aRVvUr+
WBeC7Hug8UJnC7SaaT98lKFmMXgLRhbwj4BP0RIED4Tot5x3mXW3iAs5bHoGJHBnsdVWibc2irh0
qrEOdPxN4IQ4qOIRZwSC0xAiNQ0PrN1fi2Ss4FWuOUr8RRXDxECAK6ES3hfwJu+Jgh3QIUT1myW7
Gq5QW5CioOHXP/Loy98khE5d4NV3RM+gSUWhxg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
PMIzeiT2U59Fi6TdqczCUuMONhCcrwV9QIFjPArofx7UwpTxE7G4Sh76CyUePEP+crhUwxM3RePS
3ZofA0yrKUH2VFtg7L4hyUBW7vsMHwVDOxD4ZI6hJMvYgjkJ+vLMmc7Z6xecA7A1VrEVZrj34JwM
5fdf5XuT+KOUoAHftId8SLrAyuiCZrfJUJpZJ+sssU6YwKZTV7Mg3asGASblaoboUCT6TpOIOm58
U439Pz1LyhMOpyisq0wSXWrQMXjkd0dnvRC1eumEA7vhWFV/fgroVwoqb+Hyl307LD+lAIH9o4vC
rEIqW/GT71Dq4qawSc8f/BjiSwbELxMTjIr62+HIA5kuLFecFZ2OMgwn+/na9cJ/952+SbUoTf0P
o0QypeEaZAO4957nvSyXieyA8gze6my1GvI9//qmd3XdcDHLSSgxFcBgEYaUToFLywVhgm0CtXnQ
Cv+4DO8iZpsz9ZvaePTVUbVW+7anejBFjsDxsOjT02auLuYBig1q4IinPqMAaBj3hSaa8YhKut+0
w7YEMEWUQ0sz/6jADir42ugoglqXfEUcJryuRqKojcDInkaUuvfbaKNYgn43sQRF2xXNYEmUbb67
aPUJm2rK59gbPi3hXTVs10PsBI7Y7dmBqjKoG4fTQFYuCYkjSALoY8obI7AUZ0gwWVUzRjhSHfgN
BgjKFO/ETZxK7FV39UFuRkVW8XtCTnLDJCvvqmsx3q1tQ/3UCJTnrcsWay6tpcAPWHqaoDiQ+TfS
PqPjkUi73/U1RT1MzKZwQBLBVMqqAcLW9HFQF4k8VT8jByVE6wyrlzVD4nHzDacDnOeFiRBtEUxO
SXHL3LbVXZ1EHIIhu3RMde7+2to8dVjOzEvltvulMtKWoSFlJDdllD+we77mzj1ktld50W7V9lAO
qrbQ8/A07MmZBddB3ffBvTOhERTB4PyLlohH4egfWL5c4Afmy1/P8F+SNKMgsAtrOcLYMKOpD6Dn
6PkvwaFDNnpcL5I3tPPhi4MhB9RxxWZLkecC2xOGWGWkwmHkN80XiR4Ssl5f/jwOQ4sqW8tdgIDM
f5BcmMK0KmDt0E+7dOSE92E4RkbHR4ualVPPDYWUhOZZWKPn8uebirj2invyAF9QVQxHDKhDZnWH
ar3QbdZE6qJfAXvAR6bNrRIvPJpqwBacLx13RuIUS+IPRVRBDkEeNuXAB4G2gxtZxKR6GhMQXy0b
WHuemuRHHK4NuwbkkZOwvj15dUp0o+LhRkvBo4EkOSnkdZBpnJvogODV5xc8v2tu2ntvxVflZMb2
UmAGym20DnEVBhmHz+xdgxoiNf2i191xmgs7pgqzsFrVFDzaMR4lpJ5zMoi1O6oCgkZlxYN3Ll4s
FgqADFNVKWs8GvcIwDE2bfXjapD3qJ5U2b77zlcvw928lQ5F4Hy5UbLdr+uMSjXX0AaMFplOC+Uh
oEw2TziyFL3HI0qwiFfILfPSmu1xVmsGlGKghU0URA+PEB2yVA1iV0GggPzxFgXggVYYBezD8QOG
xVPPT/cU7xT7eujAwk+oVl1pFIJRe+8KSR4IL5sHJ4w4HVOxm1EYeNcjP+AOh4LdccocSUU4zctP
GUKkNBIVwa+4Z0svXY7iTdndVF9DSdJno1Yt/Rz3XIqxhFl/g7hNgS4oz9+F6ZqkGZ1bFIdfal8K
96SYR4ynBlveDVY7s2jLCTtJoIbkCEJVBiSI4tLJGxV4J28tPtKag6GDyuxHNWqrchcVqEAfZYzr
wq2raJAsvB0SCA8qf17C6rHL0vAy+CGefoP+V8yXDJbPxzyzTmokUhOPJTrzB72zVf9yOR7adkyE
vWPCxb4c3UmoXu7yTQj18hHvcjzTuz81MPMDXM+HRv46rKRQGMHDpVBw4cIvesdURLa/ad+lnghS
qKdig2WGIy2nYeAkAAgebJAU0Ux3GSwBnhS67NVyOi/FI7KM0QE6LClfsTm8uKNge9yUNf3/rXFp
Ezr5hSiPCkpbz1Nnq0rCrPVlD/+o4n5XGb6HPApLoNu86ZFATDiRkHYJHn8Hh0m+UBy+uW3deHbL
EKuh59p9t7ocsNXS1FOc2EnOrpkxvPlq6LR2EfDw8vB0Ma1CZusIx4Ud90mM9oa8ltgs4F8S4t6h
DP+fSI+filv6zymss6l+6MT2L9j69DULZf0UYJGOSY4pSTr0nQQ4KvBJ2hG45F9uV6YHyTogiB5d
7M+O3TcOpU3oywJkoJ66AFrDAUGc7RmRi6GhAHgi1UFxY3RmyM18qCISfj9ESqIOqqZ2oYy8GeeS
/klU9i1TPxM8/ogF9zO3vy44Y4awxvnnjBV3LnAKfgAK008jddAMkr4qA5OT8lAj+e5ZUU9x5hP6
cxp1+/z8pc2Za9zO4yonMk3a1CgznBY2kUkSu5mPd82DN5SHdqS8PDmvHBYbcywOr/d5A7CGXigO
1EEMI3ZthLc1lPMdHHVpfGc+deRagZNOB3rKLtMunBkwEt9TP5KR6GhKs0yffA/++LGC0yXm69D7
s14TZONkOcThFY1S+bRcfcgiB6jNpOoRrUTSLz14Z6WDP9+RAcNqTciYLdH3vQXxLowJMb9eWdqC
VpyJl2q8+obfTUo0bovzyi8CxK+dgozBVAszVhhi5rwHMP6r8gFUAaXDUKQiahgoA81dUJ0CEm9X
07ARVQm7M3bHgPfeFhLFRd/aBPWIW021ZOdIFFqad3oQWDsZ3P3VRkF0h9uVi1XEZbPuvEIsNeJd
tskS69pZVV7HMV4W6bYY9qD8oHEbhEluBcxjJGrL9mYjhFady/nWaW/BGrKM7rbAzI+nUILSH0HZ
mgrGxP1ahn3CBJuglM8bYCDfebdi4RzWEUC45352lLud9Pd7EN8GJpIJMu2IJrQ32NNcsRRt8igC
5+7LO7o47evVw0q2Xcj/dYPQEPNqJftk2yAJUpQLyOBBhkalkw/cSZAhQr8EShx//PVnDfPVbYo4
yFnJ8O3jkIBJj+WCP0HUT9R8k2v1nx52PsqxCxAjo0NrAcTe3vmz5yK4rV+1sO5LAAyDYWypV5jL
EQonaKVAthPwtRdvXAwTvNawtTB1u8Dz/2hyqhDtIjl1FNOfXGfR8yXFZpQ2plBTYaWRwfINA0qB
8cIwdY9OtYXIA6mOeXp05o9CoH/Zh0IrgNTL6ZqFa971hcOaZHZWlYWsKbRm+pcuMx3RrMSPpYb9
TE6wYQBBKRkGrtIlg3D8cjYjH39jF/79QI6ZUhhWsSSYVLN3XPlcZHxPiwQ6ukkAkGqmCH0MsSc/
RzKenw5q2jRLbERs/qBWtwKAD8v79EpvxZe73wbMcMikxoGgWEITBxdtv8uUBst9J1K9+FVc1zcQ
Fo9tEyvybuQRR9PjYZi7yc5JSKavX1/91aNxrh5xX0jkZS/QvTO0PV3WUyMoUWHahtQ6tWvzFwDm
ZTmAt82BuofVIDqKSacoOE1GgRLJRaf3P+4VWCmCcQNywnI7OmMhFztsIF1yV0EeGNQX4Zw1QtnN
ILU6JSz2n6DISwUTBuimuMh53me2IklOdQSW6f8IrLIwKrYkTFS75tFtEL+gJihBmk1QAxBlBJNK
8fOrDeEuCnF7Kr1pDgRQIA6Graxro9hSphTe3l5B53BY1hhD6l5S9kdaKSY+MBLVGDQ+ZG0wGX4Y
rN3Amd4hBE7kBnV6jFLmREkbNFVnIxYGruUD0vKelJU+GhTiqL5dIUroZ9C573jV9ei5bayB0EB+
YUYaRSl1h1cKue8NiK8ZCdunJEW5RWoUYiiPdANJV5xJMQs8pBThnUU2EprFmyanhqXkHF1Kc3GD
JDh2mAFs8fpU8q4ineCsZYA5cZKueO2VMb1+S33BrcgXo75+7ayQVSr6DK57z67fZ5YwJkgVmTXC
WTagVmr5Zl9qO/IjxnmzM4Foj3bIMlp6uzBZ5fx7EREFjctiRhrl/pKfHgsPXU7hq9xMEUzkXaU4
DtpQNecXiaUwNWTt1w/wRqSGgnwZpAyY5MCH0PJGiGIfK8EuBF3auMh38kMpjLk+/uDgl02pUf/8
qSYW+MvtKtuGHnuO508XQG2isiYztGDwea1JObkj865V9fzGD7T2IvxbNyuTOkbwXOuynchsl54n
IFhDcHd0ntzI2HRgfhDsIGFsWShARlGb+PU3zupBlHe6EzqldCTahkCfq1hYLXvWR8Vf8U1kxSDT
u6/PzYIIfFrsLd4PDNIth874lou9cTMRPmS/z/JMqimrX+mVxeiYSawAjD/jrpz6nXJdDCEfLl6F
Xchkh8Caq/5fCtanr5HYmz+wACnav3vPmnH8q6RMVZGLD03XVPe5DpPl2GVu4N7DYaF8I8CVJGC9
cJFZ4JgW/eq+vRe2nDqq/hLMNuSbk1vWmlR37xAXNsi3Agvu5cYhJA6M9yT+VyMXgZAtm9FJZ7rX
J9F8HyanL1xq8ASuwFJ3JAGY2kJ3M7SjLFFVBdAnIdMjlGUNy6wytr7w+CMXQMw6XrkSodunTUx/
ehE0Nw+7Ol/tZantO6rhs7S5nAabGEopO7aoUNo8eiNeIF9CnoDcn9npegCxBwI02087wM5Q3WeS
ACB/x1n00w4hiAoNrP2yyUOP34Cl98vbSuzQjK+sL6mc0UFt8sOeVasbP5hOVbvJf90JGQQgIxGD
efr3eqo6e960NWlIIftHmH4SkuCTEC9oyrS+Rw9zd82Xuh/t5bJ4mfBG/loOhk4ZszQA+a75QJ6q
ZQqrdB1hDcXS7lpR3GtN9+SdAZw9DG9M/U0cGJsmK1eptbd0V3oe+i2+CpglvwRoKTJDXfYnB4aS
i4iFIMjrTikMxYi5swCcQ+tDYrXPDIwuoaATxzT99yeCbhQNKtSHSUt9hokFSJRw6McOvhP0cESl
KH4Tk6dZnmhI8sIWEFh3RMKPQkbCRSDk5RgGWvVeOluvB6v5Nv1a/q86OlSMCxicy0DMH1KX7pKO
04B0WYNNBS/k3m2bvoYs6EwsPcxYmGNuzis57WvVBMzwi/Hsm16FE0QQcPAm+lmj20nOOnxZLeAt
KsBa8RVU9Jzph3kk9UI18NASyrKtdBtKDP0wLGddoSkuP2pRfgwlffBlD0BskwE2FZmvfQOntf8h
UziDScePeRgX51BJ27RsWnPCxqfsFpCOsfeQPjFMGhU7MC+i4MPfscFJKGg9U0zrl8lFNoDN8iel
oL9lCyuAXGhvSh8ggwOUAKdV/eFvdMJaHCZ5oW6DX7N+9pHFu1+E+sqxnGCilwguVnYBq6tGerkb
aGNKDqRyh4v9XqHwYBLmsi7fM/PQt323wl4UdsvEp/p9km2ejLKyHeVCbcACr6yygxERjWcjFCVe
2hR1NDsTzj09Mpv61dQc1POboFwb/5i0gGy4MHNjl2kO9z6IzRD8yBbyFECJEjmdUmQLWXHA36Yp
xwgbYqhKzrPEHDqLfLiRmVZZG3/1bgIcIqcFNBb+fBKdePwQQcgYkMV4ECX9lbFKuA6VvMzowVX8
oDxZ/V9OIrceoYzWH1o1bYGpeF+o5kizMGmdwOeuAEurTS1m/TO1FLvR4Al7UwpRGoSIM/tWHrIe
/2jKehPgZf6O2vyptuabR5qiINI0wcYK9wDKFB/7m1Mu95mZdS11gPQS3PU++ek6PECrO4ZEhOkE
xHCq56a9nTgUR774zopQg2u/6XfdHftppBZL/EQR0UT2KYEbrIHZDUDJJiz5M8+eBT5TTEvu9IST
9lWUYM/dxU3Fma42HXVnFxyFueMOBm2FA+dxB45bsZ4IzoRrxuVZP81Xd3xiB/ggxnSkCDhg4MZ0
8oieRn251c96WDmZMJI7NDouT3Nbgt66oOWvlnjfCQ1JnbIkiP5xlli3jWmvK+VhmqR/Iuh1WyeY
YiprexCkeNaTiu6Z7OlgdyVL24LhEE6a860mDuTfMIxg0+Q89ekpXux3kngW13PBLaYnbAhA5q/k
dKwuRdzZLk8JbTTsUllo50qPBUtDxwnRa6iROoUlvjqETPOmvDH+ekHArGjybmqXIwhGB7I49teY
gcEkQ0jj5Go/d2N2voyED4ZhejpjjCiJGP4uxCAA6JU3mt2DSZGC+Cq7JkJKnCLJEfa4B0KjJdy9
NEvFqSdxmZyT8X1OhumMHRGzSGXn9VoTJrHQ0tuffe5nZiF5ozeLGIJdrm64fN0ELYsmRsEAkF2X
ONJIM7Gst76HTtFrRKHtBSCzqLW5XHMwjRo+oviECz+rTjX9+HcneFcecSKldZI0FfYiFWhFlSAs
xpzxI8/Hhypuhb4X1aPNzfzmyEM9HRw8otvHviFOCxz5252F8uH/4D0TgmnPXBNVm3hDzhF/MkrB
vbWIvr5jB98/T/q333z/7fpYb7EdXXYjjGXs0k4DlLppC58gw67pBDxgfd8If3EfN7+A9xzbqC4o
cgey9p0xaYw7H6kDDsFob/CmtQQ4UMprIcKXqxUzhNha/xeLk5ugWd1fz6s1Wf3QzSBOeGVpM8vI
odfZ72s97zIUHN8A93zJFiPOwetgy/qUcNvEsyTCydSbccNmHJ10HZvgTg3nJ47Xod5QdCyHbhc9
FMFuv7K836uztmUcnOytWJdhqYntcU4bt6kjOhmyYj+fO0tFTnd3uFpgaabnkZkYi0pUwBNJH8ln
F9+FGpujNqFGp7Ke9Ky3N49oi6Eb0tdnQLK9eYUNLnDwpwdskwHKljOEs7psIVs3D5luAJ0RzDHW
oDyDPPKwV/Gblwu7hQXW1SDimDGPmihfO5C8Cou50Al70WrBgcGdW95QaSl3xeGilYE5DUAkchpE
9vRJyBXN1tOFW39LzoA4098LQINCJOiXsoClMHJ4XgBRxtwlK3blC8mInKH40doKh/W7/SgNNRnx
05aFfm0woSCB4YAZvQlcIUtqdmpgIH8ec41YbHFsgVZYhpmgw3i1U1RGtdntv1QH+aotnlPe36WT
8IJSQCH3AwC+mk+BDL0ilVye1wd0EEvT9AIS9dk2lUTbsYXNhBYeaMLn5+im8IWdAr8OByalx6vf
HjDKEvS7Do+M8ZF8b5y5NpfUQfH3iHf8+3BgArllHyL45JU/j5E1CzshLb+j+uCCfxueU8xEETFa
iTGgqhlDs/Nl2p/nLhenxgAfuqHP6BL69sJPRZrBk1L2BfgP9K0PJUJk7bo50ZpY4NPkv/6BMUUq
CYZZ7D/n3C8IEQCdhgPR+/F6HFqcq5xopkysF8p/B2XqAytkjU4oZczfl/PjliwYTTBpFUjikjIv
qTO5crPlh4YiRJoHlMYxyjO1ngQ8sr6dqt29K7/FwI+L3DPPduzA6BTN9dXkpEgrIEZIBafgXYvd
vRMo6hvYkmknllr+254ClmqA6NUc7zsQzxUiZUWn1mY5PXiTIh7CEmm6xJ1x6gQl28h8YwEXF786
G5Lk37GmkvZkIaVuNVtRi0dn0pRXgfU+gPKPjkxntZf6kvaTz9Cet8k35GwJu1fQe2cqhdFmoDpM
GOIA1THAIaYWjNjJmb7sRWMfSskqI0chJHvRDleyJPgJWBjZb6P2mKIvdrD7r9z5szQJaGs8o5ed
kgV7l9kItRGKkUAlofp44u7v0Nr34fUubBzkfkN/5K0D8TtGOH8oMYWLb+S8Uz1J6P9NGtmvQjeu
j6t3BdCwuRL/FWyVbSYOC3zpUuBzB0A34i9LP2nJJJNIg79wg9hwkwe/cKjyWVk2f23fiV50ZhRs
4TPnsxCGsgvRcEqR+CwMf0JGcshgMnY+kTdHKAKQccqPBeSKV29LLQ+MrfQcfYE/OJNUx8jHQ1HX
wSz6ARcYvavZjvBEx5dPJ4upP7HU3G2J4kX8tKhVsqbsWFWPrTfFEzOoSbAo1g8Wjo+67JRF55qA
Cty3QoQS+vwL59h6piNP7aJACMkCthyv4tJr6v0he9hn/YHcW/IBkCEYq5U7agPEvCHmeaeTmC4Z
VAnhU/xWZaXF5iv9+hKsv4/eEvXoiFfj+V8pa5h9/e54r65zfCH3CHFtOyjBgHcxoL3XWloIQhQC
CDFuCjBPntFbnEeKezZ1Vs50c5Y06hvPOYCieGlrPcX4GfQ122zn4qCkxAWzl5QknCVY4CSiOUJ7
OgyUn6f3VF9okWuWJAG1wp+XG5PpJcCt8YFhxXp1h2gzdSfjwWRvjFtoIfVyoi4CMEdsz830uEb1
6sdJleDkEjM5nQB6kJhm/5yW2433jhGVjIJw7Hj7KDzTwPaCNLQ8u7vtT1L7BY+WFEvWi28FF32Q
6JVtMoWlcnQUtcG0x/ICDahjRKsZ1NjsXMOWVoNDTn8W5u5XiuQigFX35xq54bFZ9g4fiRpJ+QsD
B8NA5nzxqLc+UbW2r4jpNMaDfBep20OIu0ugVuLGCYmhtHggO581OLhfUioeFyt5AGqfhge1e6gf
sLKoInAnUQIQcbnfgcrdb2UMX1pL29TqEVeFnk8jhv3dbsnt1os/fQBB/IrdKiUgd6LetrKWKBy3
CNDCZZn4HQzgyyk2x9ScKhPsA++U7sTjtYTGc9T76vBrJ2Q8rtwNny+xhC5P8F0Uw8tAZPzk6AKa
OUhru7SX1Q1WjhI6A2jGffTLi5d7d70hA28X5RpzIou9dVfKOQe7ePx7o04H8OLIN/z5hG3oFSxA
a8c27KSRFqQE2nq0B5nLKBX6lT/RCxYURlHdNMFe3isYPQRk3UcmqXUe8gRb6e7Nsael8JZYamby
BqrRZ7CllxgOUOEBQLLQNT1PwapYr6qgs/T4hSmoxxNucHyM5IijKxQw0sh1XmR50q2ZS/qgdFcu
U1ihrb4MWKueVuu6AyoLDiQ3SMbWBIJAtTHc5h7E2+GDICQvI8a09Pg15rp8k+s75VnPy8l4H+XC
DbKmdVCtnLJCMHW7eBqBKrR3i7jZ/Ub03GP7mDLS/YQ521Typ0bFbmRGASmUrJCLm/O4wus7+3ZU
1TyJR/fy52DDasDAIGfpYPAcAZByMpZxmL69DqiKxRmsOfpJF2oCtt6uOGBfZ4z2wzeccuW4bKky
JodfCWAazwoghWHKzIMGEyUiqp5ifOSGDWK9egcKqqBQdDilaHoc7vCtPLln1pZSZ82J+EjQNPCd
DrbnYwBsl0WsiIBpHR72Uc7vVPuRConq9Xns3sgqymeHbrWCRyeYQ2sLYqlWoC7KGxBzbaEPO+wy
sKSPGC2KDPRSdECbdi1NcrS/r16EbelOM/o/wAuHWZW5DAaKsOsbiA87pAR+Nbft4ZqpZhFZhYl1
clHM6Nkejv3Jg2zaBlOk/IJC/1Kqc+gE5CzK7wdDL8MIFG/Go7GvweFIVLbnS2Y2tnQ4dpeCZrpT
LwNFtirAcZDGGHqXQ8W381KZRr3SSIWP81KoGBX7XjMJuU3zTSXLk3F76JM2u25mcoQ16rfAO1C9
LRe+v8oCjHBKpg+7KFkw/PgSQbn1P8AVJtf90mV4wt4W6nQbO4KYphu4kOWAanuA2BGN+jk5INGx
8EYhl/tarNbVsQ3HZFg3bHjJzP8XV63IugP04l0Op5RZiBC1hQBqH/eyRj+nypL2GlFhQ2YLsFXL
poW3bsEKHb66qidjhRK+y77S3IopKkARv7ogQ0WC3/Gf0b0pzrPQEQwCJm+tLpa+9HQPsxlQ2a2n
dsIZDBxj7piykgiIcwFZwvEHMfKrcGAsX1KjBe1mgPq2uvKqPCU+3EmcpB86L6rRqE3KBvTEmIYN
JLooaBI9OERy2cRRiH/40hBi1jqqc30D2/DkkcUppaUaHMwWTUbtTSzrO0pB9pZE2VYDED0a05ZT
q/H5Dd+EnWGr147i3XY2HAyBRxJ6o2Ry2UsLEMo9movqTdZeDxffLS6IEL0ydBTvW2OJzkoLBWJu
iHyQrx4Irn9WtNfYgd5KRZx8i1YCvN6rHcmAv/oalTB4DwePSuCPTsc01+NPfrdTyiXU2lZ6D5mF
LsGNy97XeLS3HENz6g1i+JxyBC2WFIhr/fcdBnNS7vObNmPxBMxE2kxJgO/HSTYK93TV0udunGma
oNpG/d7zjADm7UUgjJl9rMdLD8lehfFCvpW2JqKq3mBnqC7xP5YkX0c6QQhJU1EZyjFV/COCN5lh
XW+Uf2+y3Q916/84cABD2b3kz8rpSvXqPFHXMeF6xq1ugz7jzh+gtaE11MgoNLN8hTvGp54GFxwI
T5ED5m9NjYpFKQ9jj15LlIfVnVs3RZR+Ln5kWlWMdis525XQu4VyVBjBTnwc+G2F9pPLPvXvgs5z
WeOc9iQdZhLUjLVOV0NaerJDr0rRWY7OP/Dwv5Df8/kiM3u0MPDPuxH+NaDl27WRJm0RBmVOzBe3
NrK+EwzxoO5QpXq/FvAjh6X/QlO+inDZLkmsXygTJ4fAci1C0LtZ2S5xcXqO1lU61rDr8ZJcjAzv
EUWvveMBUNRUweiSatlUO9zayhut1LfldWObbFWh5qCzY3QQgkvcA3fJkNoCfknCIYhYDikFNdbW
XcltCNa0DSZUC7eh2J8dTLyJ8qe4HWW+00l66mLmyb+oEJ87Lm9rx7b9ZfIQ/fahb9JynhTCJi/A
9uM+Wc+fBNwNt+T4QVR2B0t9jO2Pkx9cAlX1qnBlChLzylv5he2PeuuApUQE5JbdE9+jZjc6PJdy
JkWkJ1NHr51mwzrDjshI89vwONgYQiNa5jsxilWjnfoC7eOxGlshqSmQ7KZJahFdigr8/MAjr5GO
AlRYMPcGv3P6M0cIRsEAgmo9ZoP05Yztejl7VdOvlJUzLjZqsVpLtTfdqIg7p/3/4CZreKyiCoiw
u6ceUoa1XooialfmK3gxYrqN1a/5mPtmhfVPJAONC+Smr8rsvKTwoo7uHYXre5SgEZyPAERs1pGi
cPuGzEJkC/orr5Lc+URYLWN+Dp9eQ5UMs622DcOanj8eMRAeFYGcrMptcYf1TfzDmb20MRo0l/dy
FFQgJrvU/ABw4v8ddixhf76F4hMuqoLMd86R+jern6LqLfL+lcfAF9WOmjcFUuzazNH6zSchfKm6
`protect end_protected
