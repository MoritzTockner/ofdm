-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Mut2mHnNuEXuOyQ+8Ldv2xfqS0SmrTo/GDWbGXwXlNVrNT+8jhRYl3gCnCEoWMxIcMVp8BG7BO32
5/1gznllGWM5Pq8Gr8uhXUW8pVQAlZMsCS0W5g/LlzzuRkuEc7G7Wl2awMdGDT7lz089HVZnHJdp
fAXTT2uwZm1RlLP+KSyv1nUnHOJqdaSPSxQIsYWHUCZbKTNZa81EpTIEZBV132kN8niKwu5AjdXT
oq1SW1MvwUNtdQII5BCY8+zVS0gZkTqkj90GtU47TkcvktFR1+lKH6IQ/4MxoBHRxM6pwHXf3h9b
OJouxatQyjWNKhH59BqCphWP81V+tthTMllLRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
4xU8bWE99RGf+NoANtkCb8NjtI9KnJAc3aaPy9LbL/fHAzNrm/7r0LaYS3RYrvAP/8NEI/5UB57H
gyXJ/OXEECQaUkrSJ2f/5d5JEJ/2NhZhQzxE/IpMzUJ0zqlHBbaos5RYbEqu4a5/wkLxbZN53EA6
6bEe2w76TVHS6+MZdd/nwT1NWsUOdJm9SVPbkhI+1Vwj18qESA6ZAOSnu+yfZmeFiXfxVIYV/MXF
DDa66ujq633Ot7PiI1MhvzAyQl63acLsvT/3LvPUtX9Y8I/0d15xqBS7NA0GlDtAWr1Go1oAYxC9
+oyhzqhu8IDfK8b1fmJQhG7igWNOtH1LRm6CoBUFycQc5EjOqFQZosKM5itaBfxxowvUsd3AhkKB
VyMSuEQ5GuN1gQSLFPpU48vaohQf5r3mriQXvGbDkPlBRgzYny1HgTWtxFB0F3bc1Md4j+FoAYb3
q/l7gcGJXoRQ01jENAq8l5PPhqbo611rQOAabwhc3XbwK5uYe1m1RBEgBmbiZ/XN2HWDcoUA8Rj4
Jy5BiZh+iQgW8CSe2ejw7x9y8VD02BJmcDVAuQ14ArriACUlQyf3csvDDW9G3R+difhy1MC/7MKL
3Q+Y53KYAVHoFDlEoDSykmva41eBEHkj7/D9AMzamZvWA2UZAXgppmD/DKmn+f6zwpXlQxybE9gH
DFTkxZu5CxIdivpSx9I40UmoCYoIDGqj5rEZXiqgTy/OKQud05VDoP91ZfJnaulBBCMmGgPXyaKf
KVugh5sjt2ngV9DT2abb3VDZpZUgEd+LyBeiUAbiH+bSlwNvFivUhJH8NM++oMTxCFPJpRH4JGof
ucYgNKjTuQ9/smsZIxLPcufr09hL13o9GiQ59BZo78Duh6Ee/DQsgslSPCIjP6es2Hvl+mZf2thb
xij3kpXDwE8EJTj1eSuLbFjZD+3B0TmAiN0KnZaNv4snSA/lURud0ex4jwGWwokGeRIDXyLFnsCM
SAM4Y/OCUpJ3xDVH2A8tYu2PwM4WatqPxRB7ywG8pxa+4B9SswQ85XSbSAeALkmSfjesm9R08nNS
D8RFK6c7Glf6lx2XdKWFnuYFMg5A+qf5H7MI1x0fisx6tF1XP4MSDYD9ZHKkxpb5LgJlAWBSaP0s
522YxJBTTF87sGD+3ARfeuBCDO4HSBICGEGMBzs/mBHqBKUIOSpdm2QOeaE0IDQmMCwNmpn2QhZ/
pXrls9NmWnMxi2AJcAAKHmKqMUMaq7vrxjrhQE+NnImD6abiYV0Pku7/YKSjtqRzdQLbw6LJiGCF
FhN/Jazn78i3MBBdDGRV57HNpDxFVSAA2IvSO3HvFfChx0OjLvTCrUvCpXZ6FwxWdCTh2Wb9CM0V
Q7zb/N9putHD3YwVtPZ17fADS6otTDISDfqJ7ZGezZQq0chSJtOQ8OXX1rbyOt9KJoFhugJxX2la
LF3ODNqsXT0RNFWI90Nc1Q689nDiZgNs2qUm3CT9zYA2WvqAnFkWnodR/O/3fKrr5X52ASMcFEFv
GnfBx/LY5TjLJgLHxdFOEBTtRbb7Fv5GkdDtuXWQ68dzukCqpyEm+OKpOCALA3GgkX4x1FlrrjpP
RKbzdCDPio648dxlaBvBGhc7j0jC+DMUrc2KwtJbVQ3wjQ5X8nIb5DSEtueRP+8rmA3jggIB6/LH
P3YnhYire97tTAtBqGVg+DG6ga+LReXS/epShj3msA2i4w+MgCtBgBNQ4pktt3X6m6j7qEbYZw7b
6coS1bNOLomowJ0FfAWJ2bcsdkZQOMAPd3oXtLqTf5q9ktDH8vG1/NmygwX+FCbKhz1IvZLwdQ2s
B0CukWiQyHnSuYBrrxZDiykY59E6nlD/s1qxKLJdYdVxOhblSEIgBXQ+a+rXOrTzAwiZH/ZdnrIn
IV0T7qa9ko7IhvaT840JrU/B7NhS/sVwN4TA7FhLA+VfkCpxxB8t6QyhZmS69WpnI01qcIGBgMpC
KRB/Oi4cswdtqfKAYT2VmYC16eTd3iN0rE8M9ZBZ9a1b14mzLuGJqan9ACi4dOs4r6zKkK6WQKQR
zYTktsItGWHj1RVzCvqLxvc3eqwQZNyvUmhr6pXtE4iegxLqBaz7YC0yGKpoTBcNrg0dotnIt+s9
IGmQumRIotLx78jGnrsnQSqMbXHZtfSE8pDcpNnayPORur8L1rQK/fT1R7c+E6Tab/rlMyWB72T3
DB3dG2XTiIbmthF4/aswWD4TYFU8KFVJS5IwD9D9RW91XcrXJQ27wPxdbhkJKYidVz6vqC+gg44T
h3rlNcWvz5Paek92kudVwCSkbqMal0k52ovF7x81u/jMttAON1vPDS2ai3wu+vhNFHCe3ejg6j13
VGdkDz+ya51N/kATa5eoIeDBQbeuKr24Wpk8Kn7vasrJeza2swnXL4eLlITbvRmfNXbRzhw7EW2e
FlYEG107oAI3YFmxQAG+UnYP3lXWQhkhWRHCY1/VGK1nG8uxb5HniGJCKT9FSAEsaS/kWnjvvnev
Pi0bX19j+C2EuHUzshk0mhxNMy6wAfR18nVUVUV3eLdx3wZq8qne/asIJlbN7kCXw1ysUcEkvIh2
1KMdJT6nxqGOv7dvIACdEuKf6UaFU73MfWlheH0mljo4xQhicqvoqbMS4qr8FqyVF526xrKP9wei
9uBLdmLG3C+DZzRc/+NR9YtUfGENWK3fq6ojVJvD+tv4alR6//o4yvcq6GHFrqcxvk+CJJO6FxMR
8mhXSAHKaTldiL9Kt6j1+eHlJvVugyMn3B6G79KmRcXUTRFJnF7vhx8DVX2r2I7ypx1eG/2xQgv0
L8dsnrIlhC1v8JxOmEa9997ch6lr6ExAumrShog+0Kimh1RfPnvtKHvRuzL35lsHz6gwXGVJxI3g
O9SMLcyydjDVc9WWsicFj55c3yu+2FSpGMvT18gAkB29L1niHzoFec6k4lLBLZrUspcjp8Lsp/bX
/WBbL/VCLf33G7hqhDYhNtj0ipnLBYUL+C3sDZcF2kx1uyEEEMoTs5g+m/Z5bWngYLuTCXBW9bqo
qmjiy1vux2qptUZIGmCcc6MMyRzSm9wkSew9jsENTob0RLgfJoD+ZO+aIC1h7O9nuZggFNxNhuJn
TgTG8qk+nGfuQKUmKHIT1VnhT3QhvhE9EIlXt4tJfFUFAU1LXvZezXEp0l/b9iCHl4BRLuiym4gg
oprrcvna5YZVVVI0Wq6joYhaswacETQU8DFl14P8FLhtMDLIuog39TraFjov5th5Pzo2TzrZNQER
b/UXittzG7QiLg0qK7WtANbIZcpyc2XBGGOjEIYcBeUBwvwrE7GFEmo9FCrGRll/Ft6rrixqBqd7
kQipEcVHG7I3DvEMAdQm15mG7uos1Sik8XMWR7S/w/yTc0Ty+CCG2KT5SjgVTF4ogdwdUrV0ZSRs
zBfb97PcYTgHL3/FslWDjXMaSx236iO+JphQCMCY//N3JPnwAisfPofKnsyKWV7S6gzk4n5ipM5g
fydbt+b8QXZ1QBxOc790oEMKZxDyWzSODWdyGCh8iF1cJ4aSXKXdb++U6DZKUThZ9a1sPlqat8xd
x7PgGHnFjw1oSEHZ/7yoo86gw/uVAyEgpRv7L+hyaMnL39nzkcFi8Zj9hnL2jn4BsPog9DF2diP3
/6ZUo4ymq64vLvWKumLgFtyIDuxM1oN7DKb/sg8Ofaj3jfz5OP7Tc/svWL/HaYhRCWf/jnDofrZw
L8WQ/A18RI8r0x6A3k+k3+RNZ7dDL8Lp1wFEqeXZC9t4cClMMyoTeoNAXYotTrP99NMNziOtcjHl
kd2VQ5ixgIidsV1sAa8Oz7iNi/sm9dvLC0N17r3w/9QjvSYVPOfRLABJpdKGXOaUuARnr0iEUbv+
baiBIvQP5FPiq/XL4iWFzyRaJBEfgmuJpNWCKeTbLf3sgGIaCP8jE4nIgqEo9eWQlNimtZNSkB27
D5WGeRqDCoupdzh2W0JskPH2XpRmVlvHJiIBghukCGA85qAgi9doluXNvsomYit8hGCIBIvezUCD
ROi8rDJpC3CTXtju5Htd+JPpxagsgMdTlPBmM/rEwIDT46MHg5CshDEH1BVTCX4MFkvcjIquRy/+
yMwLP53JndsVdoZ9N6UbYPE50bA9Iv5PkCiCmmgXiC4dj1Dp6NFedH7ZS3rXV9lAvQfce6ciam2F
38YUwA/Uyuh0IF62Nw7aXGJxd44WQDf6HPqzbevUeEpmiqLTcA1jawVI4T7XWDNDvsaKot2CNKFs
dpZxV0eUXLHZZVRblIZqaGLeu4NrNwokDMZAMGm3w8tsrGyEean2ahez8NcFFLwNJFTw6heW6iSm
1qp5FplxImj9oGslTqbIqumyEvkePftaCIRYm8NDo1VnXmxJbO1mpN+4iT6at7HllzpfPBVRn9RY
JxPoqSDFDF5A7PwZc+WNmomqR6WICPLTqLbkJ1c3L61W14lClNDQoI0cvnC5JdGDC4F6iXAuzdkK
FlzLws1W3fHIjjTbbOpIvXclTGqQkhSneEUHm7NDBF1c1XEtkV/+WBEYBSZe1rjMXuuFlZPor2IZ
o7pCm2qSoUikwxc1Pf4tR4yhyWyfT4FGzzqtT+BZlqTAGyYxPXFlk4WQ409iyGyEUK3KHtOcv96p
cx/RDf3mlo9/q8KUGE3nV9FaeOd2lmNfYUB8x68vEoed0/A0mRTCxNY4yKaBcw0XST5LRu9QXj6G
rPuJCB79eUN7qZsUWihJvfIfY4uGxEXOf/e+UjL2XJmYI8f+oDiRiNAsq+P4NUanVuIAl8Xq1kPS
C8fRQvs2lPCkF84LECpxoR1G0YhFhkp/TiPxs8Pdt0bO0AU3nGS6GPWXNARz023mDvWuOX0P1MfN
sWqezTFHBc0ZHLRKStvnc9eOon/lC4X0A+sQDjvRZC/Xs365bKgW2j9Z4rpR1T5G6UlaTyk0Esri
nfOcQNeVymbHO5wnzXwYT+9/yjbL/vGY8okC7i1H7ciDoy4A2EMDwQhAFVvh6BAc4M/iSbXEv7cz
RvafUXrBkC7syLiPIXBWos08R+mpyLGqqXSOB6lMhG7zTrcxwa0DJOWUzVDeftc6IpYACWDC0hyX
W89cwBCliz95NcFeb8RERPallSjk3tuCIWjynHjGRDsLbnbCHBDAyinoC1SZgjMWoF6GhGqx3Qnc
IEBllOXJl5yae437noSXlY2to1T6uswDmtxu6l8kbmxL1miKKVHvN+aqvXINKdNa7AXJ8kAvhd6F
owfmU1OjH6BOgUIOqTPgk4dPLJIXqXmgxzErsJHHKpePKWvq4elxO1/gp/wz4DfvdNaIrrK+k4sf
EKq+c/oRD6Fvl8GVtyUKSn4xHl2y/anONsEj8p7ndOoIUjqzSgfKuL0oGIp8W3g/OX0gXG070ONz
0Mm/+GNfiQjBJEkhSuoXmMMaht/7le420nB46Ri1CiXKMrCHhbamoHfVE1qiURV+rrzi0tsO71cb
e1nbngOFP2AV2sRIu/ZxvQUsHVu0OR9oyZO9Q4iFzG+ytp0uCIjocolXaTNAeqQXuvI2wacpwVoU
eT7goX6ESEgpNcSEnEScYI8g//pj+4L2o38Qywv/3FHorL1Rk0yGT9sTD7JDiMqteoHe+ErL0vHU
41vVHet3y6z/18CaB7aeRZegDEdHto2L/ct4smuPf0IMmxTolH21z2Mkj0c/KekQWWpx/ieS2EHj
5begdKeWlLKLirWgUTlRT3q/Kg+sT7TnEv5QjYPu7iej5TJSKIbj9J4CIeXSGFFpQUtLf6nj3l1v
X5UxiBV8Ebti5Gf2GTXUarq18CHA7QHlZyOsjJjtLmOyGcyzaoNJ4yWWFKgY2VLHaRn9GJ4J1HmA
7YB79VdwSleuHiOLE5aMZgsyOG2pZcjgjW2w87jAwn+EaTx19vZeWGbEMLNb9tssZMC6oVJeOZNZ
9aj8ejWJm3rawBrL7OUTDTu7Ns2rKV7INMxf+qdf3smiefLV8EzQraUXOQR9Fq2pVobm7zbIiOoO
CBbauK2ZKnFrGaiz7DLvglm7QnJBbnwspNaU/WBtIK79H8ucE4xVkoOT7OH2IwiIS6vM2nlUNhUc
rwO1yinCkM/EeDcz7cuTomc2GNtsBg6RSNJJo68yO+rHT5qR3vDcGJKsu6BDEzngY9QLaKQaJ8QG
frn4+0GbfMX/e3AzrDA3lApU0PuFDo2PdhDYY36f8er2EzrQ8dzFNSucWGg5TF1HO/HmcuNVHG/8
7zRPww5hABQrf/SCs5pOmRy4e52fiqNXy9wkvUQDbG2JyjdllyjptRXnh5GBrHlpnJcDsowRp8JY
rPTGuKIgdSsXGG+p62HOODZpmU8Vizq2Mu8H3KW781mGB6D5rElc1gWwIjjuFrxOWi9PkIXRBOue
AkaUYhryTP3GGw3zwF+HrplEFuTjgDJlO2nLpHKmiAk3eJYo0l6eo338yh/D/kaxp9Ac3s9lWV4h
XqvW9hiR25sf9e8T6UDYVBZRCBL+syfWIxEXyDByoZ6+D3pqAk/Cv9q27Pld6SV/uc7db1v3U9Sm
LL3ZOpQ5cyC12gAXfmAyLOC8oS7j3xcn9G3/iPat/BXQoFWRNpryKvGYArJrw3zE5jaoxg8WQhZ4
ZxqcHUsUUhrpNBoDHqq5I/EBqamqQ/Hieyqsj3TEhtmzpkaHwcoURugvVob4tKKugPtLdz9CrXq3
rR0gpjICMHqMRFwZaeu5eJRIphHsDwjWSGJdEAitdTzVcrdINUVblP8mvXSikLWL8nz43bph61W+
F2UjOsFOgwZRwoww+oPZTdCLWAQstSTHyiQ7KiVrcsFDULIsUd26IVqmgzNOSm5mQmGdpxnT/VOJ
pqWQ9t5WfRtEUJtXN3SvFZJUom0KrYdWAvyJg4UbYwXjcwn+KsadLGGkCgGB1xF8qsNw/dKRAJ7Z
CJ7C9chU2TWErNi294pv3FEirrrEtDk8sMUDsScPeMgp/3sI1dTpQkEvzpPlaE9gfOvi8yGpowGk
s/+6z36Kg4eJg1uDOuPwzmRuuu7+Y+aT2pi0O+ZDfGiDmw/QNeGGqTAjj2HsNbZnOU+cZ+zIq0nV
WOBVkH0ZPd1tt9Dfz3PFyuoJPs9tQNIEEmhTsOZGcUooot4skqyjnkaIeqsa3RA8y/3deXtC2Z8y
MeDm9qmGNydKgmlco6uuO8SlqtktZW6ZAkqbH2vGfe1Axa5ul81VVOWfAhtz3JrCrxe29feLobRJ
rEcm2K6vx29ggD1LtsXeRS/C9IfdAb1g+me9wBSrGlkNeQhCeNG04UUR1LUyY2hP4dNSzyvWVOXP
DyBq+q4Gr5abpc1IKH2N7ZGSfEk+mm4F8SgP+S46yXl3xXC5NkrUQ4ififdrgBWJDzIMq1Fsr8c2
ulKDaGJp1+CS5XIRiYajdJrWM92LNX291Avv7bIDfhKB/nwhp9kl6rRwF63x4kWp4csKOozjYnfd
eyD3JoGDREXJM9cm4fLwYU4d2hcgLimABOpa8UdwLbabFjFq93jz46OV7qomc05H8qDIcVmiVAkZ
6HjxtsncR8DauTR4m0JzkMT5nzEjT0IYIrh5mDxYdva1WC/ynaoaPAU8H3coJrlZoQlrtKClAvM5
r+joE2tBT13rmC6zQhKA2ADHB8sM3kLxKpnd0NuRc6HTEitWIkf2I1b5IicwbnKzc+lKtMEXnN14
J7vhktufycWp5f58kHt8DU8w7JeHVfK0aFzYeh2wsewS5yerv7wsLFo6jDzL6/hIO9hC7uRUEpVE
PFohc2ZBzrJUTs7homcTnvQ9pqzyDd8WGn+yY9nThZ0pMyCRY31tEoi0OT9XXcdDOcaQwdcNP+VI
Gb0xMbPwhtDr0ayROSpETk/2sDL/K9JDdR9b0x5CwX6qwirMFdfFp8EKwervYdTRdFKhicfgCMLz
1sZahX0AILwbYag5aVmB8JlQ2lYumuBOlUhF5IzjHzxrinWz+ZNWh5HsGKsnLcYb+7RcH6QkMG7h
1vkGU8muobeI5qumxQ/z7CuCPgVka6NTviqFnCWOhKakQwDIf3lBx/nqpmZDH0Wel7myRXis2Bdu
Z0OSaNcElW+zZij6Hhn2rrEEm7OlQd1jreOEFzY1+mthuPj3FGcDZo7tiX2Divnt6CMKD/V4Fgk2
N6IfpzFZ6mGruSYsX4DtCmosmFk5HwnIFW+mOTz9KCQMiSA81RKvkcLJGlRt7MeuZ1E8AYphV47q
YH9nSInXw834uAcioq1pC+JS09d7Hgta42XOsQWF1CMxr5d51ebUe7d3t4/Sg5b25ZoRmkJnhua5
HvyWX3CSIerTLBevjJNTW+RRK3ZwSouap4+rBsRcagBiicegRR+CIfxXlrznErrmes03qrsqLoQE
nYoHALytBlzF/EabLJfs/GgNcgcaQoE8S9PncQcfg6OvoL/s9F2LWsPHCs/3+dx2eur0JvmnrC54
yLtq1vZwuChVsrmiDWFPvfmYWVAnaXs4lS+oGgpCcEh1bMxO3MfFU9szTraPAyatiRCBNyKtytWY
bRUlZJxK5O+/DYWcFRteE3UIdl87f1p5BlzYd4IpsbUvz+Nqkd6DQGPWJoP5GPk6VZEZas7IICEy
VEiKPOJmed+i+nCT+shnl3jRnPI5x3g9B/nS3aBDXWq4VsSZrD4TyBTBiROEPbDYJS4O6kJaWxKT
SB4cGAibXCsPjZlxrXXMJDg1DTVI6J4x3d1PRrNc85udu9Qy0VgqqbuaGsX+s/xx+t9AyyobUsJq
cRneNRPDSpxagsSF5ml9Ui2/3C7fseAfvOg/u/IFsnxCLcpkk0/ExISzEWGdvlfhq32jYH5kPbD5
oNc1uh8WyfQoLKC33Q4m9HbwBNiWDMvFIXg7ECa4rQruslAi/ycXLdQ4GcYI0F1l32RbNhFTa0yP
G49kQIPwIWXQy2ZqcAhkgaYKVjCrpEsIgPphQaFaWiKXV7tImegFdmrBFG8G0D1EDibe/KjAg24r
wEquahAdEHJhaLiiV1qqQDd+gXTxuAggBLAhi+OxZAuSeAskByr8zU4QM/X1rLxS8yws4AukuGSl
oppilURMnPw1ohAXILEMo1Yp97lRS/VLGWX/sO8wKZowksifyOghkyE4PiPsVSrbEznN5TR+f6ih
7EgS+xjCCzTtsFIe1hnrUoroPs8+Or+FuqnIOt5w/N0TxrcDGoRIMtjnMcSxMv7nFxXl5kRXZb0H
uSFoYvbWFCK/HX3CPUrmiI75PO0LXgkJzooGzhJqzmJlWAyp5Dr4jLMV73MDktqLn3ySpKLFcGM3
FO/nlwR+fICnsTL3zzlsnrFyOEy6OpeiBi2B/DugMSEK31lXDxami9XlTzmQvgrH4vM1TFl5VjNN
Bv6ZCL2Zk+uZeiU7LE5jP9fHRZB04ZMoyxcCTamL9qDbvJBtwpKF71SDKgD1NZXvRPxeXpoJLaGR
G/CGjfJmd66GiaQkDK5p0Z4HPXhsIOWL4ZE4aJLrLw8ebFyB7CTKC5SqbjlSZwH05dm7cUtY/640
WRUI47UOUylGLaB8vlo1ua5s8qgg7ecJJurMnrv5Lumt3DERsXpYCQJOpUkxqQP8vc6StzJBFtBm
MgoerDW4qNKGBErsiAYHxLrwwEUAAc2ruMmgiL9hWYqdvyBtux6UGfq+s1c1m4m5CLc+5+Hf38aW
S35wOIhKN10+xVu+tTCbHosmx5FsmlLUk6BEPz+Ad4hHA7YJlkJuOrD77yDKtmEBTsO7iD9PCR5e
tHE79jkF7/pxpFFUZXFDA81f/uyQWdyPHmUJraip6sju16mJjbvkoXIUBRPatVRsyj7RTTah1WyE
Fli5jAvsaIPnr4f08PNWbUl/rVScNoZZLpjFyYq6fSeNL2uuUCTCNuNI8NZ75xK5c8xx4XzT2pSE
QARVb6INDfprfmcD30dufy+k030phw8VWdZhHy1mer6xKHQCbmGwo/ZiojesXhe+aAbiqicxjvlf
Pbetmwt46QF2TwQId+bamNo5J6JtFYcwxA2iU0InM96Ly2BEjU5ZknjOlJ0R4FTQt3mJgTKFzmhi
fnfgaeasszZL9Bc14XYS6ltd3N50xC0AxsnT3Kc+V45eS4YLzHx5xRa84V67XuUK4sLqzqKZPuxp
oNCYs+0Or4E348OU9109v3CJ+VKx7ucxBk9u4g0jwi5OY7nDvXYxnsJqQvpWa0IlfjT0KqpGX/5b
CxlZkU/RGU6j5O3Y5KgVZsNHuHt1VrD7VvUlTAnWDbSJsphCQ8bUoAzxigtbk5VRLi4PliVuCNFb
gaQypg286WqVxqT9Vm/Vhx5LqpmRieuFQ79SjUV1sX2l2Bfl7hLq9OsgAEwY77ym5vhS6SVB+Y35
NQwFw6ajK81UOc+U6sf3NEE72tDQO0WaNzmWWztxckVYBA9yMu4N7FNTHFt0lTTx6hehxyq79JUc
s0houvzQ5qodpgTHqhN3AwGaxh4ZkyENznrEi0iFlfA+Z+LQJ/ihxraZLNc1etAYayIAM04BN5I/
vAsFbf8HcmUETL3LlsxzqjFz+zEOvkZe3zqkkO6bpcAGvN0tXz3ev2tKjJcfrU7/wWIoh7eU5oql
UIiCvjmrkc6eMS0R3A==
`protect end_protected
