-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iMt69RozzLxTjSeNcy6nPn/8xcHpivihWL5cxSt7xAIy1WPgg3c6kRTZfqUKnLEY5yMETDIgifeP
xQNaF6HPooqg+h5fQnDXhTaMRxdGOQtuNJxeattFb15M0Q0IVWRKzsNGHnbsBB7gZ1zw7inBIOZu
qVR5EzxxseKVNJfPe34farCrqLEjBENjDNKsIXZyCgKdLyFDw15FvIJEG+hm0KjskBpwGMReXdmJ
uGEXQWMpNLOsJZDKUL9xdh941sMxDLjnjTJP/o+wAKt9eBvydZrU5w10AN2ritn5J+a0sn3YCEH+
3k/x1m69RLgJiPiYgLVNthsc94tJqdL1Q7xbTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
p1ttWNMyu6vw9U/VB9CPSG572vAnnmPJmKIihIFUSBF2Sxi+cIPifFN2PQYq9JvYAvAc0E3dj8In
AgXS4qTlLLGLyemZBfyh7bsonZ6imfa2xjHEqsKJoO9wpFzug3Pyw7c0EPVDbUwBWIf7vwvvsNDp
53sHyNZQoNQFZ6E0a+X8HthwBSxjktEDs7KhbOjqY+xi+I8kcatgsMgZtI3jmEHHaFFY2bmoW2/n
ge+UzT1BpU9ppXfn7bSeXCoTf9xEEETMH+XW4Trzr+hNhTRy06MBs677n47aw1Gn+uU8sVjYi9ia
Gaa1Zgg1UiLeoCKAQRq9ekaWqko10DKcYMOtycEhCXTcBEEXEdzYCpvcZho04y5ITHyLIuMqJWCe
MjDkjQs+kFr+NnI5dofuOZ4C4hcbB+nnK57Pvn5gxnoLx2OH9QZa83YAvDs0SaHfvRG3CFDrbBQc
fG2COntuP2UDTnSn6o3r1/DaC9zsqRBb5GKW2i9dpObxYNgpHescG0/b5pDtL4B5QCdojFvApJ3J
bwcEEk6H0aNim0dJsRwVQSXc6sIUy93OBw0CHby0IXaELOkEQzPBwpr5i1/dRii6MsoOar19rWIO
iRZN4czd+9shq6d00M6L18OtHeB7nbfttfpRh5osFsgXWRBtDLYlzUhYvBQ3YQcblo7c04mMFILo
nWsm3GGBHnlCL7egwJfxBUeC/c6SmGEMd5QyaokcSatszpquklHjYge793P7O6+lACiUgO2gy2dx
YwDYvsd+faIY3UBptc3NtfA913Z5RIsyGMVOnx6+BX/GCRHabtZ0sXVNGQwXH5PPFGrN8CeDqGrK
/BP0TiZ5aCgb9fsNU9X+qPTCOYcjwGRntFgNJV3mqxfbF1ciC/nIbC4ODoiOjkh0WVN0NCXwiK0g
gD+cgxEAFUZvMGg0RJO1bdVhwlQYlbz1vl2g3R62AN7fLlx/8Kv6N9cxg8Dz1JrV7pel6AD7L3D+
l7rRemkQwuULVPGvSEKTso+zRQp9SgFWsJGkjm1xd9XAiJoUmjsK/ySQ2sj1ZqrHCLWJwmaBbzUs
4DuGDzvZ0NY8LfFw1XqXYpfIr7Dyv3S7igD1j3Wlztaqv0NRnVT9U5u3iovZydong7lpinYHHgOg
oR5NPPR9ZH/un0g0aGebukL9GvHdUlVANcZQF1hOyHvT44UXqzXsn21lT0mi5hNx2Ny2OcgtBbZq
sGIe4uPRNpMwSxwE8QRPisBRo0o2k5U9JAdwJYJBgEQh0fqQfN2H4P2sx8fNdsTGimCVYIJlTlUX
/mJZeyYrJpNLY68q4XDke/5Vr8X6z7QjIJNHZqPeUel6nPBuPuf/bIdcS+5WzSANIibKpXSEBvzB
8z9Ed7evRsOy43z6bVYTqOtsEhM5MfrPUYB+4/GT1/P4AdV+8kLapQTJ4WxwMMNK1MxHZDukSxFh
3r33TLjPKlRQSS+6FXCYDeRV7tNkJQSCHD0pnaoX93KUzmyZtj1EmJbKyoDI6AZAsXPkXpGcSS3Y
ZWXF2q+jdIKsyaCe868QAvnvyv+ypZ9pX0hPw/0hFIOXh4amxZnRgS1MDGF4+S47g9SxBy/NLvYK
mOCO8iqTVsQQzqQn9J+UDfOMe734izdExjj+VrzShadjOebUEhZYCqM7vw/TpdhPVK4T2nXfhtx3
NEDj4Dj1Qa+795eQOxoTHIH6/96VEJ/y7yRaEm7fBjOLIvSNtN/fONeBpgS3b1lJRYWRRlTRNcKB
pRAfFkLcV6qRzAH360F2HAkFJQbbS5ZN6q898aw8NLLMR8MwfvVT9Dy8e33TxcZQe8rtUO5WjHb7
N2HLm9EK3kyZ/wpc9jeo659hy3ufR3i705DY/tkQK69G1H2UNVzhQ40Q9OKBRvyPcVNFy3ZRwg+F
pGcO+gLfEfXjbPQAhsTttXmrwYRp/4wky9MAKljUl9BttL9fh0mz9EjTL1py9XbSZmIIfdiiM7a6
uS8aoLh3n8tgB8eh1yWvNv+ylFszFsEUdWc1tuwAb3dgA2hQo/Iy+HLfHjjL6x/GM1byE6dVT1Sa
ORlvXyal9mJ0a9EdkgaMsLuHFrg5ThyTg5APGh8kms9FPPQx0DQKg98optWc0Jk2ey3qyLToBgoX
p1Fl7+S/EoIiFOb7K6/uvsnZyIDXDx3PYR4G9LkJ3XWkR9LPoQI5LpgvWPyfpNdlmpZiGWv3Z1rT
ApEBfX1FjEYROXPJtwQD2KIW/SuWaKB8/LFcfrJ+96JKdaRRWbEIzsNAg5zoNLpEC4/ogWGAOcRb
gwcnNYWsQCLctUL22H/uizlZjFcr/Cx3/S7dl53i3neg3LZIcXs9NFba/h1Kjx9KGRClAGI6VNfX
OIZ5Wt/mpTHGjkGgkCKC/iMkZ1DEVNd7rtZNLOXJk/AfHojeMva762BHjqlvd9BLxq71eWoVMoTZ
eKzD3OSzBB8dLIeUYyNiFz1UpUa6zl/+sFst8esgQWjVCdGO4xE3gGKHz0ZH9ff+ePcSz1TgHRrr
tq4lv4ob4+uyRUMSOkyZLig0649hS/T4IWX6o9TkW2TEp8wy8jJ+h3o3kAzKQCZPgkJG17wTTv5P
swFL/2Gbczqzi0EGsOtvaWu27JHBa5QvDNNPWCFERFo/vyFdhWmGB0NwohY0+PLyVR8k4My/K4wT
MOjAEacQooCuKkqrz6LarAH0iODHML9rrOdkCJsH2p7QiJ2Z+7YMD/R6PXdd77F7q/BxkQn2ZVL9
HcS3+v6YaFqXkXqRt/7KKDjLcCPvrSAwnPqCaYTaYXqtsyJh5XD4iJXtl9ZvRbF2gJy7ZEg6WyQB
2/qcYeh9mMHxI/VIbVE+b9nK5iMKn76zjYVFsq7Ae8Pf3YLcrivfKQa6DEpYa8TAIS9pDN1xWUQQ
oYvhjdSDoFPPLDUqn6U/8iJIln6I8QBLvuxw6pM2t2ES/wi3aIU0NX9y35zrUwnrrHK0UCrHNcw8
OBX1nzgkl1l29OYz8V2aSK0X9fq+JH2E7nGJaN5FI/tfe2NxylJIHDL5tutGUcgKreOCd6aqc4VL
hYe3nYkmnjaHe8lL0MpA0FKThzYGd2sU7DjKWmzkf/+3aJvu+vFkn7ioJ0u25RKSBE7RKJ0c0ptH
ph/5dJBvj/NafGwOVKxbGMtdMXcRNw3Qu0LSQ760/Nr9mjdfLkoDrtfxuo7RVjX/D+BENdw+9b8W
ZPIBNMZqNrkgt+rk4OuPeuZVSUe6AGjRszzbb3AS2zwnDBq0Lekoxu8sDPNWb1ZXon9XK8MSGdLT
W4uo5x7MBA4KnPA0G3SBKN2SVJPr4AIGyf4qvTjKT2uzyrmNCYBV7LkXjTB8FBX3JBS8F9nKixt5
EHL2J/EeyeC+7VcCpggdMiDLMRQHvVKgkOddmkOYQl6PptMxVyjaC1VDJDfC3RFadVAoAVYGP3xw
yWCvPZ1/WgUaUKJB2V0jJgnw1631dSybqjxMLP4qwxhuiBus9t4QhUU7Hzux8ykqeb/ZIXdNs+j9
UDMqEHFYTF+xjV5nwxQZZFSNbUQBcplkEdQpYjzuZQvvqzT+Yp3VlmZpsLnfxqheyH5ke9IL+IeI
gu2eiX7QhTllDOrhnMqw0tk/H2AQSjYUu6WnNU5ZAeslzE7/duaRYziqvNj0NQkGhp+jO/AvVn/z
OG2k/IypqMUJ3HSN+rY9TH1TqnlNAD3o/GcSkiYf9bpFB3xQXt6N9A8ENmw3psJrWymHdVSnA90Z
DEtjLWl+Pr0kOmF518Rvk5IIgLkoU+mO66nvVxzqLWG8y+HngElFi9ywwUpFHgc9dof1NxA/AJsA
N8e9Ua53KvwKIALjR7m2An0VDJ7SCEuT672eH8b/ybCgSxPGQSIoZX6gSQVWsRaSKnZMpROhcgTy
GuPL4Afu++BjKJjkjdwuzxdJLkFlehp0JYxd8lJFmV7XmDv7/4inrRfemCy4SAey8xzR6gbk86zx
rImp/pP3LIQDfhpZAjJSKLErz+KLGJm7Y/ny3GbCY4qRUD7Qrmr6MDpwhYR/55O8Xj8kfn6QjSvb
SLAj/VWxtBVxAZW4lW787fmYc7Y1JcwB6M/+AtMf4cnRdvQRXKswXrsrdnyflpt2BVtWBRB83/XM
pQ79lZTC/UmdOcLaMLUz/s6zcNIFBlZnEaFxm6gIGroUZ0aE9zQBPu3COKk1Hfk2eqZAX1ek6xLf
91vQAX6PQwVwMUJAKe5bDs7z4oaGMM4b8BcTZaOdwiar5UY11cOCe+aguuSXSYZP/Jb/rcGlZTTU
+SOUaJXHyJftdLITGvflD+4pCDo0fkC4Ju1Mw5GHaivKmgub96Jn4G2a5WYIRw/cUU+tAqcszFhb
v4G/EKYmoa29sj5yjF77d+utHkqWtjJaUxsopUZtY0PEbCtr1VQpRYkM7Q8563Kx6GUF8xRNf8Bc
Xf5pabBOlxL7lvip0Ja43AGZf6jrABPj46KjljTyq2TfVNkOw/PU1XR2YfD3E/4hq9FN/JbIw8n3
q2RcFAORvF73kEOhq6kwnu0F+hnaS4o4GgSBFiFtZtgI5JTpNr3gh/+xHSaw+qOJmppJbABvpw2M
SXxMG9bO4ppoB4jq/7GIshNT/XF+bGDs1YZjhztu3XGQNsKkEOQt8bWplaWvezupiPbQ+VY2Gm8K
rUEjmQ2bVowdY+5SX8cTDaQQeWClukir6tIolclwKiHovryvq+plVPUEhjYl1LsyVFLpB10Pzm3O
QK6g2WDcNB/Dtn3V9rq9L6C5iOHbYY6X5kzkZRsy0H3wZsJspbjyFdP0XwI5ydidaBNMXjJf5SWI
uphP/hvGeSpcG2Eb+DLXL+WlD1U/Br0KXCVdo9lin6Ifj6gnXks/l1uWiQ4Ys64Aofl7eW11SfMc
od6ihNItF8rYCxTGULL+RgdhFVIHqqfsV6TcscGELuAZGM6s515rLwXs28IBezDdV8rKqhnmBUIx
bvLeFEpo24L7Mo6V+O4qRhp0DuHPvBjHrQiIQA5ELJYj/8a2qEsXlNb6/XPf7ff1rT71DzMCs9QF
IMEhC7mNLXSoRQcVAITs9RGkgI9My3h17OweA++9oWQYGFyQCG7kFF+18T0WOUhdOOPHTMdfak57
KUU+2oPXdyFBEHNCe5L6hYzC8LVEOUhQxr/h2QG5SdBUMiel5Foh7tDLxcwu70vx73vGyycc0xII
5uOCcCCXRgo8rIhI+tcpnHJ3Ps6tCURwN0LMwWJnVOojZx9dFWKn/FoHGgrpKzyQ+FUdSLWP3nyK
rHHIc/s/B4cfHj5idlYmncNv7YgNk3ySYamYWo4tBseoesRVVN04MqgmYF1naGd1j50LqS0flooX
J8g0rRXfj7OqZ5EaBo4t7XGtai0HwdF3EjeW0s+iXwnceMypIFkCRNHEM0CjHFLl4Mr4HWe5my48
sgkGwiRJokYbw9to/LQ3isnWQNxaXCc/3aCWI4M61zufpG0NwCBldRk4kKmV46gGwAAVT2jwcHwA
sVzZhYFiNRfQ36AY73Rdy0i15Sy1oWAERAe+QztLRLR038Yujal+nilZEdQ1kbq7VUjX+xYV5ml+
Ws7WmOlw/ZnUBwZbzeoPc0jlX2wZhDW9a/eh3leR9si2GhtmREtYu37YrErxd4oIqjQI/yao4gUV
o+9Iy1Kt7TUGEQmkLSyptoMwHi6bnO2Wq6pq8d3MxV4yVTC5mWDbZBvl86ybQjuvVCXMuWCuaocl
Avta1NOgSvDIp6Tgqfb+0eaf8wsCwBspCtH+tnk7nkMGHAQXZoGuxg7/VP+yGndx1xLS69Hzunax
ttuZnzxPANv0fR3QbXlWzxdni4pY38ohwpuEpuV1ArEgkbSxzucqgSZEIIShNJgQVGaMV1VykRpi
Ik4M8Kuz7uY31hjESPD+3ze0Cl3qq8Dqx445uVy1WGQecbarhjnl004naM7mpiA++kj6G8bAJ2YL
BgvxdOEjdsT9hjai4NYSDLB3I3eQfwNOtdIpmT0qY33RSErWirZUvO9YU3v5WHwGbBysczc9pMqh
Iy4BNw917sST9j0CkOxBRTKLQpWUG9j/5ZyxUT4nUdJGZHo3QfgXFn66aX93e7+FdKimjjgdK3t2
o3TLSfZTlvQ45aRkl52BCahNP17Zgh0aqqcqr6HFL2prOEknuzFi5ohrcXwze9K0xfTj4BZCoR9m
JTBAsrYme5qdtw09Rh4U/zHRwB4ZnCkswZFCoinrG6F9eZuFG39WSOOivhMKXmtSVn9VrVOpP/b7
b1Pcltz7BZACAcIAR8fJ6urp/Ou4sfWlUrI5HtjW+lC9DdK5Gw4JZHZmv4CkGVEPu6UMiFfADZnD
xZ/zcP6Cc6EzUE6U3cIKHrTFJxdfBDydmHJFu4HY+8Mrs4++viQVeIQK3vg2iMd/eoyXOXJjh7rx
9KhIicNTY5BU0rUqXo/H2wJJcWrYss02Z6PrM8vh7HToeOx+ePByaK3i0uwXAbxzcGxGgWiagsae
nKJ2n2hha59r6H9QBZtHkXqgTD47AaWVkulBKMs0QAHtz7oJWwgq2IUKViAJ/lv+dPDA394XUvk3
tkWc/35t6LeGBvoFT1ROg5WsoRunU45Hx8J68fkaHQs78EJdAS4Oq5F5bK1fsmAtm9kJNO7S5+5k
0IJC1VpFW7N+Di6DDqys3sXDDVjck3PZzGfcVI3Rt5380v1VWCZRkNRYfY0MvRGtyWWRq4aRhAff
NH5bWuhe3GqT1SNg588MqIPEtbqEcxvA0gMnTf+tC+0HS+9mT3M3PL0e/v0uw3iZ0nklrq0/JKZ2
sc7J4hPtI8ojZ+A/tVQ3HLSZnqQ2Uc4fpXvSGC3pXJshG7UD8epTM8NkpxUcAx7ByhJRVJRwSH9v
pp3uViAgCGhXT+HtDbnsUqIhwMD5balmqVqPlSNaTEHGxKRvV8JqQwrtCl1lrNrdnQJkdzv0pfQ+
X33Bf3xdxu0xs0r38fWxhUHnBtvEmwqOUWv555CEvMkFctZF2z9go21lq1Tj1bwplA90ymrodx7h
Krvx5YfZnlgEnqApOyzxbuvnsnO/8aw6qT8ydfZN4tqN6X6JzzWK84cmt/nkw5SYCz7ovFwRi7v8
hWtk6QqNK68WGNY6USSLf3LqlaO7gvCSx0EObULAtZ08bFcbWXWhdaxlvYAegJ8W7MDu88MKWKv2
d+3qMJS5TBGEzbVIJKrb2lrPMaR/PFUdpgZGj30HeCiVDY4AzZhlzw0jTahuSxtgCSBFrKu2vD2w
q1Q36L0q4EOeXF2O3nRYYNmM0p7xBLBjA1iB/Gno1dQGYtOgE9Vba6HFwMu31qbEezBNKgW2zyQj
2GJFMkCvQxgDjsCD+YxyzSuqGeSQ1zTtHWdP0ADBPytddQ6o7trKrdNAiBUJ+aw+exg4StGPoxhp
pxqFIQv1FCq4YF751WcnIFK3EoGpPZDVka4u43bqESPuIuwPqoBfhRxaBml8Rl6bnBXRng4wYeKA
z0F2knvoh89kNNP5en645u2aREOZhI4vjnvNQKPu57fSFIIhNlujFqjmhZYr6AmdYaqNp2Rw+uI/
MUaF6Xkr/nr/OeDLxT6uASW7wdBF+Bk+xVJQbqw5gMPRiaOmijWt7kSv9tkSFugR7S+0ZKY5vTj1
5KoeMfJ6ug8OmREu0xA5e9foYFKpPWSvFAiXq4/tDG+FPhZ2PwUOwWZZ5GKkxqhk7RHMpZfKDjlh
Wf2idBw7uc719s1SGBioectdWOxaZEi0NyMd8+gCzE9Fem5aHJcHz8tgUKtC6ct/J2I22B1Bp6Dr
M5rA6Z2d521p4OxjEXqvY5qq4vyGtqXJiWtB3tmlDbjmZYGmruppIIPW3xS+aZW7Tc+CfTV+BE+/
K5bSPbVGnakjgi6iCsgXv8ohc35FfBJ6jDLpbdGebgSJ8SBJnDUU6wPVg6KxCwWszpMCuwn+lIZn
VJ+zMv0sTpRuvd6IKF5K3HiRh3Xdf3IVbamZbY2sVI9wYFgRYUkqemOwkjLndhCdcobIFjvQ+PFO
mjLHNw0v4buZQzC5uQBC1rE9jT1uZ+dMw/Q3OTIoujjXQhkjyf9vEncl1kXmqf43LJscUrfK7SX1
4Y2jjP2eKU4iEn76EmzaAR4AxILpnknAf1hhcbxaPD3ojF3lu3xTZG+yTBhEVq54SVBxyW5CX2lD
e3XBELzmluqeV8aYbMxzvp6HSabPSs/2uZZrcFN2tbeHjZOKwlGWPjRWPjW9dDnHJPq4/xyZF44J
E5kEGkmygViSJMCzRCRGB4L+k3hinCcVlSmV+N/lHNmb1az+Qp4R7gKGKCIjWd8jit9igE34srYp
zNZ+YgGuaCJGKacRvissoHTHTBq4b5EdmUae8aGvwvKZIRkqYjpKqXZttGXIU+V1hQtgEHONvxTF
Bowm0ckfsh//ap4WioTSgC2bckED4aK+YnGfCwNqrCUNFPZ9/3oZhiUF7/iUohIRD3+yj3VW5IgN
69eBN9gRnrK7Kyn63Mav7AVIoZ0BeFTimtdlL13dJ60IjDcoua9ZkgClesjEb7g1ctdvVhGUInV+
0YgUYqOABYlnSeYpIdgnu053wZzifxDoDIORgCB5w0/7DOD6dlvnkee/Aj/a1wLzLPUsicDDZqCP
Amv7Vg1H+LZMw9Db0hfpTZK9bHXMdyoO2FCJ4XX2MsOZvc++5tOhPkEcQNnOPOPZP1DqR7vg/hN7
aYvkiaJNhhv/tHTONDWM5zXJmK/jfxqbRLnDENRJK6S4SsgaENe16ruPk3c94REH84uOk5XIBBrF
ScIefAa88p9tYz9U40IrGBui2rIhrNPpDwdS5o1wpKdMOA5atPKao8ep4V29to75wZvimT095QfC
QFN40R6HWys1Y/CEJ1BQlmX8TTgreAGNjNHN6OB/RHTLd0V8FPrgMvpdkj/j4dZj+NjCzj/5ZlGl
wU6pDxR8K0KqBbGcTm0gMNhaI328gdjWan+OMbbZrcoF6NeDQuo+qQQ+EMT9l+CLURyMA7p38vdS
xiUJ8iv3NxzrFaeFHBiVTTKdHAb3Fa3E+9lCbsm5/EXhsrNJ8oym3zxlU1kXy1OL0ATf5MLkAtPW
UvMd3WsdPDQID3eqnaxtJUND5tDfyE0ib/wywCDmk1Jwe9Gdh/4Lyr3W9UY2zFTmYTcheNEgK96l
Dy0qFi+FlqGTne/yYjkNtT0d8ggmaOrUdy23ZRXxLaVmTZeaHUJ8xTiEbGYN0cMMUQiMuZhdEV01
5l4yGcmeN5vrZtCesz4J5Ooi/WAG5AYLZEQm2wpCCwLK3A2sF8TzG9Ief8vtVyCU1yRq06P+VrV8
HwMC+nTjS6Zp4AeMUX0Va7MPdsK2PpWiljGqPRuukO6YSsXJKe2DjwAUCm7o0s+QP3cqQ6p4S8Ls
NpBz+obxZH1nkrdveRxxLmw4px+yyzVhUXElriPxwW1NEbXvKELD5LC5p9VZWCb8EoytGCe/Ol4N
wlh/JovRF+itKXsCLHOCLHzdQDp0UVYusP1Oz46CyJSy1COIRYKoo+fCuy0LsjgUr5qW9lGNNY0q
bMyqojrIotrJEaat0hSDVdslpGw2pKTEpV2r9JemGGdFZITKFBbQD1eFZPIiKRRsK5DYdjpZMBId
6IHiW9sBBRDVGeN/QLqkLRt4u+2LidU6UTQ/oRXBWI8PnCufTPlOnNkLX7NQUw14h+4NgclhJLKF
YppeRCbkM0cDo7u0rcPjx2wbVUGZ05Q/s29ksZPDztRFzQJLx6m8f4KWRm7JDaTY4HNS+zP806Z7
9pEZlTGESL8ozhTLtjvZh+/22fHzjGYr4nOjW3og6Pu9g+Hq68KUNq49tYV6KzHrq3S2CKDqTYqj
207fZI3QhECyfsrSL8nC6Z1WPY2KecieNuH7lV7Qgi5ORh9bzSAmBkBycO1KzHN6jRVCDOCv0tSs
BsyLjPxcysIogpzl4cbk3nmEL8f/QfAw1lRdv8FUhO2ro7PPUPtBs4bJgJzJeBr9iO+Snur9rsaS
PPYbCNa5dlIipK6ChjsxwlRoCwPJp21AxTB7NisiL9ODd6KnZGgjnf+nOmO057CvNVne8LICTWg+
D1W3aL/h/KS8fC+sX75qMiRRL06CYaCIVKddthK3UFalcPpf169uOjf8jy5qvTTvXAs5rV7hwcCq
2xCbhCKnmVhbMN5XDU8TQNCywHfZJ+X+wdGFMczDhtesXrh64k/E08lKEdKCzksH/B560fFg2wcU
xDAUexIiNMZCrxI3co6LtVGfD1802tvhhwUfTAQB/YjjYbByN0MTBaGetkUHM/RmDBE7wcCWzHay
j1eczFPw7QOCaQddkEcWoDsQV2ICxiT2fFppgyk6tCz4k5MDaHRb6tyPyuJxz+GmvriF/5ajHt2D
H/Cf2fNNfikjKcLnAgjPnFKgCWE1kBMNer436qMPptbZbrC4oOpJtinvYNAU/O1/BQhUFh6xMmpW
BLpPf8wdj7bwcxPBv5McSYO0H5xy4rkhiPhk+ysiyzrs3Ki0K+3XPVQczZjBvv1ThFuRvBQoScVK
tPhy/u+bf3f3+9B1Bwg5famWhZNlj9SootTCeE84S9H8zeZsEPC9vW4WsHahf/4VSpwiPiDchVZA
m8d9DLUSiI8q44o34MSVTUG6UmsPrpGpI4m77kOvHGYk8wZKW369NQXov4Qk06Qsg0j6T6Sbpjuc
TuxqMKFRX+pRS0U/Vj6nPZsTnZJw1rY5hGUzxgNNmIDMYehO/h4pjVF2jBJHDsTwPky++U9oyJDz
UU2MXvla6rd28BfZ8RBi7qk/2JYmeeBAGYxYu5x4ZInbvr+3sNY9h1CeFwb3PVEd/3OISnw5V3Hn
5xtFyUHSs6Z6PpdHexnmQuan3xJN7o9BEonKmWLVJNqBOrluB+ybM2MFGiufDtfvOYrD4npe4lxF
9zBBgKZgvGSjsxd1X6/H36B9gbx7c5P12/wIlyhM+D28sc1RVO3r3Ed3qRcBWGS+Mg4larGCelOH
eQJby7A3VnuvZ5qHWegZwCVUM1ube4X4HlRy5vJdzHCUJhai7GZMjfto2xby3zCydOwrLfOEQbm1
eDgcjr7Ed+5ZLNDqFXf9o+yOGFHzqb8q46zPSfj3lZv5u3HBphXPC4QYRBmh4QB486xTgM2GEzKY
8Qkz/3SoHe/szHFICvUlKshe2Pci8VWsmMddgdbRPtpK2nNrFBf+2+diLVzFkkRnE9y/IY2Ku5ea
RqV2L5IhWbxvQLFl83RbcAHZyYGlZ/rYsfPZtPrWnAL6tAtgwjDp/doxBDuebL1ULP6grYhz4Qbv
Gjcdu72ziwZRsaKj2fF8C1aK1W7mWoXfOJYD8vs8wjcsi2xq/bWbB3Hzgy1V3uj2Vmyt1N9ZqWK+
HPFgY4BcYqU+LZSN1PKbRKwInzEBEw3yeFBuGrELBQSP3o6E/BkfqW0VFMjYmYHuhZs6Osb5yAiF
bWy8ciJ6bjnvqdxSHVskkPg9FVyDbe+VkoEy5Rm6jz5FM8MRmIWpCTrt/qIGf1dA7Bjg8UnTsvsh
g3qqKCCDMcBTpzzC9j9VrXAjWZ0jTQb9Wouz9nCvTGs5eC3sUpF6w+Cgfp3hSm3CGmG4IcDaZo7T
I2SqOg8h5EZHkiB8+LYmMvAiG1Xk7+kpAHaqMzVc3+nmLK+MXccVNlsbKYv627yA4IpDmk829xbg
8VsXih0co61YxGCsVJB9eZsLc/8km9j2yulfdpPkPHLFPQJ/wNteXc/AQU2jm4ln1EL3zT/YRyE9
gJ8j3uOM4quScYxNU1QGgF7IIv0eRkS1gHFBc8G6VGxol0zUukM23x/tNTFNcFSQL+wy++6TXVLP
ZMiGbaUACWXxCHJeCxen6L4oSmSsZU86mVQBX1OUkIPrnurkb8Dy9rvs3fogWPxhyH39umXXPsoX
iJOFmam4pT0RUiW5g9+87Mh00nidpHQn6U1mhxtV9TQzZOOfhigHDlbMWXpn78kQegjhpbWK2ZWp
r5oZV08hUUwG5hbwqbxCcV/nsri/xf0EbELfeNlWjisgB9SBa/wnXl+EYCjXFCDT721Wu4yr0TP3
rnB2XNzseCD7thPnoC32yMF4yJ124zlFJ+pzPsBoEa22mP5muEYXS7+FIagzoRm7uI1j1q6Q/Qb6
RJm4OA5YfPVVF38yLxZImPTOLVQcZ+kI2rNDQWMqVpjQDtBZ/tK4HG413Vx8Qc97yDejGKyJK9ba
B9TdGYAFXUyatsAEWYoSPkpmvRJgBe0szCRQi1mQtt1N3bdIiXzNEW/iaGs5Ks74pinJQTwxHsII
edp/UQgKzkY+MjUxyHy0YXruYdzBUJVUR10X4o0EJ5sElzQYspoheQEQ5x82XPslP8fOOIASPyJy
boOJ0jEygyhqp3x/zISyOHpEHV/DhJUyF7l/neKm+j5VaLStg60xk+GscyWXOXEDxRN8pWoecO66
Iz0A8kPQqoFM9CRlZGHGBfVsMLHrpPbBpt/C3Xg6YjchYlZbXSnVtIwMHl7ga850Pd43Yezv7UnN
xKaMy5gz89s3NkSNFSf4Yt6q+43uKpvYkhq8LHMzoimtM9SoYLnYfMb1rsOvgpxqfWPoJp57ZqYE
/cGbPpieP73fTl42h6G0JHTN94E3ebsVb6Nk3AfTq4iS9+DNZqUpOVoSGWdD39f2/Zdmdprv5JV0
NtLyzlykyqqosfuGfd/R5AJfvc20mKjFVnEObcIWG+BFX4tpG+4AnWBNaV+LT23Sa++KKxMfnUY1
CBw5l63KgXvx7nDS7r4hQHsWwybTrCe1oLVINK3c4krZG3j9zXVEgsLW/CdmkTs1sUE9Z9x2n4m8
MWETH2bEt0PXrh+siq7x9ACOwoUX1OpDkb4XCT7UzBL6Fywdq9CmjtU+k9ysOl3VerDt/uCSHt85
+XIhmYYRdcMnaY0oThjPyEVRnPCPPeESemllHXs763G+8ZFsvH/9pLd/fFKjlYCWN2dpJz3zlV2i
dV8TQnonZgiieqMdrdNdAYOPC9/k3kKtnBySpBJrOStfBLQ1K2HsRSnEOs0NmuHaZPS32geBl9DW
k1HHdMKEPTyf+UFtMNMtsy2EyBi1KNbqmdMkMIiqywmlDGPq4pstk8FvvEnzkWU21znKzGUMWcV1
zBCJzWXsJIJokTg4U8BNdv7UOzXX+fzHp+bB3QAv40/eHcvoWGGwvB4rY5am9yVsmuDBD5h0n3wg
VQLqdMxZI+6/G/jNFD/8eXCMj1mGAKPCPnf1c0+naeXIjGx4zKl/+LQlIdyQQFll9t+xjzgWHfnB
rXV3wK6g5cBYx8CMRrUtaGoe8iCwu1mdcMom9tgOKeWvmUrqRG3knRtW4g8a88r6HtPqbVDoceRn
J26yeKitAn0DDb9UZAV+bt5in5cNsi9i1mmkFVESkWfDMKecrSJgPv8K3U9B+Pn8fRpJWiv4e1kR
kPthsqXi+XsjjYOspXRTnkuItOMU6N++oofsFvKtJb1wWV8pRjVL/s2i5Djk87OLwNEoBHiWh8Cw
ZqgRByp1uBQJDndxs3J2E5Tr0ZvwyzSZ8PZPuEgJ2T2FAOr/SyDBsipS4KMldINjsiN0HelSrPSr
prP4zNfHj1+apJSWOsIBoxpxsBjrhHK3NxYUqjC3OJUOJj5GssyBPVuuHx49qC2dnxBxPAjURopP
koOBRf48ihawLiRWezjnWSxoMCcoP3s4OHDQvCTJoR6g7IbHgJagCm4h4Q1GbKN2MOln0jhYw2wW
WkQzPVR95Xx3/HfNpfhb8wyZ3WvJA99bGVBz98j/crAsr84P8qYloMlHDqonwWclhxLVJQjtWzre
iXwOtELRHdwEeDNdCaigGQcRswaadPZui4Z3ZN+30WGL0dVVorIMG/Fy/W014yWu6KgtjvPXRMBK
aNwhrpklEV2BJeYH+Zq0wCpNBIBNpUizyCHBERKpSliepeNVcoy1AGhCcARlQGUp1UOMaXZrBoZw
8ysgDlrM3jRLrO0iEaXVY5LyoYgezNLiP7RiUdVuCKVvEh2hk/XbmgtXv6F0k6PTek7GZoGjFCJz
bhHE5jjAiW+P8+YCNKfTm2UGEfFnJlvsYdufbchBsljo8VWQ1bnkHsgkeKukkIL5PbMZGLPvPBTn
2LyVE0esb94xydivLhfjg15wV6xPh90b61oo/pvWNEBnLebRzpW2LikkOXttzjax24KRO2Ynbcen
zEN6b8m3ezTNbjdYuU1JhnpITzsC/5I2CwfnlEfbcTakSipKXHMpiQ39ltyy43OFnZQtaTLdQ63s
vRLzhMjw9ouXI3oLo0IVYeyTpEFnuvpju5Q58UVrYbvO1/Mo6EbmLHWKow6pgihcJDAzARjQ9OX0
6P76JR7OYyEnSLK0GhpA8zsMPplLymiEA2SDofio0MTxubbXs90yHiOrQoXvCDl7mylSdjUtWOGw
rr3dlrPDcE7OsSXIU+hOQy8UQzPDsIYrQLN+gaP+1Dx5iY9lJEA3Zo4rz2FqEMuSM3XnaF8dHg3o
xlZQ+vw6DJP85v+Qxcm3uzSZQCJ4bmCmtIWSUrq+caMWC8cZ9JBQ8qBV5rs81ilIXicGsp29nZTD
sxXK0FTFHd7wgRK7Mk/lKIFmgcEzNFNuIB3/cenEsw//IKbVuEb83imIiFjjXIIaEPjMWu1n2K1w
pIxaY0BFX+XdReBKQvKOy/gB4qRyZzejkzwz/slv79v/IUz1+kZE2Gf/UcGzz1QN6dRfkTPnX8nQ
j6oefs9boLDMFtQKzNtiVG1XxZit8ibC76WL7wU9yZZ8OkPIYAuqyPMjQ9CFvTLLN1tF25VyGdSB
gV8rHcHo7506ZZ7dmYAYVkCvg6ygDqmIxqNqpsYUFMj6oCvoxzVZlwkptd1QjwIDL8GrigqZjU3r
DfLM6aPV2KRPSwXf3Q3eQiL6SI9raJ1y06S0Gb8NUR9F0cKnOyW8HBTRaYtjX5zTPpYil32PjPtp
sUhPSXs5ROrcQRF2QmBvUcIw/O9m/1DVJY/5LVT3aPg2Uu4aTIKhEW6RbxZ9gWQYzb0+MZ9v9YOd
10XVL2/Kb7xCUH48/QZpWk0JHqbu5tPfPqdj2Fnurpk7NO40B5ErAJVZpXlgsbXbNwdGED/CwzW2
8d9vX9T1huDbVIzVZtQ1o+QR/SnRlEkiF5ldt4Tjp47ta0MX10YB4tOrANwP7ogsPAkaZ9KTcAzo
gT6NBDUb/Y2h6huqwSl8E0FY5ERt0cfwXob1wJ7Q/xs/EAi7A0+MVCiMOzks3lYXtqhse/UP4lG6
f/gxD/mFwoOT1rr5mljoRShOGh5W0wOJURyKxiEEegxnNnyxEpM/V7LRjpg6ExbetgZZpwq7yCWx
Rx3Fpo+eFLCxSllFt6NYOpjftRrOsDa7CzSkBhAfXVjDy9pWVIdBBd8iGBOyyAUDHwmtW0Q+IWIY
JI4dcjhpXc1QTSiojzwRkHTkVveZhdMuZUaocQrEHoGw3e7tHlox3LV/tRshxCywYsw6KYqTOkNR
F5qwgq6bhl40WhFsMAEh5+faaFfVGHDaSvzWlHwg2W0BA9j+r8U9uGIZxT0cJBkq6EoPV8TiB5II
ryyMTkc3WUvqYF9/v4NnSK0d/cvLuy35X0WNaxDvP5/KwNzTm40/Rm1EL+2xQcF0tmMNAqnKdYVT
Rl5UBM+eaIjiTo5mOnPXr3OCirZxG988Mt6OJeJZBKUyfck9Cja5uXDx+/cGTV5OO5UwRdIQHEuw
1IM0zAIBOpFIh8hFTaQa1wtDSQ90pxl1HH4qfcAUrQNgzw9cJxmsrOGgKAULSSQz8h/sVDdmF+fn
ciZRVN36e9UAWEolFl9rJUqDHMYMGGQnvefvOtSitSXl8PeE7ySbpc56Q9ykVR1r7BoMmqSTAO53
j266+xh+8FQX1+eBasBSFmHDrlam9xD5R8GQTCgL9XwnI0d/ZY9PC6tC2yOfk81DGaHbOKKAxWbk
tCAaKG63V/Qab7JcSH52Ega/gkJxm1alwE1w9t3ZMnZROUMXFv0nCz3bF6jiWxElUAZIhO6JNDG6
7YpZDTDx7iyo5Uj/8c0LG93K0nPsV5NwpzV0R9ghqRjaeS6PPyvsG9Qqm0oPPp8jhQh1ADtaIHzV
IOiffPsseR67lFYMh1Zvmxhl96PHDfQIhTRo4KJiXwvr9/imzZHesi83tTjdXy0u4I2RZ5yanuj3
bBPkxiFSO0iVTKNO5E8SDNJx7PNaNmtT6cegPHxOjCxIk03oDwHM/XK9RBER3aT900XV21fdU41t
sUQjBS0s/ir6jpsxce0g8gOTjBNff5CNK5dW728ta7P2hfzzYtHsCM96OtAiA4d9TYsoT7poc10G
LAeY/LXuNsOxYGMyw7FzgV04RAJBCyUDzWNnB6915+s5+tdSh4qcHVBluWU4oK8GacbT6Fx83Duw
pXxKStFcZnV6qT9nBq41SgK79dMbeDUTf7pJcC7HT4Rr2MegsHeAU797U2iHZRyRBxg8S8e3IQNl
2CsHZ946ekcaeVJF17QnjfzFPpW9AAVeJGO7BXNGNP0VAHqKcZ8JW7g5JzJApJdJC2MNDozNeoxv
w4BgUY1FjkS1ymkjhsHjHymf1mfabujccfmQGW2G+91xPhoRHtwx0OWssdVXuHPFI0Ai3WYQ3hAo
0i/EztZUzuVffYBAHJSrErIC8U8RzSw+nBIH7roNAE9ij9+UNg+hnW2DyWf7WSS1gul1D5S4jdW2
FlE5GrDlq8Bn4udhYNDc3qx6mkDhNWzdB0Z15XYJzXHJsap+oSci2JSNwIwysv5LZraW46hH9kk8
Km7TVrsCQcvpzxuu8ifXGsqjVl13dbQBriXphSqk7TiVMson1BfyYcllNyBuQPzq2qG9khy7dET2
DoewezGy++urVSBslF7VyPZL7ek7kWnlkbL0s2LnXUT/b+Z4dRHZYUVOnIvWyRbAJjUjAxXn1PaO
7nmSXA6niX4LaigpOp1eE8SdJq86iomxLOVxDdChfFuuE/mJWmLo24ih4DVcIt0cBzNEsI/Q6OzO
97THUHLWEaspYaR+GS33ctXgvk9AtN7Hm1NBdYQLMO+OuHfOb/q9eu1dEh3mJrOm4ClwjxmivZdo
mZ2/iFXgaG1hiZcpP9BaPIBgKw3KZndv6i32W45b/pA7yovMHOaiHAHoBn+asGEdkmj76gFgPoWI
xsUMYPw3DaHpX0IKSkt6Ni4Oc7lzWjbyCRbxRRTisOCO3FjC8LEv+slyfULNU7UL3ozkRbv31QQG
47UdYGXzkZOwSJKLheOFGxH6ULIg1VfDGND3CfvKRlMOCJUFm8scLIDLMHIOwzeZ6moLwWRNuwYj
QsS935w3c1NZaJLqNQomH/85G1GN5i0VAPbHeSa+iSwOFWzGpZDfgQPeFyPDEQK1LlzXfBZSk/dX
AzAwl3eqEntE68ejmhyjr283II8R6eSDNvNR0t5vAf9Ljfp1FPKdiUc38TxoC4G6L6OkZaRB446s
efB1ouxFoDN/4TNh7RwB1XMS9BgpXs9SpUoMFm4RPHTyVM3I5StylIMihIi8m2mvoDyZux7WAHc5
wvNp81n3VuVdRrTp220xsHFPcKxof0vxDvwKdL/3F0UFxDKE1lqQesFaD83pZsyT5+0N5oK+bZ/C
09WFv/Kyl51ndre5Rj6YMNHUYKQu6mxip34iOqCBRTFT9DzUvcR1VP+9jeaC9Xdwow/5STMMwjFh
h0m0oSbVC0XBVELetTLPKkr5VwHVDwR/N46LBARxdp12KB3nJr4kFlMW8F5Uzije4f59S4QHknU3
snOqxg27Q+HOLYPkJSGRdmwEGJtNlhZVFnhMLnEeSEwZprv2VNfrbxS3FQrx3FL57qyiiKV/0n5I
h1+2tuemZqX9t3ZoImK03VGJCGjO9rHp9y19E52oEIKux2PMvVunoFGef5Skt1JDuUmTQdYzFl9c
FeO7PxNf7Q3tCj7iW82MhP3IXTmZshFDBm9t9KvEZnMZLu+SWwtqNrXYg0u8R65T5fMpQuoCFEOq
DCQx048yVqcJi9HEsmRDbATGPIwxNQrQTaDhRnm7LUBJ6BT6PXGBaAjYRHSd/U/xaD2Ho8MdQUz1
JcDJVsdc1K30JEO1sOk2x6SHQP059OShpuKrvztIDOjAVr67t/iGPw9qFYeK36UbC8KKfwMaWI7B
CdfMHAmHf+1gkJwGxYjBNsLpG5rapIazYmc4k39vBSpAfQLqAJzzrEi1P0wr4JNXHsLsnZHMlb69
WNJnfUxuhXJ/HTKWCNxwOmSgMKx/TZxtqNhr/Os4YztdilEvSYptlucHz8Cxlzb4VMaeDbtWJOm7
ID7DHLrrVHneVwRCMrj2xIBGT5Zj8KeIFx7kgoQ6WDPmzbk1piGNDtzmFQlDHzpH94oAliwWWr0e
gMkd1asb5SSy7y1IN7TH5QWE3qAQ/8tzBHZBehgncJ1MLVr4mgoDF+NFT+a6IStah1It7SWyeRkz
kniz75JhoVB2S/hXIHFNIbeJUrp3rxyNDLbxsje+J+h3r3gAEZ8xrGwDZ5W9oA7df+9n4/bxcZW9
tWYiJ1gUsdnbhzpXVa03kDetP6E1IIDi48Y/5UVN/ELD/bqF7mNHa1zw5lN6a15eqGAppWISW94J
i81uJ/liCSuTPLYuCjIyyWy5LobLkFVW6NlHq22I5cRByQ46GfnWdBHPLFbg5k3MPjlkl4R0jwDL
u1oEUVvlXWfgExoFZYiFmfCHI6ZD7ZSV8fSCnLqbbrpJ8b/1ZDtGsB5YwFEJVXVQgRcsZcQMhEzK
SV+FeGUyP1tefcpqD7GEGAgGOKziTLzo8nwQdUpW18ScexSavxpuU6dc50vXkkQ6ynx4eWT2Yfs5
orMML1IU7/r3idqXJHb2+UiBoPlactesUqaLq5jFsK3j6GBozu3cazIIIpXVFyI33cHFjxoqUyUh
98N16nqBHDYwTkUVPaHqJGS9+oLPFKQgTKAOsWHDO4WAGVdQrxG/QpipQUoTMjbICY3OtiN/e8nw
P1+/9SPtPe91mitbxTtl2Ljezy1CEhPafWqSOzHYLIZ0+7oxMndOlIVIIpUg0VbL3Wv5yhbBK7Va
O+72o8HbxjbUGFNsMBCP/A2rKScEEKwSZKQZk9umALkeSQCbltMs51ScbT75wb2mID8KH0I0nnev
5pWuqF5pw+w/x5YpIJ3duBEcRUMUHtX77yUs2wauCMCrNuMnaypZ6a0vEdU85NCRmk2zsnEb1gKa
VFT0fjzRp6xs+cQkLDfqGOSJiPnso73rVu9bqAA+wweqPUVrMbSXJOMlZvLNtKsgFbN3NbOsqjmh
zrz6JoU+GFPym2vvGUkTS+eLQIHc4f8UAYf7UDcYYlmkr80UruICJpXhhYj/RB0ExZzHUaFaIIbJ
dNMZIGTzUP4+OXygIa0xZ4kjVT+Bi7+7tanbRT73K3qmWV2JZZkMI4m+sEciejG1f+buTp7D4IFp
hBVK2+f5wXkeWl9cBlWseKMtT9MRT18ZG3/xXsi1mjJ/yQyU5cvEYKKuSnu7Xm4noWQBmCTsfwH0
mpxoY797J0D4XU+li30YxDyKxNCNf1sE7sw0MiLLhnodIdhH3TspEB0Vo/GWOBdWSWFaZ06dkXYz
7UstF+KFROW9qS5zuotGoMBphf3Jrf6ljkRMLaqA/8zhnAjiX/Ybk4AVXHcaXZKkXqzf0ZN6fUhj
S3UfGgg9CcLKgxnZ2EbT+7+g64Gs1N/PAJfCpfZLteuJSeNJUWCqHuV9nwQzDKHeonjnUoRWOs+1
WAsnD7xZWI1auK6nLyeZJ3s+ZgkmdEDdcTqOeZvoXDX+/tzD/SHbKIROAkSUEDdsAlDu+rch1Oh5
CUeBKcv8adD4dFd0t2Gz8HW1n7B0hFTAfvLhg9Fo3E8OizVE+9e6OA3iS4qPtT4kq5gMSbgjry6z
5+zqpKf7bc+sw2poiFauIKBO1eTCj8TTsGQEG3vpVnml/Bmlu33Pg/evrzQ/uWWTd1XZEWyc15Mr
sb9WxcPVzblr5VjGkzHuO/4h3FuTQL2eD7/KruyrZPWvLCM7UmGj8PDyHhtKQNX0RsJs9/hza1sQ
rgQoI0Kr7CirwyB0L3/xTJ1i0xixByVvJoUoIKfowKtMrfYq7jrv56U+9WPjZYy06NVH/Mm2vOZz
NxzP0jIA1sXq0+9/9j83W+JV4kiIROtIlDSDq2c4gecPmwk6uuDZM4lWsUyoCQ3erZs5ooQQP4PX
tS/8WvaOvVYGyCbwfm0N1oyTMNET3g6YNvjwmlVNt9FCWW4ubDopIvPi/xXUfsldm9jn0CiiF4qB
AtVEqkjC75hfNB/OKsAR67rxzVoRoiQxInSQhzVWgCBq6l9HJQb9fB4qpEEt0g0l99vWCiovH6Bt
PZLzRyopibPnNw2g2nu2TMj3qJ5V6LFFn2KiTGA4PPX0whdpVYxzwOGzq66t+INqxP5QVuGvi4Oc
QgdYTLmciK6x5+z88lvgmK+qSvGF8X0i8T9z+oyXxXmREieDfUAuU6PcfXOzkn1CNtmWcRSoCccf
Z3tNQ6NyFJuCQ6FkIilql6349V+XKq0jmlOeCatqxLIOJ0mEvo+XQhc27Ijrdm7VLPGJoyMLOZiw
t2aoQFRjoQf791/fSlOGNEMRVAANYJKGQGlDufCi1piCK5sRCtTv6yWCYkvET5QC/3RCvOaK3CJM
GX68toyCjsJ+4YoWB1R/Q2eCisr5g57xOQSJuKvrxAAa/PWxm6A/HZcpxDWwCK7bQ+4gPrTuUszs
TfvvzS4Wcut5PlCcCv7pPNa4YUKjQc9v9G1sMtX+RDN6aGEeyw96BrvNIxl3nS8oDpcChiFG7xgP
Kv3EkUsUnoQBLtrLB0qy+rzwf7ow3Ad7THEZTnJZMIucgNcZk1xzXJiAIZxRqnk7aYcnZBv/n0hq
KrEhcfC/WU9i4ld3yX0XWFDqIlAulDrpeS1v9RPi8+r4PF1Rf7dEh6GLLrkfOs7mqXIqXjqzo8SZ
53ErKgfCLJbRwkCfkbB9HyQhkKNkHYMixC/9P3vq1NdkiaUUxJQWRdCcYJS5MotcTTiQX/vzTlFe
/Zhbe2424hPPB7/5TndjXOYAto22+HTdQe3/P4j/NQv38bLZlokI26Uf6WW/2PPZ2lCZpNQIRHmB
+3qW8G33T5l5uiyFW6uZFYO4V0DpbSrvKPcrmfvWi4cg1Ke3eB0DC4x1nL2eftwxsrSd6IMOsDhr
rWULiYqcUUBbBl7nWSeqR6ggQ8i1p1stlGstRLGy5sM4/8vJAhATNXsMlpBF3Lf2lDN2/IU2S7uQ
361VHC+426cNgZiRYFa00MZFJj7JoF3DR9zv9fTWIcqe/23UTMPmusfh4dZdBMwKFIpkKVd7J8V5
qAN8A9YFlN+cK+AvvBMnd98vp/4M82VoWs6LtFnuA6TbkYmQ7iGpzHnD0IFzx1F6VaZPhuFcgDyw
JdynwVqncQ05Nw9KH06/LOvnCurQ2hwlfLQPJIGgzKFEleZTroSoXBgmgx331BP0NDhoBD3LlT6d
vjZvkaNt61Z7ky7Eqzyt3dXqICRPwvuTjbLCMNcd8bQXn1xEUdVCDmIL5TBrD1eER8xGQNnf2J/9
FnVg1C/KodGFV5yiOnT711rnBu4/oCORb8mFHDatF65N8kNjMrXpHt4cJOzU9G4QjDe7RYFH3UCT
2oNCmF7hM6IkFWBWz10qq8YKvEP92lPsSgvBdQTUQsDf2rrOZSS8pkMQygoo7bEElXyBxRLPMSxP
x01Zpg8Jnqx/iW4eZm/HTeI0xTi/mPMoMlziJS0uw7KBsIwH+lGn1BeHF5qZls88OjQzwkd9HEJI
p+xo8qDJc+7ZqeanbE5gUpeHtgNAM+sPPYsCKJCuSDoKAxKnIS99CuCSmgJF7dpEU4S10veOtER4
p3C6U+kBkZ5pBgjUqTc6/dvkgFM5T+tO3C64UosB8q0vIj/TCkxLPT2DzQq2p8i7kO1v/FcGvgkR
QPdSlq2uzOI4iwFFB16bD60ieavVYBIv73RCWHGqQiFc5getDbsJ0GG6/4p/of+HrapifY/xD678
lkToCodnblWNjzR/7hoE6VlaoO/x5wNV4hFxwrqlfTVcD0rNNLxUlI2GlTxG3qamA9xdlemCEryg
qWPF+XOtpmra5FbWAZcCHvbPujFNF1WmTDsZyH0kHmYLdAXr7J6vbgtyQ5fHZMwjeg0HQK/7zAyQ
J14AJQBZH+S2WVvs3b8hOTB9eDcDAcZ7SwjrpH2wdzbfMTxB6FBNYds+NQGemstIxepiGZnppFeN
O6ug1DFt/+JTOFrfhUX+X3Vs7r39w05L+J2uXGzgpjexpw6JU62+DAgs+oIrcE/Q0O4SlC08O63m
WibNoQUdMZQbRw6lGYwA5RV24msXCkaYnU8JFMNpMA8K8JZ04W1l7CNBFIBBsZjwl4ptsHGvt1a4
rXr9kQdsr4aOteXj/4G2D2Paoq4dGMeAQzt5m3A08BllPFgWb+gco6QfRU6TGlwZ11Zv919M+fgz
nAm/9JrgIuxPREjVttq1C9Zv4aETkZo5pvSzqucUR3WDyWLudGw3OpjN+gqI+966gDwqPdmJQdEE
zT+YzDgeYBBeQusqhP2cpCM0zO4QpCXyF3ydxA/nDSiLD4k76XZBA80j1e2v92o/0lWstSfPXx5Y
exnbKWNkP/RjWykWH8W2Z5UwBejXslBpI5M4BvKjYpe03GnuRRLXr+ZXlBQn0r1yJzeEp9dLap53
7pzqPbmotM7tGsO0CgsCVSyrxzpr4qcA8fY+Aw+Ncr0FZJdX+tyUGW/PQ5q0s+gKmJAK2PRqbqqH
tIcewTpyiHEiQLTeeald39dh31kxWLVPA+Ar9u60yzYcKUXEiIYNqpQIk0TBRY3aoCSgq7SNEORA
scuN/bJ0cfXSUneHERP/9QcpADGee1DzmKcVbx7lyn+G8h0q48HJBXZd8WSY99IM5vBh5NyF4HB0
WfBRPKquDSF6vp2zscYDh/pkv58kJvCdDQ2u404fwHooGQTgOCpCBwa1k829JYwkvijVq6BlgFMO
CcChWMzAlETBQRTgWob85yq3/HVS0Ry/fsRqy+hPtw0fRD7g5rrJYlRsZyzPah1IwtZK80EmAFE4
XjY9TGnB23DthW1WWYNF4MQtsFhG+DCGwGDc259LvbV7viTTjTSbsqhqOsWv9VHVjlR7aY8V7yc+
2lpXHl3FM2OWHzTw+FhD6YI3VB/r+5YzE7fwprKKaH7KTwtI5FiYEdphSUTkHGxaC0MYx5+lNo+Q
jcE6KDl+FJpyFmZJe6lwaU3xM2TGxxkEoBm/8FY+buwJXklIz2yAzdA9aQ5eX7tQdwkaRpTugu+B
OUHv6gaDRKkUwcuxsmJ0fGKic2zUQI2wBuxL214fH4dQ1QumWFNWlupDt1AxckQJ0l+uVCSpvymE
lSdthrQnNiyaYKodS4hLslVUEt182edcGMyomzTzcWmuFvXYCvvOCH/rpQ1lDbJtAuWVXxpYgFN4
bFxdWV3bvF4HAFNr8VYMHiYyIgF2a/IEyo//c1cPaoojwLqJuEu1az9VXyhnnZknKyg3wHRnA/o3
UqyZ8sqAd9BnfecXan9U8FFF05yybMWcyv/Tm+8GnBMcJIuHlypBC2V0mebgrDaMo8yT9Z+huFTi
KgTwD2cI5mK6IJ5Ft6wQ4fguVYYPXbepkA3o/drKSzKz1+FRc2Knxo/rH6VU5GdoB/T9crevVhca
t09rOogomfMWvxeayNtvvyalz2+tggmefzU4VQuW6Pr/+oe3W34B2F0Eb+FKIfU6xLrWo55kkFuR
krL5qSzNSjaMAMmLlmgG91kGACMi15mfgDzvzrKJ5/Z6jYEs8039wBMqD03ro1+jcSs35owiFgD/
5RoBwj1XefCk/cIY8nvFEzXpBXrLcFifpHt1gvAaJGwD/fjce6AhHLCr1nJgVLqQ3N91pjR41jxZ
9jrZRoYGo5rTR8d+IN6hkPpyv0uwac2JjkhORtWP2HexLHBN5MeK4zVkefvz1A63FoLIiUstYelf
GGnxtOzbIqDQ1/9SGPo5bYA8/5M/Wc8CUD2I0gAUh1uoIyfFZ8xXzfFFQkhUfqO3nzZJzipE8NYc
CYY9RbVVey096WoZMPvTLtEiN0f8wqXbkNZsE/QoYDQ7xjJtdAn+FCBoO+280HcoWwzTsLl4hluU
C3Shd1+ceWLMV/t+Kfj5iaih/X/I1V/a5MoTWcJNIc/0cqOcxc1g3nArnrRjrs/xOr/UU/eHGZiZ
q0lTS6ERA/vLquXboCotGi9pY+RAGZ5bv0M0q7yhXBIyfKPa+/FO8qXOEp5KB5atp0OBeO4H8Nn7
FMHd/kr35ZTH9ATKwBukv/jN9cF3AVKrl9v4+175GzqmJGfhO+XUrkkGdUF4PKDIDaiw4fAFFQrD
OO1ATYbAnLYMfTrgHZ/XGfWHBeR/I/HfMnEjeir8yCvqf6XhFLaDqZKt8l4Fg9U8CkbU6TRNphtQ
q9JLFCFvj4Zi1RolqiXRV8SbL6FfByH4ZE4DCy8zA/cPq7+14xtk2npeJ1AJVFzuPKpkBUSJjgpQ
XMTDodKlnbiehZytRVS+PnRzptMq4tiuieAX7gYBXfjXAqdDBF0cU7DYwMis2mjGW7PUscAPgySv
xqD0ME6JUSiO2ubplqX7If9U9JUzjWG17fEy0H4CI++hKfvRwTv0yLX2QtaU19rmO/PURDNPe+qb
Q3cWDgBcXONfUNFiig77i3azBG2R3Ss9X1zyACjJzkvoViQkN4LOxe1zjQZ0LYWOyboaEGfUAYzr
Oev/vinXbelld7J6p3nKT/14lRcH13xS5VFDcpPZoTs+Vv640xYKVoPKrgJjQjhdUwfKlBkU8FPr
EP7eELXxS6h8CjzZIYPpxYUc8wrLXXzW0jLeCzTwIls1ayucFCMCrHLkW9BU+OfWsPkHWizT16RP
UnqSKtI5yv1LPAjOILZP9UUEOXL1WvnMWYt/rXs979oZvIbDiLrjJKcD78LLlClyTQyjli9bNrQa
rgCb4GV7MQMfRIWOk1jW+6BwlD7IcICKk2G3J41Aq+S49j3sXXXF40FxFe+iYWpa5S4Vl/4u6DWk
34Sp/9+xraKAuWAgk9r8iF3jfzuZgxz+W3/MGwzjrk8M7pGTVnke76W2uR4cBerOZTJ3BAu+zK4A
96VjAOKTZhYGQHif9X9CL50Npxkyg06LCPDBt2WMyO+KmfWcJWa0B4jpRv+EK8NSPJ/up18A13d3
fiulbJs7iBocEQ1TqJ+XgraV8gP5KpXhgswqgsueL6m7Pl0+VGlIYsMgkX4EuMkWSfLxjz31SODZ
ddQJNMmwJpMML55dHrxcVe3IM7FMqK8YQxBRXKA2E5fhyfnSoLIe/J9pXO9UUnRu2rylz9Cpqhs+
xoWoziEI+5u/Re/8m38NeRJ3cgyr9EK5DIc8sf4fs+fU0Lp2p62CKps7dBYk2KkZIuqdlDNwUMbV
dcionZa4RSWvhkVKicKMCqykMw8yhw1hxL8ZME8XtldeekcoER9wAywVhz/BVrY6Ojq7BixZttm9
NbpyyKGUme/qG1oddDXadouNPf/Edt67YzIr2CrqCtn4oQb1tADB+/QwODSLRVUKsMZBEkCH0s55
S7ReH5fmASgTpoCRX1sQnbGnsYbWQ8siDGruUIWkrq7b8/oII7L2dMXl2je8o4zssElRzKVaSpNc
37OFdcA4ys0iyGfjZgnaaUVomVAAF3ZbzpagjHXaal16oob1SyCbJ6D+tcT9MUKmqCyOXaeqVmaK
XWf5dxOCOWERPTgcK+gG4o1Im77OGEBg6XsVFoOGL8NwpmAeuMBl6RI6AJfBvRlx7eIbMh80n4AD
jPkouaAilsduqRI8uYNmhTn5NywIWgkviawwoxoUB72W9FdVoTHT8QHYScEUz3OMPfZe2K2Fl5Lo
7vJVy7uIKPlFSnuSKMOFtYJXNSiD8GXCTMPetbFaBBS4lUj6+0vGlT+48Llw5im314zpJkyWCo4Q
7ngxs8hZE6KxJgbEIuQcihMQSPWe/9FegS7yRSlDp1R26TSUyEUmQEyDZad4VMDfoNTEW1zltWOp
obMOdAjmAZ6ZLT78gZ6WFgIrIZEnGtvPdylmesH6tzKRMa1HrcRBhwYO38DTr3mQegECSoyT6Wqe
QyS7munih9UkuohFs62VnkzjgA2Y0MuqchEd0zF1bkivwpPXWWBP+gyglsbzAAvOP8kDvoOG27kF
lWQ0PEnQ/ZLK/LUsV7v9x/uVXgL9UjAh1gyw5IwA7JVonvLFoSz/4XZ2mGQQAW5m4oVMjJFBecNi
C2hnAe07o5PVWWsD28usTCGQANkA6prPwFfACoyXZYWZwjdsXBBEvls1Snc6cwohMafIzh/NwkXz
pKahgn3WtE0D5pyw+4Kb4tNKg9GdAcj31VncLdPlvL8VgnBozk4qiNh8xh7YzRf6kdjz8Tusj8Tu
sY8ZTeWkbK6L4RKjMcmQmjkLbPZ/4o+dsRiFvRWQmuFzx88iEbEbcIofrbvWUkh36CcBe4sR9qwb
eygcu1DlRsCNsK/3z01YWa9Gg7bSF0NbzrMhA0ks0PvWOc3I2BXjfEPGip+MuOY+tRFh9f1L4bcl
ytB4fJZoUs+zKMOr5zVEybPAjHMjZfl+r2V0Zz1aViwwtMVTNq+hPWQ6E5apdocuWKIpKBkpvkck
oUOVajuuaUIzkXWYdugINHHx8s5+5S/Fzuy0lE8MeRCWvtMmHnTZBMP2G4Ah7L5YADbg/I22vJ2V
lS5W8mBhXZLuJ3ZtEyhNfgYgYtOk4mJ2I4oXVcDdTSHGtq9Bcr5YlAOJhuI0coHsqy8pND5vPQSy
fWIBmxkHPjqxkAwzEkZDt3VWZvWMTfV0l64JD0KnAQpZRc+z6LD21RwmXHAVWUD+fEwEuaL+lDwo
P/C9K+x/lu+dEQ65QfeYor+b961bV0cqqHyTpl/N+C8BRGq2POQBbyxcL8VVQJ4q1ciWykFOe/uc
a/kHqcnes6K3NXQtmvfxi3vFU8lmJLCbm+XygqnyGPbN5eyYRgV7giBc9nEj8vYJHj5pKUEVq/2l
kF4vt3qZsOdyabeX6hzLSqKy/hOcu3vwQIoo2mJ5RcfXfZCbsBU8eGhDc++kFuuqXvg+bqUm9Z+V
nGnRe/7wyfDnNAdrJblLSQOqMJjqksYFpLqTqJ4/79ZPFnr1rrgAN/quDfi9wbi7JIAPYS0Vlmi+
z9kbPOuzLA9wRYavALoSjGzvZfgOG+vNeiEVNyocHATAtKrhxH/Yn6Vc66P0wOz3z64ovyCv10HJ
4twATt5yIyPTnnm3Ey44uUXJpXZatlQWTa3eXJ3ZiznLbIUl2F2mfJVBNNa91ke9aAPB9yhBakMC
QY0SDgBKs8rXCU9n/5XKH47z96Szy5cf/qJ3LqDS25xV3ukVzDoYz9L3YsJvhTc5L9sLHyrihvQK
STgwDW320uWqNecZwiy03dqgINP0JYjYRIhav7dATEj0455a9Rzh/80mo+P9J/Vy19Vwx5iCQ0Kx
0kKP5pJIiSmyN1X4X60hWGc91DSdLg778S4K2wqOX9nNzyJUYNmHtAIqhdZ0u1zKVMUalJadaPO4
1YgbDt3Nd8JBUuKuTnXbT0oh8FX5VTAipOW8RlXhMg7C8v2SwGSkyQNW3jDQXgs4jNsvU5H6lhRC
5fBfNYfkqdn+UFe619F0PfYc/dWuFN7/ikYgWcsx4DUhmDEdOFWfrTTTz3gA2ihxpBdo3eaDqsWf
7ZLUDQjtXpYIzWENNe8huUA23xsIS9zhlgqHZIXb62xwp/gDsLO/b7gb3Xa/Bw0uBPcCNBs6Hyee
Iu7cqL0/p00YmQ15mLc8TNRoX41pD+42yquG8m+QiInWpP9lLeLjov6TFKf9msEwrnIecgsjwaue
UMBROfZIDpbkmKoLum0jZcZY20Hck4T3da006xE7+D1OYi/+IQ/GyhlS27t5HW3y1uJy684rvuSJ
QiiQ4rOZW5PB0urYBKsdbYaWlLENolAKryXmuM/wqfaKkAIbQKi+OyrCu4TYhuV0wOFwnEr+BKyt
KGE/QVx+bnhI8/u2QHj9aPoTkHjjH2hW712A6Q6KD+jP/OGjm1eT3rL13EOajOmJ7CBqomEUiXXi
fDZg8jBt3Vy55K6/Wi+h/9gZvh28GXepGnbb/NwkHUPTnG/X5IzjfOaL2n7JFPazoTDFnYh8CvR3
dEYGWVZt8z1Y1RrwYwiUkekjM6c4uOTl7xECpbUaSAHCiS2Nqmqymxm5QjmABusiEu3/ocA6k31k
4b3xD/FEt5KPSjSTSc5+Bj/a9NbvEWdBG8Httlldclf0967xKkIZzw20hnkyeq6RWN7FPzX8yku9
FBMp2UTzplYw3ysUQfryDrDCDv7RT+SMDKPljpBrcZiDl6l/5lORaL5xFsWYzsSgjDzdHYn2heiE
xxfklwg7xf/m+mUIGgUB/GuyHODSRH3exT1EhNEaVV/kXPatt6Of1c0pooOMCjS0XkH+fduUZebk
/nlcSfQ8D9ITjScCA+f5E9g2cgbHm9vkfElu/ULdyY2u0krKQyAMD/h6bEhwqCu5xGdroNIAnPJx
iPtj96OBCLhJYoR6WTNAnycbjoZ/1c6d2m8IBSCMQrNCCGIYhioNqNHulCGkJSg26y2xoj3XFXJP
wgZNKuYvRKndg7HbyWSuU5e5xzwxv3xg/mwkp3+qD138QgiMFkOIeiEaWlWObKekzzec2XDC6hoF
/zVhiOv/oL+PaxOVSlMCrlitqlYpoekU26tIufrjUIvLJM1ZlYpOukz1NiOY6KNJwJcRzKiBF3/n
qw0UVL5gyG9kc7uJWEJ9779u1RN6UZwmg9Bkw5ZMC40BQINh+lZva7xZ6fuZ2wMBl+C56RDbKf26
FntIbMIrDB7o1B0jacWxFgtVN7faejEuwa3ZYpWI7ObOtLh2gGql+wQbSpZ1EHxDbEbUqDorBhvL
kj9Pv120+KNjP64zNfuOpSNqSlLLxf9jMFp3DnvTPN/+54YG5rhEOahjdPfEVM2d7PvjQpC0qu6c
bIOW1uPDFmupl5DnEVjvIVomZwyfUgQRYRpnaosQFC98NSJ03uUtDllwCbnwQO0cL0mrHOGhL6xX
qmyh5Spi4JtyhCd62fYkA98+EavYKUd69NPgs8fNVu4iSyzCTt/sw2TbMkPKPCADL3Rx/BWr6cla
T2F0gk7MpSO4dAIvNIeKIkOH4wYQRWvz1cwZmcxs4h4MUF9OBRWVMHfItH5KvTRnvCp2GZtHnwhg
nuqw43KWnAYNic03dZ0cVA3Ukt9aMWeBOTIAxFhgQED/IybedgbSCVcn8o5YXwgfgcStm2MJnzyD
nv2mFxXLrb1kqVp/10xHvjG5iidHtt06wcBipVtfaUvhaggLezFJsM7RdNxKgWlnUa3xrLrMXWRJ
s+BgcPnU7YyERSQcP+33fPypkdzK5Y+LRbjKowPk6N/vNYL0TY+dyGxkPaJhHaIbxCtxAFIrLl4L
eDwWn/2P51p7HiA41n3+fLhVgcLTHaZrP/CkWSgvBMmw0tXy+yNU/ApFas2Sjk2oR0jAMLlLhc0f
0+Gb9qpB/JN+OI8iaes+EXzxw0jC2VZfTm2yI2DIgrgo9qcL7sOR9/x9j1EU+QwhSz2/6yua5vSX
aruWjwuWSCIvCqENOK9vrN3TS2O5roGsd3beiXWS0OnjF0rBJdeMWt0WUDUNJgM0TgVJxwHO0Aqj
RF5PphKGNsqYrOfSaRaA51/fBY9gQ6BU3S//FFs6UsopXiYu6Zj70O5G+JOrUY1YoJ2uu2Fzoa72
P23TlcNEfZoAC9Ws9zgtUyrjqu2poAQjATcEp0JMJMnqW5EBuFuRZhBVy5vqlyn+FFmlJwIyiDRo
Ad3OsXur8A0Uw6xsxHCO/BlE3t50wMTvolkQ1dQQGo6+Z8yUIMQAsF0aSBMT0n5F6SoOu/ZD02FA
H1fSFMCGNvIgDweIzAIbdx4lCNHgJ4iPnty3Zzadbr1k22ZXn/U1kbcMK5qiGGy8mSugK2ZwIyJQ
mu+ZYmEVflU43jRudEWFjNIsU8HWwqKepWDWJHoFXeMGaYCci7NQ+Z5SJsjbtkD7yC/VkieusSy8
T346M78l/VkwNQqThWn2rKKedA1lQMHiJogIbgAO9tADhAn8wfPMO5XUQFxA9PNHOLrw2FAo91V3
VOJa3/D8J6yIe9rnCgtbEQ10xVIUw/I8SN5FvPzcq74MSQp8U5v06rwmZxqKqKAvPbdmly4rMO0t
yHXN7/wmS0XF7jnGFHyo2Cfn6+DpAOLiklRT/WgPBXQ9UYxFnCZjaI05fkmSdlWAdynY0v4AEHF4
nNtW+RkFxCo9gR/yDAafppNWZ18fbBMJZeBX84vw12EgvQAiCCLr75H8Siy/bJE5npxCoM52sRBF
q7rlM0zapll+x7WSCSI/i+CqyDLYfze5MjwQg0gZ9t8pD9dhDTbLuAKJP9g2pLNm+vq/5ti7Tlxp
RZAA2ttU9IlePAROI6Bxldh6rHkpDb2GEHrri+iNbl4PwNWh9CuVl4IrdUIDUWmNhsvmSgqrrzUg
R5r8QnjhOlpWbKZbJ66GTAVSiFrf3gWxWWl5wR8uI1KMXIPc6Dr3AJNIvYB+fY/JNessGVub7Uea
rvl1xFDJze1Z8dCw8WEUws4PT2apI/FglbA6v4ItD+/+DSVO1chUEHaLau7Ax8ak7ONiBH1xDAMM
UvPkFrgG6YRBBEAErLTYiIW+w7tV3QarCVcppngZaPg1Y8gfe6wuPgrLaNfPeonlhbKIyg8TH2Np
Cp5p/5oND+yh78CkPkKs5n3Yk747CKd1E/jkikJiTDMmJdjJdOL9g8GSyKs559lFGAMKpHyH8xds
PuyBf2v3In/yZm5HnQUEjZLNoTNHne6lhkOorLVcvccBRnCQUvyDE909TbawXXHHOIewd6TWnK2H
gzZE1Ysc8VQ2p+AQNahYK2bYcp3QlRnU7yjFM0b8rtZgIzBaIva4XATbbvHp5BiWSEe6kFopLQ+a
txIMHKgoSYBhjg0kJuNfrw6wB166OIkZfUJr8jfNt/ZX9Pa4TMNUJkFMx/XjOjbc6XqKvsFNOpDe
UKHnejmYHA7kcjPgwvrMGorlFzIa/ir2PGsCNHD9GDlF+KHMTbaIJinoin2UMuFLsnRZ2KhDb4NB
4JPg2fZ29NZwZ+dRXdQgXMkoMLDTuvM66SLXTYaTnjDHf5kpoOPZrBO6aJb7YJkVnHaoWcY8mp1d
9eiqzRFw4+3OVS8wtnR0SdK1pOY9xJ8G8Oaw5S9jimWk1Zq8kC/JMbTkw/Bal2tPE7dPnSp2f7Z2
LiplQor/OCxhtAjmZLZts/VjrqYqMRiX6wkUmDziE9YpFHgbIS7HphdSW1sZJAO+rk/nKulTuYnE
04kr2ADYmRP9vB9tlrw9YwzjHV7Rtjjzbeh8JYEmTIjJWUrPXIew8oW7NFLomno10kTbkKtR+0ET
JskNyn6nxnvRPL0sSHXqz88BeNfkbMQQGOk3jf2K0dciLm7eZnOHIEnE6UXXshBBnxlvPzikvSkt
6oWJexA8yU2X8cbJ8TDnzC957qavjqxZ1ayoRdqOgiF39gYnZXbEDVnOrbNdufpuJl1LbsgO9Ann
dPbE4hR7mNVeqGaZeG2MkMpvL/vAS6JJi5onkOynxvkNNCqyAZDbdAOzejcYmukv90ivXORF299b
Nfw2pxuK8+X7L8F11uxWxrJ+iKRHc45x75DWNvXGOqxeU2wIP1s8BV4CFGnnZ2zhicH4VI1kICH8
ziKSmczGTB4EE7ox/6/3CIHOPP30tw5+NEFzSuj8CShWfJ9+GfbD06iYM1WPvUFhadGHY/CV5GCu
6DB//WSNifO8sxV32Aq/oQu+5XV7HuNfyVpayHOr4NECuOQiSohGjxZJISzFF9mSeVOhYIfaj6QH
VqaOES/Dtz6yZW6p4BCKIEO2gocKIlWs6czOwg5qci/7j5T13sAnQcoSAUa9XxUlJVUhHRWhXfLP
TJaYCPgti8ROYNXLIxGrnNd5wJ1pkAS0s/aKEpMrEifd9fW5yMHCn9orPb6+RlmfUFLINUfmnH33
jrcaP8COaSv6eCFtm+UvlQ0dywSy9ecKsC65cJec4jDzh/an6YDKYL0uT7XXTuHX+cjYqwbu76W4
KrnC8hFUDuMDtu/V4V03QPDONSFIb+u+PW23zdoNNoh7bEz3GXT7IwkG7ynaDuS47FeWaHxsJ8+B
VXSq/DHSjq53BxZ8T3Pogc0/QyKrQxHCrpoAtiJNUY0defuApRfoPHzSAMhHSBEvu93RYz5J7Oy2
skO0onxfZ6nV2CWi2gDPiVo9iBR1ecDwEdHaaiErv501DLfMDpj692zQvNKL1+0gBmliNYJW83Tg
fFdTH/OycxfSVXQ3ejfvSdi6ACQXBkNSfNy6xFKO8N3VLjdPeyihDqQgcBQlqweKjEeH7NOh0Spj
Zc5ubMbBY+8607YTnlUYhT6qZomQldLnJpq6CZ+/ppqRKYL4Kh80dwee0mlAOpoyiW9OS1Vdtlta
s5PoAlmqo0f/I5tlrTFH8PIwziaWAdPjXESoBNkIXjXqSGNo4OqbaXWbqfWF8uOgBl3axMomO0HH
VY5rES7PVKcrhK2i/nb8PYhAi1gg7NWG+MlN4zOEomqKtHCK21t8m38vl+bQP4n01h+8cu5IiCeZ
6aSoGU7UM0WEtLseCc7SJL0hcel90It7ijW18JAgCDSLxizwzva19H665msRVLH0ots4VytjVAu0
B3ovnOOLUx82gVzl0gBNcq05TGweScdYYbh2/I/uKf2jBKIGgnmB9Mfc2u4pZ4JWCuEscdEAboF4
/w/1fYMkfhIwJpz/XwHZgATDVVaBhfawcZr78kjH0gFT3WZZ/cAKPym25ChelP7i5JBhYSbhtKWn
XNTtOaouavb6Q+AwTO/VwbjJQacnCf1HG5nR6Nei/j1jg1+P0Nwadqk5TSbP9ZwvmZeJfgFy2BWV
Em9VQut7TmsAzTZ4TkZgzaMuKIckvHKkwIj4U/2+76b7Mt8DphEVHX1yId/kgEsJRKWNx5nPZzEC
RrtJgdIHY1ETF365N6SGAsZfkS2sTjyBLQ0bVjIheqnAtgXAhqBy2MQsGL50ATpgxAP1Xl5D60eb
Sjs9xLQPaQnclTmgD3HzVsPGevsMqZ0eAkGhmnN8qZWcTlb9lsYHCUizxnbX5vZCHkU4PRt/8s2W
DJpkxMa9CLQZRWZ4oC+OIYygN/YsithZfnw7tz4qYW97u+PBpPVVlY4fy1FJnIhQS/pzS/QM2NWm
mi/ISwag/VIU1fWyjyfIieUNjAStroddES8bzi+9xbau67DDLR1W1f4WYKdYUc6WUttzw8q1a5g5
8qI+IAei3CiuudVLZevWKYgdIkUcHTj13+P8D83Q9+M2b9JKU8RT804M+IMMC03D3NJdZt2GntxA
907RG2RHVM9YUmeBWXWO6wBzDCLUnjFKXNV6ai3yZlxDTpIPZQeesX+pKcE3bgL4D2TurWmrFE3i
6MffnrVS20tB51Gl1xpnkkMAizKZC8NQuot5dnv7gAp/XlGUDOcIfp0XDfeaZUDdqAKO9Wt5/tzY
bX3R+O8BSgUZ/1MwSOP3O9tUB7tS3x5dWgHrdLdtRCGGk69hYdHKM4ApG374aqlOwPvjkiYx15JE
Kr5UaH5Q1HhNRdw4CZ02qhq4EsHaeYgknSK7P+UHvBNYsdbxLJ9U38qKFbL9Ob+QmNGElPtFaGtc
jwcXc6BhUExj9UbtMJ2XPG4bTsEq0qboaO1cqP9mWcFRAbgj3PJEaO3IPJY226woklvNzA+L0X2Q
XY9HRrzGK0Cf+qe7jPmk1vJzG707ExyDsUCeueqLGzrzWT9U12/fhDaoBv37VRNMDBWP2XatTF0O
ukTV7RlgwclOKBBSaTBC/RLx0sBb9rvvoXx2q0s6btM6IHRPIjFN1BRHilSjm9YWNQtlLPcFe3M+
0Fm2I1L91lIVorrPlZucPiO58+cXQPL4afekLwUbDen9dfd5uYmN9Vy4ELKi4xYQRuK5YbfMznOG
VFN7HdASvAtzPd9QYQR8JGLDq6R9sVEkrcSL64U++4/5Y8jMrFh0Dpyr1epYbbkPMRS9jD+rIIhV
iLtxhxqatSqm1iKpTswUAlNE1GiA5eE8W/eqdLItjC4PbJkCT8MwTl1u73Q26KVfAfdoS19Bt6n8
wSdJ37+Po3an+HDYvHYfkyh+IvaAbfdqOXYKjdiiquY1qqtUxVV0UAwVG0HRq9ocGFArq87m2tb9
hpyEtXqq7Yju3v6a3l4xFPs1NuPfKLYw4ec4ix7fArx+3fL+XQotdVDbil73cVeS6E+QmoCIP8h5
NW9u2m41TzeuJ3oVM3Bi05ybxJ1JLcUz3Y7daT+uH+LJOWGc2fHn7X83lWd/x0uqh0GyVCO4Z05x
lhQRg9torRp/aKgfF/sLvV1rfB6Nr4N/lVKghAl5tXEu1DDQyyk3eWBtZ42rFct3XiJdK604EvDj
Cuac6bUUygpFwO3FvLAmqO1SKsthfo5aip033u/q7d4d8uxjcwJODT+aT3VIs3gnIDhwpLwd/T04
HucBF5POs39Api+ZuEJy8IunP0w25Q6trfsPqAuupp94ZjgoCNurnWCIXXoDUbI6C43+FmnfTHlV
qH/SPh8L4TwzVyGReCeETb2jUsmwXu4CSJcfigp2MS4A19hd6cIQkIQ6WvBYPfMaUMAW7cLeWZoz
PmeBfSuNPz5ayVyat4i2adjZcXItxSHot/4AUM98W4HWl9BPvT5BxXwPJiSGpI44yESH7Ax6LGWt
J5HKa0OJBMDMGeWsKKkdMlh00ByQ8ox0pkhKlGpLKEIJu+zG+FAAmN0di6gKGwKCV/wW/UGTBt93
65GxsFffDDC+xD0nFrv3pJ52KGxAxKNj1D1srmtsqiXuv/7JbwKvRGJwn5++b6wWAKj99QkaW2CM
h6hTL9G2fHfojihEfYD5WAB6VQr9X9RRqz+4if8bO2NB99Zhm4nck1BQi6UiX/EtrZcy7n1fSOop
BYpC4ebNCpnGpFheHLE1GlTvqxTkcIGTgZ7GDAk5rDkModoadMIay8LB6oWfN2Zj/EMHlu1QmDRs
u3ieNqYhCUE/7+DQD9VMCQRvRL+O+QCNTPiYIoL2EWvS5aT3HbGQwMpFy+YS0JK93rc5cQnIalj7
xR5ICR0K2YBk+5JVrqJRYVUwBikwfVO+1+eOrsyxXihtE6JuHYDkp9PoOgkrXTPzA5J6lQZuo/uw
CR/VULKPOU16KFrWywDe7dwdnHj3F/ZLFjn6DS453MZxzdScJkt5bcNiIZOrDmL0qPYCBJRv9z08
DkScYhgDBUHtAmG47smx0SBGW8FcAa2TaWDtlsti26t8kMJ+Im0q/YmXcOblbUkVR26eBDsimHQA
Gii97kBeaPwrS5OzwcVC4SRWbEAAGFDvzNkSQphX3J3Cln4GCZG/qlmHlDBeuF7RZC3JUK7wS1wG
8SQjN0Poptx+HDOD7Xb3rZrheq5kMEHUcjyl/DTKI6gjssO1PEPa+O04piMhQTu3Rm781Qa+ghJq
R0H9rydQV2Ebo4fCam4dVsHqUptH6qh3Q857t60JozBwpCBpEsETAwH8jRYu/gNp/u/Ik1WDOlGA
1PeK1r9ijWN7deVRubUhrdoylWyTcKK8sKthdvv9+vpmJ6GB14WAbiWFjZg2xh16vpUKOmoiudDw
mSVbiwxKTf+dRRhhXLLg+C+bst7auep8J/o+3+fHvNQ1pn7ZIl04PWdJy5LaK+MJPd01VNV2cKae
mBuMLWRkYPgrZvUc5XEPbhrpK83mJtAD4+IKDtPjuWNwuZsqcvyQhwvD68Lu/qn6+bK91OlHqliA
3/qhx/p1Q44P+G9Kq3BysUG2FUxYexRy3YVuek9DA5cWswmZ7cTdoGUsiUe2giDfihzQYQpjWBh8
PEAMdLVvbS9/EIGJk1jYkpa07GZNMlBqLCI5YIt/olUnFpNJhbGdSNYiOpwir6HYLbRDQ3+T9TcV
G3D2+WQJuVs3+ESuBkfWFnE3Nufso8qCwDV3yYs6TlNLFqqpJlsoJoA4z0675+5zYXgspw7HFPCl
sLYCQQjbSHk4WeTH+scFs4ic/JFoSAsn3Uu02/gaXMTSyCffj0j1UvQPlPJ8+PNQUNf2nLYgliTV
D7x2m6n61/jw0c3ovDvGeGUzuIbPwy3mr/Fj5AbkzrFI60qMA/vRhRTgKu0+KdLhlCvEzA2NsmUD
FNQWhUl0ACrdR6+nG9ikWvCUZdvVTh2FmTo9Hd8jUEIGpXWMcN1u6UqcJek/PrSdiTbMJSlZrK5U
CpguWrILw6Q1pzHITWQkCXHMtMKTPglxUbhsdrPwZ7sTV9hlnHTzWIbMlSPSLBw3hAzOqZxfmvU/
sh09B07NZR8PeWhckIWeMd45r7wn6e4PBdwIBwxTGw9AhYeaWJB6a9MlG5DIL3gcUSAjHD9MGGx6
VLwdXvJVp/7GIqdfq9CoOrDzqSSuGbP6Yra/MypK1N35FPrycNNkJXeyO2I86GzHiSU6yxudCxpu
IFaQ3jZ4qbORoPHXnYs0cAFqlqX/4ctHZz/NccqJuJ91YYvtprMEzzkMiznXoziolZkX1H+eCPLd
3GFRQuYyGDlr19oEiD7KICVbp0pEMVJtrK5UMRY/1pyc4T7BIrgn6+HRI5h2E6XeKzdKLdhysVya
LkDMK5qc6Z/JLLV3PB8yxMgjd9IBF/J+du1rmaUheahLE1LXqfbUE3zWvracv/oVOuJ03UKbGoL7
knvu3Th/bm1kguZeOiySYt+9r9GTngyomnEe/bUrkLLj65WJ4Fg0mbBlgb3229fzvZKfqlkx49P8
NYo57CVQqX+SnW2cLPiE5M77qaTpX4uBfLpnIqQeue0t7F7plisI8QkKzjHOh5dU/6nZLPojzkUk
Vc9/jmPdcXQQcZxUxua2L6z0e2mA/uaCTEwq0hrIR7kGuXDDnV3ODaRDeyxYQBZsJ1o8sTfWttwY
zCVAtg9xGwiudYeEVbamJNYMgPcpGQCunB0O6nMXU1zCUlwHs95g8wer5PVUT6mpQ6dYznnyK1Bc
9Uaob/lfSAf/HHxRO/jKb/aDOgpv6K7Q4pquMqXaqR1aow+fisZp8BJvu3icXW3gTFkcGPej4X7O
Jg6iJOkgQIe+d4zcinlpf39PtcEuablTNzibtn0S+PQUfklUC8GHFe1iVP8M42uLGasUX8P2kIhd
EHbr5lutPrs4BwppaLzVunOjwFpwsCL8xRWpoNe4QbLttkKEw6wEWSBgZSdm1DfFrPB3TZK5CroF
KRac7T6Oag2U/6aGUCbQLDn+Ua0IBqtbL6rkiP0mn8BEmUvY8mVo2bWoRHpNChrG3toJSGv+Rzj3
uQkz30OADbJPtB/aIxXXChyZ4I2flKst7SJIbnqD4iyH1zbC4rl7RL8vtOoqqXxpWF9GhJMJ67Vk
FoJBvl9FHAhp6dMUNhr5kDLpMRTp8ikFUYHu4ARPxWpVhvXqFWZ+T8FRbork8O28hkqTl63+8qLA
qHXtFpU8f4rKdc+mtjOXTKRivr2Djgf0aiT1YUscC6FFYorJJXZIaGjbjKb7SG85x9I/fHujFqSR
A2z9Vnpv5klNP+ZnQEwq1H65gnamlf14zol9aUonp2yqHoKe/Fuq9uUNnSFZeS4pvcJo0+GuIyav
4Zwo62krczBJI5pbUF+mj5yQriBosDxfTyCW+1O8QwZhhX0vvtcrtguwy9R9+SJ1K7B0RwT80pMl
EQ6C1hHsaxObg3VACQP+6WJ2a8ya2/myisoPz9rRhZyT41f3gAGicFIjfVO+av98opLXc1SleVn+
KMyMk7cMx9KZaku1/O9km2n9KmB32eZdx0AcZVXpghBmy8KYmDXlhTbAdNc6nEoPRwe7eKPLVeHP
uexzXhkhI/E4En4h9m3/4Dwqg8Z7iLd/j8R+LQ3vfP5Ls7g2S3fojeFRhzma0YM7e9bsI2IIRg9G
W8CAJdP765CYoPb/xlEVDLuqmk/STMQ3oXu4BQP7O697PBZzt46gugZxRCxqMHSw9VPJhRLDXOL2
6Rw8z5qraZNBftx8gcM8XmtbjfGTWW2EeDeleNFAjL3HYUvSKc/qUBdVgapjMM5qPg9JF0zjO65q
LrNUqdQ58mtYnUJEYtmCsGzpqKyTdHVlV+Msp0GbW8SV1OIx4e7Xyldz9AVA0GNtaTc5/hyoKmpM
Y+EZLy3Of19P8UGirKA8NLDtMqhixsUBKOvQu6DfATOc1dLoAnZvHaUZlGw5CFn9IsKsFhU2hDDq
DjJlf+VUksx2/6Uup9QBq9qyVi8i5Ic0Cd2HkAIbw+OD7OxI6uYg/H8tSngI0OL/Enypx0EPKN+8
OetYy5RLiH3Fm7fEgoXW86Ja2gf1LXPEJYPOwEtmUhtoNoBEMU3XZ0gg+UKzwF39vMOLEoyaq/4+
QwPgOb/Voi32Bt38HTvvkNqniiucWn2eORWS9Ylaaamiu0e8Mr5uNLSY4JI63LSgz6Dn4eu/KFss
iL/ScU6Eyzi4whCS1rDPFGei/zBnHwURo0qDshn2gv8nbuTfkF4yNxoIzoAp3UWpES/AJtKw4r0E
muxJ6PBdaieGW1TXBWiqbftmIfkRBC8uqcXqG3APmloSFJnM7ZfLWRgyP9lLchTJ1rDiLsGV7uXs
R2r/9iDn76RapOHLn6pEl7Ir1U6Xd3nRc3cfyDx/0jRzqHmO8JukwPyFEZWZ+mftlT1J+VqPEpB+
sm/NKbYGW94PE2C4E/5S8cPF+6NEDrsOxF1+2vhv/hI4BEgUuGYIJUwY6Hs8xVouOQtZGwoEHY7H
3tpnPie3kUBVgu2r1f8aJhdxW4kqjhbY/t6lib+4NGfyipg8O2KOvdk5L0BYFWe1PEwSpXmhL7NE
WL4V41mTDAU6QkE06/9jS7W51Ssys3mu7r95USoByGGNo839WJ5C9qiVl8qrLzG01ipFCA6mrQZF
1jG/1VzLklVkryQDFGvprD4btMIWZcQW/zgWhAPLak/6PPLvv57LxwLvj6pJvwcCizltz//XwpO/
iaUdKrz89JEdsWR3dIrqIdT2/zgbAHpUk0dQY1ouJzBzcrpZgrpUYpXm9qDUCL/J8Htf6bCoXj5Z
Tki2K2l4PuWwOaRtC+Y+Erv4U74RR2a8PQneTATTO0m8aDxKYc+SsqDsF1yAMnCm1s245m4ua/Yh
k7MGawiQYANJS2u+bo3kHj1sNM49/6y/MfklmEmWj/Kq9aA0HdFrnIC/aQ5487VAETF3D37R5Rn5
rhN4VNRGgb7tj3hiPngJWTGTZPsaN3FA7ogfCBQZGAZeIeY6vOQKS7m4Cvj0ekNDmAUJ3lL7WFnG
6dvjCPLtBLj1LKgRhb8xiWSpO/iCjwjQPeQhWpKKHuzxvqKXG9+wLJgrMxwiA+mFSsZzwcVCwTtQ
ePSbr/sK15Vk92GVyQ3s3DsgZ+2LK7yeQdNBLR1rVJdTR+eFGurZTn+xo/SwSU42tLPBlfG0nsdC
dNPIbVksXhvEvSp3EcFqKV6dC1V8fUYeRC0Ct9Rq2ndc2Xw5UXBx2pb3M2s8a5H7dw6aCSQMFqHx
RwLFFDijplwAMl1GvDzo65OjT2hwkUz15IKZIxi37oZLdN5JzAUJs33MJ41BKmUPjVNBB8mCs0dl
eBV2sb3cEkJPoxB5Ct5wuWrwzAZOHlXjsTzYpjLkOG15pgZSsbUgzAyEm0he+ThzVM/OT8He8Y6v
f/n/0K803vgK/opENUzdh80BlCyv8PaFzc+BAn3Ijerl+vpTuFjghCg02+RCahbUja3AmyAmoUHz
G203kS4Mo76v7JJNPNpqIj2SB741r1iueyC2YgR9LEo/T//jA4TTC6KZfzeAaIXYyOgiND7VzV9C
XKTKjY09GqiLv7LfC/IRaU4Q+NzYdU0EN7qdwSnreMN4TrVqzrX0BS2zDn1w9khYftIYqWA7i8D9
MQ84KSjxXfOe0VaucOT9fSm1PycRJvJGkYfvKbAY8D4Hja/SW0SFsZaoD2oyus6EljPrFRVuLAaX
kvh6Veu4wE6Zpy/cgNG8EC5cTIXRZtvPDbWlD6Rieb7zUcGZQuL203gxq9ITX6HISe97Fw0OW4Ya
SqjsRXi0GzhZ+W/byRjjzDvofEznTR6RqEQZTDKkhAC17DMjO+sfh7qhe8DgM68zO4mCXHCjgXPN
lDj35eV8UPpGrv1AQwzDi2NagRu8lAgnO6IIyPi7OoxbV/BQYg2fXwtVKuLb/CUNoCXzeJclIcN6
1QPNUa4qTlHg25OJXtWjmEzhWve5/Sq6SbZuM3hYBr8XKZ4GIj0WQiyGO1bISGlhxd9AVmeRfP56
dADdMJM4IckWZ5eD8RL/jLxuv1BBo/ItAIHR54jH8WC2LpPXnpOjofP87xHbYAMo3q7aZKQfIWEA
zfBj/2vEo2SzPGe6Q44vPclsSFG9AqYIy5DECFrOIjcYtpyX2cGYRCdCunPjPTpWwPBgA6fvPSWB
zkB9+Bpzwf93WbUaiyLXuGJLKFWbmR3e/gICvy4Q6HY7mASOtyL+8gl37BXeZG4uMKXhKYHVygaJ
ltMsuIVv+VZ/1H6Vx9vVFtdYqglRWn93Z0iXrjvOH/lcY3ypLxy5VqLCJb7mswlJkt6/8lAMRDJS
b7Dbjs5NOqqP811Dmacak7p46uOYquGTELxSpmmpv2g//5MFKMy1ODZ+CjjVHXtXc1kWouvGNtFj
Q4gcEhH7v+2zNffNHiqXahPJVgCz5O+Lyb692YRj7ll5gszbrFmKn9xbR5SexO2W/DlgKT06o+vO
yWHzCDFiGf3ytZNw4org92blvPTLF6TXbfFO+a/jjTz0rZ/ZSnZn8VUPTERIYz+BsFnzSjc0oDil
pQvHd2Ks1pS0gU4SbBXwYZEszls2REpSfNROgdcGoM9aBHWFbOyMcxGx+w1Ny4XCgy1+bIhw948W
kzPc8mS45/5LlpEgmGf04XSVnFVuuyjimEXByScyNA1OItORlkC8dCaCsecEC00CVENtTbQKCd0L
7b1I0hFGQoEstYE1KuZZu7uSGlOJa9CP+fv6JGMjucVVaO2TMwU3XEUPQRezQKXcd1wb9NvdBBe/
GAugGK34/DxO+vkhfCyyO83rPre5gnfySAvjhf+beLfCZ63hLwMTZ4kDPgYkvPr9rQZQYhyjE/3j
OaJWriUWhyik/WA+NYExmnwBz3KXRjVitJlhZ7h9FnJky/k0jAUyYNQa2Qzemx8it1eFf5p8ySYC
10svRz2q5yWiCunapt8pgmAYL18qOcnAwZ8h5LWLM+hN2k45Uj+/dAuIgF48m7DWOJtNL4DFuSxv
9UuO+v7LnZt10xyJYcfrsWXtuABZzWmjrSui63MLZXbVrtddghpNeM0xpV0e60zbmdLrnPauSGjB
h+hmO+hvNXy43UGsO0CqNE3DiCjddM5MNgrE902NPw/X6pF+yLe2aAGmdmsiIQlYcEp/PXarnSbP
MeTTX9hhtXtHRc9qbKtVFm61m1AoBrnNu6L321r/cHPH64TJqsHFa5hXnSr1myQKC1ZVERwCYPLq
bdpzR2jFamCAaLASREzP4dZtJBm+rRl4wCxjwbeftVP2Nt4yLkZg9CYK/StJp7ZV0ftuZXQf6sru
HYrTjqhHY69/q8L7Y1ajA9QLqVNOmmJrKKMyCqCH5fPue2oyhlbQPhjeSy+61fnz3VC2M+3hSo4g
M3Gx8PfyRM+EOjWIuiXXQiJYkisDUMGHCT/PeaFNde3VrxEZ0S5jf+Dl0NNU2PMp3b7gO7awXH/s
B14381FgT+zAZajq/Fn+a+P74d03lu+od4u9jnQg684VP/lfbjawmZN3pN0vl9/h6aPKGXnRs0PJ
vGKgxWaP3TVW5QYJk9Kpoiw790k7htL7HzXSRzo+8cLjS7Twu8N7z28tM9wJxbVW8rAH9N03hoOK
7tyud9yNU8Z8VH5RBQRog/xWnoS2kkbdtXkd8Yuns+vesCS3kJNPuPfCFTV+rErUJVXVWP7g140W
oE2RNxCLJm9jUwi3O3kQCkszE6yz2+PFdr3jCQ3dxe91DTla0M58kxN5I5Th0xNlwyAzDJ3w9BOz
LbiYx1h0MCP0cTsalgdU4MMmfwThnW92gEaochfNSS1sVH2kWxTmhsFTO+ImZnGsfDADpTdTj0Ft
dX2KJN0DQH4v2DOVJVQuiWcUvlW5vDd8H3Z2igBChnHDVJnxRMvVT2rT+jaEWYTITnIIT5Bci80Y
taO9/t8sQtzj/JHegqKt0XpXchEKyoRlP8engxENHfkAkWpw8Bw5iWtajPCR0JnJMoiU/b+LQ0Y+
8in190wSeJiOshYStw+vs88P+W5lhROgP/+qp6fApdwLFVtXIZov7yf66isjPgpEaDji6eFaarn/
7PjnjxSz1ZcmdzsCsx6PnxeOiiPx5iF01rLo98ibR/rlpIiCUA799zH9Wo1mv5A1oJnUUzBJwrSM
P1Vse08bK+rz69fpq3MZDh+Q+RKbAGpjQUyomB/eMuIn6BLwa556ZZA1LIjY3eTFiKks/EPkv9M7
oh91Bp0sa5qixc4iOHUp1Mrp0+rNeCDB9Upedau+2csm1Sl7olNXVR4aj72Ltmob+b8oMyvGQGtC
w/imHhh3AvAp9B10bHSQl+7lPSxVjLB59qxMaOy9cE5RM1C4FqJahUPiNVIF4UiSdpwGaw1WhPKK
NY+/VzKvAmxd6hWTMnNuhaRFEyanuHpbKReqJlMasu02mm5DiNwdD69XeeHU38XYsOQ11Bc4oLtz
LaduUXxFgSclRztGblAM/fBQAktoF0juL0Ps0rlIx87pUXTR2shwUs2Ny2nogykBsTaUXAVQU3MD
2TodRtsCSQDaPuhabt71CIupUZjfJeACjt71oFbjOy9WmQTL0WbxSo+1fASoqEHPT1+uVJgGyf4w
kN3ag5kCht/cOtO1gB/ZWzaW14v1CZpUoEP/x7SS2J/6jYd55i3K7U9xD+D37l6TjaSOeHzXjoow
6ir5pjamOWsaQ4lK/eS0Jji30yhQg38rcJvkqGdWg7omQyp3IQbpSAzWzqwU8VuuZL6ira8l2KTa
xr0yg3nW8cx5VyqVoxVJwdvgMwc7KAc6IcWNifq+ZrSFGkEGpgJdTMJnF7uMLDeGlph1MZct7qs2
Ye0FB76e0Qd2iB1iUgPvCTmURTYpnoVNTaqndlQmm4dyqgHyZXA3RfMN4QiYy5QShJ/TvJIbq2Cu
62k3gqyRagYtg/njpeB5QKrEtt1YzYXYaC4fYB/bb4aT3WmVcUzUUn3cYskxvu9V8XRXna9EQk50
SLlZj6fy/a4wzVkzrD+9sR6W54L9u96UDo7m7ggTN4R8EK7HJ9mvI/G4J7Zk4+Y56loKCUA7OVX0
mODN/GoNjxUTZwECuD//u7FtMJNw5B4IRadtsfFKjvx+t3QV2/f96zt8DNsLG3vYB7dKgoLzjH90
WHr81QC7F0lt9O2SwB14JZpv/9/qxb4uHMyOo4tAXoQLHiXrQ7LIqvrgW88AqxH10X4hjHEFRmd8
p/T5CChwVR4Zu+58bBf7gRHZJGjYAkkusuFVbIgeVFrFlZww8n6Ui8g8AusPTcN3uo7aIdYu32zJ
4hw3HIoKishUVORbiT7VuOpvKddgMgMn9zebVWVt6stPxcG7WTevdCl2I59qenSC7i8FJgCAON2F
lgq2ZzYtIDxAybnxTfgbDFVmynOtgjgER939MeQibVGsA1m6tiSrWAvdaBU+lxztlfENT4DxAV8S
nODYS4aSe6M3tHgfpbhqav4VjxVGBHfTyP5/RLYYvfqppDcDFJK1sfirOZtSTYW1QzjD/fNU6u+U
XG52EEiH5K1R0SX0aduJQBx9XM4UIWJx9Mzy8AXBuw8fuN+ck7v63TEHMRmZ2BaEwwCUg2WUBiwm
E/yiqAvYdWeyETMwpbUmoCOIeWWtSDPxDPwyPOQ9drRsfND5wEpW2g6Y9PJ5wkaoc21XGeqeNgmo
iWt7Y2uyfInkzhwTNznhf3NxEGqeDfsX+yBPQ0KvaYVyGmMzlmHHjEyjG/ecwUnQ0Pk7s86KjaxP
xJ6rTLI1oVbC5qHC+3SxjkGU1KONfnKDXct1B5N+tEYBi29zr4xj3aLKL7OoWH2gnEL39Z9s1mFy
Psf7ZVFOHc0so/pK0JFrJlg0wrbrw5xG56k3XVgN6Mo4O0S2yGyunnnXdEKIZAcB4Rorxaz3R0uF
fwLJuom0E3ziwkPXr0UWL60/5pEgThFwy44z1T2/Gyjt4LZV/K9KUZaQFKdOovNUlhvU1SiJK1KM
6nZEFHH4vwjdBhoeceR67JazRTrxSSUWOh+q8XdeZyL43RPLtcqP2GNzvZGGC0h2eTPTEwdYYBS+
/yLoIV8FXcRBVdJemTmEJzoo2Isge7STJHL3L4sHYDtmhmMwiZX81ybIDUZPyGNJSJ9UXND7TOlF
JazxMKOglrzP1OMEVry17167xVddWI56lwTATeg2TdFD3HP0SuuGtVddHhtHUXQ58UrRLa7gDjMH
R1wfrO+aRZzbKGNO50X/CMTpSe4Y/j65IvBFHSiNemMVUSXfDJu+5+4w3/Gwp2vZk6o15YeVC2Jl
5lCjUaelVtAlNPN6lKBQCu/Dk9J9ryaPSp6mtDN2N1FZ8L3x/JAsvfAIJyvT4CkDTBcbD65rhMnV
ZEP7EpxLGd8HQXpWeWTAB1SRY86j5K0Z7Bgh8ckLr8cdpIJAEvzgqEAxo5C+cN9lviRxxzU9O4JN
v8lzpE+ZR7jAFpv82QO7+CLt5QnRCobqBY2FPu5VayeSUUlOGQPM0VHAYKD+K9jkaPCZA05L5/KN
t7P7Dl+s+KG0NEvUUaG57jYp1rm2SSTm8XnlNCQIBH2/x1vcqDA0CGVaLZi0+gWPgx3gedYSfCdo
boYMU3X/+rO5HAfPOo8N98xN1nutH9JcBoB6k6ncXMW7YYiF7PvG/Fy+3x65R7dTkBvFF6ZQapuN
tssj3eIIljSLU9rtzWgIPcaGCKIGngjSlhq4gb1Dl1IkYAQCD7S+AyCVbtoZufxoTqmJ61Q7Suct
KzU408Db6F38nEe81Adc8DEzqeGTHT98lY2r2VwK2eDfi82rSYvO4vwBhbiyLXgbFyrko4qQWlXD
0KNxAuECuKcC6tlQW+TTXAJ1t6HTWQOm7osdE4SeaC81wtlaB2BWsvVdZnp/2sxtH23L1ZSKKA0J
W7Lvr+DoWTL79b9d4Q/lJ9eryy1bAJa2hkuFKND7lC134SN6fGdxLjn4wgJiT0WqxkAGE9OJ6y1H
jArNTjz01U9sP80lQrJI1lhQkreB68Rt8VxDtANq8YxPzlvdGRYgWQM6A2IcEeNpJ3kfqo490tac
BNs6qcdh75FWItnMULtIqVOgjrvxO9HmZCYWdz3i6Pfm94QwK3C7lW5qIUB5wwgy4QmiSxlYsWMN
/WiZ62SBDvrcSE+t0Cy3pLUrIdzj9LtZcYJcavs7SYkvyXktu3j6YCCalTXaCPJHQgRjBDI/7zi1
7SYk1UB6kUcURGIQqLsfNjR1fiS1gFo/CJAEQate+Vx8/IrDwUepg6Wi7Qs9CbOtrnUptuKV7/FC
jlec15mYcnR9oe1ZXZ2vsAEtBFEcdSaFnfdl4p0DGKFLCQMNkFdsq+VJbib0JRX0cXLQujysWoOg
SkwYSPjQu0zx+fksSb1ngrVcxuiQTaG8Uj3OecymyHUbCrSw2pf9X1w8wRWYw2JGp6W12V8B3mtd
oheaDmX8ndqUIMXm932jQdm1NhKIwf8N8WDZfjjjb7XmTetv7illuPFtEXIHyB8JYKo2+/6LqqPw
H1hps6wfg74NTask4Z2knGemxPLj6IO7g1d461k27lUNmS0DlLtXGw0OEfxtm3S8i34fgblYV6FO
5VuJwmA7dI6mnIpOW5Z8vb98Fa4Mc6GhThW/YaEMzhU4t5/xpY3mCNnym1sU3ISesELCj2NfxCxz
Ek9CVRBE2Z8V+uqrGkjqRdffP8UG+C+mzpu0wIpB0fFmNHxXOmhj1FKhNJeEej6PpZvvwcUYf9G2
GoqY8AQbDEWNlg/HbhZvBEpdJeJEheDchBojnzid3F/vagDOQTMIawAaMdkRQWGL+34mI+I58qNE
sNONFFzM0BGBSvrY9h8TgM92UrqWRTAILauwNCUr4haFGidS2LCkUd3hNRv9fEYcCeOPDry5n2Gi
zuJE+zhgap6BzCoc8cWHZw+FKGzPKK4d6n6oMNpH+SENhGCb+8u6fXJLBunixRz1yn4Fy6wKDtPD
yg4ge9hRh+q9b9jxFHuO9BssRECFT80tN5X8KoKTrDWFB2KlMltU/IVaDMWcXpwgwEDSrrdamBIS
eN/x9WWKpKj1B7MsdkxZuYo9bv9WwIYmT2L6ij0YwcVkkYr2Tmu53hz76uI2mXp9CeibenbuZ3K0
klAW2mromeWekbjkA4HWwMq1Cg6LNg8h0CR7Bh3Be6W+OPPKXCoilstjVhpicF9n92/jkP1kYEjU
xDhhg7B8YGscnmKi34EVGxm6CuQzpnAcOJwttFq2dGWb4Ui82m4z0gaTHh4mn81QdH5YOwtXvH3R
gHPGh98m5Sd+fkAeq6PSGkOd6V+TBL6HPl5H45Ira0aXozLg2h9oph2Mm8OPQZYaim0QpE2eFypZ
21t3Tpxwg5wmysnEirHSY41LhHwbo53c/v8Y819r9XNJq3cDsvdaFTk4srRY5/GucYz7xPShpVlI
BznHoxMrh+5DyJJzPjHMnSoXM6o+PWlywH657AKcgQk1uo9VOh2G1Vm4WLarAJfiqMGsrY3++eFh
KKvNcQrexOiK/saAikTNchyNmvm4B6q/0ZNm+6030lk23GDulioR0ZXqGxbtc3/fkh9v9n8ICdAx
YZn/WcwQSJ0hk99UtqB3nizxIiKt/Vy6qWO3DqE8b5RaBOfBrn0BVrKeX03YL4RrenzndfSJnN3z
DH8Hzt6x6jkzvGcfv72WurjtNRqpFDPGhSw8qyxzySVTuGX7dKTOBExWNE7AHXVoXTOn64P7jbMH
JBZCCuFklTV6wXMsq8AzS7K58aVXdHG/Vzm62tqAnte1a33TZIOanp+xu9wMmPPb463YJidTQctk
vCcN+NP595uRa7nXzPm4jyDvSI/Ig5p53dLS6pL4loODZnBzQSBcq9k0FSzk+Q83oq+QAW2rz0wG
Kf/d0bSQC9yVUqyWTf+2fiRby0QEhb3Q45DH5LHMvXAGJYJl6a6HhfPmEScxGEg78Lnz3R8Cc4bx
INx51MIgPKJXy8bDdFWmO6yRH8uSoDn8LP1wTIv98ff7+Qdub3XPe4uVyyrxB6k+1VFaL6pnl5xm
JFfdZS2s2mBdD1AhkpMfB5pMLnQsLkUuXaYCoiMrjle3uVk7ZziTCX9PbJgIwHzAXQdiBjF85OCF
yPj3LOpGaTMS7NBGdFQ3BA+4cZr7tRKafRihM4CNtCeNAXMoRBwAnxHbLu7RjBVVe3DKRgyvBiLl
w1eAKj1AdxWAOduC4T6i+S2lQCKB8mczXQnYXqZX5+FoJEJ8XyVvl23LSIXKTSoiZK7hsVPmJuc4
TXfkTbHpXA9W/xc8/+ODmDMK2RIoamAQISBl+Q+5Ei8f4K+WMMInWwS+FMWurheKwjkfvwJhIF6J
2ekNHUhyIf+CLG6c2NdgzQ84jtviDqBufwHZEOsO7iT4QluKNZ+2B4wmzlJSRD7mou/0kg0rRrav
Z/IdTDfogz/b8lxmkkRk/BotBECOWkfpZ/fcjrcZl1rWNVHSQ8dHCSLSE9xgvg3BTPJX+WBZsf1i
MnNa+pDHUXSeMbZcMlbh0fGN+FeWARlahtVgudagatiope42lNh5VRbdgPp0RW8hAgbdT0FoFALw
syP0eqBO0MDoUA56e3HUPW5ihgqsUmy/iDQl+oeLvQJjbNwf0svYf0gIOKtgjxGBKgg8uXBpttug
LAcKPw9XvSpTFqqkJb09eoEKtr+NZxV0tY1G2aK1KQuk+92xUBqwkpAvu7qthJKWNK/i6+mxCCY4
1IwSxydNe47W2RpqBf0fWq4Sy8jhwlE4XKGSvIq3zXpWZThhvz2cBt+Ik455k8FpK8dEgmjmR/gm
zzv/iFFYLbzS47sg5TzLFva4zv3tTDm9KM8SL+wUlyVK53FHlUxLpgPlr2y+e3B0l5EQ3xPSW7Ob
h055IJ+CPbDojs+teJ0RW3c+h2yeSUQMFznbzTUY26j7S6ddv5KsazHvL/Sjj8tYcjVolcoOo/pR
kR2i26LQ3/mqIMuZtvKNAgo/dQEDo2kgqxvMj9zVzkZDBrxKqmoEZ1qhdih07X8CwYZMV+XzbwV/
9zoyBMWQDHXQ5w7mGHqNWZMm0yqKSC327KaIYOgEZeh1pVxEYaXSc6OIE5X1wv+zJ1xxvtUz4DKd
pXSG5TsU7kg1nfarJT3etlpC5ssODBxB3rASXK3UAmoHRRU6Blmva/EJNijxwvoNyMSdkKBNYD6N
i4HPK/AFuc7e0dJLPcUXa2iXnmsY9BvAsyO3Rlpo6uBj4M+ThrU2flzgZiY0qR3KGjloBsaf2h1r
fTS72QgfFqdCylEtwusC+iv8PMygBZFmVYg7zfnOcJSL4hfBH5WcYlGJa3r/SY7EABj05nMNPCKY
Y24+3LfdALuJ4l7ARP//31oqqt1C1k1FqXKpoAD5xWtxU22i1dzB5kwgL0lgxPBVNqMAG5EC+Pgo
UP6D5h8TRZ93dfT+zPJnkYDCV8/hX2uleKyBXAiJwu60NemiVTM8dTuIPVO18qx8aYiXYENOnD+j
w2OHsRTR+nGIJ6cly4xVGHj92B3yso9cJIRCXrOSLNJ+k3Vl2H51TaSPD3KIBKq8+wFwEiOnAWiD
tFq423Ie3iMyvEW1OPubEUFqJ22HiMJ60HB4YD1CIqvwJfqfHFWo5Sv8Lu1uz/J9J2N2DFq1elnr
hYoQi7TciaUvol9Wpha/RV0bEDKlDidE/VmOtCCP+PJvkl/K1DQfDrbAKXVvWE14uZRWqy7+wKF4
gsNnh80Ggmiob+mTCXMTv1P4faCs/wQC4pNpzO8qQJgc9+2UY6sNsdolMg51pAKp1ISukwvUrkCc
wkgXhhyikkMuzTuMsW4Am92va4qdi3EzO4Tb391s2ciMWzPRdUuzJokYADqUDrTY1hvZiMVFoREb
JsflsW+JcFuKnPROzZoSsrjBBjj4ghZHkoKME7v4TVdy6K8yuQILxx+UtY2di9iePicA4Y9oOg4S
PFfvZSRYKHhaio7z7n0QpblnPiDxkjG9o9r4XJLs8VfxFF9euJRy/g28A9lv1WIvLmbIryXzM5aI
cFi8GVzon2NY7HFJ/6s6H+LhOU/e6kIzSn3CNAX9Y7SOLexuXujeEDVS9PcWJm9Gkq6QlsoQ5Scg
zU642sdfBPvhokrbnFIbFiQSEX1av4ApXo+Yl2is53mtDC+tNytjChrQooHTBeRbhibjyrVZeUdf
7LlAbfdd7NpcFoU9H16ILsMvsFHqF++CVODIwlTk2c/rUH8H5coKvByeiXBUugDc97WZILTmBEFB
L3MZD68VjCD2ZH4LV+vu9wuwmz5LtVpZORDeJiIwT/nr2H1h6mH5KenqkYCUNzujJTnLkjJu/e0g
qzKS8mLmvaRMxyln8f7rhxOSJSatHAPSSy6wt1rJnb5gcibUydc9u2hQWtVoxFYfsq1TOoudI3pA
1fsmurknzmrBMXXjMFcnVAp2WxoqV9lLmH/i78WAs64XLgyuluLkFGO+zB7oyJLv6Kvtr0lQrj0F
S2K7A44fXZlMTIhr4I/2Opbph4nwK1GxW6jvfGbwj6+c4HOFYj5rhy3gzcf9Mj3CblKwTTvfUlT5
hGJjhWy4OJU2Xb+s8ZO+YHr2BVYbRxe9yWU7OwVKEYHEFjjsDpfRY8R+e22hLhRpDR85DCuO5nLK
tzedtxTEA1R/i/2wyXxxwh3L39kPHtBZtFimmaT+032PjXgg5R07/hW01vSKPM36qxOyvbN+3TTT
VAt8PCGRomsIKtZdRg9mrk3aWKBMMs1MkUAhHueOOTJ0cXgwokFaNF/fKMVb+QHoT6ROE/gYWycL
dEdfTr6zUdy5q6T5AHy3Kww9ir90nUVXvpaFu5/6F6llBKfLVLr99F4GsXt9P7S09zYWCcKKRZtp
uTgbFchuNOb8hKBjl/P+ZS8cvyxlhgGNoqHwg63/aZtHqpJXuMchJOLNmp0YIcvSnBZ9ZjopS+QI
QDCibD3GF5++dVKCcpk+M0u1ftJk9ZcHfYGDJabGkD271hxan6gC6oPRpL6emhbF5OhN7e+hW2E9
Pk6yja8K52lTrstJYaDHp2TTkwxnoWykZPabIaY8XmGBJGxCyq9i7DA1O/JjqlVG+B/Sg5YqEn33
xGbAV3i4PARm5RSo3Wd3YNUS7Td0IrEIw+pzNLnNtOaY3mGjwypTvXfn2HvnqVvrkFCEpWYI95uC
OUHpb9FlyaZxrdm4KX4m07uw4O+xqdFrPr04JpWcrx++LsZjIrxtJUPtQQPVeUpKr8IcbwuTGR46
UnJK4EzhYKuajnHvBoNdJ+rrRF9DihG8m+2CHDw1KH5aopQHFK+HgvBIdGJkJOPlN42RL30kp0S2
y77Gi7NgtLKFGG16j+fJcZf/uDdnJtoOPRxDRdK+k3NcDOzyn/SGhDqBPgQ6DNkrbl8mmO6+n1WP
ZPAve5qvLd/AW3YSUETrnNzse1cd3fjGra/N/AIHki8kSKVWsv+V91pXeDZNinsPYEp+1dRP2sB7
iVrBU+Np82NQ74n+wFBelveoLyQlRczEeIJlrkKiSLK4z631DfelzixF1j+NkEM29BldRiiP8aqw
vzLSNpY0W4VJcM9nTuq9/xoEIDrpKvOiO3A7sGMj/djxUnItcv8aDktj42kCET3U47xJMMN7E1gN
ptIy2xGLuKC0iu3ndCu+v4rbLch+JxBrQEQ3qys91AFIhXet6GBeVvR197KlLrYFvTvKW5YgZ1ID
qXstG8t0IYS0ox+zRnPiSyVFAmOvXRNMuC6b9GAeiJiZkSe+KL7XXVk9dAwl6gy/E4LZJkv7vzZp
e4uWosIWf7VGiJagraLalnt9ljtxvu2Hkkf3PjdNn8tbBchcn59ESMAn1aIVMBp7P3wq9zv/7OgN
PNM8Sn9TIv5tH+lYbbHZBrHQFLnjpblcFBuwWEIN5BIi68Nr05sZMskKZdWtKuu8S1kJDGIISMUs
exXULbmcRt7XDrqWgAAhjTSWvONo3GNjYwCz/VoXhufn1Ypdtn4HfnoURd+t7D0VYR7Xj7pXzcVM
rJI4q+NExgX9zDRdVLpZjBAsT06jNmopLhMHjASzgwjjo7GpytaVfisXhNb5+i34QLSj9l4xBNKW
0h2H+uAWPA1KdkeVFt/eSw6jCk5/dMp50mhObr44GzBB/rHdu7ezvbPfOJs2IGXNVofdG8KsYfIW
zVPcFDDYvwakot5rArsgsEqzTPwuyJFeYEBxy3LLCleATAxWpQv1bzWzrzqNqKY8Qs7Q7OG+FFnq
B244rSTIm99q1Nt/N4rO4+z/nwlpx64KGAIKgW7bDQYM31pA3iuvdMNVLRmKzVekYCWVOHAYMyAi
BNWdCQJ0W2a3SwYeN0ORaTXUhBpr8I98mVwzFodOoJRPRIBvWbg+QJb2BQ+uSZm7g13hf/YInf/L
tfxKWtOQDfAVC0aWP2IThvzJvhw+r6AlYzVoQ9Nl1HLncktOiC7bSMp/8XbFTEu6/51X4mfsnUtk
Mqtq6djw1eG0SwdidBh4J9/6tjVolYABvZVt0cg9xUzX72PLsCddhbYI7l5RwlO2miR+gIFUuNeO
/UVadVKweTdbCOdt8tgGsqeedJWYa8TuYFPTMfSC3sWB1Uv+ce96YqR+Ws2gPVjfZ2OLiml+f8hg
N73aKzH00q9kaP0ciduqrvo6xcQdQPGIDya6ssnOQXGcPxc8UShb5rPSWQvxsSOrFuwISr2IxZzk
TnC9wO/WZO0F676n+0yx2axmnEgFqfVG13x9qUkjpTcbNYJqMHCZ+OARbWyVZZkY71kOT4RYibj6
sDoO7cEywWy0a55m/WygZ0O/QGNugRKv0/ny0rR6fFt4lF5MW/wtYPVUwzZ9nztBdjqKl594QCb8
Zw3EfMJXTcs8sLwxvpCZ3H8/byn0cmqhmpEBQSjVNNjlPZ7r6cjiBFjhIK29151RO+yYbceCeZGC
nihUFpZ9laiOf+k5RCJCznLTpdc6632bcMQaWSI4uGK7GjB6FhxCnHdKTZxW3hLyCxgSiGqh0BGJ
2qXjkAW/W/i7OTGNAgxAFpORmlFWwU2DOViEmfB00f0LfAQSWiCV34zNkbBMjWgJ4Jf2cg72HjXY
RVH0uLIIbJVsazy0wDhlqMeXGYDqyW4ibGzRcUhsCX26OGYUOANF/YD1TBH2bbebdzQc11lEXwJA
xN8wpOl/ONLdHwxdAq5VZ5CPr4euy9IH3XUpwVOzSxcO5Trxu8qfCQG4p4CrqqKi5HcoFcRr5Usv
LRgYr5XDsTt4y43PbCm3ZwTRPavIUSX1u59s8PHrX/f+jKQFYWdKyKxkwgndQHEQUamyXbrA3VYc
FOzfp+oa8Ta15z18I1cEOUcsbDiK2BGEnCFx1CR7v2vURK4olRtOGY3R+cvWWftut9kqKpo9MUkh
D4bUnHN7wWR3YENYvYUuHfasrYjhCpQhY5NByMJsgGdDbhLcnQ+hPHB+YHgSZDOqJTBB6xlvtTUc
0oW84ZVyb7woTQFG/CiCzfCCR9wdb0B8Qr0/Bk91o8WYRP2yNrHWipNUZm6xt4NpUa9ZIHhzyX/r
oMh/zt2DAcgXW1mvFX9CjNleJk8ee3kTHtwqhElBfmoVPXzbrUQzoA8Ig2yIW8EeWxMcOFLVDXcC
0ulwpapD8mlCaj6jNylyr1S8IbuzpChbQWnxlBOjEybjus2Ho8iNjhLcLys84/wQcSsU1QjByQjs
rN/Ec9nangaR6qvgdKj23KRyt32UE7XKKYzXsa31V0iybiWyV6dVijTzacTWbFACNDSQCY1w/YIO
l2pnf3hztCyvU9fLw8Q/1tM7hc3Nu+lJe1MjD8oLL+xvqlhNpOKvzhjkyIiLcz8vMwmVdtfYC9p1
k464DLxZdiXTwmpjgdiwqP0p8Vt3gaTQF8TfTQLY9pUy2N4gfKX4qzPMuwaar8UMmn2OctdbKb2i
8ftnal8OKEVhfCU+ZvWDb8xUNnsnxtskaGgQ7UI6kMrO+wDiXTFcR9RLn26qOwT7lTHOZNSvc7dO
YjADAeK9AQQ4GBBi7W1bZaxMu8HPxXqWARXILn5EnF+tmw0DGvAPZFIzPkSr7bjJEhV64e61J2aE
w2mMETDWSIdq2lJ+yi84KtfUWtIK7AmR/O+mjOrFFV8iOy1keZNbg/M4x1EYIGzPSzxCPLEyOjqL
xj8EY+sQxqd9g3PIMlJ/nlqBwpLYS/Mou3luTGfnVYyNFqYOZjnMZ81HUQgTBAczXyJk9qs7/CFI
fYzdwhE96RlKVVsBoWsAsF8Msi2APkTbQ2tnQiyKg3Uj/aYlME0p5yLTiFJX+O1xec7iANDUokE8
cBYuDMts+9Nd1YmxsfD9Vb2166ItKOeL2uGu+fjuWUnnaQD42y2+gUnivaH/KRAVuKgEVWdVEKw1
YSF63shTN/XoRiQfH/YwhsQ41ijFeL9CbBr+TbN8iKb/VhrUk7KdeOsjz3bn5dYrnWkAzabK/Yc4
JGEm7NbDvrFL7964ik9stf23so8GwdBcG4SsDpLhp3uUh4sJXqZbtmvLHIOWTOZGS76DN/Y15/ok
ueDY6yG5MUEGwe+XjEZkCI+IONymlnBYlmeJnCmoPU/iQv0W05fXru+YJ4VqmdZ7Iiy0FZdrltY/
6DwTXK3NOdedVuY9nz21/kJ95dp70cxpPSv1/dSVfY74r9iouCuXbRjMOflNj02/RpOth7c/0ru/
HPyigzPw3lsk602i/rJe43Ve+SMgFPwAx2aLP9qKKuIoQn/lObyGyxEQ3kVYQs9HDIw0chubOVtz
948lYjScSsWx+AFMOjhFVF3/XReOsJSSxNVTdAHqXM3Ex88Kz3Y33MvNAjcN9bk1/rtJwGmzua/V
60yrD6Q8ktasrR5AsrUZ/51QfWm/eKfvADzMo4h+7FXBvEDDhGfY7aSBY4aNPbF9B9bC55YvdEQe
ulc4G0a0NoQz/RSVuSKqDo9Orf1pAhUKfa1sPK7CP8feAUPc0zWcCAcRFyTCrmJnOrjSaAFr/Ny6
E7M6OoenvxegSBFOQtrohMSHumKUd4+tBaHKT/nrPnFjZhLWVAPuVmOGKX0Wg/ujrK4h06trxHxW
F5JTvvd6vdGn095SZHUpi/IF2DwUoPapPrnxaf1HAKpuQxTqhCgEyZa7UOn91NIMawxvLCRf9rwC
991n1WSZZFVj2kbNvmgpArP+ZpSd1jfzMe9Vi5SMzayCEimtrq3+7r1mvpwE3fSZtcC1wGHE/0m4
5LSfFYBwLLdJ/pJuAR0Bxxrn9qHddZat+USeHLMgLktVLsfSV5f5HYklwp1KTFwbClCy4J4df7NY
4heK1iDQH85do7EPNl/B5Ga2wr3a87MbcB6DE0D4FTJ3Q6IhCXXv/kvWlkA5qcEaWbKVqkPoQcAI
YbFGG9ZOhXtoHF9viSK+gDueY8PfTqlQwgWCe4/Hrmkprm2Mkgj/k513i8RbYsUXd9dN2mRVt5+m
zRsWDVIBA0WypgojwPhbqNpjKm7fA3kahuUJKUUstEyk+h2VfA6W/1qoO1/ODNmi4tV51pjXShMY
oMAJivQQxCqY/kXABBYLMomZ+6wZf/eBu5DXdbg9KnFiwR3btoSLo+nyVSmIbr4SRFcv5HzDQL+l
c8ImcZfb/iW2uBY4maa51x1bzlgWXFnZE9gg9SboSZXt/M0Xm+n2yVAVxYEElhssUzeFCYoiTlY7
3FY4UcBg8V5yDA6YpHtxlWrQJ2E/FWrPLL1Y7RP6SaJzDWSKpPV/ihmuAD8oGj1g0Ue9opeQQAP/
Etqdt61n9RvyMmrBsnhbKEtP6SNm+Kt/49+faCaJwutntj5pNmS6E4fcx8+4hOO++EyWjj3UPy64
lhRW3IZG4auLA2QDiLzrz9iXSWvnkhG5/6cH3yYMdxCjPX2iZ/vqR9egSjA76dr625U/2JLxguqN
ZJO+cmYimgtjT9Vm4/rTL9RpU4blgd9L9LQ65R43xebpvw0r2zxX+LiOq9yhBrZ5JTSFV/iGFPyK
Xf9xB+59KjJACVIiIQCVkMRIbV2pgD5b4kATavRExAFTaOHDbADJxuqejYY1fpibXWR0LLhlcebj
+JGoURzr5LgPaPxrpBxTFZs+O8yYtglcKKpCI4M+nhStuS6Ahw/ncwAz/CkqU5vueniHSyO/Hjet
n80u750UCmlgzlSpxopWKRexdXX87wtjZYL6RSsMSt9EZG2S8Lo9KIzivooygDEqMy70GR9wBpfU
WHnDJ9DlYbI8g6x1bRDWFgQHvAPiPNMW048jC/GPb3ALit3HC18BsYtL9ynMISxO24nCMdktptzj
M6yhjoQGXd1P9gyY1N6UnzJ9r3OYeHlcD4Bf7L1EEwjGwlNixr0fGKnTIaUpmYhM6s0Dw5vImNe4
8Vjafhmdq5cdEDmcFE3Mr68n0Oe5n9OTtGdZSD1jYLLijK5gLi1JFxGfO9kcJKX3L+Oyz1l35SAW
FltjpGvtX6GjerH49LA/pn5jlOhvU/Z0pCF9uIpEvkJ3GaVK3y7eBhlSwytYAaeZ2qt3cTsVl0VI
52sJ+ssLvMXxnOGK1W8dLpR8s6Ssyk768XmZ5h+bowHPqMv8zImt/wnJGpeuxLD3UM5xLfQk7Xi8
3zcN1ZHhK9j05pywahfguxvXfOfyMw1QGObSI8HZAlfgx+kSIgFZOYC1ELJQmeqdX7iaJXRm+m3i
dkKw1REbT8KeXDvSH6U6fmIwaf+Sk+BJuPmPbKMXOx7iGTVzG8DRkKHNgOx1VQdfiTSUNzJ9Salu
m3HPawf9Z/M/tSWeLdYTijoT/PIDCzmgQonIfexMPpCmHD2SzmzAYPIwaHa7D4YqhjXCdM/V9ggd
vBlsTBR25S8T1LmUrvfvbgmePzn4FCaIEqhZK3e+Un+a8Gt/mvXjzvPcVAtiHKss0e6l/W3Cj9se
cvGAqkok0Q5s4fkBYI1ZqS4wNU1pDl5eK7TP4DSVMV6WnMoIgmkWbnUzYGw721QWsrdj1S0TmRAp
H9XDecb8KTHoE3C400/aeAiDTPSYjqgnJNhySU/sQJgN59BaYOPFA919/VQ3OtR1nI9TSXGJf3C2
DncpCa0ch5ENDIy7QLfB6ImB83ANwux3Id6zn2iznJ+/JO5jkF3+KGTMwj4V3lBiuGzW/U9HGSTY
W1uEkXaY5qXDzXuLEiJQtMKfY+2xEWI/0B6pQ2rdZ457wy9L09qFRYKnsHUOdErV1CwZZYTZoorP
NXYcBD+9kpNRfkms88/ayj4FO3m+kCzVTvjQYTB2xD+rbO64t6igge6axTq4ZDYdXRwq3gz40xUp
/n/xCAu0TqZgAuCvggBnnRumfIUwgQfgsYrzDmNxxeXd33rLm40p3HQDkywsVKT3e5qIS1ziQ99r
a9Lf7vJZMbZCgUbUUBToNJiodRAfuffrJmqxC8tA1CgLzBxbrk7ATPs3JQ5YiYANalp6BmB+i1uK
njXYy4N7yLWZCGW550yd6E/+AD6lcZ0QJDoY4K1xXgaX3+6hyQNr83TPw2/VAjUnusywc2e/WiZ2
0zVfUpI9U9vYy3wHYtOhZDcc7J4Kpj6ZSC8hHWOrfBI0CQEC9B4y4peChK/Bhz9/St5TjCWdiPjY
vWrKFKhFrcsa8mnD+Tgodzsa9EHSMKcurvosCBkQsKfAA0wtbpBz3k+A4pzD7J6Cv6o5ECoOazTI
n10CiFyJNypZ7s8MPSjpZl2pwIgFE6FPakE9V5LCO56xfIDHsUBnsuW+Q4YeJkKT+bLqeG6EMjBB
1EfBvc6K87PqFeCCtN/bmT4XYfsmfHiwJol9g4xfhnMNSyK7CCXcRbJmZ6i0zm3FnStWb+870QZf
PTtgRlKEi/V8qa6ZkJLOK66oXLcxys52BCJO7Pz35B4280+f7LF/1tibvidHE2hANjP7L6guMDds
OK9vvE/R6Uluju2Qn6JSa2pVaJ89RYCSD+gMJ2/a0dHHe4mvkxy2HrK/IDsrZuRoWQ+CGMs5AxqR
9JKHVtU1rKPwI2YLRuY8CedxWEZ7kGPvDg/WS1n07NJ4mIP8yRGZhGDOTmmNrgKpXb7Jq7T57O9E
kZQOfOFyYf08FyrrWvQGbBXKRXYHSioHjH8rzXSWfLBU8epOPhxZBrs8WGKD5yDBX18W47ihxHjw
2/Hsyduw/FAPRIbIvXdCZb1d7ngJBEpdw1CjaAFzVLzc3avyeikRUj76z0Pon8sYNYJbHqLEy+//
MNDnbahBCPaxLlKNU2B4FNd2lnu71/8R8v9qDZ1fczvacRRq7E+kNj0e2/hXJ9TEUkGxSGQIi3Sx
23LIFJQAbeZRNJ/1GC/edbI+Lihsw6DjaLW8ASnrkn53tTZVmCgtzGmO0IQ7Nyd3zaaQ+/vPeQp3
5bwcc0PoYdOHZQhwSz7GSB8Yslcc+2cuH9OYYMv/iwlQXVoTd8XIjArPwWjRhBm1mGEHbKRVt+BL
fmGwibtuI2Clsap0aY0b1eNikJIPcWQNeKz9yBXIf7iMe77peiY9VwHzsmk00/d1LdXE4rwDOrzB
7AX0nUZObx2bK9SaQc6udLjzKAcmr09rn97igxM6U5+kKOoBiwEkWFVQQRxNXkkzulHyCl23qfwo
96ZBoJ50AOF8jZAx/vmYUXMb3uLL8317sqErwlYiWLkkW2lyRuLTNsoH8ohGMsE57nO96jFVxblR
Fw8RG6AJ/wPFLYYY8W+gh9Gt6R/OKvC+AgDlsDwbjOY7usN/dSHP4nuoZ7gs1tcSONj/Pe7Shvdz
igfrVacbBIpkkhPkX4MDDnPTf9MXQuZxqT69xXvNvr2/G/jyd2nfUI1auJ7/ix2y3eW7ypZVM8iG
R8KXQIlgVKTO1HYxzB/966LVCRP5H9BLf0Ngw7z4OzrpMLAf/untFL4rwyJNG6uvXNTLXHuvhHEK
vB5/djdsj17sYdd23J+d8X7nF1jSZyb0K7UGa6u/FwfWAbme551jNK1BC8M1GfUZw57ujUqW6M55
gCYobmU6phH/cS+TiKgBJA3wT9IKctTlsy6FC179eJBXrH0tBekCKfeUExG01CxYPOpVaGKuZ+ka
q5CzuND5rw5gDDe87ZAytEwVtONN5c2BOYEdPiv+XDQK0C5jQGC9qbugI+D3oCr/M//XJKgvxwJH
Ho7+vpbraobqjSAyhY5FFLOd5SLujn7HjIT+PP1StQ3UCG6GoJmLVrlqaGM/MOtAcodUNtVCIPZt
om1IiW/hq3FkG45kxEzTbK9jKVOt1m4T8TJzJ/nc31m3wMVcBzsRELtVskjBXrcp3URW+TgbSvS5
L1K76WLgGDQke1k36AsiGHnaRICv1do+76NooY6myoWpSt/1V3Ga7NzKEgwQj3uNsmkoUNpDQ+Ux
MNQIMDzhiT7sPI/c7l9BhWxe4L0QQLg7vize0hCMkYlTX73oH+2+8a6tSeP/qfPwd0wMiZ/ufeen
2HqsNntBKb2PDqdDeiEXZkjlgc8MeyKxakJg5ePgjpuqC8aViF+q3Uy+I3bj77oF7mVuUUXAcYil
v+FUoyRPArej6No6hgdUqRa6CoV73gRACfJcZmAbASWlp3zHRgjUHKxDcQNigYWNQ0jBO3ldKKsg
7P7OnEM2Mt9oPLRHpYMk+I8q7I+Qur7l8yOtjkAtBEzuQp9yzimwRnAWCbxbBJmfAG44My29w/V+
7RewfV0r2rYaKqC44xJa+HO7Avg4ygNt8NQkZkEizcEpEGaGDxyZNnxnSW/1PnNza+bpU0mZI+KG
MiKdmTIxFsPuI+cwZ4+mmYpX8bIMIleMLUs4RjmJlu8htANm6LZXaLUZWxB0EFl7zJmt4ksBSCPe
hgSJrZiRODI02NSSHHjt2fuD72DsFKuvFDTNU22REwiW4/uvqO1+IZKk7pp9n7UOsxtkFZ6lv3v5
LYiy7GdbMgG/jfr0OcyrwBFTtwvP4IVs3ptE0g3Tm/uVMN72RLZRfjaloeVEHkmF60cM32WiC+eY
iqiisvgjp3u8m5+Is5uAgiarcGs7iKJ8bkYg8ORE9Qtvt5tcsS6f5T5JGXBp1jp341Q83Z+a7nWz
/G7t3fV7Q+Lh3YTJWqo2cXpSy1hJY4dQlGivgYqHJelPOX6uqVked50LM/NNtbQXv0UgXkyALUq2
UzzrQPu6N/TTvdQk48l5ZghSBdU0ffft2ONsVAEFwwmjoNhoV9AUClhkd9F2IvOX1NPVJWgiGpwk
6Dwk8X3Bg0E7wOif5Bl4pR4tgdeuhXKyWRk7wAlXfQOb8nhK9F6Bm+I7E5LoSvqJn/4H47fb3Pv+
GXrVdPfKvosJFHMNkt6MT1t9RV7FK5T2WtJH1guTBD9WFyXWjgd9JAQ3g8xuTb/daOkFkIf+T8Vw
hP5KteC8A9g6uXug5cpggOVzVSlY6D6epv6fOJsAU3m4SD9VSfgiXbWuX6em/2qPEd7+wq84RzAw
EUH3jBNtTQZcFueG4jPZuAxf93QsgbhNsBNM7f0OF8zNq4+UdSh1zICFsVw3zK8cRYuV6zJ5IUUm
iwzQLmVlMBxbsEy8YigjaoXLe8Vkpa5qW6djVR3nCc00FABYSDwbL6YXCivPKf3m9PxRNpkFQbDV
IFuLsTxdfVblEvY9XSUPxGxWtvYEyXqSAdisxG07GlQ9kAPbG+NZfF4sdxtSG1vr+xwrfyro/8R7
L0lEeEPhrKI9lHmrU/HEHtpeHUTL6+qquHkRgPjCFEcshXfaCalYoBt6bP/nHOHHhvLt5ZQp5nGL
55EMsvHDiMUCufqrSqQTeUa/pC3eWqAq6w5YvhKYalEG0AXTsJLmPuQ+LZznQUXwXOa2NeX/W+KP
zr9Bv0RaqQgOCfJ5pe013RduZLEr5Vu9kdMJB1XXxfI22+yE+SfPQcWvE1PZ4trhw0FvxC1ZH2ja
BOFB7Tjjaq7YLSeCo9IWKiXHI89XcEwT/aeyLw/ZQ8OZsr8IZrePozA7R1bHHFbRLuFRP1cr6kfG
xq1GuJl+1dQk8wYQsBRz5KxFw0ZuieSgduVYplXiMmPcJtAGeqVI//1zzy2aGTYzolKuZwxFkIjp
W5Wif1oJaya42JdK1INEgCb0KG+PBv6ff1RnsTs+62Qm36Rml0/BcXhUYQIyuLx/lnR+NgTeuPRc
jJWSzbXcJSnlzCveDA3rNd0/hfS/15wKgsVUUkcS31rnrTOsAx2+rCepFwFGfAuYcuW+M4QsPfHF
ZBzEffeYDcFnyDOj8x6JAZ41Mmj/NsBNcuHs8md3IDuPmOv1jhhU4G3zy2VxAuKtX56DvW+xeAN4
fsgNM76+8FPgDVbbE+G21vjrBTAmwGPOvUCLcN8UdmKFuIlIpsANRwRIbJvMUhXZNXFf2Pfsdg0U
sffzAya9/YoJr9LXIw2hbxJVFNWeDySAUqDrMNWHKciJwL253WFOxM9PPGY6tTZe2Gl+x20g3eNZ
ehDYScmwHhb6egLLDdUStcXhhzYzsIFs6zhvBDcsCBw/vroT0qkQ2+3eREK+5XHRduSfZoTpXxie
JqLvtPLXdJE8ljAyhNyVUAYBZ3vx0eypYBoGEHJnoXUrLtLaZe64vNlYjNfenOrD4zARpbwd0Zgw
maajDvzmFzGBI9GNnsBaZS0Fvl0s+5b9BKxmhG3eWleL6XUd4RAHuZ9ElOioi+QV2PWXrJuU9bTO
Cx0UhJH+6ipdraTb0bWq66pEBNPUoJQs4szXtu9L3a8URdegx1D3GZxpB6IT6IuR3g6ruiYpgs7X
9QYwfpdDoemeHzXuVISweLbNYs0TUl5dmre9sp+C8Z8nj0fp7nbNqcCeivHypLBTe/KhBRJpLRrO
Fjs989YVbFmMEaABmgV2UixTyaNvsz+eQb8aGIRNTUV8XXPlONgOqK6X8q6p2wnkpwx6KkoYg8UV
bMW6fjYF697e2I9KjoHqEeeYP24dLah0gg/31nkk0hdB07ebRWf1ZfVlUay7GAtk4+Jk48nRJHW7
vEWmCqM39oYmgCZrX2S5nTHJNaDN6XZxwtX/SDwaiXkUNb1I/9QgS/5eGrld8eo+tGOIeikfn+59
ik6Oa0081KnGS6v8ogR8rkUgVaf8vAtsu0siNN3vUvAkxFeArjf5C9+M3OEu3QLbGlkiKB2uRNWI
VZVSRMfgLz5ZeHGFWQzh/WExRInLHz1P52HD5sf4b3YYO65l4Fy/pGmV/iRoaXQRwn6Y+CtNfKRf
FoYJ9h2kgcjmJBvzIZ2FOZG50pSkqYCz93d2fwAxUWnwgGV1B8fCTkyQkmYtewTuy/0ql8ZC7J+4
3lgZLeLEHZNCafqxHvc2OyUJS7oCd/2uP4z1wjsqxNrjzRfJxhHEIIUD7YqC2ZsIYIrCAIlxpPIW
+vpKbgXeV5fk+jLeDmXYTa4mwDAhRQnNJf467rn6LQiOE9tTf/CxhpA3U2F/CtLta/NY3UHNrk1v
PmXNz1nN8Ah99LqawgLHrDAHwkv/YH0VF9hVEGtvXfb8wg5mocdP1dFxZgKiS92i5mk9K9ac94K2
f6l7Vxjqs4IwX2tFs0ZyiYUmCqTIxrog2M2xACEKX4jAtlZOLpdsuqpSi36Iz/1Hd+oJWgryR6fS
76JvsOCt4bDasX/bybY6MRATeIQ+hPGeV4KEa5swdfo6OAY+Vvaqr/lhhfRlGSJOxV5A/0C3e9v2
XVHXTzsvp/n77RkPoe39ZQR4L4+TKRnoIE9ykrUVZWDmnASOuWIV/FwXgUBONJdv/Hc6Z00BOzTQ
/EXToHGhAQh+7aG91agffLZyU7K1PGRPXInpZcSKzVippHA8jDriVsz1PDCbbLuxDBuop3jKoXqd
yLYcZXcSobzoWW4IO04sm0P7uBEYfYDqBTEOh5UCDVk7rszQcb39Kl25IQi6fxgFY2SMnEzSlGD8
R57oqbwDtdzetLVO/pxTlDuEsJ3/dhIroAxRy7Mi9jMnZERVJr3xrcSd/HSfcqDNih9WC/LgeL/N
ZUUgeMpUnYtkCouVrjX33xvfdwTcPqQpLsIkolhS8pSGYXncg7BV87XJjkULf1LJiiAId3+Ze2gi
e1Ka0XYet2LMQojjRJ8KKRKFgDKMyfwyswOF9zwxry6ovFlXJLBm2QZpXar+9URf+543+znwYTkt
a+fB5A0bJ6qKq52M3Xy2iwTbZnhyy8cgJLJCLHz+lJtxmdD/pkyioxpTvE40xlWsMSUN37/LXJlp
JzHzdokQwmjMRRP5dXx0d1S5ANc1zMt4rlH7hnh8rHqXgrLnCUlFj4g8IbO80Fq9eVt33eBhSQIF
k+cmAaUYRPYQUy5Psg+lfDRVcDp27vAt8ROuXo0l0fmRcnfRp/idJ9XSkiuhsK78sEvTzNRKuzPR
aJOxROuRH27CANH4HAevWTnFdvdRJGuEGjYDyuAC3mLJvLYjGChTqVZoj9oj1U2OWdozFcef+0NC
mL5xctaeSRthvb+ex8LCEux60aNwa/kPq4edQVKTftB6U88cnqKx5+TThv2b0is1mvYRfjjHYdqp
JnJk1QBnZcmRVxOXE27TZQ76icqkCC/n4/NVxP8oCATYTUmjOpw19k59w5dfMYTO7n8vMnZEdwhm
vSlr3ZHKOQAQZId+Nc5Set7rRwCxGcDwyAXqMkUz3noW8oQFEb581qHS873A+7cf4gHpnjsfJ8QO
CJ2KbDOzOtiJUIYz4iMK8LZlupFqUkCdUQaV7KL4P+iJdigBdIgCAYKkn45/GVqtg1enI+bzc499
VCIAOh0+4+O78O48gEcNAKLj/MeACW9qDJG04g/IbAMdwfwxNBcb8508pzqzqfODchr/IT/2ZQWT
wDLQ+tNhk9+7pJmieMROgda1rr5VXYZ/k7e5iw9Hoe+prPQZeFlbEMFCzU5yKkH0b4tLCHGqdO2V
OsBPBUdeTPdGqsWAAH+cHmEu5iIXgURUtT3OWeKRSotoXPw1h6p3ICXGjhqpKzdKpt/GablzcR4Z
6JKxQCgqRRik+qzOc0NQ4BsRYVwqoSdCrhO8LzPsQO8r09MZyTxbtwMeRBZ9prm6ILE0hP6HLU3b
t31F30J45rX5ZAH7Oe5yEyMOvnl2y72bd+vyQiWXAxkR7A8SUmkEKn6/0QxpmnxhXGG17fEv0hbL
HWoj03sinLx/qnfgkyBnj5ZfnxJ4W5IElRg5T+zvtAfmdFtzwfuFEmJOii8nZz/JM8bbIiI06JjI
R1VfHTl9/1vSOMdEYJSnuXGjgZ5m/fohgIs0gS6+78M9fAztChJnF7nSRd5qXI1YFGP5Y+Szaz3/
FGssnnEeSkDRvEimnW4DnHFINWZGH7+30MfhD/G1mswwol5NY4UKkNM+SIVvEdr2Imv/r4/BGcjI
sToiUWfADMH/wTU/BururBEZZpyUdKp7vAlFwc9fFPXYnC3KFtv/0UBXTiboYU8p+WjC8P16kRRZ
4CSP78RLVcsDHrGK5TaLvlZxf/Yrq7AfiseXP4k7fl+xhxbezB9Yw99/gnHANt1sE7RXjcqaJh56
ahAapjsIzKZJCMHMC3/GVH7yePcPtrjB7Om1lj7RoZR3O3PUCSlt4PWygKOj5yel9Z3lXDkByCoI
/6DR/fzhghjkA8/rHtHoC/3rdgP4oINCnOaYNYKlGkjBqGwP3EzizH9ZrsL787bUWtco06Pr5lTz
L0OCkXcd/jAqqza0vghrXDN0YH704OOcjqObQY90rTtoXkb0S63xDWHm1wgU2wR87xZsrzsAdenk
SuRhgR/VnwJn7Yrtcu/GG3KhWr3pg3FQPZL+DOTbsgQuwCzxX4p7rBPGfBBFwvsef1xbJ1QbiUCo
aWPYaCp0kyL0IDUMdpDJG91GrpFeQ8sK7ekkfi606Yeobqgbyt3g53Kt1Dk8P9FhUVMAV/oXfoO8
YW77u22Gfodkx3mw8jBMSuoEhJwCDmkoc1vf7EvQNaTyl3oabP67FznvSVbx8fr/lgVqSqP9ydIY
3G5B74+iQg0Znv6PcxDfBHUtPqVlIUH2bkRjNrUMczRbzQRN+PWDCE9VyfsC9JyX2Qmt+GM1e2C8
vQ6Lm5Bl1garOCB3RFbYN+8/1hAiK5sMDX7hXuoWzIXDQ2rz3duNPQQcvPOP+A9AED8ji8fbjYHk
afqVhPEh1aP7C0xLwmosxL2f0zyAHIBRk92wgR5s58Z4SH0z3f1ENZU1uWBwvD+xgwOW23BOZ+xj
myWKra4rVeWX5SSeCtE8cAQGeHtrE5CmlF8V5q8f4E+hj+kk2Ndz7A6O7Pay9Z2xPsaX9Hx2nu4s
6NTPalwgU9CrKurOxTYKjYOr6oPPFy3F0ZuEr9hE2SFpLCJT6ekof7pR/zhtFaqb+0Nh12DVYOyo
AgCpD5M8K+MtCq2EKOVLp9Wee5A810VLbX5srTz0lKJfJayrflMCWa8XmAGuwbOAJINrDQ0tpDwz
TaqD/8xB9PcBNvNMPdhDzs27Gm7opSoLWbsbCyjVl3uroAOQ3xBXCwXq2QkPcVwEa9P5Wrte+dr6
FaX9Bh719wzh3JXuaXG9+w/vryn+hy8gUP3pPqzojsTDb+l7VmaA3MLqPOW0vynizUbyyJMyD3CE
F2xXt834sgM4aIgfEUCtTFPxKA5ZIp78Pf7XIN2vKXEVBaQWMERxEginvigGAjGGx/VfnJ2paM88
1DXGUI/0Amw0CggktiXJ2YjuohijaHoXME4IssAYC21UEzdXYL/uyfatqYYo3O0oM5z5rj2Vkws8
JYFMV6rUQZJbry3CBXMbG7fmQ7V0+Wr5+HsVsmaPUsGRV+oWg4tIwRlU/6WUL04EBDSIonqA5z34
iU6JyiKQhcGH2WQ0NA04q4Bd8XvbDOAYwfrm6uN49o9WFuKYWSBZ0Xi3GCVGkhlwar5n9MtjGXM9
HIDYMNwoThxokDj0+RtzMRBth3ttNocJ8JiOII6FcQDyrWdlb84kRyoRJGd+folR7d1cJII/h2rx
jeIdXRNhwo3AyMj+7Jc0mwBf1yKxtifVI+Ql+tk1g3m7KbVVlI3tx+yzuVifcb5WXwGiQqqNqNWF
80rgfiONLQjrPGSQdcbZcIKsqlBxUr0TTBIXdIemjNQf/aOfr5n8sa26w13ESC33X/Zoz12Q+UtV
nS+pTpGlI8/Gh+TjGCdB3Ev6mj+6Vci/rf1ymkAmNSSsoFqIdF48azjwvB8ne21IJwEYHEEzVwxR
N9eI+YqsSKSE+UTYVnHEf6KH7oB7vubhdzVglY2IF75CAY72wDNUQENEBUqDarVrKTI9td+ZUrpV
jvwe+xS/H/P+8RPpqxAtKheaRthg6g5CmYxXC/29sF+PfAYfSp4fwIBkrUwvors0qoXUBvkCg3s+
KuvLzMLK1cJ1tcm+m9Wi2+S4uj2hKRxSZs4fUmrweRsEiZEHmB1Fg6JzP0xXTLHmC/HrJZrjIjpr
YkLNhyXD45tge1w0/0rJainl0X1TpCjYTgK99EBbrbmRdfqCWhGnfRYzKIJMGX6C3qiFpgeBhOHL
HK8GHx96u4kyNE4we5qjyS9PhlCX3cSPXf9gzcwkiigPm7qinQkaqUgFJVakcmGfOZiSgSA5meah
Cf+fdB+j/oZyc6Svv0RUSWo1bsBrAAmU1GiLT3fTMvIbRBmQBj0UihEoDPlW1fFjM/AOhbd/Cko1
/E2t8xC0J2nGneZFZPAAwnVKjex6Wmh/TRMHZ9euT3EZrmmXM98eqvQQcOOwVsR47Arx0/AMEmo0
TfXA6Rs2rU+xXU0q47hK0ZHdwUcqJeI8HfWz+CLN/I7lco+IrQxgV1oPUPj0q5eltYTkSMzdADCY
HXJNyJWBr7IWpJx4/YCoo1fZ4aXkL/nE60MKtCWs9wKoWnS1GxL/VtPU9EMp3dSK13Ec3wTFQj/q
NhabE6IKVhTTo/WDluRR7D2bKY1bWtChZGNu+To1IYtSorOc+/Q76IKs+HHiL9Nuq4/vANrNsG1H
t94/5ZBMyADHm2UJ/eQqlQ3InmAKeQo9pF5LQDiHliQkeNX8qNdsAXtmrG9WI2sW3WP7Bs6/6Lq5
NKcfhmZdrPqp+tUTQa5sbvFDDM8WNhvm9IQNAXjkXMX8l/7JnA/OxbPuX99mQbPMUVE8um1ra42a
XFZnpudDCyXIvPNw9MlSKN2mG7gHKQedSGKsTQsfOd1I+ohzEtyQs7cI2wDDocEPW6MQnmfFBcE1
fb4RstMU+8Wqz45rDPTIBQNIBPoIOiaOP2hjg1fRNwOrrk0akWY7PBPcoksa2V78oHcY77s67gEF
vYnDD4lwg8+nFvHxMRRujQww3OA2o2f8ijx5mUIWy38l65HH34KQiapF+29IttaxCXt+uLt8P/8S
Ld0YX+JCfBYNyEf+oFdzeA7OwOUkPfUhmutiQLxD7+PbIg3oESIQw+tPM4ySA3g/KOGteczobxjg
GjC1p7qTw2/k1YP/tli+qjiNYDfI3eMmudo+SDVAjoRuqSKKlHGsxsCALe2uQDeKQrjEVVQkITdD
YSYBygh7OeQm2CCrHgX82YMoWa/aVUYtMbUuQwucFVWM98p3t/FVjUcuVUaxIy5JqyeVapJLmjSD
3v3t9AT92IuhRB9ZRL29lsbwd0EEJPGdXmEkk9PGzjXH+cdYYj9UqgKe9Jhvb2PCL/VSH87EjXoL
jRitHtStl9hiDtFD+3wLRNNR3HdWaKRKBQBM9fH2C8tRFdsZVeBiBffCYWfKKKZfzzkI5xE4H1qn
78zRK/I+QyJ2aROMNylA6RrFzo+KeuZuJT2YGeNM4OgximjFPXAJC8rIPrJsOikowXeXb5skAC1V
2msckHKrIQmRFvp4W/6hb4v7r0CbAm4JdN517ho1LK5jbgRWsAWyNw1meV9F7t9XOTbrDyQTYjfU
BrfMAusOjogPtsHNJDn5HPEwJiV/e0n3NDyI6kJ8HicrEdyaa5hQ8OdkX5f0dtLrHZrGjBXYWvup
8Kb9wadYomo1q7nL5krDUYdCsLIsBfnprvL0np9Mu7Azk5dzG1XvNfjhPUYxdrOXBIWQr4E2fo1q
nr80TNH3w6xgAr/98krn8CQwfPUtNowwshRX0ksI7tDrHxLY7e5w91LOzmQpWCvpN22aOaewuUJ6
NIdSWwQXmtQr0UdM+86guRdpJkuy+pfdI3EJsJfelA8azLebuEuo9dL1GApTXiR6oGmqUTyCde8Q
x08gCixFztN3OkFuoC2KC7UwTB6mQ6OLwDE2orTa1klxXfxmcTspoxj0XAlUAKLKUax2JHkNAsKn
Uwj7o2BLj5evxILepGb8NzQjyNR0vgUpwkyBTXATmoAKbUWZeEXR5crHl5HHUzutSfHlB1L1AUoz
+LSx/tC3xbkZnCrNNtr4DTRF1y2EM0rmAnI7DiFuAubAp9daW0XLmMJtSczjmb7j4930Ng9VP05P
K2vvMyJfRA/LX5xeRB1wkKbzwI50XCs086uZgjPgdY66uN49khDKizFljsuf4AdWVgthartlxxdo
lWs+OfN7fZwydTUcLt9FiTh/5GbuuDqM16ZSIxRZ1PGoOpGUyQ33ojp/HZJym44mCVm/4pvnXBAQ
9NJczZY91P0/mBx7MYYb4q4PR3SoJAjBrCt3vSHW9BOOAYFCY9GMws1eN5mbqF1t5MkfzF3i4yQN
m1cbTraAXCm1oY2/gS/X8QndTbrWwcaFyJRXg0GCKnz6uog6tKVg8rz3obvT7eL/o64qY+UbepJ4
pnvCh9Cr3IXBq4VDdcmwQwb2587QjedPhSuy53bN1Pg1yqVe/BmD8DSV+8eURoIRgkfNCW5Adt5Q
V/Eh0P/vDOLPOEeYzScmoyqsfl5aarQ5Gmc1fD68eTVYNaQo8uFduurzxE20MDxE4QddOl/izCxU
rwPfIkuPhgWiA8kJ6mBM7/pdWuKzW4bL9Xqnv65BJBVwQib4/y7swHpc5IkuGWncweMJ0x19o4gC
iWWVdCuIDsgPiJIvTWyKYcCobZboKzzGynUA4Hp/+vpYyTqrrOOQs1RDqiwiu+KPk0J4/pZZ/N9g
zLUGhj54GDxGVc936AuCB13zJbYzTgTWRjTutnIVwWnQDPhGz0MNn0+4HOHhEIpHy9rnGea8pQek
sjXWcfAAQyRuXtmfaZ7InG1uoxCe9PXfa6LumaOvVb9Z//ymA9b/U2HV+7vHBpy3BtDEnKlAIXdy
jSTKYHCSBubDhslnBU6FqRM02Fs4OViDQnjS7MynDo/RUgd92m5Ae8VRxIawTrGBWxZXWcJ40dZB
3a0QTJzhFfcYHfms8bmEeZ0vGPZ8nyTmRFproJDQW6Mt3kT/0Qh5hb4JEjvwwstUvj/ssDZeoiwY
9rEQHL6DXQyk0kN3cxQnxdRFqrWd5uDaJPprxONu/aXZRjRAsm0yB1hKl8KNBfQuGzbSUPJrAN0A
Ywhl/FntpVbfl1N/ybfTZYxrD3h/c3hzjFxWDKE9ghOhvwHl32/G/mMH8a8hpaNeSHV6Th1l/cko
jAS2tDG30+0mW+szoqNWN2U7JlSUNYk4B53E2LxV7s134rE7hXqdx/gNYshDO/X+2ozvWcFeEa02
uhrF+p11j5GHTa4Dk6zpMwWLj9+SEMoHxzy7WAirHjzexI1tOUq1ZFUw09mG2gqxHMqxF3pCm1Th
0Hw41eVU21Hxmufw7hGhSbZulIa63tM5vAV8lP364MGb+conZpilmZMrXQa6xVppRI9VXSR5Gmla
m7h5T1qWbvF+6DbNMRggv8In82k2XKyyWEMxVb1UUCThQwGFl0ythey7WYfG7GDZd+jjtUMcyDvc
FsNRKvcML8lyXRybI+ARZB3t3wS3pbzkBt7iphcELczkKPKXFsAcN18QAQvQ/lbUgBZrDeNBm3Vd
yW4PF1hIZAuLJ/UCoIXIrW37D+gICqalA/hJrp7LiNrxRlc7iXsdZs7PECJd1Vb87Kodp7KungUu
cTyDRt+XPN47CoYyhn5hkVfaLvIzpH44zdHIuYrjT59ln3oTNKlZFVQQqojyDdMaRGm8SIajemr/
jEDz1LCHaATu2F8AS3Ny18W9ccHPPDxc5uxZUnZcD8ItZsvX7/n6FXNe3rzYPWzM7l6PezkXtlM9
aYyjusv/QfS0xA53lPvG6WRKNYHLib3PhvP2KQH245iSH5pF9xjxROCExjhjL/Vk9SITruGRafLn
G9TB5ypGWcij7TQi1Ran2mWS3opAw+TQbIJFzyolkdLO7x9pgA8cdhqefDFzlg+GfH8urLoUbku/
RQnQrgR+ArbXqvy7v+hA7EF02EON3cL6jEndeDx7s1Pg0yjcx35AMkgKQE2t99ydJpSgw2U/bJ16
sQCHhjpRtwkXuWe1UEfb0iT29NCPfps8AeZ0CuzZavtuCUqPOWGceSOGzmbayOZF7Z4K7W2w1PSm
h2DCZeM9AG+4KAU8S+kLlRZPx16zXWwBdYu8mAqzzTG1GrdKiYwxK/+g7x483RF13Og+NpEH12b9
cOwIitpj9Ns1xOEuAjpvlPkd1QvE/b1iuoipOrwdnH84oVaXEbyR5F7/8BTIXf9lXohVvDoVq4bV
R/DL72V+0MtmS/4EWuNq5E0thB2B8Ru+hEIXlnSY790QxWaxiePRH6h6gdB67xmTSmc4H8g5Zqbx
w3sHj1+vCdj2DD792h0iTh22lymmEZ5iC9ibKOM5iF94hbLrx2SPv94/IPKow6hPplGXMjEEPZNO
KcfbgZWitk+E9tbdN0s++Pj5bQLX9ONCgmgz8WX8iDB10iXF2TzpeZymWexfObU3uUn2od4ln6Io
oxhoCIWSBNhcWeZJNAuArDADjXW9o0zkoFbOxI2SlsgmU4POTVle1pWgOGF+RBQGrumyw/jBiHsA
4HUeITNldQw5jMyHs4wZaQGimGBeBphaKE4Ukr6ef/IdSOywoz/AKTyd/oB+3NkDtgJ4BVHoH0lC
uZOou3RfGpH0W5xXnQB2D5UBsy1sHzbuYY3YRTZ76Tr8rU5RtBvtyEIqgPyztMAlPA6PGFrDCj88
7q5kodBK3A2P0C1RogHmLw6+dwi+QsXxHTDR4vnc5JRjdDaTFEt97x1DDJBnz4yng63zxGTgfr9j
eo/D9PTN6HOIBuOXWvIFm2xLs6IgvxlDyg03ndWtbemcRYIPHMVo3zT2X2vkf2k++RoxnDgys9kg
TUVe+hzurTcJgT3HLT57s4aXgcIqGuj2CrC+TiL3wslO23zhUkI9iClh6JG97iJvGhxBiv9kFFQu
6TuOJv0ZXgpTVbFOeJoUsoiS7in8QEnqVYED+6q/BqN9r9kPr/ju+h7c1he3xs+owd5Ui2WXhmTi
+YGuqPgQxOhaUiCNkGwOCXE1KRnmL1mHaz+BlXizq8wWSk/Gjq4Yh88jiWSvtlYOgEtdPNt0H/Yj
4oJGI3ntdAS/kUKktv0F+mkBCFBJ2ZJiD1Lmk60ranYudtoEdEeICL3oLxVcJQQ4vOkUNcn+09Vr
WRCUCrhlp6WX46kcJizAT1IJEzXP802mDhd6WyakO7eaMeGYz+sgbvbAh9sOz513F1BfPinbHWVt
RYyZhAkKOlaXkGPoQhrc15cqmHuaF8sa/cGjOeiM66NgUmg5ezrM/ihzJ3kushOTibxDV0O4Mw+G
85IaypV+2MVLVYxJfSPcz2MsxfMt7O0dYErxfbsLdKD9I4AyCQsXBKo5AZ2BLnsyETiE2Wp8kPOY
OrH0SgoH+NqV3WjsZSyqtRqHmrXk/PbY5WFjYzlx4XPOlr+p5+vQD3hfi9Z5SMJqeiJDG5NvDxy8
uJ48FzWXQ+OcF1b8sWpgQZGoE/4SBMKeENLQDeBWYiOr+3KFm7MNT60IqgkP6wh3GqO/5whnq+uA
60HdjlbrgMTOYlNB6blrn3QBpKQBHMDR055h0/71QJuXFCnEheDH2v3AhDom6PtXi0hIJ/yTvkXI
igs8dwU8/tUaIaHd2HU1s28yGZI6p1Pi/5L+qwsL5YVFAPZ4w+X1QyqybTTAOU5/z30WDdFPA9Ua
q1OLV6CgWOUexRVEzpMqIpRH3Ej4o2+ceVQomVDbXiCh1nroDQFWyjEI14OTH2JoYdpbhrjJKiFD
n7K8isPAVX2B/fc3tQxz8ODYlb0p0vKFJUbNw6QyxkZJq+AVA2wL1Lob5Mw+I+MVtQASBLbuARGd
Wb2FzWNC3Bub4Zo0pgB0eUqlh78TIOocQXultTTgg94o47k9xPwEddfVpU4lE8o54TWeSxyPpoV8
h0b2blj8OhWVTypnGP28RtU2dapryeJosWtN8s9Ch32j/F/HCV+aWAlVcmfQEmk4FP1DhbNW5qZS
Uey2KI2WoNTkFetUaRKEjWhpSRhA1mE0wt9yM5+eY74Y+mCRcjkb4HFO85nkwo0+ecarmxr6dZgx
B97bn8Q3KnoxUqmvF81bDZOvQtuWye8mCGhfqfGen41H2iwyiUfik8+Zi4iYUqfe8ZFO/jwBDxeK
QP48V/D6QbCTglFXWV5qhxMbMkbJ7hWsODN9hI0CkgGw6QeAByO8Yv5JfJHVszyMvJ9kG82krh0L
MxdL+meAthxylTdoK32Nt5rW3Qebeesbwg1Jr9+KdfBAVtulFprQoLRRZfZGmKtFcCOh7dJc0lij
BhsyKA6Mv9a4Ex4LkDRBpn03G5RFNP+sh1U4Efb/DPjcc/+fn/9bg3HJiXQC50OFSpKisRUizcpv
AIV12ERBjOp5xr4/OdI/FhIGHZG/noK9oIUbGmbodTqQlO40TUrwexgiGXfsNRjS7/1l6zmaWVuC
D/MpacdH2vg7/+l6ijZJzBqAtE0fXrTruEhbVl6vg94zmSaLLth+GB36Bxfvzf2IahMFz7m+o9kB
TNMPnSsOoQ2bFBSzB/uUvGeZdSAyGapNUoeg2udFd0ANQZ3nJy0qrH4IWrSu8MLlxRzXlivupPTj
sN2AXm/qjN9pHhRPTht6sqcTL/qaexKR2wrps96DowXHIFfkOMP/afnJN2oQRc9RoHGtBXG7aZb7
lxFkWN1lzeaOhEp+DEDHyEimwKod1rAfOKQcwflIPpe/gbRiPBnpASkWaLWu8E1SyNeVeRx995aC
WqPhwZ5YaNCv+kw89WQiyimn6nXTdVgcrx9zFYwTY++we1HlWIFau47jatBeEGFzLD+cxt6lB09+
8eyYJmsxsKTfQpQ5vMwzK87CRHXk2d0DAFZZzy2YFKD2DPaBXk7hN4DoX+t2avC4VvtpkZ8ZWzxv
Ou7DU3kdtWmmmAY7BEsda57e7c1rTHFwJL+ugAY1//fSNHIIABa/o4MpEfaxEYbMUOYJWJuypAC5
S1fYvIw6Y5JuvgRvqTt4wfQGdXFSo3tJkKqchdYThva8Yo8R9h/WSJtkXKQTHUrkNlm+tA27X7rh
eBqy1rGKGBbCjq4s7/exV11c5Z/IRf6WtAx/lAWhedN0CAQyfn4BcxI3fZ+hRG30sObWDra3LO4E
TY7U77bzChcoQFu0cb5hpi7SAMSlWjvzqdHqOJJ1Ho6riwR/rK3DMGXPcyCu2NNvWpwU6fvg+qWt
nr+qzQOBYxWEsc21gMmFdKGP4Qg4k77uWjK2LeExkuDHdACMOVkWBCXtCk7MtwK0or/B2xSp/ESp
eu+91vbmUaBA73gHJshtKExz0Vq8wztUWqkzK+J08zxk2xhf2DRZeyXtJ90znp3eRM8OSpxCzd93
gtElpeRbEArOpx5DJSUuRGjNVmRKum0s1YqhzKnAXtncfUUhPifPUPYvKLrBlNHc7uiDD4jLqjBB
OOlgJuuV4DMyWw7BdWmpIZNlA5b8q6iDmdpCErxR/J79ZSFThB+3BwhOKG4Suvk2aqj3fyjPYojm
tA9dVLRpTG7gUCBsGx8W0YtJXMxbpoFCema1yTOSh84JrRLvIvLElb6/MiI7Jlvym/YnALUgZ+EA
RWM6YOH6qkjaaU+dxoiLHjF/ZDU8MCJflDQ0tgqIX9lhs4HAkehizXonFGjHE8aNJzDyWeIOdoo/
W9pzNYO9N6qfFeRUC2hhU5q71EQfcGhHnwuk6DnVA3l7fYaYYXdm/vu5u9+gzTkjV9E4h/Ovz+ze
HnOHPyTHLd2lShlclMK/iIsAMK50MiDbIbsWiemki/k/ErndNPhkGB1S3MBE5wVc1l6OvG/gyTod
Vglnh7XfNIkMG/C/Y47Z02qdvgt15ZlsXBAzQGZpx6UWglq7hSZmD3BXDdcKEacxxYbrjylVilkq
m8tXohMeSZU25+s/7cMNmCHXJevl10b3texehEL8HkVMWTr83FZbDcVLWg5bvxTkDOKcCPvvVJM3
/Fsbvhtz9gU6dloSaUoUhz20zqPSVhJAuQeaKqIogA/ajjGKf1k1hGyCXOERO14krZnofkzm6h+M
7XaXg/4MTNSFmyinNqxaax4iK6gGFz1mj6UTf8hbTGWpCtD9ZnzUS3/ISnylP68z3JDljN/7W9tc
c8Cz60rfYIUBiwVwpemoVqxlU7BmhMLkLplvqCekx1gpo2j2YegbYtOiWxd8OpKbFlDkLtalkl+u
xyuH8HYlr0n9jKPX7MA39OlaEYuVbhyITFWIbPHLsDWR9f8r9w5VfVpGNPf7Sdn3e9MKFNAcwtZx
T0nsPGFvXRMXRDYkkvDBiuft7XRLLK8eq6ENGh7rw3jRZtrL61B7FZVjlh2XERYwsQN2pB9G2hY4
NHN+AFbcl9SZaxO5CBcBWz2Miaa/O21pibuJszh9T2oGCjW9rH0nLgiGAPD52g9IwO388kcQgcUQ
3y0309ZF/dDeo7PeqS+36rkjiPH0FIFPY2jVZrWh5w8KYEIouwFZuI8VK5UTxuyCOz7PPsypKWxS
ZtRpQmvx+gW6/7oJLs9sLSjpScrFyvtH+u5mgs7f0AweShF4xxSDVdIJA5fdk+MylSUjHUE2BAAr
O84efpq1UKvZZlCOGF5i243Qeap7U6e8gnihq9CkwoNTGbqHXW7NtL5T0Vl2rYQxCWcxI2yGpByA
HcvBRVRPceGtzFn/lyarWKutYbSYMW93t6urUhof3u9KHpOKJPQaP+8aneoGwgLDl2tyqzjSdPhf
ZogpfhpOF6pNF+VYDS1qpMWgqdoceIUsTr6MkJwYORks775XX3xtnXNg/HhZSszubckITE2GUP0k
O0Ruv98Or7XbMo+zPM8w+J2ZY+gzDRyTJE6zwnWWezXrfW6ZgTf8TtR5VZS0Zb7huvAlAIX8YDue
ioYBgFFCCvTsTYcVxPLEtJT2A9Dfur+x/+w4ABKEUbdiEyIdXz/Nk0JpvBVc3ZZPMVMNDXmHcxcv
Vv9uaxomfbDPJ+41NfUAvUlyohEfy+S7wN25PvKKWbW4DGisLAQqNWmuJtXc8c26yMl2F6UQniRo
lP2hxJilIj8i6D1AKaqEWY7C3AoIsk8SyuRUiOiG/5fUDZJmoL/39vGxTIMd8nYvN5LhaHG8dwLV
Gyn4+b7O91OiNyjJxcrLJxoYljtE1a55uLWVPGe6gdmUftcPh8NAdmFhbBsKyvDNyVJl6+wJakD9
uxJIkMkFZ7b00G/M/ahsfkYTScR2wyrXbu9f+EB5UHpDUeK8cRhoHMuGbz9MwO4mJ6VvuLi0QqJL
SWpa4pUP2rrfOYQeG75qmc4GSYJMuKqhoYXQzrkQlF2Rdf64bZCF3jQWQr+xg+aTzdnbJ+rdS2jn
cjrFwLcDc4g5bcH1hYr92Q9jTmhf8xge/92wqV8EmtTswphnPY9ij1EUv8Z6A3oOQCx0OdI3UA3a
hNTpnMlgghsZlf7SxFc8fRIQ1VrSFpEVa9AdSC+T/GjaLlT20aTUiQTgj2XYZAEPrwF6UoUN0MB3
bGgcrPXYIuuds/BeqrgY/223itFL9qbYYiTc6NN7iBlHG97Ln/DJxLxXi0GMy9H+ewZkIsBBfaHB
u9atppFFSVDzu1Y0Hl+Z0S4kvLaylUQfW8EZvw/ALRcuI2hsP87A7Hwp97g03y2qk74JnaVlNy7L
ycLSY/71iFF/JQXgBEZeevjlvWuZMdPnq6Ps5cpBeWTxwJ2zypKdECrk7LXjFCtLD2fOmFldMFc1
DHVWbcwMqhg0Q+MVwF4lT/B4nuPwIzLn54ITTCZDSRygxO//2k2VAVdD6shoKSUTKg7oStWwVs0f
ea5pml7C634DO46+hMNNFsxFX1+HgLZ8ZEnIE2KD4/EB8jsU2hzwMa1Wl8tEFMVy/ZBZwBOZ+ni/
gVDS4Wt9JGBOGRgPRvW1Tk8tA+5nT5hjXbldakNB1O6AjgswnfNE/FUiaAoJ/dtqqUdZd8nv4QH9
tw/RJUj5yoQ4gmNo+F1All2NYp8Ny144krLWMXLaXMKLOrZ63GgTTe1E7XY5H5eAiw6xFPpQ1XuG
8cPs52WqrlyPVVcHQ7LTeTS3kFPx9vuk0UM3dEeF0j2vKS/ej0ze6jxynYwVcYbG89SMHd9rYMIg
AdZGf/+OhKNDo6mov3SuqtXKb8xIP2SwXtp9Bnld8dLdcLWEH/NKc23vFUPISDjMGmIY6qksYQOx
Yv5d5HtAlkqj9K0mkPYSjnlHg8zj9dmOklHoMPuTEen8rUPPef9yYxrzOqUKEVL9l5+nkO0TsBsy
zEQC7ZCmGI8eOMwG/fUX4H+tuA43FK0pTQlvRjmmOF9dxdKNhO8fjEWrCGYFeubqVfSlYwpP07PX
L32UnaGX+TBf0Du8FrmZMP4sIJvZWw4rdBjMfmMH5bjG08JQXZNsTg/qfguZ65X9SEihaTvb3UgG
ygPAfljXK64fVGp+QmZrDgbvfefXyIBmRp73zOd61MVAaA+SG9VIVRKxIdjcEkZMmH2k7VHJWyF3
Z4cfMFlf3IKbG9TtK1DH/BrQu+TtetNZskI/AwKDlUPmqZ6tVg9KIA5pWMBjoeH1w79nTfwmChZf
o2rc8vWlDkXn/oixKM/wxbmT112VL1sD4eMBj1JnwgmmXnOUjyCADvhnKPGwvBGFWAB6lufF4eMX
tSW9Iap4BRlNdxBRXv3jdxgpN5KqmyjroEgSuoEuN27SyBrkl+PYjNVULB/Zl1CJMFEiUSI9a7Ve
P3RbELmrJsOmd5DjZX8K8hGIj5lbxHKw8vtK2LlRJp3Kvskv9qrmu06GwCG+/JygJGpA/h/Qhihi
hy4yMMBkcmMSqx826oMUJzE9LEYbiStpPvzBWqrsFrbUlPpRYMLGuiQxZRVX3P8z7mncZPzDtkpe
SP1dJ8vS4HZSnaVozE8HEXtdrb4e9dpCDId377rvIMw3ndM8bmdgerTYKVcIEjKWZBC1hh12B3+8
7sBC8A0OTbTwJy1FQm0mYE0qzHuWk8Dcnms8SSQDfsmwT9KP1GSnFxo9Z9gS56fhq8VXnydTVq9S
5eNCqJLvWR2jjKfIg54eQ9FaLSB2pJ8WWbz4ieMHIC420gDEIZL4GmJO0eRKiEOhfkS/8divcwU2
P9N57w+O70iaDBjjTrzi54gNKeaVgSw+bD18jlQKyn8zfxPAoJevK/ChPcb0v8CtmHaxCT1wVoK0
+MhSNRFd+iuo4t3ieym++UgAz6jzeuqYc1XMMblKHXyHH8UD7v1oFJF/25RRrBJpAiaWuC0fZedR
I5ZVIxRV0ozM6/sktkvq2MfKW7am/q0rpLCCoIpRT9jD0iYKfmz6Scf5DaoGknosSZWMiXMsGnan
fLtyP7QbG83cqpeLqxyn0aEyzlvt75KOmA4ykJbne4CIcIhXb4LMunK+RHHE4RVKgl9HOXX+ReL+
QxHZBIIDBq3kOBnkKaHwqhw4ZOFp9ObiEjrItbRlhvscwTS/hYf9jZOHsUq/J94dHNcE3rA42xap
Y3BIn4TUv7HxG6jq/IhfEw4mF7bWxSe/kzP3tTb1x8sNmzen1ejuZbjT6GebQKXIhzqbhK2XnH/u
BhKhggHzzXu68RUgJ9BrbKD/S6el6jxr3YRBx3GOC+5I/+BVVbQ5Lejs6ioikPn9+uaDFdLLD6t/
+41Jsm8nt3iwtUFwfhJEsVRR/EL3jMjXxykgL7rzZfqoWOJhsffDRI/Ks0I3SFeOsoOQAv1GVgSK
RsVvi3YpTaVwPRycPNf4hcr9NT3yDBroVJihmaIuIwuDtz5XR1HJj8+g3UOuqE3LUhoLupM6ASSk
/4G6Bh8mYtT+raAH/s//Nr1Q4Bm+hkEq9j0LoHpsGI0uGqh1nA0Z15vt2zCHFRqjM7Z2nRK/vSLR
4gOVW/0qhJgXU7lK2shLh4WW1SIo1xpGRHocYrdLhmkEWRP01SiRjRFZBz2FR4aNgB51NhuGpi4E
0IexF+3+lgy6F3aV9ukf4eEm+Bg0k97q09Wmdwo9+J+/fUjtkZ0FUt4nV9MUzf3gBiP9wKB2gtyF
tB25gejKRl3u46QjetUtk95aMUjJVBAxqKsr90xBK9GAp5ycfcmpRLhdf7cgI+282R8s8M5yaLK2
KCUaqcz4yrfOsJCDLHTVAa/0P95t2JyBWZJXDCMJ3yGtUj9UHeIG6H9xFGSk/PEOi0jzZq/GnHaV
ka2PZXeK4f/fgGRiPzNUC7IpPOTfFgWW0J3kN1FUQuFVnx7xL11v9IyimDtLWZS5iN34wh2D8qnU
ReKiqF5+IfTilBmoNkVhoL06S7ESlFNe+i27LjF8IjDNlVaYQoyDQMLmrwnJXKpHPN6YlmA2h35i
GEaRVjyWrapDMrbT2cwUpU9EcNtypVe2HfWqDmPAeaDGgYUZN2NnxdT7lx2mXr/l8F7mys7Vd/sf
Frbeqza7cD3wUIkCJxCCx6SBqq/hdvVvefmU8RDyxJHouRO9k3ILYVGETx1/sVTVvyJPz6e007M9
oUdk4E5ETEauxJJojOx8EC8RuYWOoVMxQlcjE7Gjg+I/VGLUmrJbAa624GDHB/sQs5GIQCL5CAgg
88IlNe4/eoVQH4txE6bwHdHpQ1WMxvZ9FdVx0KVrk22J65uUdpvmPO4NQ+Ip4JNaRSQrrsfeDeYj
TYJBnNhcM0hikQVq6pej0OltNCO7ZXpepE5Kg7bLQXQJyYhFuTv4RfRRqqq5+/AdrIxGpxfKcEIg
SExQ3+baCJW9zVUuSfg6MPyK98JAVgyQUC0QgsIYk0oWrvww2tFTmDMpjMTnUzDQGZz1HHAsDN5q
7QOOCG/KYxvrkauLm8+TymbCy9pAm9yigZZGMRN0/NcAuK9y8Lf6yT5q2qnZxdzVJGFP/aVZd7jY
MRwGjVvjk/53ThtcKY49SU0dX1mXquFDmE0rMCldMI3aIF4Prp4osJULk4m4eiUo066ago58n1wQ
CoXE9tpNWeiyVakhab6nmaCLJwiUZNi1NI8O6VIi9VWRx9RjTu6wKbL+UQP/TSZzWw7GVsCZ+fmj
Rph2l7IdaqzYK3eHI3+V44CXhBmwTNB133JKKb+mHtd/KqnHyNUkfzwkI4WffmHAXPuvZ65SKfvt
8WKRN8/9nHDO71beRX8bTjLXg28ztyV6gYikzoota3mOVWmckpkrIpnGfTo3nkeLQxDBJqBAsEnW
6TOfO3BD+t4eRw8+LT4kXjVIMrhNxzsBjKrAFdBCCU/0HVs2YWGa0NNdELCUlaL1iayqG4UNRzKY
UcmHHxE5K5XnT0aPz3tHQbyzHLaCeVhGEDI0eP0KA4bpqSfpj/uu58ayPpxQoggCIQbANnxuefsT
/T/3nsi7pk/d6tdky4F/zu8re8PGMoj+wtGR/pOPasaNyjhR5Wg7KG60+PX6C3tUi4hXW9uczYDS
pOYEOjC3qXnbPtUhoHlTH6hxnBoYvmuUigqY6aQ27rqtBZlfh6GI9BiWBxUCQUkTEodYQCkRkzzJ
SapUVIiwEDViea+8Tz5E2NjexCJPIKYP43iTBtzjQX7NCfncYZ7I38TjIUFuW2wc89RgLuFaRfuD
mejUH/lvPFsukBoOE/BW4fJLfOQRbgz9CctS6/Tl12Dy8fDRm3BRVQguY/sIKVim5v2D+/eiY6fS
6aYNIpFVm9esjbFQj2kKvdbJDnU+T3tKoWUdt8rgE3/zehtJb7opy/loA02sSQXQYgSt6UqmMivl
tIk+Pm0e5Tuuz3Y8silhH83IYodzno5XWrHzEvIj7N0TKWQslu4u8Dk2kko9jnmHqGax1NqLzBMz
rCNJDfyGHZhgLh9XqwY3Lb5RT1U4XRt6XG+iMlpFvzmM7/vEQk6AYmSV8DPrHoSW8Vva1gGlbLGx
VnhMkXB5/v12A+VuGR0QG52KwDavJecnhwKR6lnhAkJQ4xXTgvAZs4aTbjTFMdIUxGSYl3cHAKZn
IjfJO3CeLGa00yZVkL0B8WOxHmGpQDJIJTPXJBOAc52FAUqbeGnQYjsJHaFEkzMrDK6IFPtKPzzw
pF5J8c5ZBLlNFGnMw/xcdROGI/TA6lADFYz+6QRYg67rXDRV3/HEas30QhS/88ebRG5JIq8kvKNq
kaVyyc7GDZTE/IP/IFJk4aKyyri58CYGZEVFvoY+QTOqG/gzgSE6qiH3E1l2n/0b0FNQMGJ0S6up
9hywExl04DWyK+6V3EmU4vRRG17Vgg9WOa5hHbJmOq7uQj4eNPraSqHy+f34FuQU8vRWNTbDhneW
+4VYwCTNqTztExzIPaF5Lrn7GQc72C6qbyhRoq4RsdTsLBxE3kr4H8UnXZRSQtdhzSxF/d0VCTeT
TtRc0EAr4uA/eLY06NAAw37rnyl5WyhUxnea4RZ3e5ucVrIdOXxitUoEnHKrl8QrvLLjY2bNud4E
lfH/QfGzStYhV0aG7ngI2ixO2FLBJuNW50QozW92jXrm6wQpkX8b+3EB6zcq3JoqSLObskVp8UCH
/yRQ42rGzPvxcgbfx5XTlnXPuw1PdQPX43BMhuoEZufwb6k+L4C4vs4qV2qnbmplBcjGC3HJ9O5H
pW5UfcnL8wHjbT7nJnYtLwFD4x8l9aTXh6u0iqLBm1VzP2gadLhCJOFuV9hbQSq6nQrOPmNNZz6p
WlsmtAvLgjRFQ1swwPvvwUDOj2gVxhm1ESwedkyPh+SsU7qZajV4h1jnIXwU5bsz2Qo7W1dpk6W/
soo2hrzGnHrK6XlJ80IaDSnZPpg/6Q76OJhz9niYSu8B19kIaCvvN3DreWuG+sreo54ppCQpRZSW
EYoKOdT0iHvub34g/HCSQ0nEkugILAXgB9SzQHYpR8Xg+PNhuQLz7WA/e49fhlFx228DQ3Cb38dc
T6IDiP3vqoPwkpl5OHtgteqZusJOKAfniyKS7YAYh335WXPG++5t4jMGFo2c+w41oaMXom+j9sDO
zUopR1mlku1tYyt051E8g4+rxrznWx56pzC7grX+hT85/KlMlKA3Zo9xBsvFp//K+UDa25Li3JLF
br+DsNjRvR/oFO48v/9QE8xrMrZP7dlMU9aoDCyCq8QJHRpWKQrEpz+rADwbGbYwIcn52B9LG2EC
kLSOMS9OTAvTc823Vwb3K7aOkXPYFRUbf6yIYfjkh6j3TG6uKnxNedIHS6DNxSBkbGa630lrkDej
UiEi7HwiIHsm9UeP8XFczfCiCl3DVEffswFH+n+sOD0LoKCN4o0msWqejoEgZTUjMvXCfkZFeLOP
87+h1+i+zOsqycJUxZPZJMtOgUFsCtbiAXaxlOUzTTSc7eCCMZl3xGvfMjznxkDwqfdUEXn4ahmI
RJZVUxjAeUW9UJw2GiPpkBYwi+IgiWF8iqnJ/5fLKqVVV3BbOu5B4H590BNG6manRoBmUsR54GTP
iMQl0rFiaA9DU9UCXY8uMXnMCCMuX4u21nvANivI2pG2htcJmLk1Z8p4u4fVW+icAjFRJEnfGtcd
M3uz85ClTq3PhpV70HTrOKWSKKC3wb+qDLtb+8u3xPu1/TwstO5HtoWLEnuMmE1jnFFONIVQu2+w
RpX9pigR5Wix5SSIQ/lV9OV2LyyxOfFMTTW28s5zKeWyzmDd0aJRBh7A46jfygED//k/HsgsI6J3
xZ1cjIDUeiKtYTAE32niQ9UCeBKT8HfASS3lc7j8fzA+M74bHaQan2YgdoH0Z9JUoOwpowy81FxO
IXmm6XUwweKmJKeHKmw4CHbiOZ0uOS5J+okhkZVRppKzOH5Yxf02BVe7t5X9ZfmmKRIQJJq/znRn
GFxZiEf+ZhALvD3lzHJbcl0V8IszIpo3cF9seok1HW55eAJZwSf8r1hKGVpbhd90l4X7XoOvixHn
pv0wMSv8whXA2ffRv/73XVy1dVvptr778zkP5FW2gPbusMM8u+ujIysk++ehdpL2+EUt6HWHIasj
aFNAi1Xe5o1GQls6o4MIxy6bbabbqY/fAqUBp0pz3wD60ZFRDSNi18YnxhPAW1NiQ4HT7ZZliUht
JXmws2O+CQAUXKDWzYUAQJFW06lXWWckF5PuEqhTQL0l5l169kpoq/xcC5xG5LrElZLRR2NnI9vO
weMzCnrQB1B8aEk9jeDdz29krFFhXQfX5om1DCXLcuXDfSpPZkducmABJB7sfUo3eWtdBex/ebuB
O5I52L/NHx0N29zIiYJUTDpNDxrU+5VpCISNfz0WG8qu5yGjJUX+2w3SDnxJtnuFhELpk8Yj3W3H
/hiQQEn9bQWK/jknZpv3APdpxfHeNgyHr+bqcgCRuBJx7cfE7HdEhyrsS+DCkboJ2W6T7b6Qyzvc
SJKUUEpIYOM7rURUUlvbKKveXVtUrNl3yEVtDsulWUcfiyK+hJ4oLr9EmZ/d8MX8BUFyhiPThbQc
/EIfJYsK1O8qmYSMzOkR4IM5Sjl1CsnC2rKfWkUnmeznlwP3m91NMCCDZmkr/3oHoPi29kojUFuM
4yiy/2gZ7D9ynbNp7IxycqP5ul10YDCi3rj+Zjhd79CkCjR0ZyiwoWOVQOLU4c1rlCvji9vTp0x2
FYVJRj8Mm05YOII5wnUc6GT9Us3HrPymWG9vpcALvdKC9Yzt5Xv1vjvevd+7pvC/BnsmNid/xXZ5
Wq0mv8mp3TMrmllaPKaLWKzDGjHgbR/PMp7RvKLd2Go1n4cLJOPNAdc3YqhMurrtdbMo/IwP/U5H
7+LYeLH5tNDTmm9OpVuFoK2wU7Z1YHuCCjeoSIIbzvHmz4Xc1kF+W9evjSOEygjNxVu/W74Ei+v2
/+WoAQUHZLVxZmPPXsrp0HtJNPMoLvn2o8Mszk9k8o30RREZ9p0WsH1WKJ7DU6qoyvRsk/5WhpFW
Pt4tKTN8oPWKzzzVt5iOWe6b7Oqk5F+CAQtKZGWhZ+6zMFQ5ds60dlTP4UrUAIoqlDd0YlpBY58i
RzdHWkRvL7bmIaXEO4ZjTcm1uOcEysI314j5vxmvyJo+wXLomnAqXug3oAOTsziBOhUFM8/I6fG/
XPb0Xz7lZXXOIc6VAvbYuHG9D89UkNhGzamXMHqTlCUrpvDXOG8uw/rpiBhl/m20xbhr+PaGfcfa
kiwoyV7b9mDCzpkj9A+KnVGm6dZynhMhH8JJtcknXWhnbK0zFDU9N7Hh/sLUU5B44kv4FcE7sgZt
0O/Lr72R9kYl+EyUAdMhGIqhh6HeD3f6ICQ2faGpdgJ0QA+OaG9VRXNO+C3Jyp+VJKVUs3LUEa9v
qOUm1toYKKBHA7ZedsPXGfbttvLJaedcFy1aN3DkDC3PdjdUS4whAWX1MTrwP64lKf0EfK6eIQQ2
IzSbHmN6j53+JlNL0lzc+ya/4O7F/yADTaaNrbHWcgL59OJ0jRbokoLqjvw7WG1YgtNghYdbS1/R
Eu1Pwo92il7Y3a63FxjRrjNYeRyaBe0CSQNUWuw4ALT+Fwvin/0jOgySAMBHCGR8p52Bx6ey7M2P
ouOPRrLQsTiSl6c6EUxoeDFAbE2isTHKDwznR4/x1/rN62I+JyQarpd0RsJsg50Rbe8qLBGsNUi1
ze0tZeRQ37dKZXBEz0OHbhnPostTvDZxCRsnynO2mP5wWr/FNpK07Qai4miKCu0+NPtxwZp8Ztno
Z9NFavQAlwTzYaJeqRJaTPSV6pRHd4mK1j4VDvlAOWRMt9PZA27o6XN8JlXDM3qJ8fDSKx8VNLt4
sX+yNH1PKsaG7vv5M+0nf4jwHa9PXHUAUEt1mn1sjx6lbU+M03e28sDuYs1Kb6tPe4/ZjvPXIjD5
oLUCK1WBnGYEF7rVzbKjerp3ZP/HkdXSSh/knWlBo8wGQPXRa/l1kCqZgJ9bxsQMay/Ev3F81UcN
xOsx4bCQ6Ph5wURSBNecuHqaN9B/IfE7IyByERMtUgovT1ZPmrFrkybUXYRWDzRSf1H0X9LnBXBo
h92jPmZp2d0OAfOlWG2v71p/lM2M2c0uBaRHFFHqBIyvU1arXEoTcPFqDyHwCKCP7dfuAmgGXxSw
mBWlEmXmO9X7wKHGw3HYjsAoHsejv8dCR4AI6/XXxqmxJ0NoZI6Oy2eUXQlay54OW9DW97x0SUhw
0aVfIFBus9BErwquSZKv0dpFtG5LjK+JGCG4Vq3rOoYcYVxnU2PlsdQiagNvCSJIUJ7at+0vC8w0
ZTwCxwDoPt/fo9jNO/iheo75duSA7m2jjaEZdco87kcjPXakpranFarDBdOFXNd/mjCqM5pJpRC3
AOXRsa2inCzWpfErj6piS6fPxAmzoVVyjFHCLr/i2//Ra7RqeJivGNXyqzWJ1pnggMZhPJpNqxmw
VwqCBteknvSIXx2rFw/qpzIpyl1dHLfJPuwL9AVifrOqlzesY8E3xoFf7aNpD9cmJtTnJvUBmWwG
ERkrcj6/rPQ0aVhtLkxT9UJ/Mlu6S4tBRkv6LjSCBpsxL2oTrfZltQFVzL+clVN4VUYmM5ZurHCM
gCAE6BGC6ZrKKja3uLmbQIEYyOCX5UH7LOE8nEYFcCrPKHvoNVd/13jQyx1tjE6T6xKEvTU3p+45
6jPa3VbmXRahzo2CYbYo5/weqbBFk/J9qHSk0sFFZKb5oV4ZkaXr1A21VT/EaQV++lLzxHB92QoO
gorkby2gbbHqggFeMnHowXPoOhQLECPXQINV8txkd7ZAn0UUPuKUChs2m66oLEGhYuDxjbds6FVL
npXYwoz4YTCd0WAvpyHQrkcuiDs7kj0BtD1lxzSQk/KS+Q67AADkIewWaaEeS2C4WpSzMD+DLvl1
DSjTiBNJpsyDIxpTruA1Kz5t9CyAKtmnTqiQfumb0HgbA9V7wLwf/zV0ABUmA0UIKCq6oncfKPXz
oGxAtWCDdLq10jdxt1lOAg5dAysJiR4/Hqew27lpfdj35JSETu4muKUEyPu4+8TzhJYTQM8nFpEz
Nh3XiHgg+iPtdi6sJD31ScN6o1he1OgIKD7I5s8tJbLcCgabJk0dzJiUTQrIOTK39mX7Xk7NZGUD
6mZNw0VIZ6dIkEWYK82D76t4i1rJ3EUikvCdou8iFXjRstcbEzmFu4cdhh1ohp61KVykGdZMgpSo
bJWMybSsQYmN2ZQoFpeYP7BDNcUgSCic5HZm+1NN9F4pArLeoZk2rO85aOzjJyzbnp57slfaU9bb
QtczxPsPjCUVWYjFjooqTljZUe18WZBZ+uHqQ8tBJM2UrPSWiK0QD23KBf96VNg4y1LbO8uzxg8n
STgpJEtqhF9ozsC2AMSr/FT2KXa1zHzvr/hgKP8XxkcCoTE61eIIEpTjSlq8n8szdhWLqCYcB1dS
krpdV1f/uInWtw+K2GM/t4Lz1a6/DwemCW3IPITAdSVE6NvXR+G+Q31+OETaIoVmkUYo6aGLSECQ
nQ2/XHItWMeWoqcx0v4qiOaX6k3tsPNQpNNySlyGlpTq5N/P2bNnOxpsQs7j2XWYfGYiuDhfVHMG
SmJPGUEZoVY1sjwaFuoVqPJFSnJN/O2uKJef20gN4zGRRXYsrf4yUnBTKkWYjahUDOkiHVtKu9Py
sy7QgF27i5OT8CxkmrNtf/1UEZKDOpMum6tHZpBuYA2iQx1oLcFuYOOVqGkQ7yFdtrNLVzSlparG
4BqVRBJCC0hcnZjg5/MKBp3hnturwxdYnH8uTSzWN6ojW21QK5k42mh9td3y1JUzIo9/wNTDn06V
rpHvIhzNIXGz3NxywdlYKDhALGJgDMc5pnayCPR6AyYppWh3qX51V1g72RoEI1jTndCAv1A5zlUy
HW089WI6Md1a8lA7dCLUE5/kiH0LabsPyUnFdIpsSoDIEU443b1aXkoQPxclfm+rqnMPj388TwRy
4wZgfp7dgiaogcbuUj+ZtXWVb7TBW5fMfbDHx3zCX6jUXnrTSSIZ1E1/orEpCcngdChF/Ka0mxHX
FZZaRn6zt18JyHFle2hO/wD9TUAOtMZYtLwqRirb+aJbvhgAfkLUI/xrN5C9Pi6ICWw3MbCqJmL1
Jo0COGjL4G/sYHW23Y474AeG0ur3j/1662jkfSBYQxpzKFHkaNTp7zXqEQUQ183FGjDI3AKjnZYD
XVsmqburpwNvYe1bu62No5Pyo2jZGXRIUC3VyCj2t+ObWPl9XTxflAR+WnVFDGLWrSQLpq6XwL+F
vGnLdj+uNybzRy6Z1tX3Jet0jZpqVHrOGq93EYE+VQOw/hIpxzjsaV46oBJgN3sS75Q9va41DtsT
DJIZ6quzrhy464SDR41srAS1yCpjteBNIolRhP7bCqf7dAu6dOzvgC9HTRG42yA8/pQIY5WfLznJ
OHM2LHtmNzcNQWZNTkfu7R6pXExATAky183oq+LklyL3YGhGDSGASD14BA87XnzTB/UEHd4bBy6X
dVuljJ7hGYblondPZNv+FCXDj5aeEgKP0QWXB5aM8VeLJkzylrRl60+M3CJQg2Wuhu9bcvR7BUDx
P/dYXbhmjaaaiZv8zIU3dy8mbeqUL1zwYnFAvCMS3pqcfDrr8ahm9+Y9Hx9sZq1Av9MakoGwmf7T
J6hAefbHQKfVDuPpuAc16MYmBlgwtg08z49l4qJ6bcxHnnRsMW25r4XoHx2B9VaJLSdk2UpBV8Zv
kQvo9NH91l5oda4Ku3DAbk3PjOZDnWkWPwg3TnE+pM+XtYVvPKMQA3prf15ppDC77aLkYtQ7HSCL
zEakQnVlNWVn0XkUqfWa0BEuhn43TGPwmr7iSChkd0xKcdC2VfWtry7bUP4DhjuIGDTwTluYOUSX
TBrG65BSfw5g48IlA174hnXfkJn82TmOtSGWZ0kCmbDXQuAobsajFwBrrqM9DaLYx54wgSg2c7EK
etigeaAHreFAJJflh5xeR5uV6wn6vVVjC9BmAy4FKgJ0L9EqZ9XX+FWv3y0sAh1jHynSyrvor2oS
fMxQt46wT6Eybj0ii6DHn6OPbt8VaXOniqReq+JshPAEBY2lVAD4QW59C6ztEyJi28Ol6v+3QaBL
nujjFfkO5bVXZ/1vC2v5pzFh5YLT/Krz5o3DrKhRHpURu5eQTUT3dt+Kpb0agwDDMHQZS1TRukYy
uK5Vx6In/QYIfRDaxK1dej9a6qSNdmdDh1BsrUEDUEZA2E7cfMwcDxdePOWiD1DNL65pJJEq+vVd
l3E2fbW94bq556fdqQelT9dVI8mf9ma+cKVUkC4gARPtwFRKOTGzm1g3sWahXyJXpmevhr6zCTzv
r/D9qyc3O6bcsjzPZ8BheDiGSSbTcSkpfyXoHYzcurBSc9+uHnko/r2cYZLWpDYrcmYrB+set0wr
AGR9HmRXAU7ME52e246PsfLIijO344Seue5i80p87xC4puPKT4ke/6PGGInJBcqxZZizzoCmCxkR
TCiOn4DgrrhYam2yzjPhsXbCWjmga5Cqlv/ni24t3YnU8SkOplvT5HdPTc+r2A1wR5xBKdgRIgA3
6veo3H+st5gUCS4TdKGqwMVYo0dM/tLBXByPQpaG7m+mgmljbDb8Bb5NV0W6ZYBZHIdpLof3AfjG
RbjQF+2dybTY99Y6BbFhgj7u/FpvWt84dnJhiTxAwxOzT5c0OR3PJGZWs+bvJVpHPBkqxbnR1e25
6393lcZromGbrrmUraTz/sAsmtPRI+oGhRjnlr8SXhFyXoVEQ/i70QOyWwcxlsRQu4YjeOIbDMpj
G4h4eRR4oLTQSJMgRDXUvqbMAE3vpdA7aYE+ldT+ZS4CoJ7cyrcJ0braqMw+rUyV+pxfTxdstc2J
cKWcOvA4cI6GmL9Lf8ubfGETlKZaKAnZBtpZLK1mFLqUJ+aAL+tKY6P/rfm8ezUCj7Y5B8RLbcWS
SFA5bsJ9VgK/T28kANEGDWvj8fzMm4BwZyoIxgJZfDWIvAm7k7RNE/0pzpb+9+5UAv6zvTekElan
KBOnsuDeka32W2qdMuPM9bRSlWgiU3FxtOhD4Pd8Tg8q+0SAeW+7EfUGzluwg+bk4p0UJEwQNQwj
78zL6M9E7CMmeOPdZ9a3SuJKHYMQFABlQE5ftvcV1ZrvJijmCBzODItKyT/JtmaI3aUhPpvC5Zig
gHEQZGn0ZQgLrdl1ulzkhRi/tXn6c0Z77J1e1kSHK6+uA7n6jDIJgYusiVTbdV4eLZowfT4EBSzG
TDL6+BeVxAV1D/ytji4m2RVe+5GA+4OKU41s2EWJdiZBX9WCY0Rpm4T/MXSHVWTxYdvlkDboM71a
DthoTCs8L64ZXkDMTY3yFY/eXrDWzpgExGqdivbSI0BRql8VcdL9zcUoKbY/TQXSndldBGU4YNTj
f114z92wN/qkG/YDe9/rxLhn6PiOehuQbjSr8UdNEl9RI1VEcINZwnpKmgSPcL8xRJSF53UJyBIS
LnDHEbxdWWM5ee8zM+uBRDx50vOS8gboHeNz2JikJoOh/EOoko2MSelot/PfAMiWBOwjsVpa2n4l
Dfhc7LPYocfd6ls0QACHHkNkCyTNlm178r6bYJRqV35sE+pYWbdWmoc+KamwTpNT9FWcJE2qFluL
cWvi9sEnP0MOOxC7TLBuJNXjbYCR7lZtXwqp3RgfY6MbNt5EEllZmKo9jmmN7Ftql4aTGafyQ9yw
YDilgeLUIMF+BrPjSKgc4uldKgcr4L1Q5t9LUZs9L+xDOeFp5Nmu+2K01aHnIMTHJcmf4RRUM9Bg
HhrmNfMmSx0ZFdNOlOwQgUaVGTOJvuwrk+7/EyNeCBWKZozqZRvzXYerR/3rPRMlo7w/VV1FD68z
tFet61wdZ3ULWJiTvrY/wTeKiN6IosbuC++u+4HgUt5PRq1aVHfH+BhvzifxcfFec2UUdoDGDR1k
ytohISZQDkY/ZioiymT6x2avjPJJS8TCmTkewGsaewMuE2A1ye3ERvxQqmlAuskYwD+TG8dDGAVG
9aQirJ2NZFl44s7Bxu6LbY8yEBiLh2ZlSh40pE0ipruSkogIykh+pm6xaAeRJeC0jC8/uP3KC7r8
eFsVeeWabgFr5pcsTOq8MN6a1IxFx8E1GNXhhcQhiGIg0WpHZSd+5ddoMBWKQfBWqQnVnes9rdCy
ZRcdAfBprPt4/R7J+wpWOjVo8n5VKGUDE+Iv/YKqxAVXoyQvvt+TQDj46unA+AmYUZ/a9vrNZkKm
kzSdqCn1wY+hZWmEc5BEpeqwm7rVDcY4ee+8zaz1bxaDjzxdd6LGQ3JqQShSpJX2JBY/L/4z+OWG
S07vxJbwBVe9dhtYwOjMdgS2goM7CbTB8p3T6wtx7l1YIRLVtOSDBzrta2opulrk1xMJyjTZ00Pm
MtiUyhI+vLuftnT9tVESihA7sV+z6M3O7CN9f/jt/ZRJQ13/0xB5IzF6dR49niE9PoCrA1cLhu4m
Frq1wWoyMmIOgiPbwJTCazd2UfSWCl9IdPimzWRh6+yPqazqo6ZMbFpYdho3ciOUAOwX+MeMfXAR
1fnvHjeK33akZPHbe+iVQvgHyfuqZedEmq+s0oHJhfTrmm96HaO/MKGxeulhQLndKO6q581qyBHx
Gz/vHeoqXG0LbpB/0vtA2Z5oGFooohse/YfNSQ1ISRUJywphKgV8TypvTbX2qDML1UdJMQYqeHpc
0qlwaXDsLufO6IH4POof1whqGd9ob4qGHPwaIbI7ZRCm1pw129elOxMUr0RVxhGuOiFmzfIi8Xex
oHjOhC5LGq2zdSwoa73LnX1i+FT2W1ZAxuG+0O15NViKbIWdsxFasLLi2jqSouxRMJBSn5O35iBr
vAFvNw7SnK3Mg/9PFRLsy05vCFw5Wihp3DztwJIMgZV5kiYirY13MmobOI/Aubz7/kCoQ31ZOdtz
UXg/hB5dTEQY5jYH17mdW81pSCkIx/Y1QRIHnP3H5fsE1miloj8MZUeKx0T7h+NQ1QU6Cei06oCV
foeearfyg2lb60eiAlNw/Kca8RDqhpnLw1TqWWh5Qz2Ys0aK+Ag+OIzQ3TairE+icVQh+G3vWaGH
/aLOBE4WQ3RoG4h85AawZMAiAfDkapXKMLX3+/Oue3KvyXgJDCgJqNmBuxBB4216ZdLtgkOLzfOA
XBAvMHcZSZ1TsGgmpVQSyGUk+JvGHadvFalziM9TclQRfQPb5jFo1yNumDXAzu310Bthm9BxQ+lc
dY4YHGdIyc5r/Hg9WrpNdLAtiUJ0OZQqJkvon2WyPrUI2kk+HmbXqFl35YeVv51O9YzYz+fIxnNh
JhBLqHJyWbVeQyXd5GwFmMwQcwkCitt3KcKYW8FOaWqhZsOsLIn0oGKqRot4jQgXyuw4an7kpPEY
vE16uwGq9970/QBVHrtC7VuLkN4bP1WlKHaRew7p0p7YX/gxO8H/mRocOT6Phsr1Hrt3I5hMhfJS
ZWygsX0/ywbiNgI9GRd4r1+oDobyRfV1Cgs+VQs2/KTcbsx0OcAcQogRdInpR/qiqXulEkKKZB+K
0hTOcpjJVBw/ewK8YCziqXCGWeg1FiPwZf3s2xzzaNN5iyi7pou3gyzFdfuaI1D5JLnx6TRbuUVB
AfeyTXOhOMjnZciVjBvLIvdRj7c1ltAI1TC5OHommHB/6BDJpCwvgsxkimrXYwGNRfDYa5LbOX0h
5aQ2YdGVkE14K38f6oepX+8OPDtV12xqgaY3f+k1IOp/yMT7hjP9ji1yiJ8nM53UBp+nOH+owuql
h3MtP6wdfe3rjm26bx2zhLvyIDmElx9RDi3mpV4HavchL+kBAQvltHUTBWShEUepGuyGpQbCo0JE
klA8T9HzHFQFexujY+AtvEJct/BQVJ6l+I1HItBvG/Fns3e6D+m1fW1l65Pr+vd2NpEuyNbTb3Ub
aev6Z2q5fJBmQQge9PXqM4yCMiWOvxx+j94c2ZHAOgzCICs/pzLsedLwQXvgvi8fYegmQdPRCmkh
j0/UU5JbLQ5Jgap21NEA8/vRDZemXz/8rfw1Gv1nTnVWY54nbt5zNLmd6reAqsXBDtTAntyVj1SD
QmGvxCDUS3Bv5K/Vz96peSN/dfsId5crI+5fZoHY0NRQnRFrodpxHZdiGYrpBqncEYQ2S5BhQI+Z
nJY0iMFeVD2qbxax9z7pRff+RsGIhMYQe/RHGnICWi+PqLdMP8r/y/0+cyh62uP7NcWNXnS5lM+5
6H328RHWmXiXvL9Z7SS0zyAnvFQTJNlv0yW3fpY9pzi1qb8nRlJF5Uwn9ehE956inlGF+SGQ2bHt
1Y8iVZr0Kt5/ad2QgGXCgPggAj2MDwXkVpX02disCSbohdQwniVYY8lCuPivo6+5gdgq/ponZ+Cb
NNeS232AS/7oJs9VQSiRV/95kR7+V6FfmA1nWI9MikEmKAWAOEOrjM18eEkqv3M8h4LTytspWRqW
k4kCW+W7bEW/RxK5WztofX8RfUMB5HyHDhwlfcuLl7rFpD/2n6/SccV6a0Tl9mSlQp0LQ4Gdbikl
swnsNjs+hACLOxkOu+wgi9eXZDtLOd/NQC68coRoiUJPJm8TnjGD4Sf/RbExDFaTHVrHtMNeQtHS
slGYZ18wWcA/eiIYUtaV3jCq9F0wQMYt9TFCPlUmliSVAw5JakmmgjoQprC4AZFP71ZS9BFP3i3D
g2+Sg1IJ4iKOXcvJcZ+sPJWPO8MvsUwOm67C5ro3TCxJs5fjieJJXblteQXLWaOOie7KuNYrBQ2+
zqcflkxb/cqIhNCqeUmOpVI3XLUtPjb+bTyWcFjeQWqdST/FMOQGFPCLA+vexFW6UBuM5Mv489vI
YV9lb6tk0qkyYUjwecFy/6Pl97hKVXJdx3txp+Buin187LlEautU7bxnDWSrZj+wbQ14xecZlmm0
p4jGJI7UbWRcPmgkBGJBE09Zw1tkIg/OIERp5VMUqOWF+Jl7+DlZVTefpxTiD8kEIInxOiv214sx
UL+SVxF7xI+4ajwYpn2CNHwEFAlAE9lLJoUmhzWH/YQ+TajYOgZaUjCqQ47ABbUq8oTSKYnZCVtC
Wf9rBFp3Zg0xbsxbM4EMBtgYjGXrHZZaUvLdqpE+xAityk4gbAUnRwfNKe+VmIF1fi02112b6xgb
ZWl0e8fibea0uPqVEguhUUhzh4MW/RrpdMj+WZdInk96CHbtkNG8UnsfC7ygS/aMFu0ASYDU/e73
cRtm7yNKs58OUWYiZ9CwyBW6Exi0htm6gIEtmjoPDe0TfwIyJqwwqoCHtJZaaj+CPhZ436DrA4tD
FiNRQuFZk4YseM3n6cYifHxTtwdewkojfhPVNsFUwP5ueTr+HPZPoYti7keGkVySdmn3vayviNj/
LVS8oH+lsrTlVDQY9ooF15E/y5wfQLu4NT/VptpASStpWGjtw84MnDQQVVAN3Hcai2JCmRI4ZZIM
sqOKgIXNmKrqQgUeARkeEv5wxdhJt/s6+cyPzFTlLlN9SwqzikML3g3e8PP3JUES3M2GqsAg7sN6
g4ufYn8VbvnCUrH6Qx1thsYPYEYVU5SKl6gVDfeRuebAmSG4i7TLQ4EuxFTEzBsAf86/uz2sJiS9
BPBr8xvivnsO2iMt1z+ZPE+8mKsLkyFeCAcVsXBUaEVrmlX+wYEwFSpjkPNMqdOgpwXDVXtSAIcx
ZFXh280i8p7n9YeHmCwl+fGL9LJxM8c4uAHrYFQyeCPX/WsNyMKo5cuebERtJfuiL2QsHRD0Bhfp
bvXIvOFnKGxlIq3M6x6m/DZlUBSYVQbD+W3ivLClKZ/QugMgNoExIJzVvwk4CwiPDs7+ADSFh5Rh
/5GDFklmm+cHzOdFjV1gAB9IGive5miAwf2KDmV8fkKw77lgWfh7BXtRp50/LKnR4DqynW/faNf6
dBK7jbFnqECPGVqUNDSOTLP5Kh3EbdTBBxFzvHnEraCM4zxU6ceecalL8dYm6bvQFW3ENXnBPfKC
+/b16RlQcGlwkuBCr41wdPMv9zHMlqR6vVOiUFvrfSmq9DRBCU+rbzRnNBSm83lv8z/OriYKRns/
lAs7q+yYhcmTPMfbU77eJecD8HHwAAPnyIJFvXkS1Pk+0M66eyGzoFz/2p2UybPYe4I6Yhs7KljW
4VSd66l5j5nSEUpG0ROpIs9T8hQPGZyHsbBq6bwgMx21OVZiGrZUB61PGW9dMJ8ayGf09efAPQla
jWv6jcJn0rXavt0kpCbLa2zpMw0l42GjU0hn35UQYmuqurUtc4pkDTFcKQ+0l8EyzyOlSgEhz3lG
9S1kYnuYqv7g80EArPg2hTra/iyZAXrmRSgQsCIin9BIBuyB5yuMf/8LeX9qThpHiHtkhtPNsuO6
wlSZddEZFwmYXSSsf3eTyBWrxIC90YLeveQy13ENS0et80PYtape1skK14vXICwNlULZ40SXW4dz
tCer/TIz3t4Nlz5xIr7tUffyb+LK0EMb7TdFPJhgg+Fh9LmORieZ2g8IkhVZE5+1gGIYLeZe0KJu
RDPANzGdhr9w/HLENqtXAgiU7HIAeZEVZ9okOrOHeTdOE+T1mjsV7prXPPG/I+2ObFTr61s2BIpT
T6buoLRNETP1+gonngQtgTxVr0LaeDB+0bg+GUZF2vlVEH8EPyVSCV1P3EWVdWUfRPmdbY8GiK3w
CGsU+iA0vDqQ/j0azoknz2hti1ZZcY0ts/KOw0I+iDn/MWki9jkDExu2KzA/jUPstwrECmpJXuCx
F6oj0sCw6r++KRXDf+/GuIGWRsGhTgkefO3hqAGYSYbh0nJ1SCBF/aWKiCfc9cX3Az2zAoaGWiSv
Ij341obDVXu8Sei0U7LEZvbFtagRh8B0SHus+d5pClLJ4eFJbBfGNiuDIGuJyXcXRq9k6yqkLjbs
2nM2J6tfEKkC6FGumBAT8HaJAkx1Nkkxk7r8GdI4bGSjhG41IjW63g+lc43z8ocOFyBzHE/SmBN4
JygPdE2jDnZBytX+AZxGaEuhliuOCPCRZoI+Pw6YlIKea4aA5wFJqNiiTBHQVdH59VS6uN+jWst6
2E8Y57z/8IbsNYcYQaQ3ewpu+244ttBKZhnjO9P65sE+CsmH7bpQfgWpPdU09KWR0Ye0r53Tvhuq
6d9vXGkf57FNc5Ot5MKcmyiJ3hjHLUIgaRuKvDyflau4auUspL9swXhXAkmOcoo9T1/yzf/LJenX
O2Mf/qesFKL8rEUEeCRKsrrrR1oc+jHq3WkG+OftdvgwixkZ5+fIwNeVXDqrSQroDxCEIvBvbjmX
S0s/Wd2DNuGjdTnzQuAa0pjQ+AOxi9Bll7UeuOXCM0D0vFVVBTQEtENd8p9Y7US2oPYUBsHsNJnG
YtF8P3CDUA2YdEV8ROKS/7vuJvESIvdKp9zqMUOc68nrmuaYq5/8x5a64u9Ui3RuWbNaTrTx6eny
vWCvU98oVYuuHiYA5xy/gW3FtId3+oCpdoTG0bdvab7V9W2aNIDVzma7o8K/DPLnpybi+tblAwnh
JCkH7hAAZU+SQ8p5KIiroSfwvwoNwt6QvYILDeQcFBFvyWqEHbVQ4B01+DhSJ6/2ENNcGCN0BeHZ
pUDmv8p1mQGce8++ZvwfCCXx7RCW6zM4t9NM2YKufFCtJajhpEVBimxIxwTpQGoiD7KKCqn9Earc
3gbUZy1A49SPZi8cVXX6dP9S2nEmSjX0jc9i+5ro0eE9ZbmZPw9gf3ZdQyaSxEg+foTh58G5aGe4
hZ1Xvh/1XEDPvKN2E44BYef/T04YmLr4XKyD5lZ2calrsXCBlX1+6Wyvr5qWAk2gAv1JEXpmRuTI
lXyXnmZimyOsoEJDjExOm8ouUqFbjSUJYtCKy1OdQPm2Ae1l4isO/GPElz2woZ5aQuQdFrYMFMWk
AZfTf4cverXCWeWYrG/yC3DJME3n/Hom8N5aIDTXYIw6TsLCYuWjOASHlfRHdEH2S9UR2dzI80jo
Daga/2y1Wy+Z88CECaybjYo09EFU+8+CxkRc2wik0McZRziK6IZVw0YlZbKz1+KJFQwZSI1/3LB3
N3NvkBcf95aPKovOeiR7qGPiEYMYoxUhc2jhW/+AOomqiH4tqoeNZ8d/635WqBNyEJkKLQ/UnUvT
6fSwU3TbOymWQTmnurpGrZ/MXZgk/+pVd9tLk3zHbM0LDe06aX4iVZfoTQFEAjQRrkHE9tNpEDs7
x2+LIudWTshb7o4xoYunrLbVfegEQauyendIVcpfjK1hb1bdhhqwjz4+l7gI4OB/r7WQrxhRc3cX
H0V+GjcU6Jdkn+cs19c10UlfgA+ZI3f+6BXxEUwTS/ofZZGjGUgeB8VO9OY8aSnhwbkEQidHFhjL
51pStp8KW5X2fIDZvy4Fo9f1J255ZY3f8ojnn0xjYkr0pEmitHrJ5LYe6p/YR+V5GGZ7kW5GFyy3
ll8t7czzZGC1vgk1A47JJ2D+HbBltOTGb4X+B4kY8ChhXbPtJDJTyXOeO07doFCHgE30zoy77P7P
esTWxycDluELGuGV4VBPrYNllqfhbb8mmfdMzAkV6XoQMPAXEU+7GefCc2aPKGoa6PC+XsCj0ymk
Wx5cjKLyDG1GYAiwhX/RnKM60gK7BaDPIxHgoAhZ2tZUH97PfXo83+xZ5KgBhqCTd5GreRCaQBtt
0mbJaVZYYBX61s7RW5r0ZywZnvUb0ZE2HjNUNIce53afu0ltQ9UjiwTItJixo0c71mJEjRxEbPDn
wM/yaCgOZS8zOhM6eRq9wtX794PM/zGqnXOyvj0+BF4yWy2RcR8cMNBPlSthAezXpK8lzGBtRYIN
mHoug7UTjlVrFHz2UlPrc0G0Yf14MIiiuCkY89uFab6L152i6u7ZWPaWXRBiQybInSGXsVERr4eZ
o2MgZaa9MrygHgEiTwIMXy4WFr5po1QgUHecca6sMIdnRSHZWwTBl/LEvlG1KmhZ6guawxjiYqvz
UxUH8D7G9NwhVo7P0zGtmwI6ODUhXhI4XSz2Q8aoM6YGkegW1lOH2MV+RrWf7tIpDBVamyRWbXnY
ChEpfW1okq5AP1nv2c7RlxhXc2WWSkJJVa/HhdrCTKg7m0RZt/hjkD6/Dsp29/U66I3fTJTqBWcz
WDjXQU+wDgmFEkj+iSdxmlkUWoHAqBp7CyPP38WyVlhMyO6PSESVm53+InlxpRV3wsp8WbU44GEc
k3bUbPNwM4tKg0/tJNHJN+OwVXHVJXBbVLnjVb+4QDtMylpUWNhz23DXugwEcqVw9y8vEQ5I2YD4
874JqkAqRmhmG/rmclwBTiIA4Vwk1hvidp+2LachkhsgW5x3/WQdE/Bpd/qQvqX18XT1iNa1Za/Q
nLGeCzRjiyxvRTQ1Y8uux39Puh8HHepPnT74tQrRUwsjB1FLlbVfQ9MQ/IWs1O8SbCgmMKxAVgrB
JWM8iiVLBQdmCiqjWq695GFwwJpL+ktBWH3qNUlzV5yUlp76TxzBHTq2XGff+dxvOonrPE4lAZDS
grcyhK4Q2WvkfmSHd54DZA1jDiH9My6W865cZcqopIeW7R6WH1bUpjG/ZEBUBr/OT+bEQuUCUxxd
SZSaUuErwZCOH0mQHegcWs2z9jaYVVcBXUtLDlTcDE05NUdiZ3REk+LhpOPrb69g8yIiemmN0D87
JBkotUhSX1T+wUqNuBDdY/CWitBEXsLDYxiqb/9zKq57tjnfmh5sToiTw26B7zaKPrHw3bI37zLG
U5TBygjm+HGUPQurWPt7B9HUvyC3bS937UfzeVqHO5LsIIal5Iv7yKqylwAqzLXUYekux17yQtcx
gHyolhAv72ZFngKxBz9KwZ12i6O7wHKWdkb3Y8BYk5TvWCCrRifIwO1D+ybAK7lyzLA5Q/9XSuKW
KjTnXvkCfuj7lZe2GmgLyQZqqhhBsv6iVCCoyxfLn1IY6X+BwF0BqbOnKktMX9MLVjJcBpe/Fsvv
keMYsosLSJ/+C6CI5nJYvJl/WtDIrYeLugMAg2BK1je3MnD2zHtPJnc/h8NQTBUBh0DES3rWT6OK
HdKExEjMDtFgjnM5H1pmRLj8pnPM/LsxNEK7bKz+zFxg1NmH0EIJvmfuueeOvHgQy/SsGY0He9AV
l/KPT5Pkl3Sg4sDylDhijxG6HfdFdeCLDZQ2v/SmbC9Q3q1N6dcuKBKaOhHLL+p6y/ywBBIKz600
oZKtNXIy+de5pXa6w9v5Lue3n4g1hWzfTqnWXnVOJvfcVw5sjlEs35/Yev2ui55UFznlV0OPXgKI
mYkgDjawn6VgHXOI5Ou+q5/Ryphi5+l51nuk6DISKPfnvAjRlWHYO8zfO5lOyYdQ3B43QiFyi7Ey
PGUlr2oinz56mPl9yRoxBb8H8C/u4HeYTZOz3STkoTRn69sd5/GlVttQRqzz1EoNG1Z9cFuNuKpd
oM6WuC1bmvgtJRKMG/pn6wPzvljpsYOXsqaV11vFJMrPl0YN6vw/QGd/8OHxQ0BbQWaQsApdYaGv
QriT45C0IrFuvJNVnNToDhBC5wPN/BmGpASVWyBYgmLi3K8VMBQZmj2pJWf8lWcnymYDgf3LhT72
KQC2kNDkq9EmF4Gpf75mGZ5RpnT+E2h7Dk/LlgRXihRxbrA3NVDFPMgQJ0KtAVaKYUDsB71kAmrq
WcZKsMn9jZzh2dGzSZGYCA19ApC3I92eIURwcNtnCAb/frR8N1JmeNYahfzZljPIRzTzmpbmckjY
MYZYZAckkqI3EQ/YlZsMzvgQLUjAcNQHjQu7nnQt/q3kwdv4tcPxW9Ndi+w07bImJiJjMsAF5JWw
qolpVZNtn+y+3SQvZlYvUZ1Gp00/t3q8/BQiSeMZqOnaO0xeoK9Je+N0VEKuvK8RvMaaYuY/KQXG
CdDOfNtncLnVoMmCus4hHBQW8R7N+dZkXAMYPUN92jlPzE+nbnQO7KWOQmYt1w6LeDyxnzzAd4nF
pTWerdefOmrs6o/YVlA3bC3EKBbzvL3XAzc+znI9l+7lm0oF7v9+rtXsYoFYKtpRT9NmQjNs5aJt
WfUO2+osKJxTbBKnZxnyTzUitcehRaS6I7yueri72czALogx7tXlpB9wa3VKwBN5kvkt9hmknbOy
IuQZn/Tb3z+W/gZlyctJfu7ENomc0UdhApPgwOMzl6eyvnDiSt8z7xz/96fa5uE9BiYGn5mgUqB6
howUjXAMGwIZSbr9FRwE+tLs39xLb9by3npGQ3wZiEcJ/pvntfD7yZ9/S5+xF1HTPouLmnWCnoW0
GnENEkzw2uwRNqVdWobGFz9ka/dWF4LepMRby3IsAmlaiABLUVexi8ax9Y5SxtbzjTNrDXo75wwt
BNmHGFRnT4c1cUHBp1TlkudBRR5N+1GF9NX+sAlywWD+Z3t9vWWMKw/bnB89lzlUqa/Uc1cx2K7T
ce68h8d/kR3sOdUy3qw0JLNQi7mCrj6aJvI8N1R1+7wWmYtKWBIEyJ9VXF9jiurS5EdZji/9zqhY
2EvSiTPVom2bIMJgTWS6SxciRzERAmAxflhRiHXgAU5IhivjEkEWnqBxlWkUQjIC4TcRxG5mjI36
qda697Xp/t/j0IMoJUXfZoS9MSAgoK7JwsAsYr1+emHaUPULSQUW2OSuN195Fsh516NCOqqoR4A6
W2g/Sm80eyegHSk/+6UiuX717YFuGdI07f4i6dWHgqcN0ALL6nRxQ6cN815MZ10q59TgvQQlUBH1
HDc1uouMd8QVkCodcG+sf0panjfcMwxX+P4EFpPz0lp0cZyW79Dp9vugD7DYVwYCnExquLtAiJkQ
3sopUDcC33TIswXc9TohTrEFrj6BS3SKDEPHw6wep27dpS29M+oIf/yfSLB+D9uj3+zQgfaBk9Th
bBLku0+Fc5e0KC9jg8xsNjRhbeNxpfPccDu7fCvGgM8s7gW3PKJlvyI17/+V4dX9AFFcLVI93950
L6fq/vE+n5AOdSSPWhKDlM1Wm5WlTtUzp9LMmnZXK9XYCRUSl7U/2wzx456NQAgm1vmtqZYhPQno
OA2nh+38ou4hjOCi/QkgVqyxcfO/vgAkPo+1eGLBoJ3EEYV20UMsTAs7UhPPAvEMtKSvimZGk73M
RQVCPD7Zf6on51yNvYPEzGZVdyQkBzN6TlsnU0bugyhnZC3SNDUjZFaHz+43fIZUa5REOp0xfQwc
vxL2AUgFGRB5F81F034Slt8PEnw9hAp41jKB/qq0n6/wHA4wkShSpYT3nWWYc2AwuVNZYYLrsSnL
bCR1z1F0aYvxyIBICKqtGBDkIKn89uXDQTG5Q8bk669A1rjyY5OPSLnS7qUIChHvOuu/oNtgjZPA
oBTgrbGb48JPnASGu2kuUuUvhz1kQ5bkgVvC/zqCJk367nc3vNoELD07uLPQ07rlMQFHK7T+o7et
XIoUu9EEkTUQdc1qcmzdhoD32kAN0+B7n/+6rWBK/My9VPda052a2Oeh5gFDUQt+iptZzfSLx/nq
huX/QT/1ifkTazm87WfpeQ4usf22Gsf+RyykaVOBgcG02R7wHXT88pkzcKemdtwkhmhu0lRECAFN
h17L6omgLo+OHgBNk3mL68gJrHNEtAXI9THYGT+v3r9ZpV2KwxMUxbVz78X5spxj2JhCLLQdrJBt
OddkA+yb953lVtvAYy8td0q/W0B6p50ZGklLxuXN9TQdFLoFD0Yt9oy75tzOh8zO+JVqxKGlAjTs
jJ9Awb97qL2u8LfDMXyt0OQb9jtySwWxJVYgZHkIfg6GRglAN2dnla1LhYjm05QljVvQLpPogVaR
GE1yfIO4LBdBi/GjGPqQgOaJvvM35ooe/ovA6J78eQ5aow8p7EVn+5dT0h3ZlrENxLq8nYI+tWEB
tTbc3rBpdymuSvaZaW1nOa5lJLvGDOHGIrz3jysZQXI3UxC32RYbIlZVFI4F9nGRV6Ylg0y8bJoG
I8/1aBqHDxiXT7NGD7fngkBl/CA1JNXYboURYN9/fe4qwDyU2vIeoItinlPCKCNmXD3bihHkcT2F
LqHPGP70gBFhPz0jsMRGy9n4AaHDNKD9S9Rd+dt4nXbUVikv3yIWfxg0/lmvfLggxAahib8A7Zlz
gUaos+P8p8RrbI5x8a1PIYcu/SXPqzXBv1bDa0OFw3lFDe8KZ9l3UgOjg3dyDBXTRQbMvsQ6hg40
HhEhE7R3nGZca7iJYWGmRXS97a7rfkkyyZFXL50ACvc83MzsYi01i2oDj48YlcAutmDzTe2+31rQ
LMwW45kYEWbJxWU9XJovI0KkdSwS/SogsfI/+nL5p5HsYhkDWHQI4898Fa3KrFfKtjeTHQU0/GAW
qQLgE1kp9KLp3j/jayLCAtOGBby7O7wM7j+dWz92MUwVBDBubfa6fqqHpd1vgL79iKGPtpWu4Unn
hILfs+cukG1XMgWQm88dkWiu8TLAO9LxvaEUfyaq35VjwZGOyGSbBl65hk0715bttLVVZlfXEp6p
tR28qFq3qMGzVewhaWdOdAA3vNPsVscT167h7Q86yWvvutIqJJYXrL90WK+rIpQn9mkI2O3N4PUt
u3KM1xJyfR1CCd8HdZwZPiWoU5xIP0p8ZsvcnWELeofDTaHUwSBOI/ydtkABVllV/cIwHa+uz1ih
lB/p/rKBTGOanWUuoZZblLlOpq1ktZNs6spRHnp5PJk9EOQ54wc70zGDTZZRGxQfeQFjo5osZSPb
IRFXQLNEK67RjJaN6BWOv5PD8p94jS+ypmmj39y6DSsTyg5iUHGikH5bgAIUWbcYh+lZmYkNnBsB
jgHoBd838EEc1JxEFVl6yFXnIQkCvK3swKoXfleZFXo8bUT4KruiyU2HH//8P7VJQEHgquwd9xQX
h+993En0WTEyPQ9gSgFsvCpmyjDvhjZDa64Fq19M2/1RsDCaFoSLY4VZYjDBl3N9ZPQQ3rRCvvW2
dcwXXh9rwFBZaB+ExOfkedMXbD9wpg/zQ88ziBIHlnZSILJETRh9s2VJ1IQwAgJpAZozFw1mWalV
WEAgsYXYYiNEIgDcMGw4K4VKclFj8t2UFJDXXfx2amvOtJ0meelr1dMU5Po067Dx8X1Zq6tiGeu3
noUxKhNfCseNRcZ8A25Pj2Z9KlUdkt6h6i4+BO/ES9paPnu+AHVW565gcvW/Ys7rLghKteyZKdc6
jN57wSZHguvHBEtQFj97F1dcqve9YtXQOKOZsWmyCCv4qtgvqhIG1yp+tdpBcM5wxPAlaGtnT93h
a6SwwCywr7OZ4Qr4qNmZ/mZ/7+crLOPxyXMKrDo1yfIRHu1hZsY5s07EQNoXtvuCwB7jxa1/SLg6
87MSQoABcbnN2qQoi75q7qppxcVFtdB66T8NoBEZOLXcqKfI5T76HCqWQuq+NHTa4KosGdrsgi4Y
LBwDJUQ22Y2RP99xEt0xtH8AK0GdPti1iCsYbhIL0cQ52L287t7Hl5uah5zDtgVVcWCdKyP1ovcj
GtX77udQPkwsUSpCs6t2wo2OGLMTTcsAKRYofZkOescWZnmj4jNXDQond3kKgg3t8DsjAmBs6hqB
pr/WuQJlA0JrqhRgyy2dB5E7NnQwThAaeph6qy4YYpIlqFtsgSmCGWZqjGMxzZM+GrpDkJXh10of
qd/BUVh5nPMv5hZEd0AUBOJXHJFX9rCFUnksKds2nyGcgZtZ6Q62IUrVCr4pUvkcE9zzocNur/gm
upgwOy+1PwzM03TGarerxY+qASiyVyxVx4DbU2IsXIVMqlRLrgalt03pu6o9Bx9GvSkzABGONtnu
BLrpauhA8HbOFZEbF1b0SYz6b1J1jbKYiWeigc+ptiE45fUbZGC0hpASA8in4LA/Gu4xQ5dQYfPo
XBhdYaS4ZVVCBDlFeSmJweLBaLYWwgFsVjZiPpEzzUAzuWY4XXQrHuLBWiE2/m9VVxMiqe/1IEYj
3Az/s26zCYFOU28pcqJdZODnMARUygdYkV95mrZnTS8tEzCIr5aPnn3vZljr8Wv/SHTU9vV8LPpC
iWltlZJMEosefcJUYKi3Yc/JQ2BbLaD9F1MGMxzJ47nlpr8XrwSHutJwKOrFQ4e66KP0zy/22ZiU
yd0DxDGkg4Hmwr0+gpmfbkw/1aaK+iwEgwn1tI0IssVmsUer/8QtxNY504t/oXHGE63tEFKyqKp+
te5MWwVELrj0edQaImViC9ICLTBYkJTj8E2+/3gxIUV5sUD9H0bKkp0MZWL2J+iz3LapNcJ6ngYk
kqnf+tblYl81LhC9ITMEItBLxlVpJIb/pbRlDacE+t9Sysfgw4Z1zIvGr4Usbf+FLE38BQZlBNlJ
EvJZPZvy5oozsUGP/qcqP8QpaWuo54UmBL9U8BTwHuJ5fVsxdW3/IRxOosK8VphUAvI20HoH9Qt5
Y+lemi8ZN2hDUk7nbRNSbyFh66qvlbNlGKLE2jnh83Lnxz61/c4O6SzV0YTiHn2EFcW0AdemGXuy
Ao74z83+B8BWVbPE7HWh3YKMn5AjeEk5H8OA6GaJFJCma828KLOFZkTRp0tXt+mb5l2i+QRQgJPW
OXDuM10nWdSKQaJedQqzzuTxP50WJaJm47t5f1yRiivLPHIZNCxw+ZBadMtKhPmPzsK2mdp2IMMx
coZORnCjD+NgNLfCRSQC32fAdK5tqf/3daKzZ6aDLkQBy5g+x9/dIgBz62+TA/QSO/kwedpX7hto
ofUjmZnwXgenefN6wZucTewwqg0X1rPrMCmOOA0sWksz/mFCRBSZdzaNUkOQL/8ThIfdZtofRZy7
rjd0iJ5Mpz5xulVvT8N2t22LR3Br4IN1lmdV4Hhr9QNZqCJ0WGDPV9SjU0ngwBzChedPjuiU2PXA
qYo2HL3Fsd8l55Wo3xRztDpBE5Bo4249/awLxIgkX+L7AlGp4IY93vC5AuQoI0Rp99a1OA5eGw5Y
IDchrVjwNKtt7mgwXcL4T5XkuQnLTnOQsI940116MkSiLN9VIAcErZQUpm1nkzelZtm7ISe5URXj
GnRqkcCwIyIcUNK5SY4W+F9rLS5t5hRKb/HZn3R/TYLm6wLgdr/EQxT98ojJ5xF41bQve7UTpt5S
U9BJs/slFEgbrSZsX1tFPACFGaZdl3/zfDEvtnKfZKnMoAR+mM/jK+1b7YjjW8ee32M8to0xC3Dh
JGLTN7sicgE5oK3SC4V7PMMfOOgJR6c9ETa/w3gdodGsBfWzm5YNs6XO1TqEaVuvKgOEokKXo3sd
AnGawdPKqnd3rFwThHUKhCQ6BIcvM0LWJ+Iv2tsQRZZAjGFs2OECINM5wk8e+FRB3Sb084USOiQo
qsTZVKKNdOeSG6h13VHCkG1PT+b5R3YvpcLKK4bku+6+ULKkXUWpFjrHVqORCTQ2LZHme9JltGzK
DjuSikrqWjsO1e+gtjFQ0rPmCuSDibHW3xyI4yp+dVRj/Vk3TnasDlAEWQI4zK0djaVBjue4uYG8
G4buhIVc/MT5LCyYyFlvsKzMVuI8uGUyBlIIOt72pROOfXoHCtKy18lJlDmVZKwfqgERYyrsx95j
CYNH5nNC4Ak/RdckHkuRaGyOs6TyyNqILCfxUZ9iPOJHH/iLvWbpk0xYVgjT6PI/rL+sOT86obC5
U+BYaUMX3Vd82cyQI5W/zR9wZuTYI1CPWVPdLdTCe2EmeKWdQRFVugnggGS+uBf2gOYXiyzYvKrl
nthvs6WW4m/VvWkzEjr/Aq5lMJCZg55ltMXDrjEbCfaN+dKbdUj1WEKc5nqQdKQGBaF8frF4uIah
qmKOgqoF5RJWl+HuVCnUscwbCQrZSaAzrtFhZzWz0kZZMihNG0OHIZgPt+vXE60CBxPCKKzPSWSm
n4b7zPK2ipm904+bvqwxgId3SBQzcrQfXcTi/u9xZJD4kWytuSwxFPQvDsOtIUivr6hVHkrtHJ/w
W9t/w0+/rucXU6RjqjfLkftFFWfF+YqndtBT6pSNDTocW96+zHCfm+NKhzdw2co7gUWJ6l2VU6w4
r4+q0DxMWynS56pW07GJX/9lY8BT4QUMWvFPkcrVC9OKCHQFLqV5Kk55TTsAblbo0qS+innyv+hn
y4xZo4oSAD+xyfjza1FwJPsQlwhkuEL5ZgZ93erHKtsSwvoF49A+HDtA6b+LkqrwOhFCFS5IDzc6
5QXlswfrAK4nigJEwlWsQVzLhvo0sFbqdM+a549cfP4kU84qUaIWGkeSuf0nQS9JG+UYryB2kxCN
kTzw9Pg5EOxvv6wfAFzGCe7ATLL0ds+uKBKI28Cpf2aPHr6uNMhiekXQ3gBFlHZhg4Vl/j92//Bv
/rYNeTN9706KdqMPscB9Z6MUlduo17T1s5oqqUusmnMprrXtMmYCGk40JVmtujMg6v36mm+wajwC
jggYTOyySculmd0oE5SU+BBUcOhODmy0pmj0gkWLBgSYQZBZztPuSJMaQeBf6L7os+g+jjKHBb6d
p/+Ev/e6kpm2KbYnDKjfq5A3bujbUfUR9/aoeeYLfj9tYuCkdTmov4oL2FG4r89qITbTqWvUM2YB
3NnKb5DmVwt1NzOazYCJA8XjwOjQLrbbUAX9uSQL40hEo9Oiw7FAo4xjU1Td58TXBMeOuT/HEljn
/O6jb7DVfh8MZbxiD4hJXi+rFKj71AgrX89kVA5OzWPCqdIwT5Vx8bIJY6Ek+zX8+h8vqrNpUPjp
b2ku/+rpTs7cxNdyLGXHBvKhD2tHr746XJztIbGh9qlcPU9YU9Hww91utdaYHVGkDu25YQFzYBR8
dYBtsTLyK9dQSAT5QXBh8TG3gBcnOFPLjPD4u4M60+2/MAXlpqKrkfAJ+jpJkfJL4YH0fLt+zP1/
gP2qtd0CiqTf470jw7TlERfyW4fuKH1k4zj/L96XpakOyx7wJZ6Hg4jUdGEFV4R+FEN0tAUwWhJp
s9+VvzDzVabh+TPrwKIR9+/JPmRRhd1mbc0h6r1A0Qbm1tkgpgeWHBiwOB/YifGsedstyKuTRuzN
ZJIbaJ524Iy0PCrHUL/FEtkI1NUfj/jdAKPJ9o9hQul1pOsgQSxubutl/3nnCLw2BtxFs2+RgZnt
bW/JEV8gd+Tj9bsoBDehhyFAUBrUjS1/p0yYFxejbt1hjVlivlGx3sMDOfq6tZIn2OgK7/aSSGbx
jbI7LgDWa3lE0I48KppLXNWJYTGclcPzchFRj3Ew2+rjGIya/mHr4GOK07GE3zvZUSI2WEOSlSIH
wIndAT17x2PlcpbJQm9VkOFU8SE8n6YceTfmhjdWiyV/OcWVrOkJkJFahPbVNZtzi28FiP4sxucz
a5Qof6E5JPEs70VGpkwyb6Nvn0TlqwE9lFZPxM1SFiYgoDvs37MycopNPbuzt6kwTE8jzbX6SBFB
I23EI42srozw6lm7x8VsSjUQ/ZycmLBNGZAonJvbnPivCXiT5IdzNmFWCdl08sn/0zvAar9iaN/x
ZdWBmm6huvr+PKHpPXpRXgQiuA0hzKG4dTfFvqmoJa0XErw+6tymSRPc1eerbNPNZ/ey7dQVUJ3f
nlo+DTYJLqfeR+M+u5SU9CDS7js0n0zAxuDWCUnDZ8KyLimPEydNIYubzNg7MGH31vnbRWPTHErz
lJVrAlWCttgAbUwAg+HWi5pyoGYJbtck8Qg6zzh0CRemEV2C7R5lkbcRX4c06wNkcRiCp3yv2Vek
W9b+/p54UmW16xAu0+BRPg52NKMSUpLk5MjadBRalC3pgl3cjSU6pwVRXsg7Bu6EU2tNxGRrNvva
55wyIvOV95yVBHzOqa/YtHWgH5Na6Uzg2/341Y1/vktiJPN6US4jRpX20V+VC/Cko7MViJs8lmPn
t5YdQIqSddLRG8kKnZlL/PX+bHBkANorhHe2GQx48x/fakPSMF3FFr8nwNlM3VYwD+h79M75wq5u
tSypjlDaXxhexbbmCSyu8wx6o9jPSsqIh4eCqSS9Kws2BgiSaVMKZK914swZ2FNvjwGo7QLhWm3u
htcYI3XNxcXdaxqAH30ou58i+tNcjVzkZ4exFQL48mgEnhKAwnewM0fn1VGi+ywFSSGNKFOunNOw
oxyjqM6kF2+llgxPNEXFTXO2UenXRhD0sWx3YP62+9NO2+DYXk/YQ7jCYlXyD4OTrd0lUE8eDS7P
nPUuSp39bgZLhpjh2B9Pk6jIrIRkZhPBRueC1zmtSp7yqjr2YrUOOtU5q4kOS7X16xnZzrKPk+Rp
LyDdEraAc6nL6yrSgbZ3J2LlZWM+m1ODR2UmRqgyrhdOLJ06N5WorGvZECmCge/KoynVSGCC5kSY
IcRFo1NdNmLqpSbsMim1YhCO/HQZzvH/+ity6rfoAE55BnreQn2yR0WMIrrqqFpuOUh6TaINr8/b
wCjL4U/Y5gQxFVO4rSNXbrQ9RR53I4PjsG+7WAgXNuL8/KOK3bb185uXSjco4x9ooO2qfnOs+0bX
YcOFLmQjAHlOdPLS510FVD8VkA39XWdDYAiKm2oiY3DsAUr+cFgu3qRKlrQDYtHCcNJHVIwGIOfS
3MF4jLgCeBKq0tDjjiDvkejSWwvTzQ2hUhFeu1k6x64tGmqShIHxNG14m13e64j7LEmLZpIxoFzS
LmiqpEyh4tQoLefCOsAue3xHLFLT2D2uXAToJ3ITYQORSMnCadOy+4jSd1DVUWr89Kc+af1gBISF
bg7EVW9VX9Lf64BbSIiaWgFZjxrwEApNFfHadO9O345zY+gg1mKT4arNsqjdSHwVpzr4UGnAWtZx
j54s6KGMXfgvFyZQ1LBp0wbTXuKJeUdxti7eyr/cYWffUloHSMhkGzjaoFGP72J9wDs9Pz72jkEN
I3mncgEoup4NByDA3Izj2ZDZFtNOUjO8JsvS9d9cn86aRnsKHrJv7baw45Zho3M2HtcawpP++QMt
Gb7W4uW7Yw9LQxTZSBIbCiACtvgYHEo9fpwQmxBjNMcOCSUL6hLjmhS9DHt4mZ+yO92isOPT/Jsp
SjVj0/A09BYbnDUU9jS7ABGBXECakuQ7js9lWyVNKjf+6APryQ/qLLAgCJ56N+ueN6GXfbiorjXk
Q4piRzIetMi+t5dEJRoywQrlLFlKsIyfbF630CwtRvrqVlcIvmsTxZihOXeqhffcEBEeW7F4647B
yT8vwEUA/CmvYEUb443VNNDZKD6bnfzJck4k3okdH569tZZVEt1VAN/af1qpd9QCNdAGawb0SMwB
aPy47hpxz9bUPobYkI38qdJ7Iao9GjBS4iKhp7PEI1of4Anw6encGNlTwP4OT4GZlSJ/zQUrxqf2
oTOn9hAhVWp5bMhbHFXC9tYNoEY1rXpdfy3OKA14v1Lw9u6r2YcFWMe9khj3KmluspHR0I1yC2Hn
rDmEti+ry3vdy/Lrjj7hV3oZIhmFTZgH3D2tobmFrz0igIsrunCGf4S+YKlf+ORci4ucG3mHki4m
tQrIFtI3AvgZoyXWXT+JLQVNW6OayF6LFjuRubbin7Mx+Y+7mjtwXKPt/UsFLEt4+1yreRViotK+
H8upW47WW/puFr5uQOk04xxZGBKbRrCGhYhnqg3+uuqb/ugP0XccB5jwbps7ayaNEO2jG6Ji+33f
+iLgWm3EXfEtQu51RTrhBHU0/JC3LChz+Jl2iuuZaPahpFkluP6mu52BeHWaZy5582VOaP5vjbJK
Udg6h+34Du0aV5vW/DH5W/q9za2MDN2Fzld+ybnebBkqsvFSPi/vHFeEK1oxPyjbfRM6MnWj3zHh
JTDwIUtC4PRsHp8jhecJjRdYVXN9EuK+BxnqLjlEr5sMbUCd9YL+YGA9wWjL3iy/C9oMDKfzj4+D
2AfRwGdvk4vi84HEAzaWTD6MYdSc4zE4/YY/GxRzQdu9g92YC5ZJoIz9pj/mS/QLXgBcDzuHFYSd
DmTv9TsUsyP6peH/FqcvlVGNmTwQBpJUkablONcmAi5GAo37PFpSP56GmXZW9jl97VbYTTeycXDg
KWDCxGpKyibGuiztsbHlQFSuWROIZ7KnvICyQS+xUSg63e4FnghZvG6yFi8Ucc9z/4D6jLmkfx8B
CWBes6V3CCPzFwsteh61/KeDiqGXRB1kFOy3u9vvAfuXHNFedOFvRUQ3YNXeuOwf9HYF6U5l1Rcw
G3jqJvAb6FUcEFL2x1Yp5xlQ8n3J3krSfwkrNulKylR+8Ip0C3CUK2TVsPpMqY0Jn/sgRdEdfT1h
A5chSm8KYhSoeytT3MaDVlq3wArhtCPisdQatR7z1Az8Iibg6hHZnQ59akD1aYic+hgrti4Ixhx1
XVGoTI45J5rCFcejrjTsStO/5AepodYdGt4J0Wf6spZ88sqoYoJKx1XkGCEIsg82xdjPkNApSHbe
UA5F+dGljiHG8BoGq9t92crzFW6rODa8IUhuks8wI7EBFiQVoB7D5cmeR3iBKIy2plS1c+oWYmhP
dVlvVzdJB1LkiQ953nwsZGOX15hCM+pjRY+KrzPumCaT1RdwmMYyeuyYm91uRBarattVop58+Tch
QPgvrbBpJEBzI2Q/m7QVuHYSZysl7BMxmUlwfp7jHebW2haD7gPJdu2LZnPznW/jXc+yh4pen7XV
+eaV4tfUWYbNKa+FMxD7hS50AOtT9dOyt1ZtfqPdJWm1cuATVcP926vDtvyL3/vqHNFbeslMmHjB
V6bCOzERXfPPJCCA7sIzLnvrygGWmBNb110PQBv8BI7MibPDSnYGmwHJLdfQDkPy9ZVoojb4Z29+
etgEmn6WHIGo1tVfAYqNmTv8mMscXPSLy+EtOzWqYsT94qZ3L6Z6RS4qVv+lQiJXgWPCaU4qVTcx
3mmCsXhK7ED/iQfklhPiHrgUQCpFCSpkhVTg8axQFATCT7SBCXDGYF/yUcc5sUxF9f1RqUozEu7o
v3ZdQdLHYSUA+OZjFqJHQgtX1TM79HkmX2yXZV+pJmFv/woDDi9h5Nrgdjgpr3N0WGqA4msjkS/C
KRAq4RKz6Uzj1bhrvg4qT9ivMZoL1rJsfup0R6G0E5CraaCbwjK6Spgu29PUnxdpySS9PRur+jec
RA4LOxPeLSGvH9LmwQFNPTxc4EhQPzia4VYIt8K8C+qSzK7OOMxuFASs/DQWiR/KOhfkyer1A0g1
KvGe0VbUq+UYAyZKgL4G0GtK4ecWnFHredSC+78qyrlA4F2faKmE+QurHW5ER2EcvlztdiKUEiKc
XPpNHFNT/N/BQA9EDG1/5WMDL4l3zPozVswAcHaKlbpDF/lY/KYDcDVDhxOmz5bIT/SiTLr1u1MH
AdOJIXBB6CyuTmbkdR219YFPC5iUBJdRIiaYr/bHbzhlV2/aGIpZ5OA1xTrVjcvTAuEnO0wxdZtV
XZL14Sh/9TxMuAmEI7XZ9WwPu66WdJnV6AtoxrCs5o6WBnCxPeMkVvadk7P+DDANf8G+bmhY5H8f
aUbdf6d8TY2rCQU9EwNLWCB9rggKzmDr82mWmP+RpBjjf7LJZOsjPIhsKfFeUha+EXxVOUGLhmMq
2b8Ulku+ZEGx43xnB4GdAF4tlM8FV+KP9akw1kxm1a652AoopgGW7gNpdx3eZZue79TG8ife71MD
HoH9LenZxIaBRpoWcNdrtZlv+eMDk9HJxzB/66MXrrDftqQsK39jHZ4avbWy5Ul10f9NOhk17Lm8
Q0JPNe8jY+j2oOfOJJKcfjWyhaPO70VbWH0yDMJgiloUYlLhL+e/URrWupCFMKS925ySVhFEmJKb
IooP5SHMb5nV7In1K/Ct5KaIGCsgq4/Iiuan2Y15/4DbXj40v3FK5zDOEfsA4og+Bgc5e4j7c/2G
TXAJ4WeO0qA36MbxRgkzNPuzRd2T2phvMw7TptBAVwCjAtr/Cte/OEPxYRpVtLjNR7F0g6sH3z5Z
w5GeROZP5vkgGjG89Q8JfRrbXe0R2AYfxX0raiqURiH6vB8xxG21U5rXtR6I8FmYl7tGkdWwFEM+
Wx/mdG9Rt8HWC3dNaNk0GBen4mioUSUfFLbWZSt0X9bBqqmBZyfAeB4mVMMd3MqCtTHlNBvZ+mvA
T/LOPiXLQz2mukUucRPLiadrEwODmxk1gWcRr7WSn36E3gXFADyXnjgNoQoXa0qA4Q75veeNwNwh
DmC2PBBdDoIjEo/WfyxnP9eG8H48n8oH6d+e2kE0C8/SkGrz0mw6RIA31LBUwwC+EgYDHLQi37tZ
DXtlA+mqp3pPH8fNYgPm/S7E22qZ7gov02dPjzvmAzwsQ/qa+WkZFNMVruQhuvycj1kkpEp4/FVH
p4dYp/RLGpK/SDPeKqIzDzmNkaTbCZbZpT/z1jiORiiZIg2RVancriG0XtvN8h/WgxoFbo7GQn4n
NPtfPpqX75B4TAZ0vR8CQxwPMtzOyTyRRRRAUJXcWXCty7G5JpuNEpng3JYRYUH7yu52iMOthg8j
AaAj0023XGAupASOYksBLLRTJb1QvHrMtQd3K6cRVkcHBkwvvoI19in9uF8AK76+sw44FNJUl70Y
yByJpg+MFmzoADvr2YS3ubvL9C6SwoxJYqPsDoKGtVbJp5ifdW7V3E6gEwb+01NZ/ms+4ZpczoBS
4S8/lff/y21D1fKy0w1IXpOuK8N7SadKTtFEfJRsF6Vh6Sp4jHVEgqmTQmvW2SvvV2rua32iEMpR
H2MzxDpVaQzNep6MgODrU36cCGFvMgmwDAEbpy/R0t17rQWqs2G2g3b7HyylRKUJphnzezC3qHhN
sdnuFL4et2HgcRFNYo5/sqG1bF69p9ZXXgj49TEze/JeAktkpS0IEZ6SfQMwbTugcYvoQncxXc0t
Nn2KciIT7tJxz86obhSm+OzX4uoYr5GKTVlBA82iR3SBimHNl+KPWv84mdjjp0KtOssSmaONBWzU
fkkK+7JR157TaAfH/HwYeutbgZ+tmZqgAAJMqztHHpCRtYhFAt6BuukHqX7oks6xaXIVNe6P9QJa
hT9FJj/i0F2QASJTaGD7MAiUSVEkLjo1EFFG5X92BHfInq8iEpZNh7yDmwNanM2OoJkrY0hJwUhT
vB0P0wbMN9DKwiAPaqFZfSMdrT5Q+9iMfDNqAOptOz9hyc1eVL7ztM5N/ZT91T87xygg1xuHVNac
sTAtAn+EB421NFKhfTneQIpXRajojMV5BQmkMH63CC0HZuI0Tu50liguzoBG/Mbp9QRB3JLaZWVy
NfX99cicgLUkeZ/JyyL7UehPyKpyHsqqkq69bjKw+I77/fCht0hnOzHv+zq8bIQ/bSMezfKst/4r
6v09PAYCfh5ozb0mYWGL0q1RQAGpKIdyj8gio7CkKakLCJvbJV0eSIcMygKdO6cAPlglc21Zk5g4
qO/ZUQLrUPgxkVo0/gGcFGth3fiLX2acpyPyt5bfeg9wuKn5DDjx4uXJnbYUWQ0HN10WByf1EvaP
sjqxG3LMepQeW5oDedPH6N5v1ZkFPTNtDPG0Kbfh9D/I+M1QvLsMOX+OrtCr8XrxmdPL7CQ6h+hb
Dcp+QxI98jD4tH/f1ROgT71WSp7C8wkRwoajgYOTTl2+PobOMUUeL4oGzruHYui/gcOu2vHpya8T
Arox3nkENAqvHLLTkflwQRn0k0zpHJfKuf/c1VOx3rBzop6hcm4OG5DpOJ/TIDj2qcb5mC28OtXA
yZEbZi5NY1KCjS2GegZVxpTl8AfLHtuKMco2WdfMqg5gt7/+qcbmnqShlRt5BCQL6MpDEOqPj0uB
v6sMQUloFeycUs1zgf53+dEjYEDYCu7yYKYfBmwNTtP38E8Qtq7RSKFwkxcRw/xMJfas89vRLIwe
Lc7PyiX2O1HsdXjdhqHsniQsm4IXNDpjoK9EEsIJfEORQHNESX9OOSdSAKhvl944A/hy0xaqZbm3
S9VTFsBtwfBNVq3VN1AV8BYcHg4siPX7jz2wUYU1BMcmvyV9DwGFB7woyJDRXdtPLzDlPyWsOCC7
ThVTFG6WWgAoe3GCx3cclu9aYfy+RLTHpn1cBNDfM2G3l9UmyCTfskDKC2oioqObn8pI8UAf7KIl
nsQ7blZ59f/4ZXGse/1b7QUe/B7CnEyx+JUDZwDam/soArxcuGYVth34wi32ilm0VuP8qEgEYLrg
jxpXX/HWZKE86ctl5XOBukjALhvWWFgFXrbOF7UN1onJKD9mEgA8fsso+QJwaxiYPqsTvSdJ7Sq4
F3VoS3GwsHSo/YVo07bLSRA93TM6grd+6bgLgF82FkWP44ZSbHcH7B7WsMwPlTLu3TNZx1JOhCny
B3rHBcSzYTQs3SIFah8hDrySzqPWELV/1SecmbF1+CrvdxHLefTtoUJs6ZephQys3qhlWlQocvAI
sDoH28I5dnk05mo6NOHFQPL7lcCoQwnj1ENX/a0YKdN9EGC5qnRE0UsKLvTEWSnCrgU8djwciI+2
U+Rwy+2QR+X14ULZd6WSa4hOVFAT/ZVRKBYrcUA62o2h6ch+H6W4IZYGHAR+kY4EE6ZNkUZfpDbi
lnxSCrQMPTHxRJNdA8lCeenx620B3e3XClTU6h1CUGrixq4Mmef/5p7t3LkNSfimv0VvETFCGJ+A
ZwW/BBcVg/7qZMPYXjfjqtz0ep1SpLb05mvL/kMepxtBDwbHELZRaPv5LI+7N8MkXHV7UqBkJBHI
cjzdRSVoxD8ROfw1Axe2eAxPvXBddkpHzN9E+9nSNG6DWXW2dfWnORgM3h6iqRzuqqIA34zXhOUS
vhWn48lGfkN72O0dyZ4WMiLp9rwJoOSLoXOtpq8Tul8uADJ3eXUXUhxJwfbguWO0uPN6uOHsA4ms
fcln/qU0C99ioiKmLI4cz9p72MLU8cU3Y+38euhlUTYGptQk/7iEM9BUf1PCnnxEXR4uPjZsYh83
QqTFhiwC9aq7we7+YFHW3v62s8EoRZUcvJ5aXNVQypcWaaosIg4QUPh7GD2UPrxeZdaMfE4fMkNz
WQtU9jzL5eHL3++TO6e2FOKC/kqZKxhPMCWZgCulDranz92/iVk6nCdlY7DTFhfSEbgtPfMfS0dG
xuTFrC2C6SLyFk3IalNMWNIzeY2ItJQ3g8uqB2UKMSDXT7QXcs31cgbi/K0gsesXLk6drEZopVO3
m5c2hGjrZ+WZKec//iaa7v4J1kcY32r+iKlcJ90I0TkaoJbqXucrjpNeRNRL131WFWjbTzO0upas
24BnszK4qBTLPJ6U1RQxxbgH/98ptVrzNfpDuFt+sQ2XbBPFiXQtvyKcHqwsYIw3wBBNfXk6Btdv
8v4d9eozIOVfVjgBh0+8SSu+8obh5fCy3aSket4c07zfsOPdramvH/VAj7gCwu1pFaWyJgTC3nN7
7emOKf2uPK5a2QP8bv+YUO34sJTWNrkkVqQDrxsM7Eqzq/kdXsqVS1SKI0iyXEeDamfd1iVSHP1x
pohzEKl9R9iFa/Doqr7WI52m+TUv8nhvPksV4YZOxXqIsdtDcueUXlbSiYUKAhzcunhRx7F1cK+Y
0XyYC/yja1T5lc1AjPGYnJTeDMWx4dNU9FOHxg81VficMt2PtcXrHsOzzCA2MkbwAZsiCBsWWfYB
FLLdaIzprAYHDt/Osh62+U+ADO8q7avIQgt7HDjrrHVXkT5xSTqQfikPw5SuzYfIB55zTZXPHJB3
rnVEb7ONFXwB55XmN7yTo82myMokbkHGjSTV8WAlH5c+qRi/Ac9y4YLoiZLzljDyo55MHSBiASLf
QCB2i6dMiPNEI1qzXkCR+XqzDphaStS8yG6Gy+SyMTVvntGVtcYLMkxQNwXssBWsXPvkoNrfjpnr
QwqzQtaH1p/f+TZPGMfHYFErMFHJAwb+lKnFNrLIwxOEE8bCoUGBeLoavefIwY5chA+VRj8uo9PP
fNVpReXRAt+DV/xCX5GM+uQbHsQoylFhwNA+VvF8Icx03bR6BJSrjGKBrtMO2uTAxaO2TsBgKxHD
gXdu540Cx2IVtq3vdSwlc59EimhPzL7QKcEnQxwvkazdPehXgL1w8jD3JaxiaYrj4+zI39aavCA4
LrJ+x42KdP9ok/0bij0Iwn/SsEL5uch6zQ/YJmwqW7zq4Lzg7RKdgI5UbYiQ5t9rx7wjw0MYI/8P
FvqzigNvuBiIUSWCleGDAIMe9s2J3wCUeGnCU3MIX5ZKkv2cswyX4qMlr3MHTxSQGek3Aod1p46y
FK4gubGFeBVCLGEAn3wmONFXktVIQnkJ9Fpz68u1Y2HF8FLcweb3M/2aV7PNmGD5XemPetcLteyy
xliHtKPdvufWfFpaXY3JaigSdHUxChLyLttNa2y3FeHjnSmE4vAeXX487ni0hXuBmb/CZU7R42bd
pz8amFzT2XYRQ35wYeGU7xxOSxGh9szlnIvdnYw9Qe67xeM2fggvwtjNORJ7xZoKJwGUE8IxGyxN
md6zPpnoO2oVr1Y8XL9N8xjUO8cx3XLqqIahRkm51MGM66NHVDwXl3O+3ix1Bxy7dQ9ABa+aR2P3
Pp71UizSs74mkpxBOXhkN9CU0IsnCZTkhzDHoKZL+UnsgZE4ogGue/uV9l1pEX91zZhIgWUFQs8g
wQSAiY5HACmxhskVLRFij0NzDPi0YG2HYRRhGtpoRjvv96i+2772kOOqnqqw3TLN3czAe5fc9yKB
ZmsA1ogIZyeoQA4/k1NJlA7EVaydXmG/rZcFCKKeC/RW0NaI6gVU5G7FUfMhoEox5PeojEOQrWEN
1XR7dvnwtc3zvOD902fkIdusmJ09h/0hXL9JUPASx1zjJSzt52IiLBrsmIE+wCRjNTDTTEiaXuhS
kQfueG04k+DvAdC60nH4Gzq5zmBTTnHIAunayboy4ky4OuUOKNt8+Dyh+bDLC9VL/EXPxl29B8yi
oPFgCoMoY5GjkCOxKlyA1/y4SJWECQ4BzbLWkcfUasSxjUibAHvieOVPCvEw3woThsaj53Ke6ujR
tWS7NbsvngzLchQYY30EbgibPRTtEg3Dk424pnn5xDPFuYvBCqHS9/HmiPp5bpOLIZgOKYABFXR1
Vdnfc1ND+5vRBkwzmGQdnD7Sga7bjkO5FmZTglQ/2Jv1d6OCJJOu5AgW/hWqNuICkjebJI5OE2SK
0zLQPfIQq4XHbzVsB3G4UdTYuNzsNqOFCiJUhg0AHm3I3++lQeQQLHw/LyB+Fid2wf0+69H94RP8
taWzakyEHFiYqIKLifsL9ZuCAjosT5hSPpGTV6wRaJUSV245ka67aNLi2teX7J7pvuQ9rYdLbIdw
sBOek9txGRqWxioruveO8r+IPzsH4vbyDn87c3xcLIr4xrpZGhl3IfgVc19rPfD5NSVZApW52E8l
enNwCwnGkPpDkdXofgtFA55q390LiPGzQoGLdmsg7tokFkCb7umvbUog7WJICDnVJbHa/vh5KV7l
Zj4rltu6SFGag1IG7V7ckLMVwNVitkosQdc5JZItIl/qxrSYoPZHwGGLt8EopgLGpk4QJsskLzPh
Q0SLeYXesp8VijvHVYkWlPn15XW15rZ+gQuQGUVRGhyn94RWppByYgzqJQ5a6mwWWWJHrdMEgkZU
8sMWKT4U4+07NMEIFz9LXdPBPU6kWO9vZuIBSqaiaSv5hgo2iQ19Z/dGPkunfu9yDA9skNhs2pyw
3yyj57rtAdctnZt5BgktaCbmu9FWHl0wznxh5nQhZnZNcFf/Sccy4L6xVRBqqOP/8pgvxrPu++kK
68anGXRRmW5lHaLpB5YtPnH3SPi0WVN1BFyB0y5/j1Q+478YeB05HUgxxPoHkmkdDaxZH4rwNJBv
5eXchmHuS/VEG2Jd6Xt5DzAczRbn+YpjLuerli2i9Xf7wPuTVITyKn5uY7HKQf4VPTQfLdMHEXoR
NHr3bEArGxuYU8Nhv6Nevh2mneRD83O9+sFK9LlGYmUa9P1flM8kgEA3NCVv3lC9kpxbaCpXB8T4
ZhX1u6LmXJ+4l2a1H/UBTpgZ/3dUvMbvMdpC0sSV199EpHRRyGoSNdtDDsNaSNqXMTCcotji9xFw
hxbm6DLjNpTDX6VoRzVSGWli8BrJiceOfqV2pz8NsWzYn0PhouXIX3CD6uA59tsy52mQ09GUIl62
+9S4fGeO0iukM6y1LxbYMOAK0RIDJWFPJKBoTxiMO3vZVQ4nVEaINT5ZaZ49ENmwBjWoZy3y6emY
dCzrJVbbnuJrCfkgBChFs/kveiEgBOuBeTE32N9ncsZUjtf2zaUotaXIJ/BBvKn6T8k8U6Gw4re5
NyDOcPbD9d/EqhRkwYKBanaJT+Qa9sr8kAWQOO8ZywYsts6MIe8kpJNMTGb0SVjaoIszNYwcQPSA
BPXj52HCIRSz9uGil6CyFAiE5ndmWwVyRo9HnNaKf9xW9ur6UOhNhPNZr/M+PBKBBwo2VmNlsgOW
4nUi+t9q/KkwivhxYpWmU7RewBFqXoA44otaEPPQ06bmvebADwBWAcZBNRKxCcvo0ic1JDf7XUON
jAI+duZllaAqjeB7d/rfWU1zfrh70piT09eDwcC44PL8s5Y2/jiWyrsOMA7I+hd5D8pH2i9gIyHg
TpjMXX7vBGBUt3/xV94DpE0tZlXgenvF+nPc1eJ3C4uOX9HoNzqGN0Mc22wMGYfM5j/tYtROiRR4
bCxeVIJf0KxJpUtdWfbH50SYiEYyooR0ZOEQxyFPIEIZxrIdTnxQ9DswbSREs+PyFOcyE03Ym/8b
53AJbUuNlHN1h9cjrwk=
`protect end_protected
