-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WomZP8Z5WWtK5kLZieUEu76f6wyDHExNOGfgKY54OliPqJno1nDFxpphvX3waMTDkDOHrnrdgUUM
79aHEFVNbMLQloy0styImrgNkqFuL/HkUscgissYPftSqeBbDBakOUAGwadASKaP6v4yfPyuSif5
THcAeIscZlOAdzuas2b04y4YlFpFZhWi6+fW+TrcILkTcGw++eVmwEGKCRnE0PdAeh/WxIrqHYJm
jup3VfA41pKN4ZHzSxxf1/yvmNFlhAVElEdGb+m1gAbV6sQFyIRosi9j03+opqRvoGvOV0ef3r/+
fsIckiBHKCnWtYW2tHqJ23eBHJ//WyCJgVpTFg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
7jN6qZXftSd+utXaso1Cc0BenMafDKsYcJIaDPRihyzvJQkneCHNhMfGtg37M7ar9uD9dZzNFLGz
OntC6OzrVVFrZ5fwORc92DYBCkjyeEbhNPXd7olHUhx03v3N371lm6v2g1pMBFRWmRwoZahlsJeu
L1lK+oz98537P45S3lVhK9fILdHMlqtuZNWACr6QeGQQHoSXMcOnb7fiGOArMa+2JJyKo5RIfwTo
0PYgn95uD74KCso2KA1NS2n/X5lSYeQHLMU6zEJKDmbFuqk00kvGjRiy4xlfyn53xQf7t/OBPUFr
j9TDPTrrT7nvC5A3Y/uLlkGNtqIWABiD4xPO3SzrbWe/UFSdA+MPRJJC5NTpHTK/MUAQi7M9AyV/
tIqIMO/CcpzS9k3EmMObhV+/7mAOTLEkCXB6YH8H9APRJ1qCqSCWSckuVwc/WcEeDAEVND7n/ipj
w/4bhM21rk8c/uq0w7rt8pWEp1Elrj92TY3Ombj2awkkEworLnBqU0kivckZwWZ3tvyq4OEcBFGS
3REboq1wCUQ3AnW4Lwm3gu4S4TXb6WqyQiBIEvordZt0u385YBHmZi5AaGNBGznuLKvrySpXmmoR
Rf0cqS8L7QM50DDH4alPn8rAzc2rV1fCsUULVehpPEzcqEqt8NPgF/18tLb+vK2As1mDI4Ch9JjQ
x1KS6vSSy/ONAhF2xni8jyxtShVYupoEHJhQvWIv1JeMjU7gvNobJWoLdUtTZuWDNUDNZNMjhlsx
5xKAMmxZaHRCjLvG0J6gXjmIUIoRBH9RHHOXR1/KOHw7HxTT11BU1f5a+Ix8PTrWoLeGZzrUpj8X
4ldatRs2QAYJEIwPp67jwOJjR+LttOLE/uxE4xDF7xl6FQRQOWByV3b9EHWVAHoHOVSQY5pC5wDu
E/OP9GfN6qysBfy3ekRxjGd+RqZkjhB0ixYxoK6mdH/RQjtMJEQJ9FznCoGWo8lEB68TMbzTG0C8
FTsYrOzPkJV4sIB338OMXkhTxZ2UPmFD7G7z3qC5CteHYzO8KIZ/dZBFcGvgMQOLlb1l36ZYtUt2
ICRWhqqobcIg5BCAiaBsoLzZRnAfqnM72IlxntNNglKVukYJ/iTsOHNs6hEPRAgQDdw0ZuOkslT3
ToL4ZwKq9+Jstt92cFxSAWZep1G3coN45yYT9KYJt9Pq3hABjaOIBX1GYuG+dlA3lQJqTBLY5794
GmEzGUUQddLpKfqDn9+91yRp3l4THumQpDKiSa1cavlOmRhYu/EWozpQb7mBaE5aORjuwwgAo9OO
PoMD/GvmHQi2pLhF0XxDq4aIyoKrb4K8H9yh7sLnVnHbSa/7FnS6tiD0N8WlZOllPFik8iLjphho
RsLiPRoVN/hv2Lx9LxKqVBwjuDMg13ovpOt+wHvblF3ZlTiujbHoSq8FrwHllqYyGeHAOaFDGR7q
/xWkVDRFv3x3aBWK34nEVHzZJ75H51h77WzB34iqhICUg6Y6+gUmWB8vJNrAItoY4R+qQbuCN863
oCNTOy9RtCDA+1wdIxh5DAOKJ1uOGv2TQChRvMcRjIKBPMXwHdd/QCaIgtAyORqjRhc23oHFFE84
XpRhu4WlRYxYEkpyEcnVdBhQSQM3uWI5DJM6mDLaFGJHc0d0TOp65n3HYrgz5ZrtNMmHD8X97r/l
bAMLkEubX9AdfZcZC48GsliC20jIi3CQJZt5K8aWU52cdlNOsGqjD+d0b5CZO0XML1e8Cq2bc3IN
Q960Io8AgDCbPb7eCOV+rfK/Ntx+1UCms4wPM5QIzwURxYsW4wfWAqeO3yOu2UJ1FH5/Scdzrcc4
hSyfLrQLe9fS1mFtdKE5x5NN0GG4Xmw/C6r8fKGyqpqX9tTZnKcsiNjWYpzncBfgZVRgDO7OhcOG
IFw/COwKhIJO9VBpo1jdljnVgXVqR8PN4CWVpgPxgEFPkihkR1EtlaWYQ3lH4OSQnk3pVZPIV/1q
bm6/aAq6SZA2fW1lj3EvgR32yKe8sP13AGcTnG2jF51zdSdlE4sJgYSyd7oRQu8UilNJzqvgXSok
Q6Z+rMoet/73XNPwd39ngtznc40/FXeei/Q6Lm8GlliH9OUjd8HJTVVnvu3M3pminpM4MDTsxvDc
EfHS4xRThDM/wDutWUP3HHA3JvNelfgsTpvHJ5aDRpXe6wycEibiCBY/oNo4l1GWVrTCoydpG8uk
Qm+t1JEIOZn12k8JdwbAbI5oDa6SjhernRsx2zuynhbYXs2Ix1LHuoKht/8dKcx2/eFGvmImaAm+
8TY8BbiYUBSsqxvQCYD8IBqDnYMf7iURDKz8se76O5NsRE2iV7w9BWjboC3oQeTKlFurqQGz2zxC
O/z8VptuyDYGY8BGS1Uxf3OEmB/K1cwqPWdnA5pv1LFTGTP8dKVvIsXgRpRv+/d8WdqKHtqTMp5a
fiKyKn2hmlwvgqruOGAaFnxZb0zlCxCm1q7DPTfpBonVFlfItwOgK/dEw7unkF+MIq7ee7iBh2bc
m+jyIvqG5LWLrhUFLxJgsGaUHJCAbekALDd4GxFZ2bu8ZOljk3JHaGUTciFgpF39lZ1xgCDJ+kEW
WMZ3voBn1Uee97QYkigkdN+Fv7EYYqfxE7xhUPCazpQVxu8bnDerHPBOlKPXw7ln2jKgN/35vh00
UNdjx12B2dh+OehN3AI39qbPi0OMP7dyKuRx6//wrHGD7T/tpPr29uH5ycOct8HCkYNNItbrlme7
33rcHaJ6nqx1WoEgVeaEwUkdPjtaiQHo6jA4M7G/C3wD8Miotlpbu+DFSYoqe1MWkiWWdsUtuQXC
gcsaDSSp1CiEdZER3eudvDZYXgzTvpkII9gexuj8FW/pGk4Q6KuCWOc1ThoNSzNXX3NckEzN7C3L
AvkXF92TG4rRc4IXV0TkwCueAgQsH3zxTgQi+Xdqeh6ok63cmUe1AeXGsluQf7xuux8cQaM9Qiw2
T/kxsI9RzWEVt7bx9ZiyWY1VPRR1+pRPzdj20wzbIpghDhg8CUnhjdsC3Y4Vg+G6BrZSvWMTGFZ0
/25UxpIl3lzMiqcCtlr7Ci25dngjcA4fE8YJimNRtWTnqIy+8HCLe9sbLOqWIm1qdOBY+oZfLQDE
8xW5rdKGq8tHK7l7tl6Awoky7mb5t5BX54DtQ6feP2P4KIr8WH3HDNt2N6e28OGPw2bb2XL0KzCY
x7gq3ndGDbXuQ44h+5v1EXGdbptSKzaSqS3Qnu2Bw/xSgizTSBdty2VHeQ+3dqpfDF/mdA7gfenY
B/HevkkkEqnBcdzWXdwvDUw2r5d8rYLzbG8wh7hlv1FUPjrwaYYX6NYZAPd4lEmWyDGfS81Xyhy7
mqZp8MKIzPdjZ2QWBAVjhNCoCC5BtI6tXSpsHCmQUPOLgAImF1J/VmH2ocMVATyOHFdz+XKYuUkx
L7ja6HS5ciXGZsSXIj9xp4uuW78vgeRone/PbqPf0yaWy6QJpUW96WKvYOjVXNtH3LVevQT5b7Uf
1UUxJzKvmlPlWBz35/h1Sw2+aLb5u21xo91XTYRrrtGSs3RDbnhV894KQg6Q7GNw8cCXwfybkOtS
W/1kIo12NSDH1ScAaK01K+1+H44XM6Bfb9BGaZbow9lCLQLgMZQpilgLs0qypMRMu8MkCZHSsrSw
TPsKFOnLSMConSQlO9EXB+wFVpVom/b7baLYNgzpgmQ1IVPRPvshTt6unEOpAvhe+pbfEn96x7/p
vS0YFbBZJ86PVK7uJL+TJb026h+L0GATE4XvT6J3X2+iFbTZ2WpaTm+fJcufMlOvmFzyXmRFnu88
MGqyEjiZYeaG4NxFhTbb9l6NHeYYTH2CMVyU5ku7S8ZdnPfxsXQiIIYVJ3hQRX53gDdSrJs2+OGq
OF/xWwqyAxzY75CkdobzSle9anZHRCVJ5KH7uSkZZRc/q6XEYdWFbz2cxlEqrL8HpbAquEHxd/M2
xV7VqPuOoubsgJq/cgZjgzRCZRF1FTU23JzRpY1WjmI7+OKPEZWnZwTQPQMUSqbORXM9WrFO9aAc
ae9vR4JWzjqqhVu4/x+HJfQXwZ9Ez0jAA4XCwyl+QmOv9P5lQbeZio+raiM6EPbvFfl+0rqVgnBu
IbG1DDQC/geCDz6xG4i0iLzZ7TQn31E5zu9/fzTKsrVvXVnMo+B+6MnWDlC13zhy3/2jzNdYJ6Sa
JGVmnl+JDsgoaxiHwvZ1LPmTN1ccLEtt7xCU8rx42Rl9hDsthwzWHLzYAIktLhEQZfUQmuJjrNGe
AgfX4pFD4V4zk0Hc1xUBqZ3zkTpiW+SJuBdluWzr/4+Up30nGa/QWnziYDvhOeAcoBv5qWCzx5iZ
4XYtD3oOswFlvS1Fjl6o9zq09D1HBb5AX9RLzKWdjMuD2zEFT1i7hsDfhGJQD5C1gxTU0sFB+vJv
lwMe0/K6de1m6NCisuCPwwqWiVRmspdlqUKzUkgwltvLq2DhTW8mxkD2KlbQgRr/EwJDCvTC0mYB
g1E15sKyQXy3pR739NSTz7r7jvv/DbKgUpdtFVkylY/stgqOnPwsRYZxBo0B3EdWsXzBU1r3YxXb
Yic/yWFzJ2/1Shu3G7kY60azZf9RmSXRr96calr7o9MqG0ixmqGjUwsMEQG1vUuVbdFO9Ui8aGlw
GX4W5RNZa3OxwNx7Fs3YlvzQEDqpChJXj7Tg58HpfUlTVRTR+XLayYi2KMUEeE09ZcO4MKy+5o0b
ozipF7YJ4fpXibpiVFhAxQ19VPoI679O7WiAyKrWjNCo+X5ebewhnsa8gLJMynyfQNm2cci1dVTo
r7VUQT8kF2OLaN94t5xmFE3KrqaOM+5W9XUBUPk+sEH53uwMxLv2shr/zbQ5mMZmpHl8jJXwkJIh
jok+OF9FX2Hu5PeIOByQxR5L38h15yGKYo/Hn8+o+nYqHbphEB1Lkb20ViWYab5zwkISgwdawdNy
1DluNK6MXYkNlAuQ38PbewJgEO3+/jRbU0bhX8htkB4KOYnr5OZwYJ3K+aWHJB/QiCw/r3hdkGaD
iXhL4mYZxLmWV75T45nsmsL8OncNfmvmSBz7MrBIPRhX0l+/n7rWKSyexGDC1sK85e8/rv825lNi
/izWsn4A8+WZAtf0r0QdaKs6PCvekY76wPwJwvJXir3KBG1mCnznkBA7ThOfCLv+CTN3NHrLAWG1
zdKbpdaCUPJ1O8LMcVGh16qB4sjcvAiia2AFKRgwPmSLzwpnSVyAy89g5u9Z0T49D2kbvZtjP8xw
nG2tNmvZc+oemiPas3jeyfApXAi4oqV8PBDfkvptmnxWOHz461SeJ898GUibvvs4S7obLVER3XEw
toNYGvDp6o6GzECajRFj4giI/8qUaBbu65H70ZZpaLD2kUkRG/EL2g4m5Z+I0P6TKV1aytc/n7ry
OkVJ2XeySihJKxbYihPQFtuXegSZ0DSjE9d0VCqpUIiZ/eED7ImYuIOakoB/372k1896UDikUnsU
xZCEZzyBFtQad1LNIH2vvwF/BQc77HUnM6eOMwUyZSTagTiSCeBtVzqLtlo1EoWAhKlUnQcfbAHO
8QF4p90RgwPmUvtSTiyBQlM2+KD++E0FdTTt//lIPpM1SdNm0U3lZEF0y1LbBde5gLrv/onmlE82
PCzfV5y/i0w8KsM9y55IVv8na6DZ/4J7ILmeXalTJVBBIVaaA95qbw4sxuua+a2r9cdQaZCHSCAI
TQXViCuYySV8WPxPYpPD7hrCEoZaGd12d4ZjVEzHwf/zgecfNKokhhoCY3uOHlyfDu3ivWFmzWxq
dYLVDtFqpSu+k3Y5athsWRzUCD/ecDrUMKGyUoRaX4DTdWyzQuYoY+RZ3kWgS0uGsEobE2SQOFY8
6Cw6Z/RaXXJKruPR7YV4gR4aYCk0vy8y8RZAEzuceGPpWLNr1r0z/X4ytI7Xm7KQDQmFjWIm2eAT
vjYDrXvn4lbn8xOpdzVl3TfT/TTN6uI6riMGt+QIYOSo8yUHliP4f/95DuBpk3V5DNxmB00Z/+v9
gUaiNA6ozjN6meYZFsbcgQBdvdAciuI1yDNiD84+JuVcHd0YVi8rCPhx8SWtPLdLTKaumB0tMEPu
QaRSe/6coqZ0OASWBrPMvqQ8Jxj+BLiK8HKcSkpczPzXZb1jp6Xwc08QivumRjVlv344WYs+1Iwp
HmYpsrd2+X3vrHnUn2mjGEUBv/Up/+irUZBQizAqIh4LAoFOhBQZwHV4cfPnaegVIVfNXfpx+2kX
VuJWi6ayarexA6zWsivBYQr5uUWm9FGKDZxX0EecsBrcGfvl9B6wq/0UznazbOZfSOSyT/dDUwBR
NqcEGFBEaE9SK53IJEFC7S7Zi81wKdPW78EPeerptqE8R6zx5N8r0hOaNMWcI34mQ3kzcI9Vdegu
WStWwFOCimgipVtcSBpVxmB+LjOmF06YPYdjsqlxST9DMlQi6/Ok05705Nsdsoo4OHPaTVDLeja1
cj1X5GK3AYlPJQwc2dFYqgv+ZBHEo482dCgSAleME4dgKzipxohbR55H+OmXd6RZdtSAlwrAh087
q0vz7GGdDMsyNKAojTBYiw7lGtz7UZ65zDpftMA7cm+SnKbBlyMJruSUCHqY3JMZFjnndKj1z4z7
bshxFOBv6Volzc0VbYzj/atrie469IxUEMvn7gOL8qz/3x1ZsfexuHGwPa3HAXZYgKIr+7SjjwlS
PQkzaeBE+QwRguhYozv1/QxBr5Fg+FA8nmwIBUQWRIl1iwk2iEwOTClpt83An7Fb2j66GtUugvst
PgfxtEEYYshcq5zlFeRojO4vxhC5v+T3bpUIcy6HECDxDh1XZEOne/nu0K5o8SfOpWO+eukfgVk5
H54Uv/I2QG2w5ka4vbCz4DIGaBK6VpRpQfdlsyWczA/6qafakJ2lEoU9tlwKTXy+XIdHmttM0L6e
KJk4yxnRnshxHXaL9dACGYH7uRIKJWOLu6ylLFnLI2HMKGjNPHY167rJOlsnFMoccnz8mxpTw4NN
c15GkMbZg/xQ9e/yImgqjst7NxlZQP+AwEaJojqJYzDc4MH2AJHMY37SJP12bwUYusU1KrvtRjc8
9ZQgk1G+U+pZ8NJ2cgg2TGJv/dt9eLUOAxO6kCeQXb368kfOKwmlhYatVTeChFewouLfxZ7FAMo5
dc+xShLC/PrQATRnIamZKR2WYsXS8ohWnB+wsW2FqTFbf0Aoj+CNeJWa9MkAfWeQlTpq1hKYSpp1
gklEZtqvUMph2dqLQvs7En47JfQeKu2YlJnMnv2IqYHrD2nwoBnsr6MXtyjfm4j3bphRVjp3pwJu
NlHl9dcf2oYkdZzEVe3NyEM5YuvO8EETbPcO+QZVZ9mVHEk87RfZZ6HONE9niHg7E+qrwJkQ/MNt
ZxMVLuFGb2BNxBNUtWKFfYutjB/SjQcbH43FHOYH6BYTnI2bGazUM/iFABNYJvDYvpfMNXwfzyX3
3/pLhKXQ5ni8pv70RcHlqsi/KyEKAM4FoSREg6zBl8rpQpI25O+XkeiugATZRVTxYz0MKxzFG3kf
COePFc3VRbX9UHTyhG68+17i+iP9weinLdwNub/lWoGPRBwht4oBhqKVWOBAMdkQHg2VGbbuCcGx
CETk4UN9EolT5uz36R2eO/UJ4ZmNLlujQWMq1ffafEMnRY/5HjiHmx/kZIDvF28xYpeSN6HPpiTF
PcdElXYwDkrvOLbG3x0C+j85wziuXfSQI8XcvLNwCKu8T0xtDyoYaLlOreBI9sC+o7YVTpe/2qF9
J2RniQclu8gq6I9Vi7n3Fni0mtA33Pa1I7qkEJmXwcM6eOKob6lrbqxFPxvl2ojw15CDzsiJaefC
gU7ZAzR40r0YK64zO/ncubNc7xAq7R48Lam7RZxksKckMph0q7OEeQqMRYsxDFHTX0ijM9+DoWNC
mCf/pqjqviYmEdsEqmNF9BeCkU5v6gORKfqPh6uWITUdh2uBC8RL9Grni8gk5Qh4/M3NPWm3De+h
ZDgO+fydkwL0aoPkich9KCpE4WMLSCSuxRapQ0pLCNhOEE6EF2YnqkhPEmOs/z/xSVoDE8rO35O5
Z1YqCEZy5mvEfAL69la8tlrv+Fdj4EmuqxgxCM7QxJbPvpM6qY7PIYNd2Xs612QgIOmy/6nEbnEX
tYpfj3RRXZvDaacXOiPTCnsxvXS4E64dvrzM1RcpccBE/1doW5jH41lyqRvpiGlfeblS/wtHTyfG
AVFpN99p+dGTAGgdNDhjnyrjJKtZF5dtn8gYl47HQTgwg+Z9Pm8Y5ViEaomfQ25xb3uWeVq2ONGv
IClmFRq5w97BDdXUHe2wHTT+aO5n1HzWu3RSWxyW6rci27a2bGHG1XBd+icgb9B6stwnFUfRywxD
p8Gyi5h1SPFM4GpAQjlpyZSCDbuQpM4ujzQFJiUauFoaArDcwmyQjRJ6fqu6Nn1OiYYx1y3PVkvK
E19ftOTPahebeAG7J6UgXpmiQJHYsj1tbd75r9+WVg/eGyEDxliBs5TisBdyWst6GwhcLB02u6i6
6aTDoELFeOOLCkkn6YtaShBbfQcuhHSSh7WvOJ2B18jqlB7PxeCxyUPnEiAqSrmLol6In3Kuq/j+
GuZLu+QKfBWC5Mqc5vP8XghyUu7oL7TJc2UT2SINQrbfdACxB59KtMKBGuf/oLeA9wf6N+z0XVDi
aThxg58wuBQhlWPBf3zbMyzOqvTHUFiE9Xdsu651l1MfHwTkBfKedTqJ3RoCxdfBfBYz9wSx7riI
XGo3soSDbgjDooVifvobA+Gg954qxlcj6dtSEOwEdjmKze5F0IFSXamfergzojweL+NDtiFG6yW4
gsC0wRcLYubKCUc9ONWMDYiM9vD3LancV1+dOYfNoSg3Mb+jaEFmnzR88ZsigWXbmsvcBfw/dtAs
4g+Jif5X9ysEuUnvm0s6WRFtIjlBGSiSg7iVNJuwqe+3Lc7mlT3DU76IQSgYoEKDqs/rKdQnGnbr
2+Nvg4X5h+VkK3o2RfmORD/jG54KF17fzNL5oy7WcYInPMaNxxfD831o5JKMPaZc2FwW2dAMgl8y
A58DzMWSMQ/MFT/p1JZ0jrr+JYEU3heDXzw3Uf1poazwtxg/HBDHjnK7lyhoeLiis9EbvT2+vuTP
mHvG8uOefLLwENjEZl23z49o7FdvspqGFXPVwm5GrthqSfzElym/2qRmWXYMni2HxSfPHDTlfXRK
L2EkF30CByRC3/KVq2xhMPDsD96tHO7guh/Fw1CObPPaSpSg5M7awyBUd7x14lMkx9GFnVqa10Ww
AgTRzph+LIDz6VWS3JI02ktWz48yiisCsWhuY8ugntZqCv516iUh/dYUnJqaFD3YBPTqR5JkJSk+
FHvWBzAry8AtpgNLdkh+Q4wJC5hC+rlohU9vyuPTBSYE7Kbv1lR+Zo+ROHWiREAVKCNk5U4AFOCc
abDY2TyNENdhbP69ZRlIGKDI05xyOJJulmGdlaIrGddoAQWURNbgntHO0KvV1qv1htdCT+7ErExF
IjETO+/0zT4MqZI41LWPP18Y4VSt8oWCeBF66VlXDqh17qQhdxMGY5Y2SiEltc8BFkNhGFM9taTu
rCLuyapLCiFnegXCdxMZd/PIcLFycW0i3Db4rUQnQbvcge/xhuGDhllE0woySaQK1rppwm5zMgiG
LKp7HlC+tlnsd6g2bTt4uOqs9I8oyfYKEK6WKJhGyy4Ol6EDlaTbpnH2yvNy+x7h3nLT9B30N20g
VhmAnCwOGzvJjNBW1JdLVqbKIdicQlqZUOLVC7DSYSiCjkh1iYqDvPDfncjFONP4gZ9T3vj+34Mp
HLfuEyxWwOR2PlmjCBnwHE6uR0IVE89bspdcVqZ70DA5+0je0pYIeXT3sGeW89OuklnapxYzWZQu
VHVj7GVAXWDI3ht0tf8/sf+Ko+3cfiW1fJyZKDMsY4OXWsUVXCXkrmImiHfwkxzCGN4w+DBmpQL9
rkwHM/DrxxN+w79NC4aYX33+ngzsQH+zbwREuo6u9WDwCmcS6JN08aUfiWfV6am1WPVa5/v74ZNm
x88JWom7kJ10IrMvBUDSprD7/FD3JjYJ8YKux5rJhfrQ/satUIEm/P/Qn6TgF+km7Zzh+9Rt+xlu
g3ND6Jx8L3cWkL2YYXFaXK2sTwhIHGdhu24pO7+zeh5/R9oo1/URZYrzcIU58w+lWOV/2HfI79e0
g5WnL807ZkuhRBk0WJ/RRgHmTLAbk1vxI7yApc0K2fUQlEEyyL46g5l8qpub3KjIcmIXMbSWwz+3
pcEqWMdprd28NyFBhKuhCP3Kv0uLaijddVe7mRNgufmh8DErQMHS/vy6ekS9Ddjisv1RpUVYq83O
RIrdOcOREShypbrxSVpSX5YZGnQAEloXEddd5ajr/1QkwJ0TGodtJ4HYGAk14qpVIoKQR6Nb7RKn
/hWr1yIuOHnCBYnEwBooNaI3vPB8801WeahnweRJ0SU7IYmtDRP2UBYQROS3soPlN3KYCIG7MNVM
8WBDMA82SVNzNAcoKHq8/k8vd81JgV6o1Ye2JjOvzdHqPQuQ+pOa1f724QM+r4hzMjRu7pOp7qqC
03kZXddMF284gT+WHPBeFyAJ16112ADXgmcfRUAATqvzbzNTELlQS0L4Jxh1xF6z3zhhpx7fTzyr
qRtIiIqoInyLha0XEbfx/S7oaGmbEp01DZzgCO2tGKC/bKVr5AIc6vm7lYC+e8GW6fk8q6Pb+Q2a
4AD5MABnSuGCZnu8YDNDrzGtMathJhfhmT1QnJvZEQUVQFwHm/6H9ApBa7K+Kn9JJKNFqDSvKVXq
m8/PKO6MqBP52PDqHfUdMfc/U5NrV2PdVmx1HQ843ofR7W2jIFyKG+aSMhfZRHA9opkKv12g1q37
7mc/d5xhJjxqwY6tO8Ny7iG4fA1EUvk5P11xlZjXNJ/hGByKuYFgwKtx9cl1bpYrlD5ZkrxuU3Yi
I7GLDLlPbYmIRWmHZ/+KHGroREyh3BSGasOGq5HGHlQKFqaP7ENnKPwntPuZDourId+59Unffjnh
UUOxCwpKsgXiP0ei49YZVzG1/YnXnvc1HA8FnYGpQhA3cHAxMOb1TuYXVlBlwaUNduoiMrdwjBw+
fTIVVUXJHjO5e8tPjETd0GyKl2+feBf1Q5eE17gmJP2U81u9NaO6tzEhrm5LkR2fg79LcT42Hzlm
fh3lXcuM8QXkYQUBiQsAdnTiTwmRxL/fG23ScQWHsH3gpyZsMN4g1ItJipwCNKJj+bCFBTJtRNcr
5Tii/g7C95QzxoA5oK/QgcZqalfxtfC39iuDN2IOQBYtIiRNzzopXu6LXgQNFQCUdk4utmPK3+F5
TRp6cZ0Hu0iAElk38h16TWE50QGH0rs0kszAcrc8kKfkTDtxQ0YMyvY0hkf8eWwb23sRwfXKMPJi
mhpymHyLGek0R/lHtiMTCoJpHTYsjx4Ba3DEN9c+LINFUETFIFIpojUZZVEtmj7DoWwDqn2x0iu7
CRVMYMzFif+8KtPfX6Ag3CStVU0YRVdOjtiipOSZXJDMzbvGiUk1Z6D/RzmhhXjiFu3prk/WfShC
gs1AI7jHTZKowiejT8jOQhX00+pAchdWynK3ch9EYP6OVfu01l4LcQP9G7t7Vg+Jrviunc52xyvP
3p7wonlKdb60RowGOth9b0KbQPsdE7/cAWHy7xRVIjOq8NyGM4v6hg2vgVaRvTTcOZcrB5GMGEzk
034VmJs+nDgZYB1dlp2K3InHVgV5OzgE2IxmAusSD2JKlU9uG5N4BuvmKIkZpCP06wQtrXxKpcbT
9snovl6jTJfSzQwGKHievOKvMjr9TQzuRJdzlztC55PEUz5vPebJCC6FHtvw+1vKbAaROMxnKsc5
YCzSw5FHZMeejZaJDro5XkKd1CiYgyUbeioPV8JIY0d0EjhJRYsyPAeQsTsklv/emzi84Zq/BejQ
eBPhLBU3vckRUYzkMZ6EnHjP3zewhDl8jAuHb87AHXjiKCsMZXy7BMUQfrgHwN+l2l5VyMPjiHMI
yxpP5ceOk1x6454N90OdfIjGbIb4UM6wNR6Kn9M7QFaK5ayPL45i6ecYfWcrz6SoOYrYw4eYhL+w
yisYHqXswtGbiNDljaEM6YwT+ejuqWLGSxa5n0qfTo+sQSkrOApT3ATOWYJuJRvFT/oBoUL8S9L3
o7BbsyHJT1bK9tOyxoygFVICEkh9tYuYdPfvgFlEmppUXN11AnBkrtKVqL6ihvuP7K6HJR7rL+AZ
SaR9JBkXi9yflxhXuo90YbzddLGFCGV/r5CxpdKRrz6KtXgswWpsab1RMWpfzPv7/c+p9+ztIoXK
7t54T8beJk98KTMeu5ONTn8mImWxpY5ttP8sfiMa0K8g+kdhLBCp4spfHzGVZBfr1nuSlDnY3/48
M+7D/mHm4lRdzkLYpNcinBffRHdNWIZ1aZQ951A5MJDmGUx+07FC3yO3dI0RPtDmGNmENBJTXgLg
T/R4zeZyn16Mm0R2NOOQ1pvEg5+xXdr8UJtKkXKTW5Z9mHFNZyUx+hfsqnFFJGNhWjV9/pgJbeC+
6YBWxGkfMxh/OJIUXPbffQaxe9drUFqowLNfdzZzAAfW4bTKNmod6+wekNruaaQNHto41BWqZB33
BoWmzQexpWhDigXBRWXGNIUjTzZX93OaWarNTEBqgVMXuVaMgyDnUWSqdTox/ZRYVmzLvbBvx4yT
aj8aeAeD1XQ0oflhIjLh8MPcxq02JjdJt3vkQ3Izy4koX55kcjsoYkwYEbc6LL8GNPQdtyEwdTIa
spTTE83byx2b8XInRuc4zFRKq1fHqtJaS+F4RRMWfMyiCixWS40y1vzr6pgfeiaIguA+0dnVLpGS
pBu9ZbIejuRtUCHRLCLlUQeWbnpIKh37P0klhtUn6R4cQBKVYxk3c3zTLotfM9CGvnyyYUD5XsPh
DNfv/IYgkafxXdZ3CN+n0iWN5SoZoHGM+1XFgk87Fc87WR2nNEGg9dXkVCM10jQC3sXvUY3OKhlc
y+Z62HFhqelr+nQ32MdbVKQmNfot/62Hd2pcFpTgX0J2vZ8IdsS2iK/ArNos2W7QK2QEMNCBwCLn
HD1VRalQRmkbtS+yW9Pa/KecXiPcl6icPL7zGKKFKzBm/wyFjKKMh12iUSwsXMlxhehnAuJsCzhf
MOOCp8rZWFduDxctgf+NEP5OM64LDCPrJl6K9l5BWGprGy367sdWw+UUSVzh3CvndxvhlNJxi9z+
18BVMe+nw7DgjUpRnHIkEFAUbE2OuthgSHM+EkrePGCq5DZtdbVUvujQ5+HcA+5Xka1WM2+T6Bza
UiY6PjeHqY2KWBAvIkWZ+UzSpgRaBu0vyEtOuPgp8cSk+768gvBTGll223poByc6F+Yb2HXPW/t5
Qytdww3lMnG3B4xxVQ7jeMKS9jiUrr9FeDs/36NOkHqtrwmkCzBYNWlODGdA71Gksozwy/OUSKDt
nN9brE1ZAVuk3M8RMiNP7M/+Wo83KoinEXPWnbOkUCn/J7NBc81e506X7NvdmKeMxbXaeXKVNUEv
YLTfpmcIc2xbP0cKwdVor1fJ0sUFbcRYgP4rUGbSIuouIYkLOo5lmW/EQTmagoHaI954DXh0EkWe
YbyzlZYPfgqSMa2Cl1yEkWNJGndeeKbglg/0TJ+84nANlqH0q3WL2KyF2p0g1ihAggItq9mgSAt9
uZOhBHTCBoyj/2EXkoxG0JxGbhWFPEKdDaro0HkHyaFlrv0rF9d0hilOz7qZTm4RvcNNntK2iwD1
oWF6pz1VqNxdggRfTuQt/ZZdvF573ZJxUz5qmkg6wVH8ScPJSxRYnvGlJv3yckLvAddNYT1QauMr
TpYJgOyMNP7r0b6F7C1oBm3r5reAObJWuAk50aClHI0dZTdBBpw07+XbbKU7dBH2G3EV9CZzGBNY
vUkd4Jpd7YQhSrL1Adrhp4ZiO1ZseSn/ityyTu5790B15Qghb1K+wEl3MTT1kOl/RIiwS0vQqWRG
6jGVcXxHPRZdfDtwxfwEq8Iy+Z+HTlyt3Q/gveCcs4DNEs9zP3kigX5ppTywdbhzgcYp1LX2TPWa
Fz2fS8gNnsX+q3geoEfL6LGumpA5BE5npEg6IBY89dtWqfAISYpeZGQbIVYIy6uN1IKDNBwwM/cK
ouf/EkISMMMSOei8JK00EAQ3Gy5603OEIjNx18kfsBResrZR6y6pU6IhsN611dG6FSeEed5aKFxf
7mxaDHvoy9hoQE1TXFnA06VLR4GO3mAgu/oggh6+wnrBXIZbFJiK9I/dzojNVyEx0FS35QZe0Fez
GACVCyamMD1Pu/eIBGek0S2f5NNN6tzCKJpLKbsD99BuR+DqClF2Rzoey64XluWSdoEroiAhMfIo
dkVgKYkv5vdrkm8K4s6UrNslXfz4MRS20I0EUj4GC+CIbiYeBD+g7vG6JwXAMTy1W1NkXaZfKST0
0dVxfWNNRAs68+eEeZmu11CEnUuKQHLWMsH3KZNZPmwYl2fV60fQIMqJaV0w4cI/wub6ujyjQ+Pa
W8RimQmE/d59usOzFQb262WlO5K8UtIh5MI/+4F13fF9U+kKbD9WIadn2yMM1x7TydJZEx7qjRb3
ObWSSWGGG1PoOM8xZthv47gjioedQL/FKRhJlpBOjmJhqBMzYkG8+GRYd3448YKd7gF1dm3sBV7K
kLUNxtyix8n1xYr8rGt6nythBGM0tDEZgv/SlJtdYqAd6w4Fjs+EcPReHpaibqbcvh1oTX3hwgpQ
rgN+F2qutPqKPjC1LLiaUWdxVp4j0ifudIIpjd7yL7H9JToyiC/FuOYQcN3Y/eAtTMQ/xmBXLf1A
8WRquzpybg3mwvd2VUid3Xz4f5HrprwNIDWBFQNd2voL7lTYJU8L74A4G5IYWwTJaRbtxkncu/GM
iSwE089O2yMMWrHCC8S642ayUQXPOaP+0S6+smq0W5adV9zBoR7agWhssFn5AaWCBtGE74B5AAhA
3QCvU/MaJrRKRYXE+YRxYZkvGbF1WcV+Ws8LDyVJB2xoQAyNGGuQP0Y/Gx3/Y62M6yfKGs/AhyxT
0r5WV9jyngR1pAHRzj3R1XmNee9FpjnwhYo3jct6TtkaiAFThLqQrNQctPzXhi37SwFGjm6vQ9xD
tClDjbm2YcCbmKcm/ZEkVvnHfv6VzcY+fA1rJ9qfAlrt+e1ALnfGSxdf8k6C/WPKl6PMO3kH2c4Z
waxbyZn2H4JYbeWcQTJ1AZY9b30dCP27++X7iZwthI3GrUtff+jjnZJpxpSFGZ6yFcnSG7eFnqyX
TrV1IjHoGOU+Ei7yKQOWzpK0M0wbf3I9NkeOFgPTHCPcGwo2dlv02sBXBjC9AXXtVh2YIkPaQbJC
MoZFmt+IKNTC/jULye2OFslj/YK4G7D74KgkIkpNaAc2VRz73ctMlG3sAqltGs3Evo9VTCqdYF7I
UURyONLqpzy5t/0uuPaxARKY0fE2dH07tTMiuap7LcIRpQUT60ZvPvcGrxcp9qcsKPHDAsWL+03M
wAnaPClUZ/KR2zpfyVaETd4AwndwwAv654zRKAn6p1Ufd6QbswFKdQGesffKw+NIkNggrcs8n1eX
CSkhlBD8Xy6FZiFxzXavfw21PkQAl+isXfIzQg7IBXxShheUSxGa4GJJvKWASWDKVwA9qW8rL/7f
4Ayz0HIlGsKTJQsTfHKg33Lnt047CBuc9Gl+Z6WdG++6qSdeCYocOf3w1FOqHEkauU4s1SAHNJAO
ODoTvS9KWxihzhSu+kLdK3x0jMnjyVUyobRrlz43thNNj/POk/PA5CWPWKwaIWVcgX6Dfh25tHS0
PwSPF+0K6asDOOew/sB8bYdwEQqo2SLxzhoCG4FqAaNXemtIZAZ3rEv3KgA1GCHM98TJsuKcUOHt
f/jF/0F31HLXmvEzxXKrVPDxt12ej9UiFDx8NuLq0dG0NvN3n7t+Rx5oBZOa9SybrniygiO1/SJ0
yOmfvy19b/QS0oCRXS+LDwGyEyAsPMeOog5o8ZKkOSIXDXH2i+MOCdmQfkTgc2BsRL6WBVBgkMwC
cbKXH0fiU6JaMF8U/8V/oXnW1wB4tV/2arxi4eOSGdMTUo9VMbnjd/DmHb5gsqcuJjkbMFxkogRy
DuM4imz6LKmek1ks6dVDnc7PX1ioeh9GbywHj2goo2z5qXOI4FbsuKDW1fAWQrtjigEeBzXxy5UF
6C1WXwkDWZ13qyRY251aVELV0gASKzD9Hf1L8iuyDzEuBN7wRExYS0IyNkzp8RF5mLfFXR5n8nTy
/FoHUqU7I89/k0Pi4vs8Pa6/lUKbrYzJZymmtN/zLaTGcMebTqdSFCoanEOVZdx/7dGAUzyEO1il
1hoB6mZCXZ/fWkTqNwVKl12NxZ6J1U0WD0jgT20ss6MqDyqJRFLhnfzkenfFKeF9ymcVbwR+24qe
wTFLDZnGkQS+a6YCKS/G345AOJB5KaUQwbNktg2Uyr/tFb3XcOMFk7o+xwZQfq3Rm+bVUMUCb284
Ss7jp+0TSOJTgJ/CzZKyRUxakLFFAd2XOIdYB23HpXjeQ097Iv9D3rxdW0VMZ4/CJy7enPfXy4oV
KoVB/CA3OaCifn6UvHb6o07rwuZAaT0vsZBLCHtC6e8FXtlixZJ0Hc20PPpPLK8qKiCf8QXkxoF0
aReX4S1QwBDiglRFe2giS/yVNM15PPNgXHMp+fgOHjGfy7wq3/HKG8Q6cDdqFaiyEPt2evwGTpBl
mpFnu4P3BFztoSPHqS0qAAepJljkg9DPfBWwZg06yy8XmBnf2hiNDVUt8IxYUMkGVv+M0e6h0V+C
EXvM2RV7zAT8H8sYl8p4AovPfR4ozrheonohb+ZXN8DP42JXuzO9+rTyL8Y7O6L/TZC7vgStj/dC
kklxmnxB6od7DT29cLjCp+jkcrd4XQ4tVFUYeDpGNAOC6qf2D2cY3w2aIBzYDTOBU6ScbA9xrJzy
32cHMH20y8cStoyi7ENdLS/PCSCqFC3x04cnR4YCxIGj0okvZx9W4gj4zOwtt9Y+Zb8uPMneWr02
H5Ty1YHZz5g4iO5tx5NXF9mgbY9uBlnu9UhlYJ97tY+IDBPf/JXlKC2gAHD6eV9E/HEC3i/lcHQM
cUqjtV6C3ScMND34OhJPnQy5/08zYScyMmDJ3/+fiPM//v5rmkQJ40bJl0hWr5OOCLWBoDebuNFc
cBdGon3lBblQ2QgPdZOgfwbEhN9dxCl8QsOMER1hcBTwc07EeUBDM2px9FrM/FI4p3UyJyIXf0XZ
NARFL1qNH0Pvuw7T55m+NaMIUVHYMdLJAJ01OLog/mvM2AQHJFT2L8UFZMfhSdnSVUal11z/Mj5u
a2EI8m1HhWtryZq+Ii97V3C3owwErZtQbcj/uD9wYrGZtck/snITLECSjilTmTQEaf+HEmMktiVf
QBa4SZTBAknn1ssRiruOgOIuzcTcnQW6wh8Nu1hZbB/MtM/nUuN4cN+O2QD3kVRtZiZyjEd10a+Y
oqyrfAb6R3JdJXAkB+XB9rUHZKflYoTwt85c3GbIZeL1BYYCKk/XYn9siCz70xin6/e1Dy7BrL/0
8lZb9YVSapOwUwvYD+eltxEGVgsRuCtI3bAo57w5S3Z1Oumw+c5LZ/CDk+XCiwsxsqszgOhzkKUw
hzqrx5KSUer1t1cK/jbH5uvlY3fAdr6HDILHxnelt763qoyidLQOYE3ASHyQuVIjBm2NK3Xa4wb8
LQZOz6EWhDPCeaDMqR7J
`protect end_protected
