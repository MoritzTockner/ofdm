-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
twx+fpXsq4K9m4X8KHoAjfGNpeDel+FrFm24SX9tVzB1uYWgG1m142UJFJwNrZlyYVHu08GpqH6/
wuUr031eCxq5yt5DMKNhjPOJh5xQLEMd6M8QTZXDvlUDv05CNBc9xscleoGKedS4Sh9EQfqGMdI0
pIwyClvsxjo31nSjDfj6sL0fHlWlaUXspDElApnQMQfiQ8LaqZh2sRBgLzjWcvNDPr/ojn2uwL42
QSA2K5+AEVuR+X2t1daq4sl5NtMYNcPMrdJeUb51yfzA3WrHcnLSZFsECPSLwxt8xU4MZ9oEOk0G
mRKjSNp5seAOZSVmPjLY44wN4VmT7Ss9vUB5Aw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10336)
`protect data_block
Oqh1twQDSVsBLqY0dvfqXWp0K/1Xivm8wWlYFd9uH26qg5j3AVzNSHQ9AnBwXWPIhMXjySp3zA1L
+jTA6xxlnneIzfd3y4IuLDT5CQZFCZ0n8XKCmsVgBuZ884AIipbvAXgekfh1c9aUJ2OdUK2H77dj
UIddz0zXzaU9A+lkIIvzfrS9iXo/3FC+eF7uxVknAX/AEbz6HVbbprF2Pee6Oqo3HP/6ZXquDyoU
obQvYth2u5g5ggoEzjGfNCbPnmDTo7/xjY8pKtxJcqH8hJJDmPtdU+zzBdPQUYtvkGsnAznIkK9g
5PlFk4i0o5WCEiTpx2d3WfinXMWQ52LiQP10g+TtojkPUaCZR7nwIyUUSdX4NoVNph2MxDpzsSDE
39LoTU4Ib2i9UBn9lfdMJUih3zwUPBwrcIpfTL2ijqvpR3sVr2NzyL0Wu7b8t5A6GHq3JmKFOyAT
CMfp2wQv+Xhc13AqTVwpzDoOeNHX97rfhfWyRJicJTRSzBibDdjMmVV2hbVxj7m1ZJA83uCiMFn3
06I1F2Da6r8Zvju9/DzkCr57VD/BcNrM5lh8fnemsgVb1LUsEXrrY72eVh1/0wgzQxyrqJu6Wk8i
vLJHkigMuVA6b8wPYNnuUtzYa61oc9IvmGCMMqr/EhG+wMyaetsbmq4jhDKGn6NzdOh0clDh+ymi
JryDywHb4OwZVSgOvUwdhX44G4uIbzBnFT0uCAF0kl6Wt6yMudopL7AvUPmKfLRJND1CNfSO0o5V
HkQvazB78yQMuVYOdmYzslw/zemDq+4SsfHZvMU5o22tcpeqZzfzwXQwS7Pkj9d0yxhfK5qXpm8K
cSw7O42G8dmcW90tL9ez6oSQvyNty8LtRrajv9XQJxQg2uEaHrBb2HMf2DlfcnTG2wImPevn0d+A
Hrj0CxXMJ+w5y4tY13KCtvHodsssTs2iJ0Us7ytj3C08INQxug3GdT9QPGwOo1y7FaCRwFjgkwDm
9/JNJ4hDaalBWBOooE9bo8Uab3Hk7MdgSnWOkRsCVII+B+qedxRadMQ3SCLI2/ZVsINS8NdLS7qA
khpqrMTsDbg7aPpnBIYRFnCfZv+fIpBMdy69TjHgAPgM9ob/bKHG2b0Fact0ZMTlPurhXxCzZB+Z
dE0/F+/8EYA/JFnL+nSBryGwsdQ2KANrhD+G701A0H3mS08yxDPztkb8kIerUtM27/yCrt2mleys
SV6hFqouvs37suelNNxjzdE7fJMtDQJEjhenOlfAsiRRikOZbzc0pYvskznvDX0Rcxx1+jOP62BY
aQycPORalK6nH7vcf/6wJD5h84bnwg40jNGHu/ASw74lBc/gswA8DwXzB9fgCKg4JD3Tkp8pz3Bo
W4qkcVm89ClslgsrUkPsvpmhKsQMJgDpJvmEE58HqPWG1DL13IjuMoJvQ8PQP5xDOQwHZUpyF0R5
JvFSz7tKovikXcwIvAk8fJgbHFr51xH6s7E4YK2egXKtCgVvAQgmAonABlzDHdrEuC1+lgV0+AIp
mEF65M9o403Vl7PGxgUGcKlYJtSHMJH9P4QdRls4TsFYZ2vrQQp1QVL/nquDag+70qNewmXRbcq9
ZoXYGtj0GEd8R1k/wFyjuAGzQvHujUI82ucRZsYKuOFplUzTJf3enCbTMoF/CmdHXL9RPpZYHzjI
71A0OMiHG1clvsfCVPMyv+fb5BTqxfPGMJ4hcY7foYtX7hFWFjJOWjVb8bZiTGYkGfGgU1JATsei
rc9fxk6ielwL1p/FceWwkXs0cMw5y5/yPpcX10FKSaqFGEap3eoSewuFZlVKb2Pyxaptw/l4Hrtc
13/ko7qYMatZtEhzLjB8BUJdzvQGYEu1wlKQyb1f1gTtpP4tg4UodeLbsmF5xA2kuZQclubEzbHg
zIxfWD/8XM2jOrHQWm73bL1BTj8LEYVxuOiC/rV8TdCkmrFBd/VgSGIRP6Tmnw6MXp/WbD1r4ZWb
5sPKCE2vK7uY3TWdmN2Vz9V3X5F/NKCtG8jVMqT8i0cGJKhSYKnoVWWyWbq865xCT83kDcY4vnOH
pxQ4/iUBCpKiZNDcSpCUnWK9qtTgmBxfyChpk0giiA6wsPIjbcy4BdjLvLQioNdGS9hfChMBWT0l
BPsvr2u4AB67Xn9a0f2Znlwjlh6BJ9jxxFjjCCBJRgBFk2mrEub+PHVHj7CPNuvtP4kmTCrxJYYv
w3PH8zT86a9VQ7jMsfBNEa2Z0/oAvnddIwrvpd/+6vm2RKuz1gEY4pMgOBgjoR9Jr5uCL4l+UB4V
4fGdAwzJqSBuEODMF2q05FCsZhfkOSyczoIWV9WuXsa4zAJeK0hHZouJU3yq84LAq3VehSX5iooq
hnbCmXICvHdv5B/HMkePlaAE7aHukWeUfXUGVJh+URDnpkyYw+N6UVL+b0gIz/EHjZXcGVyZ0CEd
0oaIYQpao3hzDHEbZ1XCESMHWrZ8bUfA6gVP+/C3+K7vB8i7jOCa42P3SRlw835ugY9IhxSZLatL
7YocLKy+h6md2umahDfncz9qqFBr0m7Y/XddEBkVPEcylb44HVluZIgwsM8J2mKs2FvXMGLJ2VfF
/KVfj0DryPVcb/ojM0MmoT2pvQw4G85MkO1HSMlALRs4ju71ST6tzfQYexyBDgsH9qf7ybyP4bGZ
kMo37NMq2+W5sDtCDVTB8xxcJ65lIDlKdDmHabgjlXXihdL8FEpNE4bEhVZzUNRDEzvvno4ZNmgv
4rxAMZXUqL4E9vsFkCIJTSAsOkRr7ocnF/9kQXMhzEn5xQmKJZekDdolcJ8QtOC5gKyVbsFvi1E8
UJRxx2OsgRtWTlrwsLilq6Z4V5UDF8vLdDy+BWk7je4qiYvecZqtACqkIy98aT/kbNsh/4J32xMJ
X0ULAqTnDIBPHDkwW5g01ympne8ywW2kibj0qWHQcJnnilqNmyiffIg3fb+y0GT1fNPjF1yZpuQM
G2HntAnzBs1L6OoxukYHgnszUoXXO0oDH6vwqqKc1/4opwtV6F/T9BMoADONDXqv1ytwpJSq5IxJ
N67xdF8GotAL4xG8DeocPolHrPcziUQgjtqSA4OdamQW2BD+VOPqYwZCfFW9jXJriVfvAZIKdkZs
sOjnq+Voe+fTVEab9XaXbpsqbnaUjCekBXzUO2vSugCllcK7aKiNYZnGRvWJG1Xyrb7pf0eTTH8f
L9VQ/kDo8r44dPHGQQV4QMiHY62fBgwcwLwiYJ2ciZBnD5z4UdUCWzNt60r5UtrDW/xh3gOUJs9G
JKoWUOdGdv7Wd8BcG81CfpnqkN8m8oDt3aVovwFdoA+BNAeQuZUeJXIOcxg/mpU4pCdMG0U4anxx
2ECc3v2VKNy8WBr00SlVheFyBQsx0+VNeV7rmzweH/fQeCDLMXr4wh55Roq1WwYfsKvZu5mk3nW/
CX8UEi203g3FpixIZdAZKjCVc56BNmlUAqOHqzfvgp+nfxnZJ4ijaEIg4tiDDSHgtTj/drtVHRnb
hnyLS6RNcMhhVpmJuMQZigvGQzxwZ4z//RwRMzHT1QLfOKK6VX7BSeS1y66Tj7wXi+aWjEE7BwU6
QHIYN47kI4QrJyBOgw5LXfw9s6Skzkxn0VRXKX74ZNgc0FcA8ooCPFriHoi9DE/C1z66iXL/LRRs
FUEt5cZNgYR3caseWP3UAnRVUmRrZZP/4aurjNTwvwOuHemnKMXZgL3+kyBgqq/avRUXmW2cFHrn
YGzVF2ojdOXy2MvkoIcagWS95UMyDfeBcCjC/RzJ3eWOfJTdSJaBcrWqf0xkIUASRRiT47tiHB9n
6fiBmYFZ7nviIf4Khn0q+NfbI5NcfgXU2DDqA5l9968FijSf7tBBLBnwR9GhB1ArQpqCdWG7zRFT
P49HcK0QnlxFfgAB5xKxen8kfxTVPPZoVtEZJYnYLwCn5CEjgmkdW/pWdjsyO7HhEk43gOEHk5ZC
KDxovDQdS932A8O2GVq8EMfWq6nW7dppQ5poE9WlDUY/RkHrUNRPlIdQTPNvZ8LEAa6EwA27bR/1
px2+jGhQrN/CJIMVQzfqHjOgkwwSbMf22lLJJgNY1HLMzcn4i13H1ec2GUlP1hQeDIDeI+pOB30M
WBHKHqEFDdoMjYi53m0+oUGg3TqJsWfGpJZDrkvGYZvuYRJEkMyIjSV0DoyoFOtyBocWqDxSb8iI
pBEPuC4fGo+NsXxukq5daux6JvWtkPRbmiVbPAYFpuNGLPFDX+okwnCiNVC+2D72EIHIKoejgRaM
TEhkXLkrYx60igl1czkQbqX6jZ2U8ibBoywxZ2C2TIEqYy0X7AJ0zvE/yUaDqFf59DbkkjkM0e0L
TiCsTUdWgsEYgXA8TyrLeByPY/yplxs1aZ+CROnklFm7rYvwK51pABo81YlCJQFjyBZ7rdldswDE
1s3WbpfKusCKTGPEm5ZgGnsvEGWx5z9XQVSNcirMbKlVmknh52gpFfqQAhCZA2am39JD9qzR5Mgz
wqOAv4IzLbv8sO9P2xCVYcGQ3jgHdEwIjzLFN7d13kp/MsgeemC4GTLNn1IztUCcHuIoZSBERt9F
zdBHtjYkqZmSFo08y5+u4VwndhFeYbYWJggKM0ftxQIfQvU+Z8RFZ/3IC/dksJigWdWvtE/H1QKK
rERvTN0N9ItoQZIcUN9qfHG0QiJP/BcYbpV72vWAcDR//BMgdZItkfUiPjFY/zCYKQOjN1w4GgjY
4LBWAz1eqC/hTSp0+qFO0HaXp7Mh5fWMi3hP2Ia22fEGdhRN5BuXIb93I29/sdr+W4t9IBStMZcO
YAy1xZ0xoH+yLQT2r/0+W0nZ3OCeAy83Vvmg4jyW3JUcASjjyZN6DWEOtGkePKmCpq9BRwmVS8nQ
wN0hK8nf2J/hnWgmR56zeCBivSZp3vBTJ3MDuluaILOR6lASpXRTM/kyaWEgpBQREwNow/jda/Z3
sy3G38NIeleaEEjhBwwBDtv3tovIbRjTbIMl+hiHuTvCxgu9RszHuan6EE7EjhAvUcGIvoevmTYd
ASS19oAKuFuVSxMZBlFM6rIWYvoLAyQqI2/fMNRHGSvj5CJmBwEJd2KrRI+cv95Fyg3uVwPjokzD
m1BDLfStnkEb6XR9Oz2FOStmPmtYnE6Dk/+I2Z2DApAY8+uHgeqNz5Y3chjU6NGP2qOG1JxFsGNe
3fAk1pkI08eG3TwZPQy1B+513lvBb9kFT9FqBJZfhPTJAZGk8jpAdgR4MARc9jZXuR0hjcI1rY2X
Xg8qRSU84jcyasC47o1bJLNqvvSu/MkNF5BeKMunSyvGWkQ48txxyaBLpllkHwHCOxOnJ4bgU2iP
2xMl9ukSErX4QbUJGj5ZhqezlVaqsnTZsj9c0wF+qxvFN9TEebMwBs6PwKQwrvgZ/9d7g1wWEWNS
VWE2zflWztUW4IfJiR9xkjHqCU/4jN/RuPEhwyGtIQFfTQeaBqiLCWhySr0Yc7thHpsyFFCoJeRk
W1NDGTz+iQHqsEf/PNcJab9MJMjsyd4VcNAVBHdL5hHgjC+9aSgur4sL9uLqWsabT2PGVLKO82Yd
DZxCBMofDR+SExKuG/5C3k6MJob7KEtABdRgLnl6xiPreFhUKNjfsOrUx7J0uyb/G+DpcLhpU+rf
kS1gqtm1kt3Bkr6BDnHFnHr6YZv2fa9oWFBpPkJVfWpcKaun5Q4xlnxNdAZRHRSfU+Zf7Le8Z1Tt
ZC/7aqLk5U+awGizFCznpQYhPKyOvL7J5KJlGWZbzsYDfOgBlL0eBh7rp/MZpP0/tzdzYO6VFVpI
bo70MUiQmMhZEazTD9d71bFaPHpqq/YDqlLwb64/Nz9B5DlgmGhDEN91mj1Ky2Mu0caTX22/66Cm
968z7bVDvVfWxVmyfIMPbmrXwOKp3XvUQSXZwAAm/0pNW5rli73hAA5YLUNoFhmhItWyBQZ2BXPY
QuMV7DdsJJYwujfCwMzQgjLLkYgbRILmJyWz0lMVtfEONbGkjAEAqT9cPGps/3TabP8PCpGi5hu2
Hi6PMnDjdFKW031ZXp7iKNj1G06BY/E8pLE31SVMTlnAGrtlGcjeYp2nkqbI24vhVqkZnvRlia2q
jFZy9nFvH3N+XIuwi/dMF3Tt5smfm13QxL43cj8nJUkVLHTD04wf/CjQO1uTagTGaouRZsGu28le
9m6p13RT1nXvQcR02EdaC44mVXka1RPReqNrdNzdK0mFkYzMNA0MAVPFkdT0ACLSpB6Lp4Qlr1iE
vZCGtaULEDsExNzuhhsucVdgH8L69XhXrVi8bvD2f+TFJC9krNWILOmnLH5fxAaAwWfms+Vz8NDe
nfE30c9n5KX7lSUSQtuILEVwsBiUgU+QQEzrgxOUCq8az5JDSQkkJrMSrq69h/RVqb/rxsck3+9w
hg1wPQTWG4y7HbN/CvWbeNjlMdDTOtAqLcoA7XTqNXRiZop88h/aiaLworw+bnHDuQNjnzGIbM8q
IUgXuWSaDom90AtyBz62wmc1Zc4rH/MxsniZWTzN9B1tt8hVcKC/MmUpg/y3baPjY0r2NJmycrTj
LUc0ZbNJqqiDMyQXCHu5zx9+o9sQja5lKs4vaDLs5fGNBNlQnm3wNgrqO+SSzCAaoJvhzOfTneOq
bdeXrPbwCtadfSLdDlIbCBthn98ZUmuXDk1p8kiF+ryDhs3qI/7P7J8LyYal0BkLZF6N1V3GOcMh
Nu0ODxCyd4yRsG8ujmHWavwN/dwtdTBsvonNL0yOUb9kWD7ZMIv2naQyz8MeN2x0azFdEz5E8MIt
lmyoSwg8q2Rp3rzWcsyKHLkKT3P89CVdteSV/bzOvnJ676LK59b0kX3gJlh3+vBdtz/lqousR29b
KPpu/TCnMGg+qVKp5qJzKXkrxshMwpi884p2vHq/oliybjsfK/G7IJB2ZoyWZj/XuMPC5mc4zIPF
ZoR4SZ6DUfywiZl0uEBg+kGm8OcDmGxXhDmXnRcoo6GCLXAnKGPzJ79Fv60RTsfGw3ouVrvNmvve
Xt6T50as+IkYgCQuTlZLewiPYWCnL3YYIK42IgQlEZk4xsrvypGSQy5xbcn24x8fo1L6Ez9f5msR
r3murfM5CSEbJ+c/rtUWjqySKVlriNYcz5RJZfy09wDFZlkpQGheJfttBIFuAObRq11UgoMIlSog
DJOsko0+e8W6ywU4VZ+EUEiOPSMEpO9cr4NnuINgt9D4QcDtKJzEM1CnVRuuKkAbnINAPBWo80JL
MfK+34JSpWiG9v+QJZwUfPK4rG2fdXgkrv0G7t/SzZeGiuq69tFQ1XOd7FmYxWAI1B8ByeKGyV+x
8mf3rw7HoZZgB9gbASpEX+xKOLwL8CN23fiZkcpWAFfBj1DbDf9FMPc31sMR7HiABhlcDeaQA92Z
zRLAZuAjL5kiHqsyqGEv8lbpOrRf39ggQjYx+IkcaCROdInmGbM1zd5/1tbXOXgc4s78TCKwKHOs
pSBXz808bBMuggowpgnpWLBx5+QolweO2FslfluXaahOfMmVszFa0TC7s1z2asF9aCVz1iGSY5nv
yRCbVjGTq1YLdqHY4u7V9XFkBSgzbmOik4BX06t5MsihF1VmhTP5A5v7vxtQmCw8WCZz2AyVeaOc
P2/7TEHKoBHhxPWWNTDr3JUVnWqJNgagk0I6eIVkG/UvzKn2uas0ATlvDyZ3neDfnwmcOvCiNSjn
T9KjD7jDg7qlJHqYCw1MexQP5Gi3u6lxApAdeZE+JuxQXMfCMAc5GMBdYKdOwshn/fz2aM1mgVQk
Ka7miTpk8PtNPUMz2pad20Tu2qoq6fNFp0XG4rPMiVlcOP9hyntnf9VWrwBdh/VWEMtXQ9MYDYzT
YczilS3wtDJ+m5ueBRiu+dsdlvdxylYBd93RaUOZskUsbOX6P0bo6RQtdGmGn6M9FXGI3jRHcy++
g8aDShmpPCXdoncXYs4y7bX7QgX3rIRE3Na6VCtISFtPntTqs6NTc3NSdoIkDy7BQ447oqgXyOFl
FCog8uEcOVKIQUH/Ac25eBPtUzu0c491VaQPyEiFg7PE6i3mVVR6SxtRNrlkW6RZQwGUDVsXhxdd
253muVsmmwnbclwSWjqu3FCsdBvcZ4mrdcgPlip/OEOFoILLyQK6pzgxTYS0Xzpn7QJP8DhPVm7J
gx1+DMPLgEWsGJarmwlNS3SeWwbUzCEG7WG1cE+V4YjgW9HniqysKMUoVXDctAMiuGwmdWSQa8nM
WAQnB+MItIMWRDKM4i+RG2lLO5l+0e1kHcKhbxdMTyiT+p//8scrysqFcDeTfMPAelFJADBNVBdy
5A4/MqvDN4fl9HgIpvsagURvK1zxguxooA13cWSmIELoHkgGemiEenSPcY1ymemyk5vLY2eSjyfI
Hi6CTokbSwc0dyONiW+kYSbHnOgLUxed+XU3rq8GULGFULeeTeqlBQvU0SBQJtobT5KdmG2/6PMe
C9h7SCm5VZnbouaHc1H6gXHucN30h4CCWxSi6VZrqq4gpvb4WoMla6+Z9NKclSwNfKB6HxhD4Xou
/Y12WmO88u9hDJVJ43j0PY/Kt/IXyQ18z1J8qEospOJvqPKiBEjyO4/S2seOPUbVmgVnoh1pUkSm
JmK1GEpiB65ijubbSJ/AilXhGPDoSlyicuChJdvnjiXQ91w6300ldL2cUHr+AEgZHr+kMGK6PNus
rIgfZDHoE68f5m/XsX0d5i5vX5XONaEwtZldRcR5Vp6R8OtHk7+ck1Zd7ctovxGce1LpQ4WQhNfd
norKwkpJfahgORmFr3wQjEyigB50qnE/etUG+p/PJKd7n33kYQE1Qo4OPF4LVdOO8Y9P/2ETLfFA
S+TehlGUidVYo+hk8Esba2Emqt0RlXxDHUzxMK+JzaKGN3hpZApNPQNf/jcj29sgBZ0pB6MZszYs
zIDBu7wH4xVSBD9tcXjEbIblou5cbPWmzcl/ejoEBqVIhI4KEgvha1VfPnS/IQp4A93iS9AiZUFV
Ag0saTEQafOuWJH1cQswL4LuG4AaW6duXZYAxVWLjvmiFpAZb+mJ0EuOmjpIggW6i4uARZCF+90f
JY1L0PuRfU5JR/O4CbLSKGpy3t5yd9oPFibONbqeSVFOGSpoKFSkRd2Js9vZONJaKfP0q7MM3Cyf
PGnwjXJtsULB/Ic3P9VdgQZs5KPcrrE+RoMqmK0LIRDr4kRXzIfcjCOt6gXn0EemmHgl6RnSB31R
CCnfoNjkZaNs8URHo/C5k7hS9lg4Hr4Aw1idWddLWi+G805eDsh+SZ4prRfVcv7ilccL9RqtX8sb
cYotY3mIV9PDs9fzdJFYxkbMwb29wFyrkt4fffNVKTlIJ1Njm45Jr+SAbgLn59BAA0eD/DCluChK
Jml523x1AhbtHOEHoUX7leUvXu3FtkbuX48oMeI8mAzariJ2wLmFFiKSsOpRC8+NcuMy1iAOuXSF
YqQ1NhiTl/RmgKXPAL6FXL2EWIe2A2+2Cp8X6ikTRG5h/kfJFFKa6KiOwi9s6ob2Bb6HaD2jdo9t
uXL01V7BFuSgB4efFvqxY3yMOeT3EdOBaDN3Rjxv12uI9xio3RhNYrWHBXvAb5rmXG74jfEyTKPU
skigYzsTvOPU//GooRuQLvOaFThQjarMqcjMKEnyYj20UHe9YJgRzjN4E3APkMKN6k4+rh4GOpUn
lKa0gGTdZFMxzuSbzt5aCMjIAwc2unRiScLA3XiyWGVBXErg/cAtoEbC1LHZNM75JyFTYiqMW05e
Z7nh5LxsWLbWupCAIdIe2VbvbCQgd4D26oIC4uKUSgXgxihuL7F++DFGPuqsIywkJ/y0EdqvmeRa
ooQAU9B/3q8TRSYst1zXsAUH2uGW1Z1rYlx8BTYGX3UU6qB1ubjMuCXwnDlEurrpstA4Dg9+qV+M
v0qVR1gm337YGzhPHKanbSua+3ZploAcFaYlTAPR6qpzyWbf2E4pOvRe3ZcPxYeAzRd44yhKR+Qo
bQ8MRz7kgf0fs0RSohE1oE0qteZH0PtRubuZOXcKfQTyQwkcXIw4eS22psSAkQ0grke9RoWbA8Em
IROVrXYi+rzWr4ctiuSHfZoAyAnzviPU4/d4CBYfCJzh/KW+jdK5eb9FInOg7ZUy2BN4PWlPTZWK
xR+ZnwA95zBNdTpCyczo6VbJgJwR18GE6qrFnagZ4kTTzkShyneAnrG+CmbtSP/+m2Ho7R63+lw0
Inso6bo3x2MTTZsRvj1EDLhJGGCrMcJYd/5u4fNVwz8UDGfWsee72s1l4mAN0ZTjgwfl5WjbOIYI
gaOkH8u99lLwRsa9q94hb1XUFueNIxUJL5qM0+HCVVhpkXXRQ+lGguDSLgK2mbALcGv/d99Svfeu
RHck6+tI1nptx/AJ8/Rcb69xc99LuMWuUTXNEAHzy7QdkC+MK1Cwkw2EpIYdT8WQJzoC5kF88cOf
8izB4sqIDcbm3eUAmF/vHJO2doF6oIcg8VAXIlpInujf3mPKA0zbRC3w5MjaUi6T9cUI/wMg7NtM
RNWOQZjo47tfZ7HDz7ULWaJRnP/gcwVaCPRzaDgkgQTU9k/wzKmcPFEbBMvflRHhePF5+IB1gA2I
7ttIiSsmPF4CSKl3fRtPpVxjUjP//SFscSeSS0S3XYluUxL2YAYYo6qpZt6l8ug/zZS5QcNZsBsS
cOXCUKJ+AwYTlvr0kcsJmojG8mRGGTklptxv8+MH1ozr7fP2oz/xn+LhoeF84slTMn6DOBBTgAjc
wOqJZ/qmcf7CJN1GplDpaG5yaAPrO+SAv6ucMGYr2CAiBmbuvpEIGJvGDYS4/fHEAgdrdBEh3DZq
PGpX3kRY/kCQqIgCcNPLRniSo4S9ilmdnFfDup9lxp6ZwWPVmTxM8L3YDnYms9wxal6NGc2tvJ1+
9HGE2xA7ZmZEBv7j4FC6oNzrl9YoCQmVjFq+rpnOHXvzaQknEHlydYPXvcFY7fAwyEpouSM2jKSI
w8+JJLRNSAWjOUXbkqO0fU7gfNqatpUmO1KKFOZUNA+o6oSJMIPB2SrQsGvseA3gLCviBWiiG2YF
r+XsnsyyuKUBtVxNCkABRvcTG++LMrMrw/KL3G1vI+tTLQUC44GeKV6DpAsNtTw0KiH9xSRSGqXT
8O2in9XR9mQItC3Y1AmHi9wZudcf2wsifkq3y7E9tOZWX8XR/cI84DhDDTOq8rJ+Pv6s+YPVmmSJ
8Wrd63qCPBUatm3BzZubVqoWhFEMsj6r4+LQORyJjY5e6m5LmtwFNQbAVeLXPtrhgloOo2CEq9ow
lO4PHCX5pQ729y8VE55HR1dgsm0RkobTHr78zKeAmb4Bw3acI3irzj37LjywOPAsDUeBzrmnklnz
VvjUGyIDtRD+EX34/eJb/LCGWLaFpr5K1UMfbmHeVVPfcN3rKNR3T5r6nO5h2cel/khRWuhrNjlz
pA1xb5tmZlnMeONxJsOl9zTm6NEYDTAeWLccDHy7aAHXzdraKWfgrCqu3FHaDYlDQzZTUkdzXjoL
2NDV/FZJ2iCnqELAVuhareba9HDcHpca/AFnsN2SXUDWqIiZ7Ejwhun6zXa4g2cRtbbAjnSopjN+
L89uTkFXWzTuhyBIgpH18/sUFMAZ4/Iz1/DLGbZtA09vpqCCVZOWkbphD85Rt8coDDRGADFd5q7T
O9wr6HlCdOwQmNcZ2UGnGs+1DiXVD2REAkvqG/ddh9iA8cqNEvdratYt6kf/n7cubVb5Nq732Krn
jctgJraJSxNvRGidisvH6nXcuy9je7s+bEGA5lL49xiqrdIwB0trMR/MvcorligFZze7ELV3VZ0x
UDElrJYarfSTz0wFBic0/KeJX9XgXXSjHOUQt8HEa3h+x2D5n0n9d5FA0i2PN0qKORVYEJjrjzoS
7Y+6iawwF2w/0itpyRnC3ejLRZ7s+VVQwbhzNQyt+ZWEEAvP0X9iG3QeZohApM3qk5gLW/GJbqjI
kugGAoAEPRI5gZz/hU5HjIxBAPRC4sqk4TrrEOd9ZQ7J9J3u+erh9F/2VMQ7NdwwwqxDw1hlCAiw
p6CAAVRrB17shfEUXC5AYn8v4vEObZgACWE3E27fH9D84aKGam4ThURdh4VoThINIB1AxYOCWd9r
idQ3z+vB+ytdeamdoNnJmqYPiiafXoJyG5wPyutXWczqAxmolNChsVoz7a5xcA9xzpMTZybE7vwx
wCwMhlHb3UzPzF+NIFqrGwaiqycMC33ylAlIv7zOLEfnnOU+s2+Bvn4xVER7PMnzQjjwttqrCzS4
lOz01gseq4SGEh+LMtCv1rl2GspymmBZyVISB4wiTLOn7AcGEZ4lxu2slVmbG2URjGN9WPDANedk
fGAmMeq5uxuZagRVqbGZ2WiI9e1Sl7mUxzxfYF/I2irPNb8UFxzPyluzKH/fEXh1ChRC7SIZcS//
eJyypeO1290vnD3eDrlhGIzbb1yMmXicOKxIfdKVfBr0VIJqJw4Rdvey2pw22CIz+HNTj4CyOveQ
WHGJZp11uiDpnJiLMOrC7zKN94T4SC/osWFQ/gYqn1WublJGRPjKMo6TMmS05YAyrzD21lOL9QDD
6buJ2wIg9MG8nrBKzUwCw4VThBp3cVJwCz/Xpue4cd9C0+4q6yBvDLTUE5stDKWkS0qmvKN2W0so
RRBENOHsjxL44h6ECNyTeAZNfGK9sIqsBc3y0+xX7MkqZ6ulf2h/TtalrpLn9r/VXUlHt1djTlgg
kyvyN4fENTfQv2d6b7BhIqTh21JHrvquncPoH9wixZfz18I6EU3AbJkjXvLmXrPwNvffpq/PRtn9
e9LQGTQpqXgWRUlSFn6M9mzBrNwZ5SqULe/JhgXYyYInApjJEhbNzu8xWbZ5vATAqPRWqZLdM/a0
jE84lZce590v3JH/sdSbxz0ZeSPKwg2XHD+pnm7j+o2mCn1lviPsSIDkAfHqNxqCvGxqHJ45/z+d
e+W2yfckPa8Y/Psw4TbsG+EY5zUGDM+EQrEbtw5rlkwTFYKy0k1G2/Bfo81mLplxwtP+rhOFbV0G
WD3olaKgKmzu22f0URfoNFjcomfcA1hBqukykZEXR+qhz1PyRxpDEunxCncgBA0OUFDHbSygf37M
1MgGJ4JfQNrdthuyzB50oo0UaE8Nghefuko0oKwKdd6nxE0XJeBczrlODP6EnEcgnc6tGgXp+H7b
2OYy7JKzrRPWmI6O0WecP6k+kdFhu6gG/qM5+zptWDqOp26Amp/GgclZKdxl39KLTvxlajwb7lc9
b/kOkAfUkPW28Qpp96M2j1xDHxSBgdLkF4SSf2rCMl2JTnpFdvnMJwCx4ydKNXDnChnsGnR7fRPy
r1K00LZCdOsJgUWXelGrFJIYhZYVKfGI+w2EbzivhmQt4pvA5JAJ5IQXpL0qu7lMYRPuu1sI21E0
XRRdQN3406ZVb9N7rUclMRbs0LeRweMZN9dHtdtJeLWDNFOqalPP6Dss3pDCRnyPVxc2F1RM9sz3
QsWk2x0DkapUYlQ94GGhcS+A/eDNAIJXLJjy5Brfysx/2Y1qQjIWKeHrrWtDtF75coigCppoBL6R
AODhThPY0S73k3U1ymQuTCXxQZ8CgWutX93vqQazQwn8+fCBm1paEQy4kJxojhmmR39j9qSoR8q2
TnH9Pq85tfGzeI91Gj+y9WmFVuAyorS7ywglp19CBBAk7JprDJ8PEoyUEPPhoV1+MFZWxCv/hWgX
jBjErZKPGJYGIMnKX6MpaqqTAot+qOVFBkTGsNOScwlX4JdNX9EcKjk7kCIpc6S+z9ONFJt7GvQu
c7vVXDW/HBDpsg4grTb9iGhU1Q==
`protect end_protected
