-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
kKyIW7r4Z6d5l8kw+Juz0BrTy0naQpxxSOIvNkCEkxSVf+EmcGwCIMZ0BR5WC+9Vwj3iaR2S3rpJ
no1LTA5gnrZXsNo9ncwPYhq+5OSCVk2YFkBVinFfLAvpPFtu70wldc/6T6+bJqdUge1MDtoecPFA
nOFfSr9JRjoc7XdZjfP4FV7wRGiS2QQXSzJWkylmO+E5IfBPO7MMFU113udSASHr8yQ5skzuqotV
KNr9mL16eBMvjhvF0b4bcy5hpCZC8I03wfeadOP1i7AyPj9Xsmd41LlhS8c4zzIU+hFQ8ZakpH73
px2RIYZOC6bLP5q4VRE+zhMDyJl/wOYpYPhVAA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24768)
`protect data_block
nMBQfdWM0imNHcWSU61EQ5XkWbV8B4+8cZwpU8Fj2ydIH67ylTwm/frLka3llG8EzsMxKtZAxVmL
VYMv8vsN27Cue8ajR5tNeWIFCRkmP8aefYuiZNStCBfTOZVpboJqsHUo4UJK8tpvkN83wK6qgqO6
N1qo8kMFPvckPHOdqLtL/M+N4kPGLzzqRjyp0l2RvJsrAq9Y8QB/8oALEMnvwBZY4e6zc7myC9Gl
EiFcaPTaMVGQezSBfQEkZ2+5QoWT1W9n3q0eTvWEI+E3HmCMLl7L+Ze1Zc87OVu6RcIVTRG3xir8
8/+D7iGD9VQPyLqsmSgemW9u58XWoHQRv7hk2it3QRHruEpy9CSPMjEKjqzosBGp4dnG7pQ1a3nJ
fO0uzbd8/TPjVfw8TXTKkBPJqMFP77ye7bhO3TqGU8a7kF10MtW5wWNztD1asdxLI+WeO8k+I7kd
h/uRKxydcsRrJKmd/8yu1uelVKPTSVG1f94NyypC2jZLJASI9r+STmxR1qtNLrlFhoODnaa3GfCh
aSQ1Ij/z7pCF9BX7Id6A3cDHdz0w7gC1HfhVM59b6+JBwpghSACLQkpfb0ckBj1QjTQJ2MVf96Ai
nsR58SJYcYa+Db4bdCn08WUb4KnD+6VyhV4E7mdG51Gh5/eZnjb/TJEXd9mUOFDMIgL9u44Cjo+U
EL6kMwI3oCHnu+ZShYx86pQLgXOMjEWpTRiFAjZZ7+cNPd4G31DhIcuxnshtyLbAbA4MROrPOfMm
cUnoKVurVVLA2ZOYnYPWfaFErapwSqlbA6w6e4AAQdiIupXf/p2bgzXWXzZzw26wClo4gNx77UrF
PHTC06wGUvOVo6JWzLjdYiETR6mxsnV8xNv02q4ZTn0HCzwiVt3pUl8ZPB4WTStFBB/tokH8J/pO
BLQ3QFkuLhO2ns0goPwN5xeyz26gATcsyjmsLSslLtqztDmXvbQ9XVrXbJAF4PkDg5raC8gm4hwL
paBj88heIOWOqUpR/e21KaMP+grcuqGhECKFohQ1k95vIqY+wIgxa9BA3JAibpbd/Q+ClZngfP2t
8CJfLg69EYbICdNVHmaBYdY3PsP15xlPunGufdW/qvtJTfKIpOKpYU2gKD4aBLkoK7OBATChI3eJ
psDkG4bzJKkXMXeVzFXTWrU7PDH+YQgotZ9WG1STi57lo+GS95F2LwW/tPNroGmpn/h3ZPEvi0M5
UpaKC3mP1AaLMbMjXPfsteUam44FmI2OUSRjrCiihuIC5nK59U+Wk3W6nHQ1v4CvtCPl5EdbOnMD
J3pp4lyvTD2T6BWY5p6Tx2+Y0AVc4rKz7elB3h9tuUU5IK/v5TGFqGTanik4Oh4ekrzuBVWjQVEd
88DGix/8PIB2mMNzq1PGRD+IYtak7iwOwW9KRyPRDsAkCG8JlSMZaAqdYy8BwZreXBwlE1BaAtqO
t597wdEzRw7ipYQIC5kqktFEVMvMqubt2gFxXQlto01HOk7J9ROA+vL8k9xfL7vtsMrPDIWiod/l
AbggGzpTtdC/sdjkK1VUNtvRkoQxKmdMEB3T7gtqy7UoI2Yg2pQyr/ymO8/XxXjyPg3EnQL1X7G6
IuZErTMvzZ8VMctGZEc863brebWGOLOu/FRgrlJSdq4wz8zr2oItnyC36tBcC+g4sJEJ9YtDEqjT
o8HEf+GdLo0sERzNGqGxCs6OzxShIK/xgxoQ9wIhwVr2BWqpqHQiL+4QAkKQUuq3SN57qlXUXnnO
UAtHrHEq9kVl7F/Cj2KkxzpTJa3hJEck56EBrrlcXKvN1GOFmF6pl5uB+bzbqDW/p8SRRe2AJ8Us
fyhugNRgjMWj3OeCgW5hbKObK9/q7x7uAKBj9c+DvLC68wnJf9p2mFPOnOnc2Q4qVaYvMaRAJLBY
ioNWErrk58yMtHmdgJW8UHhOxFFnTd4gAhbAf+OSZIxwb4iMG+xvwKCbLDyq/JXdEgCtmGhm4T1C
QYkSCwHvKeqoTlobwiKCc6l/wEHKsk7dqMFeoT7sZuD7v6pscHJ9RHoWmhzpObwu8AVmwbMKe2h2
PBWSRD1vTg2Btrb73lkawqaFxB3PVGozt/AVejHK0PtTe9IXx/Krv0d6rXibQJJj3SvPzhwVL/P9
YRByJx+Bo9sOwNFjf5J+dTPSGrL2aZFKjkPXdLF7eUTq/g4eCqjLyRrO/4S+GkFgK1JfcMLt9zTt
ZokWLru+rChnXt6sY9+9TZw42Mu1NWRx6TFVYrs5WNopaSsfA5ZrilH4s50WowH1xd4WKGSInrhy
otV1afQ2LP+U3nnutAeqL0CKwP1kuFaxu5EEnL+UPiUkRw/ulAg2SxcGwm6lFpIpUlmFvRzQGuSV
4nrvA6zL/NyeEVdyeyuyUan1LDHc5gPhMvwo7awoYDnHYjPCYE/3x46dyBUjio/mBhmzMK/kGJ+T
39l2ts/g7jFeuQWI1KeBuN7wbNCzEBat6YdV5ICQyjqktg1Wm08ddaBiAx3fnNqhbwb2c43faKp5
U1iG/c0b4f4luanKb4UySasyaWLFXLeQAHcSDVq9C6J34YPQ/fTJHH8nnDjvLR29DhyKtAe2xD2W
QZGHpJT9Q6koxbAPTc4WuYm7jgxd2j4a8DN4DMTElfhSN44bo9aLvB8Rzs8P9lt3E7H0IDpn4cZN
43nbd1ag6HegtNb1cF0Msp1hoL9+Y7CqwrwUTadV7b33kynVPtaUHItzKMXBfb1h9o+rbBww/Ab1
zscC4vHT/M3Fq8vg7MSC+HauNtLpOfmXJNtILgMUv63lk+SP4+4cPJvBGJEyLLkJ9g+/eFElnLFG
kXsXHIl3MH3vaV48gWlA/RaIKHN8y0Yjb/P1svWdBzSzbu4YQhWllan5Gc51VE9UclPVBjrygZrA
FQlyHgLB+zqzeM2sFLAjvxzdIthhAPXvaLrLdQ7Dur2BcjmbcJHpc9I+gXnGE8MHWXg4e2t4kus0
UVV4Cp8OR3JqOchCrfQiY/01jpQY5nPS/FKkoK/fu2hRJPYFnbl7YmkJjkW+LwmuNOYi9QcmTEaG
Edn255D/79jQsRczE2YKtjJUswq4be773OkG9i2a/GDZRqXqT0lXVbRmPlIcH0x9NpUivTeVGDIG
yEhF3fRGpCHbZVOIuUeNbuFeuOhK18OFY96lP61mQC1Sgdxue0qdlLC7QOxFOES5MHM55akNAneE
W3nsBDktjEVLVKawaVOptCBXjTeK0neEkl8/KpzE0nOvg85yLTL0uQDm8H/1trLGO8o9PmdVuBUG
tcu96XkRy5aL5MHLJi6mNVhXGH0KkJLgzmwGCLaEubclI8zry7fZ3ur9i72eEti9yIHf42+eSrsr
CKbyQF4WOgZv/UG5ThPNLPgTg5BuOq0NbbZ52bnCZiabfzVOU/hKeFqxw4C2EXW4oTeFmkwBKTwX
S7kmG3vRXIdFxglYrrieW55QlicEm6bSC2l0M3AIF3J4X23urv23qtERtoUQEcRLI6EFLAXJekOr
je2MaI0WADHFEcebTwLxNnSEy3arlX77A1+4BxoP2GkOB2lJNunw514myB3nmGgXPlc3cJ9UcDc8
VwpIWBCOMJmwanQUMWF37lh1E3iNkmn72tWY5uX3vwuuHY4hPe/7nU+fH+m1d5aAveWR1XnimElh
MI/zqX+kf+J6ol84ULZZabpHjzFI5nYwZqsIWYL7ysVp66vYOIF//UdTTfuV6JUzMtNibprXgWQo
BRaqLQz9wUvfJH4x7hauiNp359xMm9cTEepiTOpWu6NZr1AIv+qSCmO/q82ZUg4dySGecDGJrMpv
mUnYn16QRnYN62PvI4SlLAhvPB1mMRHE9X+ZhGICXU7/p3GnJfclEghK+Aikp0xp2xAzyeoecwZW
6lufzv2scM1e2GG90fUD1VmycNW6DJZm59OBjol1lfnn0JQqxaVRW61UZTw1b50WH9xFGZycPCJo
1lYUSbGUMfXfpDHAXrytCRLc/1BJLq/O5g3GLuSbXeNSn+YLOGfZtoFPjRGuWhFlPf9/ftmBnNHQ
RD+TrXcEANfZGPG4wTEnHGiZ6oFwo8LndKg1B7kbcNKKyRdQ+sThTfXP8YR1mOTU3QaQLh5RepDw
SUzhB42X3W77KtJqEVSrIaaemX8kNG+CrFUeYeU+JBATmfVlIVCIUhNJIfmHpy4pHt264pAK72q/
/nwkVgODIwVes/v0n6QVvRfu/Xk57RzPwRkUENvc8hM22NgLa11llBk/1QJwT5iZgTJi5svfe9Rh
1acvW2qOT5WZV/916nJXNq4rQDVRp/TPs66V3pE3amSbF7sRny/U8wcktl0jdMveQhGjBhqaEdB4
ddLwKbiVdosaVeybtzUPHqDuuw22Dx8az1H/stP+VGp7iZGOnb1wAOA2A7LlfN59jX91uPHU/Rcx
HvJ7vwRRFh+Ica2BzYp0JiRZDY9CbdSPZXGVAnyd+w1FTJ+vSFMnlZSHkwn3Isk+rBnI51RfYg7r
f67tPGR0L1kOZU8hW1rYeK3/ulPVM0CtH8qiIDPP8npjSn6SiJbu847JU36rXfTdEpbM1S8/c/Hl
ZpxvoaK3FM8qN1Io0E65/UGn1MaZiFXhMuMcsnV1NlKKVsbOvq6PcPxSDhAblati9AZ/YCBTb/Hi
gYyNlZ9cDpZ5958SwKufcAtHPDU79kjSijEMtHNOcPQJUuejlDIIQAiVAhEMNI0iYMR3v4wzCQ0g
HvP9ZQLavUjeMI7ZWorqaDSgBdiScd1MEW+3WrxhS6jj5fBvv8J9SAT3c17gpu9yx1ZkpGXBV5t9
EUeiDm2B+ZwwLEUZE8qtc0a9rYildLUqgVeA/GPJ6FzUGue2sTvAstARW5TSsTbOuuBr2g0hhjcq
G9r47KyisxRGP0wC27NsZgqdHho9XoJH427tVN2ALCZVbH9WbsCN97JqXXKunHGkeaYaygzypJL9
M7iVKBFlBJ1Mp0JbQRGDKKyr7/f9do/OYxWtG2vNeIusnCDWcZDj54tKT7HabB5es8uPPx781CzS
6wIClz9mPDyUnBp+rdcXht2iEWaBVrvy5PDrvFsFIRjG+Q/gR1WocA6h0l0I4lZz6cTL37G2xplj
b9YBiQ61Ym4BE4FmDzBg2iKz29s5W6iFz4JzBYRUYoFW+6JxiPtIPrOyXIf5ZzyVPrV2gbdAE27B
gB/iABkyiA3A2nzL6wRTiB6JGBbVA2Wl6LE6ibgRBiQaET+T3QThcg37ZYWAJWAq/DuNoLwNazU0
zgoh6JK8ZpE2eZCfMXpr2C36rOymYxMvxFCzEatKaljmQQoLjWLfowZw6IqB41Mc5rMTm4oc8xA7
VxpfcO5GOG6BZq+pjTfoG0Txg0j6/XRVEY4DTqoC2FDuDIJYrJLIVWn4Am7dCFgFfSXtt2qURefw
Q9YzuwWFt2QDwsnNPy5Y7wgdaD+eEKEkUJulCFRfryDOP/dC8P/k3VR0zWNrYL/19j8UKAuGN+VG
xBzAJtiiZ9mGBQkjl4OHCCwMvccDL2nmoqSQy7bmjA6R5Ot+n9Rqs/5FAXLUUr5UVb22C4MEI+of
8A/1nFgx7ZE5KrTDhCYkRqZau+Y6lLOIesCD5utKrCJzWoCumELTm45/GjJno++CQINCaSDnvR0c
P5p9X/9lgMkSW4LlWyYfCJqfGk9l7g2vWcgi9V3iQpq9Q/QjJkaMpPiU16GOlDfPVg5/Si0U177G
nz+zd+CMW+sgoru+4Kgrbf1t+01qoJstN6LyJ+/JP154b1Z0heaxddXzGtKhnxt2owe+9l4NMi5W
F5pr680r+DQWxilLIc+13sHK7spdVbBGwbvhqZcOLndKhgnG+dN28EBUmodVHM86nzPLVFujV7WM
EEiKmgikBG2wwtV8HgDIyxuDuXLHCYlSbGDmlhcoyrSO/fwSECTQ8JiJ4nptLui9AJ+3o2v/Lr9M
4XR5PPil1h1RK+61acFg2tneswgequ/2QijeOqtZrWSxPdvKqKDS90YEnGBAWff9ROltc05PYrXl
Xb8WmVYSh+/h64uLSadG4/IPZceSU1seDDFUmZjUbNSd2ZOQETj/7Tqgs28dE5CPSjH960/ANy8M
XkANp+1NggELMWjHbTFLN+9JEZ0g/3IBNnZhsHK1/Bb/jFkXOKjtTV9DQ27Ew8UjT+N/QP44TrAB
Qfm6UH8UrP5/QMZILUJWfsruHzrd1py/3k13lLva2LJ6vNAxGhUCIiRIuMBboxdicHIy1T45p0Cf
yKhsK3tGrrsdUSa9MEG5NVlbhmnjV65uE4NKVA/lYul8wQGDxVmRE2qlT9LWqKTnalENmTUg7Pf5
EjAUwyB1xNkchLZhwf7w9DSmIVzpK5LgfS8wkO000W4flTHTKxKJtk1e5eBrmlqDFfjVx/OIRw9w
7QM0bfs8JfnLbtcezpu+CqCZ6xaYWaZjbHf0SoDLdHaZvidGmubAv/eOmLGHLW1u12AFallulL43
V1Vty7yk9bo9MkLqNYJmdSKC1qGscY7AIRZrUnRLOSiDQDsm6wxBZD9drHal0mpffow4nwqAiISU
aqKeIh7br8ImfdVHi8mEDXGS4swcW79eXz/UA27rehctuHGiYMwjBA1+4c8VtyyzGb77MR9iVcMP
EsnZwoVoSc26qA2Uvz7hfQxzh4vWaMSCd/6JDkSXMlOkAJI/m8HqBn/Zm7pl02izkMGmU3V8zd5S
4UIEjQQqu+5grh+S24X4fK8jTQijlf922bKRg1PTpaB1pIWqPAl+eWnvpimDc97/6F14u5WpYAXn
K82E09SB7EgPArt6jLvMesAq7bMJeQG17iaz3pAhJlWABHx6mDeWhWJuCNelE/ND219qc73QKZAe
2krMipE3gPMJxz9F7SbGI5oxFqVYoB5Q40utiyyOhJTzM7eQdK/G0kj/WqPFGe7ptvb9NFWVC81r
x7gTpOI9+M4YeLFxAJ4foiehmybnHCgd98OLc6Ye2YIBTqlpjM7DAT1MaS6pOsj/6zgIKN00CO6M
C2YZ/pX531tIVXYGuBBoIz0+PMORZtYglKr+pWWlhVPV8yLjqSoxYUqOolNaMJigECqx2wLttQwF
0HS+mbhM6LnovgMYKwJ79lVp+XlZSONrl97dt5nlvmL9O86tlGsuNRy3U2sMc72gHAr5bV/95St5
bSvFZesvWpIPouNLdvB1uf+tFYIebtr8zCHYU6e55wlXWpenXfKSHIEw8v8d2l/ri3/QYV74kejc
Hbgw1U9eZJef/jmm7eyj1DK8hpkFhKS3gT9iZVtWDMfiJe+Ogol73r8G73hOhApp3xa70WO+MQv/
MvAZPJneT8tashTykXRtNY6O1GXyKowMRXhpbp3ErOUHBj4d+cJTb00z7NywMkg3vvxHk7p/n1os
NwBFCz5HQRR9xh+URs06HCv8JKfzboKXpHQHrBRoEvyI2paqLuFt1srYiT7LRlYAIROk39Q9FoxK
JoE/FTLYEcJ96fdxG7/Eo++MvUvKqA0FLcZ6vUOeKRkKA41oT49QPLmou1tv7r/Ugxiyl4q0TDBB
hTnTdhZlVaSrmYay1JEbCpv1QlY7B6IglixctCvHyHpLAcxBIW8Z6XNyEbrqkw5sZqw8c+paOmM7
3Trdjs3iO1oYJXFGe7qwq6WOXzdVr65dm7TNL5fyH8Ury8wPAC7aLAwcl527QdEfxB4CcX9aDzC1
2MSSQtxGHf36XNGjF523LIrJhKHpRV17MRtzy3rFmNsm6lMNvxckSpc9nRxqaXBc6V03r3326bzt
zSSusXnRsDcPDZIl2ghTxkLWmwaro0HvMENSXK0hyluk3D6w3O0AOqIfgkBqi6laMZ6Z6HMFV6tE
cOL3ktx2cGs/x9tS8KPbobnKbQ1xkYr7bZY4TTDwYn9IGK+kF4b5xhloc/wyiDR0CvYTg6bjvYZL
9iALXJZdMhECwY1qDhXyzvWgWGUItmMsTscqb1HQmVYPsKOYoUec5D8kWu9sqbMPs6gZyZ8TnQIz
I8zlppoLF0IulpxbT+EU2Ofxt0P33Xw3/Ki3R2hDhC7X5K4SmRbmwPC2F7jWj27p9uU3YyoPAJjO
jsMk2fHZG8e8EjSmFi75wqQoXrbaGYOAWTbh0LrFikKL3EL5toNY5JtaRVK4E+NbBunqj1S+3Pwg
k6oBKOTlHh9G548oFIBGfMt2paKmnFJwktIFsqRCsTwQ+L/mwTjCUJlsZV7ysg9+VqbunLOuw+eu
K6rBOTqedZnFY/ex5/zoOVIK0Xot9SBFpeoCFNAyMhomqk8t2AibnVnFMCk0IF9uDmaTGojwtmx3
ykjHjTvR3LnlTOzlnPthrT52Wkh+xubOfZycmuSzOzJYtDUM/NFJ3hqmY0lXNXbDJrFGJRdEI+G4
ZQzLAHrNbD/uHmkNfH3UdmnoirQxMEafH5EwmBcelDQbRVNvK6WoOZkwBXH0AyTGQQsuOYM3qGrs
fu/RjZQ01kOV6GWyu4VWazAXiiRv64p7siTB/MgQYkQsK3XxQ5sNPHpewzOJGA0TSuTTDl7cRiau
ho68CKGSCtpSECWUBq6GmJqkt37T98A6mj/QeRREEIDyAJeyXa2RKhZesCVwjc+JTA4QDTlieNN8
RkRQSjNOXaQ4OYGiWDtFKMnpNy9bYXrtSNdjE8d7vKzlX4elegMNeFzPNW+kPs0s3l05l88t5zj6
MwsGneve0Ml80w3Ho9FIzMSx4F+c+4mwXzA0an9dhEbeJO83pBEpKcLqJ2WoCo/ePfZDSdiRtsR4
MWw176NTbosi1Vt3btrvmmWefyY5s8PZ2IAHx3zlQL5kY/de7UM3kUMuye6qodV3RKanKLIiNfxy
+hr603pojqqsmjQVWsmp1cI78horDbtv1cY8AJ/qAEjRAw30w9MF8oJ+dxO6E6gDkoRyHnSM4UWE
KOPtHccQOOX957tFaRxsVOS/zjtbhkXMESu0uOih4Rcoi4zbMdD8RZUZAM/B7gWC/xAsJeGvXkgm
na8FmT2ASRYGoZBW2cVHiuPOy3qrsenxnW5LXxe/VwaMicBsXM4NnuEDDhmsPF/5gpNC+GKygjs2
wgqo3Wwad2GVUAdEJNjzaykdnKh5sNqAFkjC/mMRg++wO/oL+KosNhzADE22VtVfONJ7ScvDEYfz
/aytrSfxXdYIm6DSaC8YpwPQVQqv0eq17mQlXDAndBg0BZ8SZKxxe93VqzW5dQBqU8iq7l8XDwBM
XDCa5ivxyw6rdrJZrwdJpPuTJn/Qh6TO4wJaRadyDtlyIDlwhtoawMYGOgr1n3t+7fg8iH9dhmu0
FLUHdL7t+feaDQ0exSq7M7A5DEnoFrI4Pb1gZ277ngKYxcZJLM33Cg4aQhz8llmOF20GORhamb6P
2Ca6s1QDKBEFJCUujcLvXOwRBm8Bb4yLssbluGExB5iOMUCD8RdxUmMzWbBLGbJ7gDBqCXp6pM2H
07ctonijGV2DlISM3jPdMyfInzIaEdciiZRcF4TCRHBMI44Atfz9a0r98mpuQxNIsiN/18/4R6+U
gCYYjzi/GXxP6CjzZZZf6MqxFjbWhp+QBo8ML29lvIy4iNDwIh++/rXpsL83lJHowHSIiBFiuQZK
qOeQEF+OOYVVQwGhFiIPmo9YKYO6QFnDjcMSPVkXvhK2MgLdk+1xqfjJzkWqWcCu9IDK9qMdVOCF
tQeyKMz45eUGiWLJBDLKAEUOEEQ3uRuSdCMa4ePwb//JjnCE7N/pN6cGBR9fOmX8KelXAyJOyYoz
oihKLGUeUfwZVTh3B4qkWMo+sDrbITQjlHOtBw3h3BsGFAJiZ5Aw+9SLMUG70ddhKNE2lJ342tGN
1wvgLQIcuAGla6hSCeNEm/C7vupk5LnPXSA+TsYed0AnqELd65gfFPnCvC2NsHvXVM59CK2Jmejl
jMAH68TizbumkabsJla91lEFnsdmkJsdSU855a1DP3NH/p5irrFBhAiOz8B1eDKK6psCeQQcPYoz
Ts04KuGLwT+OBRKHoMZXGCtpZm73oOj8obHpktZK150c3gGUlwn4PTivCcRxGRFDvDSlC0/XfRGs
B1qxcmiXGyexlrnXkul/P1xeBHWxQ78S4s/C6pt5FuC/9OKfE4k01Y5Ylsh3Nr/ULvKgJ54Hj1ue
jrF82ILkrGjBXDLRBgG9m8RKUdoPq9VysRKCq45VP8nIccHlQiXMwW64FBqjolbtsBQwqiiuhkV+
UUgH34I3dBQsuhUG9AAx6NpI7yEMdAVOLs4f9HR61Oa2rrlHZmFCO8N2iHxbNBsoCMKJZulKcC4r
HzCoEMlU7/cTO5gF60P5bV1IL0x03zyr7Wpb6htoymVZMeWE0H4al0Uigigb928AVPqkM6GQa9XB
Jg8kmSWBFMvVNmO1fK/DpIg3R1y0zOKhkHuPCOBN5YNtODMXuRnneERPIf+W9LN71C++sv4TVBMw
CpKjg1FjBgkiLUAB2+oRwX2wnE0TMEyLzHfH+YZbHOvT+ytHekRAySYM7RRzS2w1jsZxssV20W57
M29ltWNfuaH6tYTAoljXKQjWKwFEizeLaSGq63sRO2QAt33ylUddCpbDopJRkhrsS2Wf8HN4RPW3
Hc4Nc2q/Ombfy97clJoTW0z9Jt73WD+UrPMvSFl+W0bRGWf1GtEcbyjeiwoSeWwNqcId1acco90O
t5CW9RY+XEfS0ZpC0NWNthZ49oZSiEOt6uJYYJ8kmKE3g6UQuon07+UMHXkjHb/1ysmtpTmkJd71
6gbUb3Z8lV0CrDNPq6Y0kJGOQ2lL81lIFUnvQts/MxRLoAkhqiq0BXUVyEgCqP8cK5oZi9u8L3Ny
D1XzYQWv682M/5dT1GEq6/AYg9jRdrIPaYlD9Y4FdhAmYNjujTA/EkA2WCfav/S0J37SxyW8T5Vg
pcGS2U2ntIYEGqpzUIZUA8HENio89Or4posHlWmpUN9QzVNzvaOtdlbS4UQRikDP3+o5oOnRjJ6y
5ooMZHUwxK3ui6VR8rnx3OlYLUwAEyyrkhifb3rMunHPtCUwcOB9u5qWQ1nTtuqVw1XiuZkQE4JF
ENQccFHl5yOBcf9QcjoqHacEs3BjsGSqG8/VTojQb/5/SOGHcmaN+OFsqBqEJDaw6tQ2G0mDaoj4
7IRwoq0izf4R2ulx6lsMWzTJnDKXP2oQzCoW2O57soBkJH33ZNI/VB1O9m6h3YGkLAh/w8ryetCL
93vv97ijpx13aHZg1rfmLr1gJt2FLTyy48a2V/4uWUY7SMEJ99mrlmUrQW32U7wrHw4kXcNyPRUo
VWjft3Yqyck5JCa61nOl5RCUnrUpbWQ9a3e388Y2N1zVDs7dlQa0ABdb/LZIyJkyDttIzlkPx17d
Ep6aJXN75vdHyMPJOTaIbvKYVw52Q3JNfMM/BoA9mwpXbNJbhFlWX6bORY9tRweOwWWhVW2gRzEs
GTtEHSbPpYTMwvpo5NqWVD7D6v9cUa+Y3Q0+v0CGPzILRQkgnvULYYMUUx/R8YqMCOx/M6HPwphU
xMyNTd35ujzrZmf8DL8DtSd4jBv340Y0dhmqhNZxThL2HM+6zU5d3XIzxO8mmiu53KxLBqsB02c7
964AS+m0VoNqK4+4AHrBDZmEKZJfXdVRjZ1EFjZ8Ghwjxsj94RneF+/gQr9KhxN7zGP2wPk1aXVT
ozB5xq3beo2HpyhhpGQi1XDIytgtS8Vwdsp0X4ttyc351thdbxnDGeS8RodUYiV5sGcZ/J6hn1iR
4jPJrGllF6Cw7VOXj5uYgSmzomshIFAXRgwdcZr/R4AX79gDD7L91Mo1MBGTbDkql5LuQoFGazbI
+ftcJ9O3aD5/7dVELRFlMMsMe4rPSldkCF0az6vlwAVLnEzIHPpuZ87ppcAVeoqOOKdEvsE6APh2
HecV8ahnIMNX8jALK/vCaUkZ2t9mBb/OvyWQaj2ijR0Wfp3akRgRRN38D0+T6vGhLdJ6VYv/QLq1
gtC/0kB9YP11SmPXA1KuYjSTs9uIytgKdx1K6O2atOirXY8YQBIGnK1//HE4QIjxfwCn1SVrJeyE
dWXlOcZhmiw1Jyud6fFIvZdlP5AP5HgCwNZ9utNyeUbPT+zEVETuf8Am9XcLwm56ey+6wKzJlsZ7
arlh3kpmAOoUcIj7VOxEX/Lf2wakKnlYAxh8IfDGeqiIJFdNp38/6z+0PtmyduH3QCcsK3lwA+if
omhqtYPLNKJS1kLWfD2/LxoPVrPaLuoFlVZnPvQ9xIYjI8/XfdshgvtWvIDSFbIQ2395GXJt3gpV
H8vF5ImPGxP0mA7YNjASwY6QdOxqnxWRj5OuHW+FP6C63eF9UDZGRijf2AKXc29go2FDz+GPITi0
rpZPV04922HB4riNzLIWp55dnFV1E5Zra6LJOl90bYBzK4Kj1tZt/yLsaGnvwZMIqOomCXtGzFYP
hm8n3W/yVltcCwQk3/a41m/hs1cW31m9Zpv/HsksgDIjJK7oRX11hgsRIudzL9/w2quZZbJACoXm
QtjBd5uUrR0BSgiegaBLVP20TfB3KMLPh5EWBwmv4grjaJAX6w46zBNUblrJP54TxiI420s6Jkou
EE4CD1NDMvXZf6bH3giODPyiZuOC1cI6vUIPbah5himj2D7qYFiERvGTwYxt3k9l30q7F25oi+Rw
3v86S7TITakDBz5XcLN1Rg6be0PmLu0TFaNPl0Vjya8eibOVjdMBJdFdabINYhVFra79G17N0rwJ
fAImuOIn/fEyPZvf2NihGJf3w3UrIGsy/VuXBQVI5ctLCa/Z+do35gwlQ5+qTkEnVNs7utDrVtMv
BT+O3F4op8OUKkv2NI63D6oBNy6890UF4CcOsSiZrfRT2u+JrW75QowtZOH0EC44kSglOmvJMYaM
Ozc7RRIHXQu45LiFCb/Oi3sQWqEJkDij9D4e+at5uF3eQJ1o34SEGW1yF9jaqjf0TjQ6sR09hPrm
za+RHLrk68HDetPsb9tQ5bfygk997V76QxjFhF+ZRJQdlFX5LA+0j/hi1RDfy03fI6Y8ghpNPRcB
ZsvVoEyAkf30e6o+u4j+S78Sm1AYOxOABOTTN31y/0jpWIbW3gpQIkJqw7JBCVirv9ceeE773Km4
28Pat3UqY7gTW7rBr1jdLO7piN0YSLmytnhWc3XLWbeCP48ZMo4jW0eKUzZ4LGTtnHIcZdERlBVA
cn6D2hTqknUyWocFXX7cRhwHTYRKYKLiR/WwuIYazljL2zMdnFCfnWcqKo8iuli8WLlDw7NyToRQ
YiK4CsI0DaHGANZV0tZ6jRXhzv+Wd8IL88sU2aCnode4OTaWToJ41Y4VJ5y0GFph6vuIZU6ENmUH
EO2L/6xHhm+ym3U5h5QuzLyd9hQhJ1Fvk4U5lwGlz+8duF1MaK0WduE84sOlhTIIQ/kvoHp4ExiP
823sC9aPNXEpOPYk8MODjqHHyQEOKW8mb3oHjiqfvG/aANgrOoZoBjnMJ/RNqZs9/5djJw0gTBMI
py0CFxhu+Bnl5Mtn9flkaaJ1MFtYfHj82c2i8snavs98F4Iaqo5Qo+/fSiYCqm2/a++YU9QwlRPt
bo8O6XffgoOyYHmsFb0bG8BcHXSzTXR7WZas1/Mfihy/aeUzi6zlnPvGiBlZRC6hN7ne1TI872aW
JnV4MJgN9DEO7HoYBT7iAPGIRXFzTcRHEf+3eBarrmREq3RI/A1/IEQTLzExCNI3yvudAXhK6dkE
lgpBw8aD/sFSiLiqTlYcy5pxzn9PKpN5YEOJnyCzaGTr+RoaPaLYw6mqeuCfIgPQO688KIXMwlde
/sPt2zF71j7N5O1BMNd/PhphlvcVWCtbV0CFTmEZKMi8aCi5VSTJJumuugi2PjlByMS7iXPlJiNv
cwGpj/aqaE1INwL11XpG3q3nw5PeTxdoCPjh3AnP9sojjMSkPbhbqwbolNB3oRsFYlRw3OeFPnxD
skD2jJ49OpTBGv26KlWIgAfjZ6y6YaBNzQygY4Rpbx8JnSPoJmM5rwaoXSap1A2wmGYEk1FH0VaU
lcU4ljF1nzE3AV70oY+rjX1uWekWUfDTlhZnJ90IYgR+L29wO6rZNKm+hRPf3dpn+av7VWzttdeQ
bA/rrigqsOaByw78fh3tv6p7bEdqQIyIW2WLOJ9fdaAd0N2C5DUrFs9B+jNhVOBzBEnUX8NgoR5J
NUKL+QA7hUC2yeTY02anzLzXDDjMi1/Nm7G/nehuLKKDRBUCPF3XYQBwgk7y0VxMyh7J605taW7E
2NTGRnwt91u68+sZ6CEL2FRMLTVyreiEzcwsx6fc5YWCh97ast3LFsnZLMsibSb5/KLs3Qxpbdzb
x58T7qf1VWr4KcjehuhyphCUi1koJKCP7x4UZRRaTh0MUb+NFpAnKtRmO6CLM5xQXZ2jB5W4eUJe
tyuBUYw8FMDMFfH0tRFk/h80uHPpiFrWGfym6vpj9p9StClRppGsZTpSFbvhF4PGEQ3EA76o/rnf
cdXdJvR1l+VbHiwYJYJoPuz547R83bQwvDCK2qMcr++NRr8IRoJxbB4oVCAV4G6eOGZuB2PxX7jU
qGLwD4FfL4gFA8ZKe6OmVihxTldGVzvAxWXiMDNqP2lG/pjnTzJmHUw+R7t5WS+qs2uAgBoVIQsd
dIFXiQw11EIZKuwWF7T6xHTZgDFTEEBbYyVJUI1PfiNuHyTSZCdByUAv8OMQBqw2nchcsDLlUT2k
dNAGqf2+NYmcuVfJ873rzLd3MJ9dEndnWMODqkK+z5v+Ezt3YIZZ/5QBi0JDD32T5aKCUl7M/PbL
P0pFp9rDDKKWiTVzw/RaWwhV84sJiwbzwvHLDtYBwgdYrgD01Oid1TNMKI+y7hKNoU+C1y1GjhKI
qkNiIOgTPDylrxNLVY3zSf+pmWboKI90rw+uQZCr4amNKZU9EUSZ+RF4H8+lBfS6a4TlhB8upckI
vQaFfYVdOvrF9ZRl3FxV1i+IWIWnvVoMnZy2R6CUchd9gphCUsV5TTVx25+JlL/HxnIoqVlqz1VT
GvkzVvBsGU5Grypf7FVVCVKHPKjh14kLlBhd2nUD8dOwtTAl9wMtx3cgxie9FsHU2G6qO/FZGkbG
f6PoObIeT86clMm3TPIjOYoZ1nY67H5niEd7+8OkCgo8Jd31QZPyVctMfAqqwypvlmCUyDqM+D7M
HH3ZnMOXEQI6iNNgSVHM3YtLot94ppK0vQwbfa8iYBAKy3SzQq60wehMlPGAwZpk2l9lANhG5zcz
rB2HSDUBwHHTPQtat6BYCqs3LRVaj9Nxezs1JO10oGe3MOgBUCR6RHJJrtk1yJ9448BYMHKcjEcv
cjG6edIjpKjpduOegKFVdt8sv7xSGZTpLcVfIBMpT6V+eeN48GWPeOiSpYqyAatkhKQ45ZzmGfGB
DP55FKIcst9toDHGxKmikNxVY0OYr8ehXAESW5/c2He+ZJeGM34h5YdQ5rED7HVSPXkkkhgkUd+q
YLD0HaoAQAwV/q0TebdLKavu3bbjszjYoLiVHVu6f/BG533+PT9bmLusdmk+d+Xv97PGUfXoY9wQ
OT79F1xPlbrXk2m8jRzGb3dS6lHJEeoAWQ3EVFaM3VDULj1yu8jUl5qj1H//Po0x6pXQ7hgZh8yC
3sn7ysWd+jkhPaR/BS9Vw6unOBIKVPOQAXJDTA+c529uiuRkTllIfG6SvUohytRHDsb98ymz+i9L
w8a1gm6v7e126Zd6PX7oGqtpYYCaUQzwOpoG6jOmHMrTGJaKn+6o7CF7OrETV9fKGWCSi2Y9KqUH
CKtYT1Akje0Gvw4fTbpkuGvSNBRhnUg7piYNuaXeaBRhi3vApLp1xS3ELCzZEi/zGO3ncOEZlmKI
PPlWl+cuuRYqzkztfo7OJNdI4wAlalqbAkgomeD80doogKSdB3Cg9of8joZMKQBXag9nbWUnzNKY
9ynnJ7/nPG2wWIDybXunVo2hYRLsZd4tC7VupgGNhmmAEb8AYLtCISQgm55giwg3JFXuDfXaAMow
HS4G32DXWy7uGvS8xsQH09piXRfxM3r4rN52+D2fzNvKuYDS4IXZ10m/z0DzBByfvoCCOPd7YsQp
eu9kxaEuTdAR/LbW8yv9F/Lg8ZbmVCX98C63V7SJV3YBwJSYMzTniZhjEr08BykpZPLIolMv9Fpw
zWJvOeMyexpo7UsMWuZBoAWmHknZZJ9RttgMH9f8C9ZZ9SKvdT7L747ddeO8QNl1ngI64s10hfYx
l/YDGM5XXta42P64Sw9fTjGBNWDG9DpRjoI2xpHzVfX9vAJVTrFyEXAsCHRCqHUMAP8b0AtOJDgj
HF/MVQAr2jUBoU7oY+7JlTUblWldNLmy8ch2Yz6YWeXj99steFStsV64U1i0wq9lE1T/VNioq5TK
Ydw6UtP1U1JSs9qMsnYMkvbqT4fpEHRIMmkm+SudSV5gUmpCb78Qitf7Prq2Dl2+HbbEtxaeZXE0
FdX0BdmB7WcMEQcUlYSTeSGadB9pI2Zjb0LrzQE7UZ/CuKwBBZ0r7JyPd3eWZ3LyubLHV4Js5FkX
Pf6MbpP6VojhTepO1gFNDhUvCJWboJtvkbGmqC92WSJ/OhetBSOkrMcaC6fhX4BYr2chNw+TISI4
9WOFUJZdBackIQ7kJ9tqra4VZf8aZdKnzqBv9RjBSTuT5Isa1kxTVBjL/q7WNtctv1G+/iedVxfA
WZL9DyQhk29wL+ac+od459znaxAitxFluxZTnjUlx9Q1hRdKA3jMNd1WCHbgRZOfhO84VZ8SHsN3
alF7egvrRoPpHwYTXW3TUbaiWvNDI10MeAsP9QjrRnUMaSKaJRmLArLFW5U6NIN3gsQQPEqWTp1g
7SIrvays5fnnC1B8Wc+Tbm5AMZHLLxyC2OLEb9GDI8lyiwA7OXm1hZB5NVCqjVn5xA7bP3Jid444
29DGsdwXOdZGAIHjguWWWCDhzCXXohSJNw2oqOcRX/WMmg4dO7838qs+P/sRGbzD+U5hNKSCR8yC
eX31YVADoHrVdQzXbJ9xz+rmtfpLzI1i1zIw2RmljWeF/NUnBmRP0I/8cQEWAPP0CQyQ3Un7Mrt8
3KswGsQHQATZHEFG46F+t9fKWYPfrDV+yoZlVR20y7OHAOwLSG+VptZCkrBj4LHpnIw1M8peM6NK
9zbPK/qLAC8gtbZx1H08S0BBcJ6/Dj6e2wkuzY+PocCChEEylAtYcbdUp5YbwNZ3NRjwEK5lS34y
9Qp2FCFPLMsO8F1rKpCdWaPPWUZe2p0AJ5wNgATws+CigLtmseLWJsH6Yj5xJDWsMP0qWp9SZqnf
l525DOLZt9tBc1PmH8w/NN++jw52h/uaLJtx9HIVLRu7WihuwEPgxlap+0KeQQ3fjOJ1zWai+eA2
scWENayt7PCWQjyIg/HXV5+VWIgoYQbOOpErgjH4h+iP0RmxhWF/7Ttypcko5bzPVzsJS0BDBasE
Kx2aiffgl1E0iPR+kOlknSf3916xhBzFCUKJ2sUSkh+RexrYhWS7jgRaR37XRbgk26kuJqBV8eya
VUiUSCBW7ezh0nup7+yjLdWb4SeFQDxCHUkakjcW0dSUia9S50KhFTcj08xWHNtuJGTJMASc5BUG
L/XcWX4ip4R/3pPLOy2LjuBNf+UgCBltX4e3YLFxqV0T+7jpk9ucCHhPd3L7RX6cm5R/pl4dBjLe
a7l4zvfbh5+K64UHPLtl46UtrjYDnbEhpxd1VY/zFlztBbBhyWB03PAr79Vr8+rSCq2PupQhfkYZ
V9xEAZ48A8HoSn6INq88wqTJvTochvv0ryI1ahmYkN/B48+1tcSbv1OOj1Xb+W7lMbiAWpamszQy
0Ai+PVP9Som4Kkt+WbCZdXkPY1XsiAhlbNFuRDDt97s50VZXVIJWUP3qg/DIYIv39EJ9D66g5B1Q
zENA6XLXNWr1Y0rKb6r/le6k0Bmlans7DmTitMgtAxRil816uZheveOCiWnttb8cevvTdIDXCoJ+
e2/OT9T4eeIinGNeorHpv8/pJQu+sisuNi/daDGIiD13yKOujR06/JZQVo++x7fkR7gVuBzNEr5t
QRTXhPTJvM5BV/CPl2PwX04CaJH1mb8vQSWbzEv9bjM3H4fQ0mNw3X1ftQ/nMgCf0DCed42j9ylA
1W1nNJrH8s7tyjd7qH5pCFNHCwoGZ/34el85dFP0oz0K10diShwNfkoolndJPdFIPusjqxyHITZw
qxmDn1C4VbYxm98EJurNWv6hxhMv061iDQT621uLLR532pWyYLNORBkKIeelpPpbIqhusnwRepl4
15AjIZNoUNWAbQ2Cy+Gj+rtPJJ6g7UBp4NLtTu/9E6l7T0HoLYXvlmWfytNkA6mki+U71ESX4NGm
qVRolEvoJwzl4VTMlyGnEYKJtvv/t/kTpyItDF2A4qTcuurNXdLMQWTOswQBjHgcJc6zSX+TuwyY
jOKwytoBLIfIQaoHO0z3KPO2khxJYacKwca7qxa8i92nHU1gbr17KStafPxZraevCVJlUC/Uvbsy
lGV80SDVC7DQA/GeVsguJV8tmUhLxUr3fAnv32kcnHjHlIwEXkFSpMS7MebnsBxilzeFtigm3sPq
tqZQboN5oRISOsNjctPqgPIEZudXEW7Xs/ukbaAYFYoyyy7eJ1A4vjjXPzFOX0a4vmCqeg1e0YOC
iIwyzJGMKtkwfek+HccyJeO9ZewyzNo0lOc9N/xy9v1HjlarbkcUz68QkRMQAiM/fsPiHre5Lx+B
2QjvsOJYEd27LILGGMCX4/ZB6fyj5tGyx5DUM2ICDWm3+lZlCO9o2ZIhzB7VBXqXIcaA6VHog2Yb
0m7etWcCGHwyEWkPyHgs6IpK9qa2YDlSXPFlUzWijhqmvpvvwXVwQ3jLZIs+aHGDMaNVjTSnMJMj
F9ImxKyc0RmxMDD9SNxCH0BHOWRfeIW5x09877GyvATGuS1ZXCbrSIsbMv+DEHrbT+K9PXQSHeRm
+QweXmgBFd7Y8Qv27o2O3EjKJMTIB4Zf1C9pz2wjtMlYSbCbzoI+242pyxkSBpJ+jmbaXArIESgG
QIbQNs7LZPLRprL6fNFC8WkSTUyH1KjKHalArkSx/5Jgj1vs5MDnimIaMpMdwxZhZvaXLWJ0pqss
6vU39Uv2x33f/5CeDxPuWWKbOo30ddxjsaKQmn4sXtqGrJk73qFgay+/foWGzcZ914fXLARzlNOp
gBF7nSk0mbZnj0nl6RbKhAAaHkraZYUgky9m6oDYgrponfFMr2W+9eRlLKiO7IngTf2L2inEWdMK
D0bD5jELnmG5vfOQtlIzZ6KWuIopji/wca5Hy22K3CtkWW4Bjx9QCAvcT3sTccE8+W0jeBr2N+8g
wdbyDfT/M+gGZ8/e0iC3+B0Tg3xYxtjNX7+ERlwxnElSU0FQQ9X4fszMcxYWXT9/bDMRCJokz8SO
MPy80kWviz0jtrxGdlt1wxtaqJbHEWWTJANxb0wB1Tf1MJBeNa1rBgrJ5gHA9yzrUURUo+rADMwB
m2DRIl2Byxf67dBES75hxwNEqa8Plb8Oh2pPqs4JzlKjpfIXxhlGNz5OlyKXI9WzzJ+HtEtqDOHg
32upmCxC9BVcArDI44qfFv7P1k0Dn4zYY9WnewLDCQlxLwwzrJ6CqSu2DJHoX/yJ+IhHXBHHizC9
+sq8sEkzzodka0nsqES4ETOTW41YpGD+CA7xQmYUBORy5SbDJLxqDhET8CC16kEm4CBRG9DSLBR/
MBSTCRn1TYfpipNtride/fjGCjS/16I/3OpoyhKiFKVBkn3lhwM87nY/QEI8KKcY0Jb5QxFzev8i
Ir9pI7CVYrqIZrw5xRbAfX3RjXXICNhpcXK0mgaVbTyZ9BS2FUJX+vFwRVgsPj6jB3mmB7fh+bOG
lbTUT7LxkYs+cu3mvJohe1wuW2nyiZlcxYIUqnRtVVvllLACoQINa4izhmY3CTJyW1rs1Vkt1Y4Z
OtWjHrN0y3bEXvR2vAzRPZ4ktQrfuVVAFiPVWUn2v8lqnO9/31e9c2vpND0SGH64o7zlDtXoUgRk
q0we9KLBxu+v01o1kwyc6RBqqpAsFWuJ/YEqrwFgIhrnzQbPyqjCaeMXlRozo87ZVg8Lmwh3Au8E
L24lwgAXXn0x076KWAFFdBIqv4PKA+pW8OT3UDYykogs0KhBLILFORrbPhlt9odQIZjixCLzT2MO
s2NTDNz4MFLVTcv5anWH20F7TIwikC+G9QxpPRStxo37Qypk5gigwSMUYLEzatFn1YVGr5Xl2P3o
vHOk+EDaY7rzC3Ww3b1J6wophX0pdQ9d4ZT88OZ+iNKlgKLbweUGGJjOqp6o7G+cwlczdrxI0e5B
VFqEJN5aO1T3tofuobMXd77/qSq0mEDU7F2k0ugW35qP+gB2ume4VEse/XNfWV51CRFSU2KQqnr8
bISbHigaxPXFiTbTyB8+RzO9d6rg+GEqToBojvDC6CtCdJlrz/gie/BaUHBMJFFuUl8zwNAGVIZb
lYwjihaIiKXJXsQUWuJ2ROb4JkCh3indu8AnJ48rgORKQjb/oYV60PDOyVCUTPKG42f2NEqAO/jr
1TEDLz0AN8Bk3N84jrybgklsKuY5Cwoz/sujNcevhaDtC6D6k9ESf5RbCFVAdpPA2I5iTTNRONll
bqsy/7UuDny7liLxBV8qUhO6JCUhz0jpVdS3/siyU7gNIEmYMM1NGHHMRO3HZWc2FGfSODfgBlzB
uXCrhdiBTRB3ESEG96Pezm11QKFz3aSm9wwmFomX+OAL2pU28cqRSi6CE/NBcAOPL5UYqIpv0a9Z
2CXd3tLf6YKwsma206FYMiIklw3iQxYmQ7HYVt/6EX1Ez35r9TwSxcv5YKbbZIzhZyhhs/bBRpIK
ITxLeTywiG7cGSduI7vxdxZRKCaPh3po+F51B+67HaAwuzNBN15f++FmJAoN/vbw6O2E9DsV96iQ
koE8dtmqAH5Z4tSwCUmyCtiDVghPUt4qPX9G7J8N9U7RxsUxpTAQqwc6LmZb5OdgvNm8wa+E21iE
VnDL++hM5CJy4K8x78F4uK6NKNcxlaajVgFUoaYF8NAtzS15VI8PlPZHGANhV9KdJX1SvI4kBbBf
DORqiYYtQF0dsgw2pHt1R7rfKvM6LpaStt3c+GmWohwDqOBm3PHrPhHmB0Ri0Q+QNLvlwwQesieV
3rRiqvPl088LjTlTE6ZQKl/x2E7YzHxDnOZjtam6G+gvolwnE1MBoHSVh1CmZ7ONaZXld/u9DMA8
dh0ev9TXRRKUVTWW7t1ThA2ljUfq0jgraCrFKQCJUdQUcroSrshHyGH7gumfCJRtj7OBC2APim7v
9KvC9yTlV2KyWXFo16vIRPSk9PVMyO5JYxEIBWSAagM3t5/q70mr/cN7HhiBjWThrIgwDdAUFV7x
INwQ7Ayi7hIzWXVrN8pVGuUpFPdZEXb49CsbtqIU30MUIlkfuqFWEykpypP9oB4yGRt1kdcewDlJ
scB8kV7rrpeC2XWB56GW1VJhCMiIP+iiSEvmNggIcUwOwgQ1DxIqLmdEe9zCVG3kZqkP+uwPM2YP
ishLmJkxO/qfkKu/sTbrJJ9otYjKiEI+Q+PKfdhiTo4h8KB/J5QxKy93i/Bu57LzgSqXNxfDcJvJ
tamkNHQ13D0vGNzypz72vOB97Z20Oo3Lyyd1laueR03L89t65JBYnHjNEgtYB/fTHwrjQKryA+oQ
qKF9mXuxR6FkQeFufh4VIDSvadVCHy2qL45KZ+9dR3P94v1MQUaadF0Zu9nXws4yKrqtPPt85+OF
mPK8MWzrlGdYBMTVvc56e743xrzu9mN/5uk87nVSI6cWBsjnMowOdH2hpgd3x8cW9e67RRRWP9jZ
KgoRH3+S9bfve5Ttny1k2RM1KvuH10Pe/L6isHaz2RQjr7ki6lgsPDojb0RZjzUtOuCohXqK5oeO
V1mJhDLDPk6TNVRjoPxWEPyAd5csYEcgd+c+sysUXpaCXAqDkMlg369AOlk62FR76pRlvC8P4Y05
eRnXblCfzKHzjSpc5FwGsuaSbdggFMwjow2Nii+Z3YjXjAoOl/g4U8Qr1YixS1b8f33WOBv7Th+T
IM1zxJq02C1jux2Snr8IU0tgFBSv4yiHO6hp5KgELOiknW4zLXPrGgTHnDT2w3p+IP1dyXY6dJu0
ALe2/uQyBOQACWrWtwM6dg1Pv809HSMHJ/RpBe3NmuW191gpG9nbxojvwBCZjHpJS47SFzwkUJLP
0cCSqy1gPhzjRGfY0rjLYtH27njOoEm2tKhZIrWporsKjY6tXgW0mgvVXvDzZXe9qvQZdt0l2fe3
QeBcXUbLq6FhNRneU4fR7wPOGdBD95BibqKeDoin4fYS4O3pnlIlUF8whL2fcdKx61G+V2cBed5i
PSm97joi4FUOZb2isPYaM4+2O3g62/JIqiL4iMl0+gBuxGOu6xmeZWiqpEFC0rryQ3SIoa181nXk
jLzhIjp59cPLnDDFggIY34aXRzUz9FWMUXQM0JI3YVTsV/FZm+4qzmLDHfni0mYPbe/3qBnsT1xY
2FCPcojaK01k+nydWDeIDt/OWD2/L7gN/w+62Xfp+lkwNPWc5PvFKYnkLwAAmc6BKyoJCUNyTOqO
vgD9bGoanTDpEb52+rsS+ZRgSCU7Wl9/7zrXqGURBglqh0DjFA/yxjj9FHIqiMxFrHdJqefPGYJo
bg1HrWN2ScmqVdabQZrUEsHx2kih7DmNiEblgiv2g2L0tYumW5X17MHBIowk5r13cAas88rlLNO0
VN05WvBuH4is5+NkbjGOCclgdFkZVjZMTDvKQfDPKAEOXzI8Vpwav/8+8C1ZRteeR+sPVeqHo3Yq
dYRGlWZrzN3SPBYs3k4iXTR8NjWHrF+Aop2zgWMVNNJgRP33JOjbwmVTOkkpEOvUOsGphpEa9E7l
HzrzEkrv5PbDuOedcehzf/8Uch4qdkusgCHtxJFVWJ9zpynPSRml+4pu6ihyWWbG0D2OCH6cOmah
N44vWAGKvjpvbhl5MSSdmFjyTmUdWORzBWdf2qbsqwp8CqqvVpqjF2StUCBByYzcTC0+KY0PHqkF
/0S3aRZ+cswjTHtwaY/MkuJpNo/bEmP7oKAQz6kL/ZoohtG+0LoFLAXfkIMy/2TPxvwa1zmBTVto
5FGwmmF9g7zI1a1d5FB+jxWcWXOgpEmXcY2YrEdATaGkK1yvO/GUYEhKxlXfqPruFqF5NUvwqndx
+N5he8bQ5ipDJSr2f4+BNdMViTrmngGMFmLp7UZff7IBBc+a2Wn6r96t7hLBaVKfR1milQ6tCFkz
XUC0V32tihQFcNTOHNd2Krvo1TQnYcJE7TPLb/5e9NIJvfqyka8jedcGPzUcCIPUKK7oKE29Augc
HUBJZo5S9K7W0HAtpaqkZn2KtQiSRCE6IAqBE+rNqKW+E+JGdj0iudX5jgAbrou6+SQvD3l8eH8K
bfUfLe/iF7Aq3LiCsyo+DKQc3ZuGw9qDb5/b9IQgMEhEObXgl+RInp4oEY0KSEX0d83bufjBHcYK
XrmaVp4NWY0KSPKej4uR7mQPSs8OaKMxUKOKj3QszXCYXIGRnmnmm0BBZI27TDI9AItqExvAFK/X
0l7y1e4s60bkpwIhr3gukE7VqcEZfJwxhyzdWRx+zLZyqIf/WxrIMsdG4EEwYZiAyxFFj0wG1JjW
b6n3CpD8FHs7f4qUnv6GT8F+WTWTMhqUZJNZuq7fZ35iys7f3Z7sDWafZISXgClvFiItWCuMc++2
wIamYQHTZdEJkaIhDWH1CAn5ytl3saasWwlQb2RGZSYfOD1ZHNKXZTytCFj40Cflr3fbXisHxnLR
n5sGOxRPMCMYKbi3JSyg6sCmDx/2amtZ98tblGBi8iDHkUaL3qp9bvtE6HJrX+Nx8xX5xpjz4l9I
aTZmPpRiYDBUqnKYP0B8aS3y7C2CKZilny62MpRhhKdW5CwMw7u09/oiTXdul1GX4+9I/sZfugSm
OWqKA5xAFR73dwidXI1rM9aRvydMPx7n8if8fQwXU5g2/qF4f3YQ++brpyoRm1qGJPFWIvQGXPsh
+adZif9X+msB/aheAkesnov+LEX/ZR4AzOvE0QOaJNd+3lc4d1gQFK5d4LYkUc9gqusgzkHTSTMf
as9m6y9s3VnuPJEquQupg2XbnWrKNL/+Vyag89thuP2eXvro1O1IvgxQ8LyPm3LjjBwwu67UfPEW
LG4YmditaNCDoYXS/u4K9Ah+NjtjRr7Bmcvl0wuBV9WgKMEhhJr+4mcOZ8hZ9STiDpXeP/mePkvk
2hmRCYIaGZyUFAw36MGVfQ8gOgyaapn6iVKuUDTyzqvDLkw6eiBgWJ09uimrKJlg5sQprkKulk2X
itJVIx4WohnQ4TjFZIweszwFx/JeWIiH4l45fTiTsYyTDF3+IGK6KQyhJTYDjL/k+X4JvCOjnGoZ
5TDUL0Wg5ik6Bbre+h3sgEgOr7m2eyGCgKIODMoS5ZxQNqMsjavq/VYJTiWMS6Nbs5cUmA+lB7uZ
KHx3zHADPOP5wc0Tf5fuOOGCUW0i4c/EH4YEXFJSEN4sVJukRTgxuGeCXQM93KzFyoHTVeO6yutu
M/PuSIBrKhtZ8B2vD7RCVpkpMzu+Z7XHE7wtkyEHdYh4ScUmUrdH83LgncJSCCfPC6lm3rvIeg/E
eBtrKoBAlcjArArppSSecpq+4mrRSK6cAUogGADS/w/ZW0KEq5+j3rQBkQN/aYITMmJAvr8nwOX+
1YgLji8yNcoqfaF2W4QqaLqnMGIF6BYkEkZmOVjS8i1Bt+gvcvbdGWkNkt1sm0f+D701EllDs3LQ
CUu+Nq7Fv+Bx9ZQspb0/5WKhOdJk0D5QKEoSlH3KEvYwmcNRWcJ4Yy08XDDfJ1E6lJ9rVD57gTTD
ho7Vp4T7S851awsQxK3ZnX/awmBo0pEQhCmjR32Bi+7enLoOiPvAflTtsPdM1WDQm1n3rHUoAgcW
df/47ZfjkGXemVZTvYAkiCiCuXUn7rSGMXsHV09gZjH1P00DEsQw6W9sJqL7Qdu/GkLP5FdML9da
H3d2wUh5VL0it0gBS6tEbxyTOMop42VvGsrSlvQQnjmJ6pERuUehK6ZCiI+X+C31+LCrQN/ymApQ
DZn9V2gHVyYDN9TTApUDlqCjtlVmy/FrhmMJA3EtOQD9EPLA9t1/8WiPy6EoxOh1lDRWOHb53VoD
XJKjvNF139CsATWv0TFIagNGuWy70dmBYe6hYAXXmOBM9E2OpzT9SPe8GeEovP6wZzXHgSWFj+eH
xCDfQiJrpwiD7hfu8j7ELb39Wum619ti9x/PGMHJDzOluSMhsgY5ex+fE3iiWL5uv4Ec4ZqTM5kB
Rx9en9vuOWOU35YwDLYgxpZqVHym4XLKDgTmSD+CdxFASwm59mtuBqhkct1L6Zdy8+wKQSEPZjyf
Fx9R0IzL0vpD2HgJDyyhokSUirUhZFYXdJ4FcCJkfh95GvTzButYC6Mil8vhRlwoAVXNWRC4KVA8
fgKfw/+s/UelrqPZtJIzB08fNcdK7uAdBRQGZUllBSDR32JtFvlj9Il9d0qWIm0m+ZMoeW1P6c9h
JzJlga8En+3K+ugosCtbGPm5qlXhVJZX5EwqjAv3WQr8aMd83XBDQl1VvQsFQpHrBp8bPdo/y9CB
KmFGPSk6sTUjZEowzi13VO9nGqFcZXVQUED94J5gaNxDGP/aQbggZ+Qikq4ttl917ZbcDMpcktsP
u0+8zUg6TKR5lUgiGOIZZt7y6HNPaflHBKr5eAOhY0AM2yunx/X8psRSk5Wy0YFJRd3JY5GUxJiw
OtdkXTADOaNyoRvxZnDTk020c/JWzdBqyUidGxLoUiWk2Xj7jGLhaNmYjc8C/0RInyu62/CJxbNn
hjdM8SO6HiGl+g/Yd0lRIPDAuIlHf0MjX88WanfTBcaTNEdo1I9Zod4+47n1dDMw51/Jo3/JVwlA
SVMDCT7KD4NwmjMV0SGgZMGQ5DCFJssNi/7ahVKwpiqri70zkoN/IsXSQPAnY4PfyHu/RC2jzKHC
u9+V1vfrtcAoIMBge4RBfj2vmnD+wKEHaKW4lCy8lN8C2BHO0XQT+jD6fSIRq2kyMNb3Twv7dtio
mhgatos9gKSPIBVq2lcGLrE7a7E9HnPvOOJWf5udyTdFz7XZ4dKob0PC64dk+za5hDVk0NEHzad0
xuqREImahwZDMXoi20zb3GRsxcvTIjs0wxLEaOJ7q9/sLjV0LDlyxfOOTTfgtRcGPXf87K4FNCQJ
Rqy2J8Zgzkm38304N460O8k/ZAVsi5pxFhvjHOkZZVooNjS89gcgjo3m2TjGQi1y4GWuDu4PVDBm
MZTIZ424Rtt4Sj4hCbEFJoX46+uFIUT2obgpoghTgXkAAxejaxHCbPmEbriwhzYk+GyM8YIdx8Mp
E6XBEH8s6+TCB20+1cICy3YPqHZfb3OCwIU3HYUOGheg+tc9f1J1sj8v4beVIa6xd+FnQ2zDfuQf
c/kjqvxZl1we4fgUJv8w3GtBtvCYHjzv0ZOoVGboxXClYn9Rdm1k4ZMQDc2I17hNjWyT+1PhFcp0
mOl/M0Y+A0jcOGZz8qqhWT2pFmwlz1dlOT0Uce7yTE/y4F60MZRjXUYLeDd5/YXRkpB++BLFyDrX
C0QfAEabtcbBMJzjHCsSi0awMKQiuE7+jU+RbvT8VkLKdONAgMmOwQmR+sEi1DxIW2aFfLnREDnQ
Kc6F4L2+W0XtUxcuueTdwrB5zgNQF5xq2YO8ShKB8CHxJRzorNnpWhCkbyohaY6wjnmvOHnCUilF
dfjFj/+yXCGSfR6/gO4sjGDdN+n6nawwcXILxCcUS9V5gGm9YYLfBZ1husm/YEMw4wQ2EslmpEmD
ghRf6vhxkH4loAwpDjLAduk4dAggtQsQZcZx6imGO6jJXGDKlj7mPsVu+a/z7iBqBwiaqEVaYKtc
pgNI1mFfpiCWWmmM5K54a/6NIiYoH1AwqHINRQr2yViXIX9OpxA0xtN3I3T0swmURPnk737Sr093
RQ47R59EA4mZVQ8pnRkIAGjlc+4Fn8T38V4MSSAVQfnCWdxGGAG6Qmr1sP3JlKeZk2bQhCN45ZBs
o/TUQnmW9jmiPmMpXx2oTUlEoLexq8zEnsyGrH0YmuOYYNK098iIhsHrAxlCA1v6io8M/HCtNBkA
Q1tww4Tab3gR3GPPR8u0t1lBGI8yd0Akcc/nJru/O52gwCR1z/Ebt9gAtjydEAXnDQHi0lBwLGQg
suX7hgtGRBkBUg1Jg5zRXt0sxPNZRN/p9Y59i9w/yW4TLwaVgdr1JmnpCc1jemnJkqJ+k6SHPxBe
tOSqw44STXoNbA3Zd69Sv5mlUv+RFa64FTKoWIKGjk1RryprbTifhf9DNz5VAr0nFy27zn0dqhrk
RwT6eJd5dkVM/fouqZ9a57bNqFS4qhuyiBiua5kOvjh//Irm08d3PyUThgQEVE5+6y5TZ9nIJkMj
Sw6wQ+CpUi1mXQ1wt+MjLtDlzybDOhvBtA/LeD68jmoY5xSbTUnK+oaW2cLKX+XyO6snrgYdyxUj
Rcrj+LR1vxeX8NQFV+DHRuT5IEnIQlZ+S2oiJPEe8eE0ihzZ1bZ6DIw1kRneVhS4cV/ZlHzf1fBH
QeP4IlGUWC8j06QUT1o/jd4b5mhpDPzYw2YH2PKNJErKG8umRdSA+nxlrHuPcmP8S1p4EMRk+Ne6
VwKizlsU9HbWazQbRby1974IIG43F8t8lHo9UxEZ2XTeqrsBDqlGKTIDccM1/4I0jrmEuEqXIq8H
BB6kxfjQMxnpWLA+opeIcB2/BNLTkxpBHMtSuFDuuXt3aAbUtZUFVoPPXO85BiLW1+YyGqQooqi7
1HRUVI1xe3EcvgGMkEriZvWDehBN20Gfr6aogD90WLJDrWBXF+kmCDOF/cTVK4NosFjwAzrICi2u
DajfrOLopvwCA2R5uYoM2TJ7gF43moxnCA+R0g/Fhqi3nxqlzyuUQ/kMq8wOehR19k4RqXqbXf2J
L8bGT/j03fy+JjwXz5KhCXfVqDaf/jscHqtw13XDbXF/ZM2szio7d2Wix9gYTzK+5St+boGTub+L
14gXJqBmeFWAjUfCJth+VQlEPG1ttCC10nP5B8O6+SMkmpuTIWcfWS/j7xSCVSPCcB7mXx/khTwl
vw1REcnydsF55lc8T2K6w6kKjwEo7DMHzefZLomqjVS2qFPIdwNejPn+rRxETm1HUWvTvALv9Nu1
kjHOFxFRCCMT/Krq4x/ci98lqmrjE9sJm4aeZ+Mjb/ypmXRbnDPugxxmvyCDmV/PkoS6jWX7qkbB
19fGDtCCFIk3RefU/6i0Bi4S8mGi7nsFiwJTDirwc1DySlvT77HxcW+tHxWLyZ85tzWWpFRsamuf
YQKzNaWBO2zkcMIwweDSx5S2zHRrzRc1GPMR0lpgFrdHJNM3dDqbYupPWXHJxH1bT/5avGAAEx+Y
ofCRQ+zAXFRnoRMRHd9XYr49TsR3DqObjQ6a+6/omhTVZS1DlwnaD/JL2ZZyJDISNoosZsu/dLBb
7Bs0+S3Ra7KIGqp2VjIidgyOcyZ7Di12xAx0vZr94i4ikzoh0dekyjdxUH1FohdeMSXy8gbOJ6Hj
pALS+K3yVlEKbrxCqxZHOLUozQ4VHDLeWY8+4CWul71qHrYziBq1/mPlQtalRQgfm36CyaZxoEQs
fqvJN+ElgDNEx9RJV+em04xZCE/5Hp3otm+/9KLHISZYHv3hGh/rkqu22SKkzAJc2vEdlf0M0LDj
/XGaCM11QK2rl5mdiPs/qJA55Idp91A7pKvnGMCw6tuJkhtpOBmToTVFePpK3KsK+3kIjf9aBru0
vEzOE8WUpeit8135as1q7uy4/DYnNKmLdJM24fPlBzumQhlOv5m9hNUK/ieDv8ZCxB2yFf1G11y3
ftGarfxV8m2TUQj23JZ5xcjQmb3Nwn/kJOWgEqsxj+X/Vkyjbp3S/mWz9FSQWHEXZ/ZF8WZoxsfN
qcVlEMwmMth+7XhfBwkrHEOBmQO1CBseucFjBGJxqoKSE5izXtKKUrW8/ssfzSPduCUYULHe5Yi5
kEaX+1K7P72VXun3HSMhnxzucJaLkGesIFKXJ4x7CATt7XX27wsU45O8f+npOGPuHEB8XTyB3mNc
9RA3s8txUGRdJxGzJNVuC0mlpOsCUMA9CZXWHpt88E+I6d1ZOCvwt0xR38KmlpFC9x3SoDzoJtnO
AbAiECBAfx1VRMCo/eBLJABMI350fDA14igNXQpg+yuhxxywterwxIIRReF8Ngl/N31EhA7wv/eP
tyM1JSFg9Q0SFrf8m0vNM+oXmMwPBeBnyAux5Hh+/yPNS8eLHOd3ow/2BqYojJB/VhkigrKkInvz
JjRY4hmhd8jfXwRZuvDed1l+39EqI3YHNM50VXvarMJN4tbK0adsJ21UKQqhWwUVaNZNQ020MVa9
xHWKTNOV71AGPtcdQl2Rnh52uf1a/vn4HbfmwXDPYzaX/+p214KzBnW8ZujGAgXzct4t4HxxBR8u
6d03QkmGt0014eWAZE3rUVPTn+WvxhiaM8s2Gc9zmJuA+7YJk7ub4ThR8fdfPG1R7xHqlWYm+R0l
Ce6XV5xh7/mk7INXEZ8UC8M+fPpuWKlH17OhME83MQ5JZKikTMb0WJ6+FGosPkiO2eiJ0RaNZvJf
+coIvIFyvF6nXgXCJC8y0pkDgMTzWZ6i6AYl33uhzLRjIIlj6E4jNwhKamHAfYzdcnfHisZbBqpI
u95fnnZKeTU2XYebIgorheZPVxyocLQjJ26jUI9eKTXBYmgKr4T59rA56sUvxgK/GRsC39295G3p
2feoqrTREZ/NFC/WaFL9qpNUe8gybABCo4VDF5togH2rpWZlrzDAg0ufFIrFsZgFwqSfPxfcMDfW
bUyTaXlziJT1dteRkZ8XV5KKCup1Em7EQELfD+cRQOhbXc71+PTQD8bafjpiIiD9A/oxhMB5miFR
eg+DkNY0GlI8BjaT1MN89BbsfID8OZKUpRIGs3UgxzoWG4xYcXkjHveV9O4F47IJAQQ8SKVC52Ks
yU21xKe8QxyC4Ffr2SBwdshNNuWXS00A8w2iVfsO9HiV6Mbnb3Wuh+6XMQMs8qyRVYoymCIT9E6V
vddHZFze/dzcZ/nQidW3w2igeBZTG7YOKYM1VNHiGS9/BHoPpnlucM8kPVI/SPUB0fgxuYyO4BJw
ALdx9Sl2seKjptBDSh1fZGj8tuOSozQGyOVVcF0SZnlJ3qJOsp+hD4sMfMhFs3d6pBliAWtMVbf/
wSK8s5sETRiDcdKn6A4uEiUYnO0xw5QmgJbpR1VAabq6h8aTJEOP/9rZD58ng5t4bgUyCAV347t9
PGt1DRauxuLayT1nmZ0GwxnV8MjKnihUbucjWrTx+3f3yLrm54gWKg5efv44EEUGdluMHYprwyR1
7cNZ9iRH74RG0exjk/F9feq25Acph32Ha6ZOzQK+uUwebfqk66SApxQAS3xLrrBrXZs8d5DnM6Oy
z/bu/47h7XV8FakYIpXbPXFqy967aTONjEh2bLPxTFt4dMbLWywVrOb2+zNjgBqVnIBay+12j7xg
s8wzy6M/3/+W5xGOEnk6PJ4gJSBB+pKOA542A83TVxzQOTtNwCKEbzdcSn0OA4gPoBkRjG6EOffM
psPcQzwlPu+SeVuzBctGgQ8Gl1ziVSt4+1ZzPTmY2CziU6KiV6JrAQNdTQtTutnE7w4HazEsT4Wo
m75naVB511SVofvbL4ZMeqU6btYRnMmc177tCPaX+PPqck17Sfx85YAAkp1qvcZdbMiF8B0MxDM5
0P3VzMt4rwR015j6Xq3KIVtRyJ/1VfTRmBkrBcj7AK9/likbwX2U1j/4WUnwkRaJ//zJsYJRb2LF
RwNYIvbqn0he+BYVfT69mAT2XIYP07cPVcpbfcy4tB0ZUsQVzV2JIfaKAi1XQaNknjTE2xx0Qf8P
Z6sS4WlQYu8qThcJ3kyTyqBVD4REspUB0WOMdBTvxDtYcY1T7PUmk0QrQkeM67IOXdo6KHMvK/y7
kI6cxaNwj/jgbxhYa6LsfLvYEYc/ZOzMavUv9AO+6nyinU3VH8WafccKo/f79XbUycUE4UPxY7By
l8ma+wAOwP1wZ0+AO9t5P40jm2DAmW3wD3oCRQJm6GBBs1pGSvjL09HmO9rFwzQKTP7HCMfkQaDD
92AGjWAHbB5K0NXAaD2pR50/okYJL59DSAIRi1/IvlB7RLPJ61NokXG00NqfvPku2jg03Z8eCbnW
uQmsum6bBcdE6gvBXtGVxCgJ9i9ZlCJQSWmFHk0XZzcFDQwm7QgGNR6h7ScQa9IryG3GSlRmO3dj
0LRISokHWxU96sHIL3NFZHA890pI5ts8GNiB2qMiN8z0Ge18cIb/DiGFigxpPodhNkIBrTKtz8xr
CuAw+v7oReq/CDC4anwrHBT23UvhPLJsj5W9Gi/MvshLp2TEYcUEcY80fAQgtNs3b3pKImA5P6+W
9g1CyxBipwq2xP1R8G+VthLAZFjw6mC4ZzqKfD2f6va0NYJzz7SdxYPWSFkDc1Gw5uR2CQcgyx4x
N/v7WtrwNOUJQANTqm51/sJJQdvIsz/Oh0eI6aA3B3shYHOKoR7eFDqIarffmyA0qTkKpxsWUMQX
xlHBQ43q3KlqXyTa3CAXvVTHvgjMcHPAttwpvuAH99a4qTCO7Z4nNFYB1mCMIivEyzZvOaALilr9
d+8KTqMoD2JyyzNJegCydp2lk+7whwAtEgfcXG9Slel7bnlvWkPYASxqYfTDF1sogqgUoseEiWKE
avafVsGi7IiuXFXtozbCm8/uGkFal5sPLCtZHopTu1Bgb0+r9ZDDZY9jAyy6R3Lzcqw5F1D5BKFQ
viJtWopymKs+q20V3zFripfdbHFk2/QavyqykbVieQgmKkp3fkKoTb5efZ3NHRN5YJxNttJBXs5o
WINEJL/TloYNO+yppjWFJdrAGflPNkKRvBJcXhffFFbAnb5r46IGYW3Dqy4/fM9OZ8GsrmQ/RjiZ
dmsJkQ8mZQaqwMrMT/Nm+oG5ggl1Iz7HC7Efu8tGPDHmD/wEG91pM2En3P42zzrSiP+h5v3XhLnw
l9bcaZhvUwOCNSRITP2IZIdohMH95ZuMndr2+l3qRwk/r44D/JvugT+n9O2xiYB46/V4xFMx/PI9
ZhBboN/gHUj9/9UVGCKBlRX/P0Z6eM68yMXYOaIu6iMiuIr2rn4pEjpwZ2VoS0OJeqXurxyt74jQ
5zmPMWHCh7QUkfV9kHSGVaaVikytSETok6vLavle5d9NmnDkMicGG6eTAzj45O+OfBsGeXn43G54
2nGbiqT1AQJ5Fj8ZbucL6/WGldeqPtiKjQX482qrChMLkTkr14AcVprcaglsG6BZJFXYnTQrkGn/
dHTr/OcCHmgqG1tlVb8vrV+XRqRzX+CPoaUZ4kJ5nXYnjHihEGZF7+7af0GSt9CUCld0Zq9bFfHa
TNKHBaiML/0bgcezWR2SpocXNuGxPQX9PdttCdkEadCemkjRlnCgFkJUfm/nQcgPLVY3CJ1pch/T
qzpEAb1Q0OSddFRFpqUGPVxXre9fsueT70tlWQTxXC6Dy6/q74lV9tPlmUOTandqh0UN7lUVEgw/
6BRE0SIGpz0/LzOrh9dRCVy5/L6tUxSMyJGz+qpZr8KO/XV4uNA0452VQ73uS8/Jd5Xs5moonjm1
H+p9QZqNJJ4jcPmujZRjc/zjpQxLGgz+X6vMMxGprcWUyOVoM7+kB3zvGGHvoNMwlyoR7p2h34Y+
o6uRo0CJY6dXmUc/fm+amZjWeTZa79VkiiJoAIB8R1BBYyMhhAOcHJrR36ziXu9JcNK40RDdq2rW
Ba3f6uSTW8yWiITweZcAAmbLq12wI1AlfytsuG8kmvQOwShVyxscj7KHNAZJXLI7xPOOnf34oY9R
H4byakVBLtXwSMC5z6g41FyVZI8SJUxHTBMrS7mQjp9KAsxB0PNhcha2e7xzKzcPHNvaaF0anxmy
U+wbhtlBXQSd8YRRGAq+SJjHInxgiUsFftdNWeht
`protect end_protected
