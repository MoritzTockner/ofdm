-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LEcPDGOfenr6+eChME9MkRboWXRtz9bQg5gxlTgDeGof7HYoKxNuPvP42KvqUbfHFZF3SVaKRKct
Da6KFVeQw88W2HUdCw8SSYyB7ihVWXVF16k6LkWwx9LjsdciJpbEj7lB+lpxYbs5GopRBdk0KinF
8/eDaTd5D7Ec8oj2BCdQylb1m+1xuZaahpvEouLkyAxKsZsfdB4RRuekv6+SpA9BYjjDRV6WzPIM
0Kyi3ZGq1GIsFGssK6TqCj4bE/4txygDqgwIOUmzacmGHMOt6PUvvAcqa9DE19cCvqo8ZHAsEo/o
SC4VPfZOfke0Vuk6KbZYWbxlxbD+e6M+ePO72g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
/My/Ht/FF74CY8uyEGuJiLa5Dbj+TSEXnbGS/hAccDSpwdlclXTzRjWoNCqohc8BKqJgTSEARxcj
6wGkc4jqgbFGJsL2T+oWu01Xe5D8kkRVeNWZM58WQ+meD5+0X1y9M/VL2GTACxKaguZgOzAZAfYx
AS8excdfIilL4mkFlZ8iEYR6jQB0yj3VD/y3Vfqg9f+Yf5TarlEv4W5ZDvOD6VPiRlndAnVAVxSs
W9QRYRA4z4O8OUuFdoASF1Js9Xu7gsCpgyaUmkkS+5T5FJ5YKXGkD5ImTAgAEZZ7ivkDXMEgYuwO
6AnQ0JVy7x7QTFnJyNcsk5+CzcyinOfaK//1tgStI73tTgtZf8UhjBoxYXimRZbYiLSkz8rFtoLJ
9UnWe608314EhP7mEHSh2DlqFym5muudIarMbUZXY0G/RwrZtQvoX5qKbIL1WYbeNFqeYU5Jy7MC
Q7v7bz1FevyJMuvlJ3WScPOVpzfTshCbX8xZNymq9Izg6DrlVfxAMk9Z8zXQX8yo4r8kV+1idDmv
5i3+Kb0z+JGSXwRuUOkBQX0jCmVlBVpCRB07FFxYbVkyx5SsaI2V8ahfwpU2ufo8KcsXa3/knwTB
nZd9gmss0ldbaReZukzYllxxgBh/trKe3rTyRdqSNtfT6fnV2shTE8+heDAzhKUu18INyvpfVWHs
tCyC62Fk4tZZOyEkAAT6/8V9Y3qCXC5oyhiUomKSJSXLad8lKcAOq3r/W0tZtsgLeerk1XlXv/jm
2XS2kEld03LbGj8STC6uj5XDxHiDVGAa35kPICpHDvdEtSCCfI+hdiq40jp+hYZS0lBOGmyt6txT
MMN3szcEv5viD8u1XtaxykfDizN3bmiS83jpR1enmxFNwjMJSekKm/AKgUL0BqgeU1q927kOwWW9
Y0eEalPjyfV4Sk3TRAN3dXn5bb16BhYwwNfq7VC4Ml/1YW6g+riBoHJvP70Jm6yLNDdbUH/pFhgl
8M6w4WLqQ/tn2XKoiDxH8PF4rmobKBug8tWXXf/Nz3qrivV1NGqOjUvL2beNBwCV5ozzuFbGHUDQ
/no6pLM2XoPheKTRVV6oImVh4ouNZ9L7CoEZwDXSCuzRQVoZu8ax+zvuHw7E9fO20o2hc8ZWal8G
5J/cD+AauDIT3kb84Z/8DXWg74/fRC+G7smJx6A6XhVzVsxgsWsMazCbJtwd51CySfE8k9C5qVPj
YTD+qvL9pjjou2667/sbfrk+eB8ojhtJpNIHm81gYqZDQ5btpnKCXq4Sgbk1qnpwJEw+/srOQOCg
QSN4QcpruyO9pZCfvGZNIwWsQzDBQcWEumKENoySvH4QxyMcplPC44vHMoGdIG1KR35/pTaVNkVM
vs9jocEe+/noZFInXLIhtWJO3qclcBUgA+OVLtzf42n2YTvwtkRKYfxPzv3B/e8StNZLCarHXQik
ZFNujc/AP+n/9XtVjEXauGhoNJYAAUJt5x+MuClNxBchL6Q3RUbOosR9o9MaQ4QItSH+LQoYXghq
yBq7Wb4qwUhTXnWve0ymljSiJ3CiNfL3fSUBBqgMLLprIBZAY/85n8WEyhWIvzhX1ZNlHBN2kE8D
whWIeqZpQaew6GGawsEm+w9oBlq6MP99nQaw/4VmRWb+fmMBJwLaEm+p//pnoUUPpHZc2wMkL2mS
QYtwSVGtmvPGOBPU1vGaLUgcX/wQBZ5NWRT6E1e/tCLKanH0qnftTUu1WluTgCwjopOrPh7NagGV
E0/Xbcv11q0T2zB/n8Qj7pshdqifj/K2eBdD8vVaEVkiWVsWWB2EAmiwcKeXkPK+EmYinSoooMAU
g5mkU025V8jZgoA1JWUOYZs47IqI039jDJ80Fb+3JyfJ1edUCiCvnsqFwctS2L0sZnCS35JHTSN6
7djjjS378QB+awO2XTc+1yhGb+tOVaO0J/wJ3RpTCazM8Q25H7XB8NC9BoRXmN7eD4zhoCeztSw5
jBi+HHysvduc0BGdrUNbhR0ULmDLAFn65moag0pedqM6ucbqSX8ov4HFD7LOr7z3DhNF5G/0kJ5w
Szhmbvxr1Nhi9CJ5Kkan9DxQyRx8ZFyGVj0xKFyTxtcHtrXIBj9MVoUB5LNHHHnqjlMMexQT0DMu
hZD0cQNaOhP0ExzCYdGyedjxukU4vvlUIz835aVY56xPZgzzjf3C/9ODLyU4jG8eaJXFWmyLOgpg
85ML0KCpudpieXDSqtbZePgaCSz8UIJcDkwymw3j9MFad5cEcjLxD+ykXim5uLOWlSbVmvvZzLJa
/zYoqTAVJRk5Oi1LiEIJ016X2Nu98S+FTo53X6jvZSfuc7fPyr8+uowYO6KC9HXWyv4o98OpSjJR
coklNoDVf8Wfyn3bwhuRrlmvzlW94KhmbK7wddLvUZ7Y0zfNDaNHRGayal7ejMyl7Jb6J0W/YWAq
N9B2fsDNpHkp69knEpBTLmLvIZZv7gXeBbTZ/nOVoCd3dLh1V4PYED3O1GsgP6GBb0AwoIg16p1K
n0s6gIMtCkIK4R/Lemd8c31ccs+V7DlJCB5uQsCia5to7StS+rAsbIa7jJ1w4HN4iWrD6wO13z45
N3I986g1/Z+DBhVm7ItTVVBQnmyFQUq83BHUlnhyOodNOm9H5Y4RF8/nmXdm1jReku6cRGO70BEP
esYS6yoORA4E01exwADcQNr++76Zlr2PlQFZ+F63m6CLrAp7Wl25jbWPzh+34mIVwztrwprteX0e
ljyFV4NpStvehgGg3JuSDfnanJVrO0ReUarGjTP+uDxAhDsC9DwggkeebeT39yyS1sabvXZDu6Xt
wKPUpvsc7/ziig74/7no8H1cpR2ORwMnQk8/zMd+wC28wRgu/UdlGdR7ns1Dg2rfxesjg9H3RkRE
2zua5hK9gS+NCbY9uEs3BExNDzszENhQ0+0GGidFdxQXNPMXfvGiJPWzn4E68nqQrELEkr1XEhhj
xoukc/taYfBeGseoxIeNySjmEwsSOwljTzeq1PGUdwW1yCS5FUkqrPhWCF69vtREfvhERBJWeNHT
QA2xN3X1+JrIadUlDMVswo+ocs+D6TYs/Rm4zS7BUsVjP+Sr4zRsONEq2Q+BYCICfYifIvoPppbL
4yBhkTwfY6DGfHIGbOMZl6NcVDqS4q6rHqufNxx29YD5Xzj3NjxFhsLFm4RWJTx09iLCpdARj8Xg
wXKRZGsavz6wGstE0mJzVp3SDdUpBhue7VLgsl5VE2NMAE3Fv0JQ6jQDhV/3mhYgKax5HSAVCpNR
2MYtpcSPlL8QutL8o+p/frcriz5NdxyYMy78ht0rYGOPw2SQ9mhFMFp/MMiisWBiA/OgBT33ccXS
v2IKlL4t67ObFPKCV1cjFKOnUC+wWsOH9CUDRZN5wdPDX2/tKGfvn7lAjeM6Sswo6HGN54FA2Mk6
LaTgDfi9Gin/ZOKojLw46kb0RRkDevgXFXll1U+4Cdbc1WUFw1CfIfWuDFiZK2xThdhFD7atQIx1
9XClilAxzDOc0XgBX6ZF79bi0KHKRYt6WXgemMQLUbqsckheAJXrgi+IiBsrPTDm8U5UBmrMrjUh
AfqpG8NdXvcA0ikImoRye4d+a8cN+VwS0RI7SFaexRw8b29koekv/p5lb6WKRVl4wnqDLQx/f9PE
XV0poTKoAsH9Ek/iablL4rvmRpWmxeCSDI++KLMdN8XO9ZkSmP9GNmqXygNyclAZl7hWJZWMD7R8
RIN7fCyeIbbqlpHlp7AKmJQjxfL8jqZZWgZ5oGoXE9kTDdRhDriTWkgTJFyjacPeMgVk3EXon7JK
BIFqDUH140Er/HR3NPc+uN8r4nsGm6Z/Ei9aStOywJ0dLbamSEcKCS6SpJ+CN5CzsZjUMzJ/x8tA
1PKfi4eUkA4qz1AFkkx/4BjJnJ5esd4kgjr5WzJUwWnpmdndQwO+QC9PMxgF7Kaqr5f5ZKwP5H2o
34rbk9FZ2GceVaQBaIZy1gOdkufEWC6ZybUrFJ0HvHlzqvorByt+2WQl1TTGDE57CMvxskpSxg52
LwMdammh0ibFYEb9YlnTYZBYvUHZZLFEw4sX+zLZ8ZOqGNTHm7TVOroZ71KO+tbACethXmDGQhKS
vMZY1AEfY2jdR+U+bIc05nbPsfPMqlWeht9Zq5ilPX/kkwJkgkzzcwj/y0WS9eZ4Oh0B1Nf4Gww5
pVzY3XvovtAVsyvJ19bhIKskbM1mD8pZe4lhFNrtf/QfRgDX88hxsotSyyNUZn9r9FTZ/tdYzvFI
3pxnHDnIsoOOowUG33u5RUU7yLcwhcv6Oc2VeRKChOAMq2fFw8RMiFsDnAf7ScJ3TsucMGuwYh/5
VnmZd7qVdxdt0RELGNgYoe36KDFAa9OIr0++1a/bpSf8TwuOeUC25Q+uNZw25sBcVkvb2BrYfV1+
VEmqW8SG2Mpmu7EOX86d2VNSQyMRTqfZxWnhd9SZQqhdQqGWJMKtkRfbB0qSKbFTiuz0MZ7ZShxE
b+e7WJre4dI4JEHW0LiSY2oyvaCbQ+0AYS3vmHKjZdHnkALTrSG+VESTvDVqtIXitzJOI2Bj15zo
u0BC4b13GCGnSicq8oT9fK91fcKZE743ohKitrhZgODc4ThFiNdYVki6iiZBwohxqrv/5GYb5aoG
rhqrKqdjh/v+CqlvcrcLcAEYdx/Vrr7j/FZBoykECNyjjARa+6zoGFFoi9ip630lkreSfkqQQBsR
yKTgISfGbPRm2w3Fl7BrbrorfOocectULDOgxzpZS/e+GuMZELdH3k4quBffWtI5oimUYv7DMaeu
oe1eru4CQIMB98QBapf63b8Scb3+m0zVExhVcx7aVa9ya7AQVGSKFv0l44b7A918S+O5j+D/mqrw
l0+4Pxixbtf63R7nfpOZWVE45L1ZL2HAcPWVZyFfhaVZGXxZBfcKdhP1T3pcqXfccS2J8W5JLzvC
Vk9rwUZiw8tihZnUzZAqm7IHWczwZLf85GpVsxmCw/hGxO5cARM9qwXnLrD9p2cApSIiQP6thA2i
wQL3HolGdmylDeVeaEZpNBHU+FS2LESJEuVuUKChgV6oKmfEAi5sZIuyqynZHwJLL9bIsI7i6bFc
KLcFBvlNFYOt5l9w/mTxB74NoDBEzXd1/yi4dESzsqDb5NJrS129gYMvu7uY9bPRoYZ7lZnupQdJ
8aKrV+pO7DInFxttUNcn7JG/spkpYcMQ515modUDvGNwm6vYsJTgakG0rR2UrnZuZTsOjf9s7pTP
XBHTKhDku4grtAO8JgwTqmN9zVw3Od0NwgD/JFHV5w/tqBWVG61tNQ70JO/phjnTLdvAP3hjhyEf
xZn7THF9i5V2JzcVV5XQBEtNEAHNPSXYtDFqE0J0HbHlLmSs5P5KgPt8ncpaBpyIgNznXTXGaNVX
qq+wCxh/KbNmVhvpBr9hUzNtRxe8Kto/5AI6FRwTtd7RpPnZC4kFjBZuReSz+RkSaX2Ghtd6112K
NEhRfpFAWha/kk6n+0HzTKydDaJhK6M1nQqGmwKjs6IiXGMMfJ1BYj3YoqlAAGrZamUPaLJXr4/H
5vx/zJTow3ZA+RhA16vU701mANaC6ujLXXUBugRL+IRTP1CVa2niPSgnQtmXa+hUczoeMO5fhntb
+vCgUNPSPufdP5XZbP/f9Q3xpde2M342aPyRA/dzKBVQ6YSGZSl+fq8CygWRbbLo8rfsurMECcaH
EmC6qnM2iwQP/FGIagPdsmeaaKJbHa3zvn0gQUAgNNw3WC9mEpQOzuTSQv5A/deWLmS1U0DNqf9N
3vr/lxqbZGbp0LzFwMWxN8HI8WqXpYjLA3K2BA0Vhdr+Ebt8jF4H6WDXgkmL83kkpbyG4JVgG62m
69PehvhdsdZB/a3ZQtEGAQosDpWWGEaAhOyPU3+tbHM5mbB9Msowh94mAUkoaOAEZ2SpaAkL7a7v
GOnQATHsUmkL/IV1SzcHB9LFqdynQYB4HfJeYuZ9sYoSYYbadTRB05ad+AWUEatVGYo+xLwdaaEd
E0JTUypmAuuVvPhBggYnyJGdt2evDfyYMB2nvnZqXpwOyXBUnyoC7QhG7g7yggEeRa2LTVEZkFpq
kVaHSKlEPsjOAghrz1uRZQ6yxwTwAxXvxNLkUMDR2Fck1vAjUvNWy7IeqnPcuGg3djcwC7tM3AIF
1qwc2pBq885gSRVaqZNO1xwLBJZKYmzEO7mCptWGT6SLjA5LaawPX+sTgosbZjZ2osI403uXH9tT
GFEkke5GlsGxzTC64k5NQkpzukwxmdesSdBuWbJGYXNI/aYRjK8KJILJio5LIHcn1t6Cub47F9YW
8fYpuxOIgplIuz81ANVci35yQ6Th18/yb3B2BHHTXH5KNrGfCOJay+pJO5pJtl0UwUvL0JRLgeG9
dGGcbpYQzreR9y9CzeE4AFe5gac46rF7+3L69h4RTwC93U+e8mw8rxEZZkgRa4wyeqb2ZRAJcbX/
VgtmSp/Y6Xm/O6+E02VOBIStnVafH4JCOvx3BNsNrnYeafdQLdaP9kSMawtwc34+UFQH9TSPnhp9
VKZ8i2VjzIHiX9nUDOfi+1H3qkWd4bpTYKu0IsbgUcUNU0t+QNaliqzmbNYktDZBU/u578BqMSBm
/KDDS+C8mUZvx7gMLRQwuok2rWDkxOwD86g+Dkf9DdlJjCJWjypWCZ/Ys+kzkguvWvFFuSXipMEm
ZJgJi11c+LJg4GNqe5rCJQ7t9m2Xo370N5nQBOyNN5LkF6tEUO7/IHR8++EfSXszfz9RgZGW4ZJe
/0ARrzq9AbSZa/CBk2ye0kPr7MyN7ATbZ7+ZrEWFPD72MWYzXhXIcBVxhF/w3hRIOFocRBcl8NJq
xDoeTzrbmwtCRJqB7utszVo37JBOxLTqxoBhWrAp4ve3iSAQOdRckFBn/heHkdzvqMYB7JXC9ck1
P9RrnTmvelcZKqYM8bh8lm9qBP4Ayt0BlBmbtbU1++jXHoijx621L0ocTqthCr0SP+AxOdXB46UF
TjAplP1EdAuSHvuWdl2PDGbndX+3GRDiqlTwNGnS7xahCjCD9gfS345bb/w6azrkX69pZnhwHqox
Xp3ofoagh34eNp3vBM+QHFIGtZCLgUIHqioQa2+vKFwaav0raRESubYCdtuIxuR7pxKGbJqFXsR+
aoMvHGOKsEW/9Q5Q5k/4VmSzu5+6fNAi5xjZEHdBfHSP3uoMGnXzLLpcbEUmkXVDv/1YT9JuXKa4
/WzMSn4JAVJISlQlLJtFKSy2LwZI8eleN2b95nKvtLO5xZtG57K9p4LD/cYA5B84gDE6rnWYd0Sh
MCQmosRR+7uMKwk24cHINdMSd2/WIy0Ziwqr96sZYoSaIg+wBuXLb6zpoGhKB6+2yIyQ9kc/lEzy
mB3eEDTp7aYRcJxHmUFBuJEbrSiUtbOYED7LjM0iMTU1Kw+vnAX7J8ccIPbKxBHgcwcrFBuO1SEJ
bU3h6HbGi4SuN5W0YmpHrKqmg+8NtFYN2Zdaxp05EblfcYD5fRjHCy06XVOrM44A3ttthpSgiTqS
iNYftwfLpKr3JmiFDdpupbNtRTXxncJurLhsvhqjc4U+RSKot8op1wNUZ7G48hWz5oMtBNb9M855
U5kgb9mbYnhRVsXz6QOAUGLNo3E/ChDaC/m9SQcYUWZOz5gfkxOc9Ibud4hMfEPJoOjVAoXFwP7l
bltkUw6UPoZNPHefb9It3sIgiR2NE/lvc3rNj0t27fFEKk0ewya0+wY3Q0FIM6Q/t3WEir3LSVGg
SwxwRmPVPfVsG9VGiDxwaXgx99/Jw51QzJqb7C36XOwLR4D7NT/M/nUlZ/6XtG1F3mlg5DEN8nPY
4TJwiJPO6faNdphhYTLIQmrmQ53oWR1LMJL49k7sanSxoAXDGm1Ou2J61mNW+shGQDjOzkqzj8CU
Q/K7P10azZ7FgM6HCmK2QnvUmkK5/FcLmsu5QdxFmaGBz+QCaVzrcuwxSO09hdgXUnwR+9tqXbBj
8p7UiWcWlVVaYvZJGHFabfkYASP16POUEKtxuqoxthG3sZZ/ShH4ptmRtnvhQhDuGMUNpOj9TCRt
vZOy4numSY6S/0e089a//I+k5lAv4yTI2jvSKoPICksWiVB79eJK7WSf+t9DAxaOTQXLIeJqf+RE
DFU1uIajLl+ph6TUuKO09LbwpKbfiHcBLLvN5NTgWKih+wB10RcZHxu1zUj7/6K2WhJm3DUZJ1yG
dDdkJQSy+9SNsSlGR7VMWFZciYEj//gkV2vPPz5KV1uC+k1m5q2eXuuGa2Hsq2YmxjoiDy/Cjdnc
+mzk14x36doTABlpD/Im5gE6PmQePlcru3gxcggaxgnFiYk/VdXFj+lJIVk+fDlZdIXA7Y/S1WCt
J9zZYodLtKbfcnCU5qNgFdfjsLA2bCf/MDtRFM6jwF6RpD0Ojd7cOcec4WDlRNA5l1S8BNniFmU3
1zKqYK0kpbe1hl/B4MkpQZ95J/74Fan8oXs7UlMbG8oOlN5kDUF2FppgKmEdiB47Reci8gEq699r
GShyhxXf2jBcEsS95g3uS6I+OCbAWPeIS6t49JBmNdk66grjVxgLVxPWWcFbIPUmDY/tmZF+uTWP
jKfou2U+qLul2KdXBl7AjXMRq2/1bc9RlLhgnkfViKtrSCvqX2OzAbLjpEakvkkbPwi4PrOURGO2
+4Qx4OzSxPBuYSyEyQdiKRQLyxD0Ubwy4gtYY4rhWIcFhzlBbV7mJqOhhPVNRNLfkmXiQJQlGtLW
CMrFUAsI31AH8jl6qkq3fv9xyLpPWexEWJlkYh95f6KF3iSh1gIPkoYsxi9e0q9pXKIGxdO4atkm
C7KhNfJS+fsvx5jsu7YFSAANrsCtGNhwp0xx7fJaUhE2+1EzNj/10qyKy0xCw56VtnwGgBH8Wf2B
XcqP23+JiePFo42n78URxQP4f/hCVonFtRN3vYv204/VNfiMcq933aP86sxpoITEzWhPN9GP5c65
OJ1qJ2DDcnUe+fkBrUFZpVRAqfsJxpdAnJ9tKjmMFXE8IJoyYAilXyI0z3F7gjBuuKlZLyyNNjjH
0eNYiwkUPtNmM8OvAxE99tdLCXQDxvM/vbSNAN06P2NrgJl7zX04zZO3y9acLYRjsqVgI0yVZLY5
VC5h2ybHFHuT6HMbE69axb+Iuq9+gZxXs6clDO/gneGe5tkja7Pj5ddjP8lseIXL2T6NNa/5Upe/
P33q2Q57/1rMZJ4hmeqm8+WfUADmCIrBBU7JheDQS9iA6KEHblAmsC5Mn9rgJcQSBjH/M2D3xUzi
VfzgyuEaoGNVOwqjbVucj+ByGJjy1IMGkKhthhjHjH6BwN/NfT5KgTq5132aEs5ou6x6PRl+C4rW
ZFCuQxDJZutMoYJChXwQ4hbQ8Qj0aWCWRNHYuO4uTTX4m5J39s5kwjPYm8lSCOOSCIJkJXRKzc/K
63ufCFIvBlBS5IaBMoGQyENCdjVcRz4SNz+nf6Kcq2uYxdF4E245Ofx7Lzqp3Wzc74czsjMAG9XA
p5LDBdzXbBbAP6tA+PEyv3l7BqPuk7zdv7QHdihF12C8ufIYcoP32CYI9Qdb+w5/3+dbUMxxC0hB
Nm/W585Oqi6qXhWloR5/67gDY7kpzfPz8jRlCT7EAryN3PqQqn9SnSnKD54aYwsj94BicmtgQS5k
hDGtlcwMUo6RlCvJJd5uRcklRiJepHdxuEQHp/GkSn8MtAsCgen9ENlnmhqjaEMKbbvaMSX/seFu
erpGrW4yLSsoCsqFQg9osm5dA2i2aSPEyJn7Kvos4AP7ufoq90KhZJUj+IKmrqX+XmTrJrAYZZpZ
dEfMm8BjftYTUm6Ea4gbeVmKTnAL4wm7x/CbhSsMartvtTeSEaJDSKJ/QuOTRCJ+DbcgHtDcFaFM
TdauCtYywscu83OTweTTpcw+i0GnGFklfTpTvyczgIoaqq9dvc6LoZdQXzVuqa2g4cb7sOb6d6/G
aKVZtUQC/SXgJxTLRVq5MlG/rWaJSfAaI6DIUMXJgZ6QUpA8uJ7o+ftlD2K3MaTqbnaNrpf1h5o/
Sd1DCK4wZ9xcchnw2tfjJ9FIhVNs2afvPnOjgQHIlITsu4C64Gq2hZ78opSqJGIcUgrQjeVc1syn
DRoiAmOFz6I/eeKpgfgxzo+0ixZHN/PkkHv8F2V5Ai9awlyFvgw4Zg7SWKUGqQfLN/w+pefgkizn
hyi/rkIIlWU4K1OrL4WkeUcw5tLJuLRQMDgwBqJ0TzFD4RV1GjkjjvU0EaezT1Rtu404GMZ/7Jaf
mwT6D+kH3aqEBu6G5tsW6Zgo1I0VJij9dAsIyXh3cuQPch9N2Cxk6y1Zu5CRhSKA9YnPMKMS83Db
jViOLuQUiyv5MPcNK3zUBr+LYc7igF8WYGsFb65ejt5ho0QI8UV+/7fPNhfDPaOGXD4zfW1LBxU8
57pereghonqOwL0rMniergCvCJ6d0UsOiFXeomJAnt8J7IVldn4NbmlL6OxC0PKAiLTYVhgpP3pL
mHkVtepua4JwnP+iWnSQEehF8MmeQ2MVXt4iY1KUCnwQffDu8JPtSk8htFLfD0T9Sp7apfuDSvnX
OTHA/5RLLuHomG5FGXf4Bqt1WzX7SKxn4+TZxtipfoPZsLkkKEKOUPGt0lZl/M2S+YxP4K7EfNWd
Xbl3LHOqgL2lbeUU64zwsBbdKenGxukQHiWP6VrZaoTgMoaOWTZhPCYTQh+k+0LbAa/1Ot8Mdlgs
FGQXPPuNIwuh6cegxz2Mhi5vfZ3R/6uC2zur6XX6U2lBpq97kNZgnW4kulPkqNv3qZJoFUZedE4L
/x0tp1ZV+KdWjRMgHNByTWISs4AVW9EY72tKTFRiZE/n1Unpkr9KRnpdZ/47DG9nVfmhy95XxgwV
Pnw2uacE/4L09IGI5vJmH74UgwXUKWtiKY9HyOAJl6c7caNoOwocY9FSu7o/Gg4H8PiFHTyZhlbG
l/cV2ZWtdyglpVE3SoKPbEKIqaTm6TCiDtjd6vf4uwhDKsiJWwA3ThdNWTJrFGvI93/xKyOVtnYq
/z2HynJFtGv4VceSnupTFkfsByHVUW/oWXiNakSyUV+4++O3uUqDpmtx0ydaukrH4TV1Sa0Zvcgp
WUx/Pi40d3tOCOsBROjgA0iVp5TuQFe7TS+V0WDIiiUHKxRakZGx4Z9PvFhIb5J9GfMV+CF2Re0/
TDSFXgFdKQc5Rr7syEfsvx3uRLNK55DWxIP/Y2zQG/+2jF50HmDRA5mWWA7sTyKO+ZQsiFI33uXe
E4zDDzkLM0MuNRIsDEibW0DhNStcMzUim+N5oi80hjli0yE0VCvOc+1rW7eSnJBGPzEGI7RyJUIU
W+PYcdP2WVrXe5P7lHCicrNi3ZzSXgcSrCw21g6TdrwwUW6THvguTT+RxyMb16ALa/zw9bxWAhvV
9oGJbG3/tCdiW9pOh5j8OIwP4Yl1F8/MhA+Y5mGBITXjh222YQ27Jww/iRH1tjI5Vl4ENt2KjYld
8jvaRDcbDe0wzEbJ/Otm6SNSjtO+DEp9KiBDCJ8ClcJO1Hu9nyvW/IIymu4n23Wmpv7l0KEL3BSB
SPck/gyc/rlDwRuBz40Q+ECL4QDQnxlbrgJbghdoDnM5rekYQ/nZE1lANqMfTtN4otvfhPPXeIhW
IwILCSBtaSBUqOd67eUv5dbCJWhDJPoP0bHz7pWKUFj1FipHMCs3RYx31x5W9M8Nok9W+LYq4Aee
eho1OxzLtUj9c/upFx1WDwAQBn1xODmJijQWmsrzIWdj0iI/yhuVtpGkdcmcjxemmM9HgdlZc22y
EJ8XqrsiSBvAfzhKg6qs1iZ5pfWC50/c0h8BEDOKxYK6k1f9cjZILhowlc8vwZkG+fPj0TAteSkY
9Y9EuAOmANZrGCGkdHPjsBSP/FzOljR4LtYjcPYzpjLofFBY3a0HomGgOhNoSNmIn8JDXyjh6NtB
+6Rm+rO5BNKdWXoN/7/j5oWc3uTJCzRfP+i/gRuxgVadYOEwlA5Jj8nJEmId21wc5bkYCB61dWju
CRHYedu928zMMhKCsDQwg6ZMshHt9sh6JwcjwtFUGYMEaCgA0tTvOpGDhuIBTi1U+4Cr9JfEHp5E
PBZB0ptf+IGedo4QRaWyVPdjXpjdqix0VMzsUaunM7EVTxhJwyh/fjUljiS34Nznpm5xsQPsLPbN
k5Ws1TR3PA/ja+WZ3U/ciwAix/UOwbMOk1anr8NvHlm/56jDRM1nvfrc3UqalO1PiXcBj2aqUcTq
JUwW7z/5h/ca3DbgXvdvmk/1KG+dk5H6lyaTSmTMkx0Lz5X7t+PRNh0KsF99gcNLPSMXBLdQb3/k
s+gsie85CAgmLmqmaIVjnwsH1hI8z6rNduHp6wERprlnZDBebdN0t68Oau1hWGJPwkm1jFdIfyEK
kGy6A54QiNNzmZUupkwcQyjGsSzKTCZOyVTLfrlR5OYfSCnku0bN+v3zyFTI9QPRRKc+8ySAG6Bo
ypGePRd36L6vvULMMCfXAIVO7D2zCXfBqjQUXDjVSWF8Ne9a500BnYuGCD6LXPdxq+EvdwJ1caA0
9FyKMB60WUOCDBiggj67pQ6CgPmMAYKikUD/yk7S+p1Y9oeP/0ZhCpwjiXsFV1QP7ToX2QSEz8i0
fUhOxCit+RDQypQRiVozveWMnAU7UY0r0Mv3OsI0rWE+goDoQDcHWm9b9pTcylADUaU6o/fZ9wBX
2xUaZ9Mb0DQbJ3BHVwk5SoT+zZOJkC9t+xoZPN0oiOQqwMAerVTlpGCaKVuqHOxK8eZxH0UISDxJ
E+w0G08HSE/dcicVPMVb+GC02gpr7YimTTzx2bel4ANies6uXX8wg6eoa6jMKlI3NK1vOL3VWBIj
9T55mdQ01zJ1ix/xHVVAKZGDF273ynm4v0FYK1N9lmLaWW/RTZMTbBl2VekW1pgK93wF7QmQnXJk
z6tZ+9S6Ftc0SYCf0SvHhJdO5td+koMQzgI2bRpzXW/k0uSByzbOKCg32Z4ZOhLlOY66VHqLupiJ
b2VYqVl+Bg+idJ2lELEXs7+69osISVpaZRyWEkfXbQWh4+fSN54vQRQ/H6Hf3IgH8E5daSzNR8gP
P9ltWcRJJCHLNv7ZusxiOhgm8FILxn+CN2w4cLvvmnijKdAq9aw0rv41xFh/IW1hWAudmWB2RfQA
RYtdKT30NPSgRCGIZq6kc1dniWWR36t/EHK16LXyazd/pSykfPahAKEdKOvcKAqLqVfRh99b8phS
HDh/ofjkFuprGiJkX57ePdNHSEeBAbivRrOE6QpcRAOLz7NKDo/wXKu0R9jA9T6LadlBkk7luvwm
qkCR5dB6ymjuuAiy9RHNUcrRHCyVxYDP+DdADDmFTblgTG8KxbGqEFZoyUAfx96JndzorFdCbdvy
HRim5RrxG0oySuHGQbMpfRCR9JW6zSM4KcHAy4U1R7EY8CrO0XiNxvVd7MsLUR1unQd0jr4cAVyw
sHibAa7Q6wDK8l15mFPlAj4f+azWKmrkzyiHUHICpIe9kpmQsN96O/PNjY+21IMI/oHiBLtw6FD0
dLaAT2ye2C0mxqA7m8h4Bk7hByDCEtzRyUyKsRMNdXzybvCYC1OnTyYtl4pqECVcZlkFKxdrcbue
B2xp5ONgPsG+TO1YeUKMCVchL7563Kg7ChiZyv9Rnl2GiiY8gZkIxupmG7D31UZ/UsqJ9mfx+Umt
Gix3iMiD1VJuePy0a8USTNNeR2AMcAjyivVIHOHoPpMYxOlUZdJwYs2cJw6hx5d4AH2U6FWvq3Eq
VZBTPoyltUL/SUOsEuWGDdm1DOoRXSNqvRy7jORhfUUDI0XOaDloRp1iG6Quhrz3R6VyHOa8Ar2m
xy2Kt9w410c0c25XtF0j2eBRvI+3eT8sO7D0Qv0TmekMfNsl28gqmZPAq0JjBrTni7Y752tO3hVB
e59JWS0sZsglVMgS5c/7IC81b4ohwh16xw70ayrWcyIUyEsFgqezfxoS1p6lxaBN1aY/O8i55tQp
+PgiZFyju7sefu9D+bG8/hKzQchDbHSTNvy+9kGFsrMSaedfH7WLdf47ctwKDCTeDT4uDrCWu+lu
yFFdwoEF6FSAZOm8LUnz2mR5ZQRwo5BDPB3K5psnNSf3oxGjUhkf0mNtMGVqVYByt8Lfjgwnit/b
5z0Xt3IIB6sVYjNols5dnh+80Lf2G99UNhheRiND6F2EMU2wGvK+p3r4NatzLFSn35JdhQlw9r9+
iitlR4Y/0bM7dR6NkuDgr53mB/pkQbNOs5VNSx+neWpLzLC09DXY1l22kumCMO/eEJ6SW/GEh9B+
JzsgA3cOgVwJjQbFyEs/2sJYS+TFuxGv0X49xHEZ/Iv+/ffYHEP/XvFzZiTShIUp6tXAYq7A6X1F
HrSIOjlJ0EcRxYlvy2YUtVH/ZWzDZ6CFFA8aH6AeVhf+Z/pWIybUCHcGcrZ2AX99omK90ijmflR+
y7Qe3n6JJlSw4xXCDEb5qmwS0S0opu/niztHRvDOTeQo+Or0M1pUo6QuOxL0IDuBBLliPCalgab1
FQXtWS5GSy3aZTyXUmDAH1Huo0C41d8gnycJ6UQdmpAKBVRod7xQ1Qj3UxTAZ7oE3k+nDT9LEDeG
I1w4YeiQz9OKGt7be13CmKSAl7H8wdoptogc0zgpV1ovk5npLpwgDSEgUUmreuicJDHrhF/9vxZd
qcRdCVvlq1LEwAQ36eyG7g5GfSJiAlrIcDwhCg6QRcHBsJqgKHSs2B0rlIcV/aFVIWrChwaPVpgy
8iI5jI6RBmrf+XKIU6BhcPkXIaiI3mO21jHKSHvvRHPVpHf1SIuSBF0A48ExCy5tgQzmEGZgovDJ
764Vr9SxiR7n6gr5M48U+hUDppAYGhW/s9ElgduvA03DMKLAHCFqXCAckUMh7BkZDSNRp1N42Kj+
a6O+a4eSghfyFjCOhRdzugaizd2K+nJhzZ02IwB8OAXsiLnuSf6VvXcooSU5qipwRQLLuQeCsUai
yS9P8NcyneX//qlSGl1b+r9hN0k+jZyul9bQNudi9Z3AwGirigutfmBfLM1zvSuJg05cJg9GpwkB
10Z4AuZJ/nf9iHvajs+uegxe2TbTrOTFCYCBCxS/EJN4duKXz2ikCUWKhVjCg/wmoS4QEbo5d/nn
0g/3aJgP9ixIX2eqGR7/Vq69j6dlLXpl891NY+ePQB2L5KG4zYJHJs4AiK+UUVCfC6nt23PL0YrS
UFfOOEH/SwipEUmI21tyl5dKlVXhtcl1Y8aMfh//+1cCEYXU1J6cHZRnRmUCy8gWstnuMnFc4lme
iYtY4djgiQlcIdtyynWImMpwsHllcpzaZtgeWppp6Vlte1O79pNabm+vONRyo564z5JJ1JsOSQ/p
LhPm/ZiQsNMBKAitQ/gBX2bLvPS7980GhiOaIabX1qsf47fmV1T8CHVMbYgT8dTQ8nsQc3Esijh0
I1Jyh1qm0HoIR8Yhwxjv9w+jsbuDjJ556ovKrJ+W8EepU30Pjn2XFgMUALAXaAlaJ+RlfMQJXT/b
WCKrxY6sJtNez/Dv2YdRdED/FXhIfLsFp4rY/ZYQG+7XGr2R7NWd1DQFayUjDSwjdJ2XvgCZ1CDw
EBfzQotXmZlyUAOlD+5Poyln73GtsrvgCarIMBliu7MEnM5f/bRWSgoWRKGHOPl6H/yAUq9aVNGG
jfmHUUI7GK5Wa9LcKEXGKStsZgs3h79TJDk9TpeXHhvG5ueFrmWW2uOP2sFJhvNTaVKgm4TPlFvt
XZhxq+kfC9VemId+FEtw9jkwJXGkEt+FDx2WYtnN2Z/SnJxQez02QVK5j6E+SUO496EbaehGrAux
sQe6m6Fokm+omC3E7466JsFjwOcWGikv8cgokQ67SJYC7S7hudz+oFUSWreILxGReZ38U+B/3gf9
JeULQ0eOKwkf+Ocw+m9yL3ZcaZvA30SudMDSCj03MCPEnqEQsUqsZ7dgRkVSqvADvsg45C7sp+sB
t8pqkRi3LRZ/HN6N68tbmaXugkaRoEU2+9TVcl1CG2QsQgkzJheD3NOE5FjADXWpNMg9XwqQp4pu
Y81aHVLCpkWw8NXAwlR03tDgWIISGR3+lZEDczV51YHHN7ztHrhkixaSUissAfVQHWLpUXllrVP4
3ntF5uckM26slp3kTwuy4BxEhByEbg5fIsDHxjwoT6RzHwKp0ydMYOK/waHPxImkZ+0fxJya7z/I
JgGiC3inCGEH0OGN+iOxiofPDm1aVM/hQJnli6JmFqk24BjxO6J9ibXt40Sc525BBNYeJpl6pGgn
xOvBBc4wHG/tnN8Emg9BecrKt4eit2r2DmNueMioY7P03X4S9IQonYl0oBB5cvBWjRZO42Qf8reF
AFkhgYF97tYOUHKDuMeMXCrjIBLhb0MXITG7d9KrpBRCSNTMhZFegWPozQgtmliL8X3OPDQcMsfR
wbNjEhovzsNkxhnhg7DrGf5fRV78drmexiwD3hbiZ+WJXyvfjnJy486d0tAXha9cYvmmE/XtffCk
NcgvA3KbLTIzvWCe/kLC7gnjF4YTXK9MUk7zgyp/I2gWrnPXxwoP/aZOoxam5QEIK84KZdnCn6Kx
auI/v9S8hnAdfmagb6jRlJ3sH7wAAQkR1Dss7LZ53khlzTdLXhSj84F7ZDhqa7xJh+lHcVUqcqZp
CK1Vs7APX9+NwTBKwGrba4cjmY1DR+rJapmqw0u5XV0i3SsacpbrgT+pWrWvw3QrFL5JoU4BL/wk
DIzA34L6US7ekU/hBRV3BBKKQiWmhYww28HXBqrbha9wCYJnTiVHdgd+klxosBGits1IbHItWlDR
NcBvaQV8lrq4mU6fXVYzL+cv1lzo1mMJcR1Qd2On9jVVMbsyQLjG59j9qMozWPiFz7P0BEGkN6/S
N9/QucmDGDiHY2+MTJJg9BRkYGMmO0+vMFiHwq8ZTH87EzQ+hSzedI+SAa+mFKYz5uQhOlRviq0r
Ovc2/08btgYTqeZduBRyh0X/uQpQwMD6bFWmbmICoLZUwfTWaKPLAn5jsiPaL4CIeSBzpqzdwlHb
O3gma0D8z0kzsnhGa/9qTqTdSIYqR+hTKxvX4rSZEDRgAE5mI+THpMDeDDawpBt7hhzs9T+DDot7
Dhc0DFsj8eeaw/Uuz1+qqB/ITTkZPc7lB3MxJIfMCHyWXtts53129ZdeeBCSwYnFBpeLPJSf2zkf
V+4EblNFohK/GdQUi+tWVO1E+ld0IUNjXTjpqDrCcceQYljcqR4IXIi7FFcE54Znr/8ktpgZXB5k
GwGbJ3Q3QA9kS+tgBAWBMreTFj2ykbz8wvchGg/2ZAnN1xIZSIbApMJEB1ImWmvf/nDOPrivar8H
YnGmu+izAvj83IPsCtwvsDnsTXxfDnm5SHULV//5kdMBTa+7bA5s+6ieCR5A1yledWi/dv79c5VU
Wc8KLOjiXO8A2AiTa10N+AgjbbShcssxaTZ0x9zd1SqJOsN5+1vFscsE8+OCZxn8pdXsqTx/iTDD
kBzaktTwKoyn9FQtZEua0sjNhBNqLyjNvvHNIVTjtZyWK0cJ1Dg9xlNlbKSnWSIxQSV4i988X87w
hg/d+5WZ7CdFpQ2fWvXwt4vXrvqs29dA19uVHA1t8v5ypnL7He02oC8F/1eWt0chasQFPJ5nYTOh
jEdrIbgKUlgw/xNAtMH5tSggJXXC1xyUgwp/j3JL/iJp0DrBhCSZRQ+Xeh+tYzWj92vvLGozwdRz
xG/e5vUZct763p25tZMU9+86ckxJnCwnsmG+Uue8GKfmY665JAv1YqgFFFoTVmUs8Ob8GnoLD4T8
EpVDd9UdtzadpV81l1VxG/gOf8RqM1KCL8qTjRwVYoitJQSCEURs+4/ZsODuEeTkIm4yupMAV5cu
/OEr2K+gnql2td27m2i/K2Ntgqq+eKUqvnwlCO58GttjMpJ17RPiyZ+EDwCaeKiSBo+0tdFDngY8
054QopSgsmiUJ/hS4FbO9qKkOasuABDY+OoRIwsjUJgHvwqnF1sBUNlY/OWKwUVeXL3YT5gDn4QJ
JUQu5GJK0sMYtZMX7eKvpLve2JiCQSRRsIMbbhpVKZlMXvriGuZ7nRJS3Jmb0pnnkFh4PU76HXg7
wBVo9tjWcl1Kvj2kOuhEkfOfa3qImtDXGDhJT5kgj7Q6N3uIj5tbp4KXTAHxt4IFOhVSTIi2iY38
Evfn4k2+a90+AFIWcmQrmxHgGZhDYIA20L24bA0NKXV2a2PeCEUUVWqgO/ES5SwMJMo7/AhXYNYa
dhFOT46RqI2dbEOt29dt6axb96JU/4WAVWkV5huypU31Q2JpIHMMmGTCByt8pvitanOFWplFyf7k
aZxS/IMY0aECu/pCePqCJ22YhBk4P7s6yg60RCXjj/mgGsoJMHIxosRR3Ve7cQGeLTpTakwN5Yxh
C9Bw3FWpyPoUuu5iuDN4ILmRKBQ+MVmrVKMgy6Xn2qGLTO5vI0Ai2Cd838sGVHsvoROlrcdApgp/
bX6r6afOYl4Q8OTlSvEg+Hacl2LGEY/hP+LbxO515oU3HjqalUEhhWLD5GjtzLIs7HTcwLdBrqU5
A+jQ57PiV0kDeJQ5anKmvKk5vwp2Pg6lk5jnTZwC4YsO1+3yPyvstaLO8S/bbmpcIo7FfGa0BHFm
OKTO3sqosOH0VP3cZczrJKegYRJS4/CYX5hLRXKA2df4FIfaRVOlcAw8WhDa9q0PICvOLHxyECw0
MlRH31lkY8QMgXd0NGcrPoGd7J9yfUM5wisF2ifDpYZ3mq/C2LhqJTt48/Aqp3ju2/ug3XT1/Xwy
RL+Z4wf+c7NuYs3vBC7TpoV4kLSKq9cgoVnudx1ykK8lId0dSsT4XYdTcn27bNlRIv4wS5B44RGJ
j9zByFFhrxPDqGKfW7Ov0syz6b8Zp7NSNT52e83BKK025aih9sW4ZP2Voa2fXqoVceIogf81yD9s
dEtS3D/srgI563yxGM18+4UL37QPRvSnGC/pPs9kpJRxGjenHrx/78P3Hy3DuYdmBq9Z5lividV8
YPB3iXeWOcOXhy7sczNhKY1gQ7tQMXMpaFyai1VckGJ6UtV2p1n6OXLKA60kGEJhHRgikSgiKcUo
TXOpIjNQ+7QQvZOosm/23JGHw7O4zclPeGpAX3neypwL6UGCFopa01/GW+x7ccsnkkmmOHg3NrnC
QOuYRl/CrmGjKK2bS3z41vG9KEtLTti6KFB5hqufUqnj/OiMJMfXwk/CpQP11qNYzf7BH5eSsiKR
3JHD5YzoIWAu0X/GRET0Gwiu3WJaDw5oo8qCITj6iORx4ofQ1Fay6dPOdbxSXX5+t27N3S25tUbG
APiDeMoPK/wjsQIRvo0poXzOOilSk0JlPgIzogsPa1PVZ2Ro3vspkiu/ufqG5VWkwM1T9gyYtY0K
M36bmg/36OOPXYPywD7WHyvzSl89lD5ZyQY4aFt/3f9YnWPgBtPfts+4FgzZsVgIIOhY/EpAj+of
1Ahu6fi/Zg7NGq3JE6zlp+BbEA7sZA/5Uen/pZKUE8C2kBxOQ84z7td7KTrteqroJy75Kq5xYWzA
Kqa6ITPuUKOPVeK/QHkjV1wGBmcFEl0mokDf9/hql0JW0NiDAZtLm2PpIApyVkehzygZbFKAVv+M
z/LeSdmzLbGS6I/7qHGJwlIgG8RtLLeSMN9K/XlsIrUwNm87Ggmlgky/4Yg0h63LGBst6dnmNMKU
U4mf2tgV3wC1s/4BXSgmzYR8NvMAH11QoSPFuaaATIq1O5/pRofUgia80RSSAkWEBXlRrTFvdzUw
ahmStIuIVJnL0oTBZNRpuEyt5UBVuz1G3BefHeizdo/0/PSFlBqI4BH4qmfTPAIOjHaj1tlHjTj7
v2dibcFgvBU6qM1qcsEcQ5v8Gk1syeNZLCpnmo+X944Dv3OE9zDAZMOjLzvlQ/UY8ntaB1GN8RD+
icACTDd1mzkRrrBxd6xkjHt9kiZdIXrCDiMgQxAJNUH3IFfEfyYLF+arWDMiZ+h8zfl2sl7a89+j
h/WDAuJB1o0VJS4tVtvHtdY1gAiEtWbWrBiP1mHBt7DdZs6Hc4Zwbc8LoClTY8nWDI3b2cS7eZKk
3D9VJRnAbk198w92mCSbOZCrg2DXq6rQSrfvxl4weWkFEEQ7unlYLmNT/lfHO7178VEA2dd2WwqZ
yxzn/crMV8KIyxthd8ilVb+BcfMWKPn/WjksVXNWPnJjTk58wHn1sNFBKeC1qQdbKfQ5rgm6KTmP
HKeqkgG87gpEGObaY6laMJztFzL82eyEebxzO0rlhNKfuW4OZC2y2zeNOww/btr9+4c2m4hIscGN
42VnLvbgs8jXi8tt39b/eR4j3tuSz2ZSeNcwhV0BdlT7c14HBn9HAS0nyqEiF9uGBfVXhbhLkNWx
sLRDTbL3iieOw3dFvExTbT3hwbk9wF4vshPC33T/owXwe/+3HoxorY7wRQdkZafZqVCW0PGAtjfK
3UAGoHdV0wSfaKz06WIiW3phzYQy7CRMG/OG6Gm5W+KXXhrbpg2O1e2/bVQHU3dN8aUlLlsSgYVL
MqswS0to8fIFME1DW8aUCFGfd29s5kodxWxWKkuyChPoFQ0lTav+o848gXt4A2J9v0jCf7lljQ9n
GCjZBeRs3u+hafjDs7YGl6kjSFDqxvaSJTSiKvLEYQ8IdmOY4XQKPHjlQwP0sNSFqEA+2bW9+EyJ
1oWrPkc2edxe2nHmWJb7Ou0EosRrC26nu/pIk3HrtM629Evvr9PPmVTErhPaZrocD+/yl5quXh/m
6UGJOQvLYRinsaUZjs/wov/9pYJRY8Ts285wMH16wGWeoOgqpShWdeHaySffcvQhSdNlQBEJ0JO5
WV6A8Hq2mynYSBILHTNY1mnRlqw7uKrkaBKZ9VjGpoV+GDen0ZK7zzpeE9hHkOfy3twqbaPzjff5
Lq/E0QyV32W/J8KrX7waFFpaTMScFUes8L8v9vlwc30uapXaKCdYV3rjSZgdhwUKOOonghyD7rpX
D6fsyzHoTMESu3wpEaOIwWDDHrkjYU4q2YTpxhLENz+4Xi8wfBpW3T8Qfm4JFa4l/LHD2SCqIscv
HLxAxpxnIAEojmJlaCmIynPEBXRc8WCP3hJmJ7zUk0BLJ1jLtxf0roTDtEgk3rriyXRGkdqWKfiD
DyJGBcKhw5yabv3AxPBpeMmQy8MN+b0Z8MUWSivzM/NlKlXt6pWx/jm0UNWK9HQBiWRdLM7eiVhp
LbuRTSZMYJIuWh67vmhKmCezyteeH7nFSIlRG4cJHUdzgSqY8srKIxb3OlKIc4PUUJmI3LBufFOG
mj048mU812kGpzebbW9clYn8zxqzOTbfU1OKf0LH6NVytGSCjtd6O+KZYpoccpOrco0luJCJwWaB
EiSwhyKbADV2M+nNZfMyXVK1QHSSUrPKMrlOvBFasV1eWj2wMHWoKo+4+vTcbkU0j4vz6Q/P8/Bc
wEfkkfjpWWLHj/0k9RitPQcLK5vmabVXANAAUiilqb28s1564pFT2gqyVldXu6bHBvcGIiyWL7o5
NkH4vMr9iNsb9Ge7ravLSjpepOCosKLBiexMwUpMu1+fvrkgCU5LTYuGmYl/kcqIDHJzaZovrEcF
IPc6f+etoSS36T+Vf7BJ7qO1Pa4GxOf8iX5DpyhrkjYjt6hhTuO0kXXElii5hxhY/0sVu7GYn8tg
pW7fm16sLrT2FNSNu1GMmiR46doPzSyoLlBELOl6DYis7CCeBJyvqpBfX6NJ7L7RN9nU8ZmhVtwL
mCvWS8UNUEV+bVIXx4CcSYzAZpVvvG6X5tvKX0gTkZnkYhIL2dx9SAbPQdUN5UJCVxFj3Qst4nPW
i0viQJS0a6FhBeC4429d7albX0vxnxP+b3fArk1hrR4hm2+Io0oYWEzQlZIi0WiVyDl5uj+OhxsW
y96i0P9SxkxHXG6PIrREWruSgjXhbKV4nSApiLOv9ipA+Y2L6+zXd097qv97rU/p/xXFhJywBKrg
9+8DzZV/d2lZDqlzuuRJksZZ8r/2EwsnI6XYTBqFi0TiHHXlgpGgu4nFWbgX0gRs6xg03gCzaUX2
qnzkQwiNMkda+UjlrQ22D19vwwODqthhJuWDmdLQ3lBEVXy9/GUH4Z0qROmZCoDgiAZDHB5sFUvM
V8zeqJAx4YrWd8oGNWQan4E/kO1v72qVIjqxm/Y3wUOV/EDb/1VAv1O8dKjzDo8DHg+Kt6+iEVzR
Ns3NCum9F6vK4VtT+Y9RZzPNnfByFBd8spueuxC7sJWk0dBjHPINsQkk+UpCR/C9uVVnINTEZC+g
sjgrIBZPGKTcw4coW+VtMqE/28KDPY7CfuIrwwhhl29N75DhSs3rIn2FSSPPIJq/cjG9WKE4fQHZ
bvBzKLkSIiWaFGCcbtKdRpoc9nNH5oLPgY99tiyx4dGZEFsoNa1/9LOjQ5dfX3P+AcrrRM0zw/4H
wTRS/Zsg0iksGZPeeEF+ikSAfjO3UVLFO7uA8iQ2V/EQKzrqYzLTrRb4Web+1OjVZ//eFNHa5hXj
UC86kip6gtkGz3paed2G5Sl9xTsi+2PYhLYABBJ23RCGeLFODamiL/xzZq3gRycB+3+i2jZOq1QF
4kbjhXm8HE0fV/IO/zYahzdt8VLE59S3FdUDdKVWRQl3I63I129VCkq6vc3nNQGASbHpBaYGYOtN
BxlBHhYzDmaAUdxakrEqUB3bu32tIXndMWtwonY/DZ26PA3RAcuPG2iRGDB+9Xv3/4t//szJpp+2
6DQ8G++Z7bnYA4gd4lKyK026nOv09V5Bqz0L9DTxcHujVFw4Kg4U4mwaJ6mx0oTiR3TCOuUVv+RA
rwD1EQ4ea/5KjJgjjhfnxpPBPKrh122EZMpjaBVlW3POiaUpWKGXQrIqcX3dGs+lmveOf2eqcrro
WksmNBuT5MLi17ZDRGUpoN0ZLDJECX1CD/B3Jvc8gAjqGsQip7vS2QDYzvqjeOwrSwnR4FOquEmR
z0eeTVwMOxik1wnCu+WjvMf6dygXysT0lPuZHGjlKKkRJINqaYmL9Krq5OUx/jdjuDIkFDfsWz5G
mUEbLC48yW9WxPOsc2AJMB7QMgw5eb1VWgSrKW+o1MYjwy/sd8fX9gVXfwjH1XZ/wmJfzT47nTYI
lXZm9mABBiEu1ygRZT49tSozwYF11OYAo23Ii8cVpZ7sxf0EXzEfCDH0L+2fX8DrB4OUBqi3c8Ia
FhldCM+vtqOWSiY+OBI5g1W70geExYanZoEG8BLST0TbFRlpQNnItPRjkHVUlh1enwABT4tAleqC
zQibSfgVkjSeBohHgL49rRsQAzsD2UuygpuBii6AfIm+jn7dfsnvdh7Lo5vozzRNBvGSWGHjTgwN
2voAbhv+ZJWASrh9Ql1WYRSgh9/LlN1pb3TOE2liZPQUt+xZ+euWtiLuYgvhPAZGsd9/RKyS0u4S
O5sQZnkAsiJ03TrUmVBr3LRI2vViR/O6TT8kpi8wfeXXRv4TFcFHBSd8+tgNStYtgzBsFXNAa9WX
SUI1mnLrRzhXS8HUj3HZPnkeFKW8riQ0nMY8RoAZ4ir07ULyu4OryKpaEesmDgwnryVKQY7flOAa
NXCnfrpC54DckJJEUx/jTQK7jjvRKeeSoCPWZqyNAsYr98jlrIKj8iIuxX9tfoXupeYNMdqqkIMm
ySfJKpM6/d7Q6vK8VHOJd9hltffcbxH1S4Wr/l7vxtqlTmJb6ovJBOsGwBxH3sxGuVmmZom5sOYA
S8N/ge3UUuY1uUF0pkVQuzm8mG9HSAWxJt4ruD+tpFxj7dGjJSZBfbwl32GCpDkb274e7IGIJQ6t
nZ+xfDBNoycDMJ2J+RQxJAhEs9Ogr+Xph+HJgmM09NQFZEovFL4peiFGFHSS0juTGXRyBi3pPKEv
8g0OrCRUc4ldtdSbXvauvWT+UiSuPWa+jAq1R091w6GaqGJeE1GfidMkaZMYwJURx85lkpwpM53T
ZAqmgzceL7l54z+Yevkf80M1Zos1SNYzH2d9hAcMbGnelARAAeEzXzwDbXRRySSSF7qTmBBHAX43
XUB0MoNCaG7PyzOU9PqbXJ++hnYwJ3JUh698FQ2Lt7rIFr6PstxhtR0UyvaYDg343n8WuRpy+emF
674h0dgZYViypHDGKKExpMUY6dugbGsJeTBdnlZcsGB7A94/4ZtkLILMJj3pExMlN6JaUmYsM74s
0kuMIVqhgn3deXbHWJdDoeWFjDV2LQIdz7iNlGm7U06hx6+HGtMNN/oUozX1LBy/92Opx75WnaDv
yQHMZyiXVS3oDQeLFVdgJIx5mJoGWBEzq+HEOJJgmGCT30+kfCZj6iW8Y6misrPfOTteTfvG2LFB
Iuy6CwrkLdUrtY5dVk/QTZKZu0ruJBYIt/zcwxJ8M1RMqweSldXjbZEIsr2HlNzL7hUkGEfFl6Hl
cw0/bScyy5FeznK06fi5i+e+HDW8718+X/nkA94kB7mwjN1kTd3BJ+D7KUVKtfJXETXg3oaRLONL
Y3Hy27hEJD7DpfMMdwW6Ko96qsRmXwWuIWqJhMFQAH7ul0osWTsahlm06defeilQcBvNnGK1yLVn
PFz4VyMIxFlB8JUsDxN+M/Q6q/T9ZB1O5NLIqSvLYSN5Navt7z5DUhdRf+MwEK8XSEYgSbmTrE7a
REhC7x1WUIOZdEvPRvGso9BOCzLfF5BJgeBlCzK/G60e/CQAG1e04yJ0vFreBgAXgmlDqa3RXhmz
fVoIr+23LczcvdnruKDCQdQkIIvULP5zBYKnFKQkqBfm/GB8VQHyMgL2DCfisw8Liiu95/W22hZJ
tz53lZ5WCZ0RmqzJxI7/eTSq0VlG53qDuSvfqMyr7NK5D+1SnQ2Km2NiDcyPCXTHhFRjMZVlZ4+O
lKOhBhuxojIzbe2m2XyrBRQrmumC2UuwFbeQO16VOdNRexBzQlTUt7ith4FkR1uGS4Mil77ckG4N
KffhAE0YX+7ul6Q5E7oXnQeW6w+Wx94vE5DJEPSxO7P/wcVLCUgG73tmaV3EVz1SRPisGX67PAhU
ZEXjuKB2kmTeTxUQeOBc1Nf60le/0Y2ehsTwyrntOatmd+SubjWLQ9MaoS+h1UUVKVyIPodebrMt
BbuWGEupt6ko1YEv7r5maWqt5i8eT6snGXW80IxpV3WIB51BSidkzquo50sJnPr/dfBlNnTBlWwj
4truubQPl4WQs5ABrmDVEn0JqThZi6s2kgxKa88t3gl++WehrhGvoqIuzhBE2AMfS5FAfyaXte29
BYIezulCCHGj86Rf/JJroDPG0Uie/I0CdtDhG5qTe4yiei10sOYkNJDPj2W8ybKV1B8ihCWx0rb/
ZyXDw3Z+UaCFSA3FtEDHUrjH4HTWv6KK43VpKKGze/29PZj2u4AZlk0clN3S18mYvoerkhFq0ns8
r0TQS2m4mNEjr5dydhdT9NUKa801sZJqoe7FTtKVORgZ5xeK9y+rg4+Wi1Y/AAsFI00kXD8h9Z2Z
egiBAJEUgCNO4Hsb9ctWmKPpgkertD3f4gaVXBOjDpOrNYdwYpyx7zNXBjAg5Vc24XwmwbtyikzD
Zoo9bSvwn5RiBWob8lNOSkjKPypYFhGDJIvD8PQwtdTdKy8MWNw8F7tUtn8pL4+MNmYasinxg1Qc
EMRjkTuwKyzaczCljudw0bey/iKbA1xXMfD4txEjIOmRz08LA3jC3c9cdRrCA0CZYZJi1/hN7BR3
PZY3zRs0hCQWrswKtQf26q0Kf/tTR8Tpw6D8Ipy4d89DV/6/BjpaquKyDEXlIO9+lEQ3Fn4Q5wSO
ED9bdbWCVgXhcSniGeKDyE9wJMvEwLr/XOVPkahQO9UjydNoMBnZO1fDtRoJmVYBJMrfEeBdSLMT
p0Vlh8+e6r6ibSY4ho/0MV2GPp1doFfpxUjnKtUIjI1FG72USrS0V0PVBOogDtQIb2DDnnrVWvOH
wNgdzcS/ivqO8ew7P82r+UaSlTKen5Smj5vo2EaWIbgECu0O1+Y0FHrZLdU3DQgo+dhnJ5b5ez7F
427LDMuTQRKL+DIK526ZoNK4Gm7u1FD0vRLEKt3vB40sJ3uAfD4TqGb4mhO/Fh7+bnKXWIhJMXHf
cjcSMGqq3gDscL2Pcnwm3C+m+dohgmepnDr1Y9wpWDG2kxZDxTsQtfBu09NHvFGmR5yriwYRsOBd
9LzOKmKb6ZSCS5mXCUdHPudAJ0AHIblSnPwaWUzpY8e6LsI1PsfjTKGWGTwk1lqfkzgSLOoPwA+o
nUY+Jvse3oQ/ss1351/salN4X7DdFQ9cEEkUB0cltiPjxiBvjZgGaFM2ZLrg0NdhSMLJHNxl03EK
IcURkalzBmTWL7tTKN0fj0ArLSHwzSQB8OeKpp6aKNqSigX2GW/F90fFkBZvnhXU7iDxgkG4YO+R
WT2VhyzRb2un4S2tyl/es1W5hvM+9NE+xNAfSvIdsTZAZuAe8R+DN1djcW1ls4m7S5YYvIHBfGHJ
9JLi4cTsaTDl82bdOLOFdAVVYoxe+n2ltgoWBKBhElkIPaYOFnCT8w9mCVCtuwm7GCMkSSKjN0jA
3jmHnRfT+DMyVv7btXOzQdIJ17GAqviDbmufASycuPZm+bESaGIKgS2zj1VBQMLGGJyG1US/q27g
NFPxc+lVL9wDgTrJrp30TtjD62u3r9rh+y8nO9xeLx66f0qxe8h3Ijzl+2kK4d3ATZbJVBcJEzR7
NDMdrReB1Vxds31iv2aC8nio/9O2RlXzN0JVKYmidy/6WtlkRxbEbWTXQ9FHftdzl8V8r1+hka+S
R5GHptDRKLvM2IyGbL1WqluhKj3PNnZmUOSm80kisdIWeXDCBMhafPVHA9cwVcEpyiKm4mnt6WVY
2JY6hRLE1H/ceYcMGwrJs24AMwaH6crpAhqmyoBWUrFv44srs5aJk5OX5df4EFGGJtqSwLkRWlly
zOBye7/gp5LCvJgMeHI42GYnClrUPvjCHUuU8f0l633HXUHo2r5o7lsBMcHucGIbCK2KDZopFQIR
hWPVk1oSw+RWhh6Yu0763fnmSgTifnTNFjdbDOMB8hIJ2qhd3eRS13c8dB/H0muKBUsl2Q9KIS9e
0mgvA+ECK8AUe1FJuGmGZt43IJoNUjdrLqDXIlOfsQwcAqbTSri9jqjx1tjgI05Te3cv2aDKnm2V
V+JYcAf/r1q5MW1vmdk6xpugTbmFH24Rs3+awjkrKIqRXmfxHrBRLvjNiypGoxWoKGuSN3teB7nz
OcXRKqmuPHV+hrch7OV8yjNJQKvyEBvJChvyqNlDygkQaTuj0hctY0mButpu1O2118ZJlfS5ZcYZ
G8Gl+Hi2Qxe97YuJm8W6HusiSVV+zjkA11Knday8/oA76lVczNb4cTQeyC6iEnPiN1vqe7ScB4BX
uWlPjy2mfIFiKbk77BRtyX4lUxNotfH9o7uB7wtxnXf1V8/fDbUMrmEI4qWOd/t06ks3Ff7vYZAN
aYmeo9c7dyWMRxwUr1+jypVkG88rDNftXJKwwasxcFw5Kl39qZV6DEPzKPngV9cDHKPzsnQZvkqA
eN/s1M7PTUGDAQMmkz1S4WiV+R8TfsyF+EfELzftGwloJaj97x0OH8KHcTxDFH8nsju1AIsf0FZO
dTeu+dFshNOMySvJ7KZD/nkIUm9A+fV/dGvgxIf5sa1wkVPcSQyztF/6EXRVArrjQCyiTTXJX0VB
Lxtd5hyhZf0f0bOXP4c5y6HVdxGq0ZyrNF5t6MQKnbv4CGVraVaEKwlpYANGe+QjITyq19M2uqWF
p7Hq0RJjleMLWGMqzMysVclc8fYpbiTzl4DIrTROd1QrXkT5J1aMgB/Nmn/GMch3vvOE6PrGF69x
Fe/oxoMnv8WJtk+RYOq0c1ju57lsoG3kkPmpPJFhlq1Uw0/LDa8Mu4xnVmoja5snIYujD08Gj9TD
mwulcU1qiGcb0WVGPdVYluVCyipWDAFkdbmGvwGm+nD/MZeW2NRVqoscY+oQf81boBqktiLmlv0Z
dqB/mNkL3Z9fpTW37bl94FYyU663ynxDufoWWp9+1Ab1WoV1LgYv+4FLLG/TlGuGK0LGn5rCArmz
KzHbf/ADV48VB3hWVgeaNcaot/CE7z9zcXl5NQkphcFAJlWGzHeJodbRXyjDiQ6E4ONTbJT9bDzm
dPkncMRbeBv+mp7yKrdE0CNBDAU9eE24DSi1bQK94gzuzp6sdMI1oLYRsSJn31QjrRdisZcoXU+s
xRbhXfIqrVTGEhUzD9hxqxbnk4mb4MTAaEF3pAbOSgQXylxLejqZy5dQITHvpjZuMFAHUwwSUtJJ
Y76EFotkf9GzLxa1lTiUfv8HhwbVUhIEZtsMHnuQfrWlN2J2zDHmFdAorDsPW/fwwk48aQXbLUNW
Fr68fdjPYNeYmv6lZ7lYyHwUSgBRpX/2aGiZDRgND8Qp+5Mxk1T3SYs9dpWLhAb0ughWBT+KUW9p
/ageYdMi8Xm4evqmAT5FIY0YgCCJ47DVUQYIYNKy/6Q6YH/IXN/lBZf/5pr5ipWzl1+eajVfel3v
PcE/4QfinjQKlK5vqFzqLExL4AvTAaANZYd4xgm2t6VkpTvapDx1m0qF99R/reV8zWKoX3AE2dP0
PqXI4y5JEydnzTpjx08juYGwiAa9jefOXCkgXWfbeVRr2tq3QuiG4J8CRZxT2btj7o0TKU4ZLzcQ
cCee2SxLE2GeirzOlmm7t+cohdOk1dlkG8QNJ2Y0644dwfbg0ujMOAsjlSLhWKEO76L6tBgJavHR
kh1464fWpwVXoHXEQ8y8iBhAMtPut7e5puQUY4RCI6+c+Dst3AfAedH6MbH5TIH/sk4SfS5bMTRl
T6Ay3oYEIwGxh6Jg2bz+eok5v6aixNS6KbX5xL1taaEep04GpIvTGyaIyy75z84wGJDINm/aFLTL
amYMbjLO7NwzFMYJvJljmZivFxmbqCTTG6RtdQsXbz5u2CL/kMsjAJWXLXa5Ntt53A+ia8YIOynl
eVkM7I3MPAMdtxooe3EeFk5JgChyoGS9DXNpSwZj4i7WcBWUQYA6Qxoa+RR828ZpcXHbwNdfYcsY
HERVrRg18HnSXzih2MWv1KRX8TVXTqeIcrwcTT7vr+5uxAethATeBujaavuZw69C1dqz5mPpObfw
ROHY4QYiNaHY4m/qrvxijS+WvulowSJyi+a4exAMCAfOxUi+VAW26q9/RZRcewwskHqwkqemXNw9
OPOG3fTSQ2miWBazYXLR/h6WgYJBnBvNV+cxFuPPBnrpUhqVh1HdCg6by1j+5HyfKXymxfvHoaHD
3atGc/VeblbinCNCyIh167OfIJZjVCpxDsWyGyHhniMXlMIrG4hMWtWwFHX5CBDytdYa4UvM0Wcj
OtBRwGKW0T7ktCxidVLbbODYdhNBRZ/Qv8QS9z3c3KU2R+za97WReOVm2vrh6COiF7X+Ye6MoctP
3tZzwu509DHHP7nzy9mtAxNV1YXou7zzyPQ04LHrR5k+aJlCLvLzJ8Z9+xT4wFO7IKAF9Mjhe7tP
WXG+q3oxdMCZ70DOYSy0x4zdVzlw8MCHLqVeWCAXWZK0p7cuOCgAe24PlsDIRQcT6njFUnW1RMZu
wI2+NFWsHPGdyYcxc7E+DAG6S6QbzgVotbf2qWemd1IFmzLE6AzyLwcLckGnI7AHJv5li7ZPZqEg
1Caixw222l3hFiyIitTE73/GnR6jn/aFmW2YEpk5aS3PJ40gfrTtY6nnIp4to5myLPuO6E5FR23O
IVwhduLx/PudFk98D7PrpYhXgY6y8+vv47yKMqzsIPZx2n4F3oWpkc8iR8zWIe4ckIePtl/sr1kX
z13VLw4xiJuthICRM1AbV7z3r3FZNhYQ1425FIfYMDr4gnbwPOq2NgZ8iIpxVQ/iqjtdQlmp7rmP
H0XJsosCINB3497GbSeQTS/L6VKsOc4uKU4gKujg1diW5ECU0e9Z+WRpDE0Mgs+rZOIVGPJKNo9a
MaaBANvT5ZjRSZboz7kh6FP+34ZtQkY5gk+PVOkEmiXXFxSUV0D7uRO3+gtLrNsDMGt6badNUkW1
wFO9niSBvpbekTcug3m9+ZYKTzmj0FOsVsWtUkA2qoqZqgxaCU1A0jd1uq/oV0BCbTDIs/mBBcdr
aO3Y4pSykxjrQYG5GO+iFU5CTmv+NL4PjFOTEhkRpEz8xEQU5XfIdFucbK0DEJ/IYahSkD99NtNO
Yvy/H/kFhe8fFdNnz+0k41irNcYEPOtgxzD0O2ZFNwP4CDcxvz3gDZ16/jKG+EFxTguXLhXwsltA
b2zfiHkyFzylGhiV5ytWAk5L8KRX5ImWi4apl2+8hREbgCIBr0iezicadM8NaBFmUMDN0XI4RowR
Bvu7v4u2hxgUz36ZreHxaX231VorMgkZMMzudZV09Z7vK3VJvucJUPXEXAXOJ5QAaa1hQFRIJHK8
JLnJafgx0EmCWk9L2SSqUfqf+kH+LqwU2FHe8+34hqzVJotKfV1GaBKiz1qvDkCVzrsHfmUG0W0Y
2fkqU+N4tnRv9m4UzkYJw+ByLth6/buVLMcFrPz0qz0ifPIkRRasNWELcVpt4PTFOAutPSgeTTUl
Q5d29zJxIQf7vPqS40GXGoqLUIBqBpl5lgPeltelySbe7eftkkJNrqaDwN4kPfmFBmmGCiqNfV1Q
1+Bd8TEa4qqKHF+Ojunpk1fkpNM2lEg3n8x//+4BiMl2HjojCV3zOyvHOwNkyhKP6Ri+17r49Rcj
+H+C3HyuZ9wUJQ5mtEnh5yv00pBPD7IEpiS+lnCxvEvTauwExeN54vm+v7LS5BSP1LCM0eoM8isJ
L+DihHGHc2vBdNroePIzdvly2Evl5aAztQ50ZBgn6i4niU1u0CcBjzw0IHMPzZO2zsEHcX+T8wNx
MINQ8uo2kuv7cr1JZ6rhVpTH4uYChfmlG3Szx/b9y0//bQ86ayw7qvQvQdiuibMMdkgnEsnpGgcR
iLvftpkSF1X7qADyQjldb34pypkkXy8Uvj8unbKAuyfy5TSqOMcEJCGGUyk9CNXSzWtJChus99pI
AyumkKYMIyvDrFLbgW1Qgc4a32hbSy7xWIftAfTdhdEmfzddR8MTWcqtVC7sSQPLX62yBBES096h
33yff+Tr8GAnPugAlHwUIAa75GfbSsl6kcrYlej+ixKK0MGLUKyKQi2h4zoSxQQIcdXieSiN7uNh
UG0WqvNln//wHTJkZkeP9H1+5WSd1of+eonwehN3U5TBxCI+NHY0o9jkCGYQmt3gjOv748JRqShd
99xM+5lZRph/kr4RZhTVzFfxCu6L8PjodxhGYWPxAw7zAag6t7NetkKeEsr3q98OmWOBEVm+l5RN
UV584seWJ+j53ESdLSO/zzGvZ0Gk8mvBWl3qX04yY6/Li5aWbjD8pHwOwTzP9NgWKAoTZnTxRDFO
4m6RWRfMuP1MOmMWcSKNOBeMwPk1nq7NPSedPNNaAl0UGKe0cwYhTykuvlA+7sCRa9KEDfItnqNQ
MPlaJIYRbV6f6qSRyBwcVj/zdQXqHhhmSneJQz0w/1hMx/XTv/6Ej+ZN8ihEeQiPF2aU/FpIvwNu
mU1GCKgvF64Erj7xsA9ahz9K+rLWvSU5m1gm3MvBaB9zu5Cb57sbPp1l0upAJXbtjB+xzX4rSDlZ
MSVG90QNKNwazPlXqxtzd/t5tpCkKQzL31MgBsIuSVpw1BAsJshJzPn2LvYBOJCCR4M9BCT4xBSj
ha3IAyBUMroc2IbZHoDoK25//gBJMKvDBQi/fTwP5cD77Hkps0H6z4cc8xRXO0hnDkjRpgic0vuh
u0S6WYpI+hc1xSmH7STtsNwYbsLbIHvc1tib+VbKpGh7bIvL0dBROh38c900GMoV1XrFaSiZgB0c
HSoNJBZi2W11JTCsLuf8JAvMhY75bwsSBcRfWBnzJl/BrvGq7VW0oh3DtLg7t+0L0zDZvSE0Wy7m
rRHWokZrPwvDYs6Bl5PG3T0RZJCcxt/ha2OrIVWoo+Xfk1/qi/Qnn2E8nIFD7qItaogsc5gehhO2
b6B9FE2fg+rkYks2TVn7HLTFQZn3j4/tkQ5cFrJ0OYsBcBShHmCpMI8zLsekmiaI80xWTD9kR9zv
Yc2lcZhJ5bzsWhu+L54a545kFuC63U80nyPGpeTR/IACw7Bnz5lx1zkCBbxRJ1mcjl3RisR53Dqk
eFRa0W9aXXYe8nEApT+HTrhy6m/bE44XGWuuxur3DIdvs7OAHUYcjBHAP+5w5UKiLkQ9hkZjgrJt
TxfNuNm6cPs1KXOqo1xVTIhvfb3iKF9l4BQcNBY5TE00BiR4YatLEp+uxNved9XLXDQtR89LkvvT
mypGjDmJnjEZDz4tiocG1mqkv2UgmlWbHej9peRKjE2J1z1UL9IOKSiRU2HhlBEcLQ3me9wo27li
Pp6pmx0pNiLlLui4hPDkTJT4MHpCOCXNqzVgC6jsAInMnfyD2g8tEjYA+eLgunnCAasunzhk3AkN
1HV5RkkpU9U3MaZb8wfTMJesZn1vM7n6lhMFJjHSzTz8c0vkZRdLjUs8kufv+19sceVgta8h9PQ8
DJp62nHQ9cPZzh7INxeXFvBcZank2EpSoZnVulQsbzRc67dSMAxVc1aeXoDzymjZtrPBgIwEIGle
plwmnDNCLsZ3HoyZD3eCB4MQ6kcH4h3KtiJcS0WFHP9wPNWkNog9y1Lvr+aJMlwYUv0RIDckvn/0
WV+c1ik0nxeIM08EwPm9r47bJ4iBHBsag8UlZU7gSOR66FpfENDFVUagwOAHpTg4fjlhHZYUw/kl
G6gHQgEYrQ/E0dpeSSaNEKP3uj87JW6/LrlZ4nWt2dKhB9a+KBBhVQv17erbbkuuv39soHtKPD75
4bQ+sEC6l8+CRNrBaX9Vd5dAuU3D87KwKNwoT0qLomRhIYjLm/GrZdRUszDvG2Sn6s2O5PwS7dP+
clVlNv+4PVEnc6pJ5K4HWSIOyImd/Cd+svdoIOyCzl3cZpsQHi0YRMMUEOPPjSzUWq2uWbnd8lPg
Il0HXG7ckbIG6q6my68wTYJlR0N4Gs8rtLV/9C9GBoOh6GEOv+HzAQ+v5axvtvUKhfOK6ZM6YA0f
0mecN9sIzsyytgVVBBonzhdO9orN28zVhqNjqDBw6TvhNmmqi4kABXwa5G+wfByOa9OHfhURVRLm
G3Fqt/oXa1X4c51y0gwNmAPT66uLi4qJLHfzfViM3ZbsNJViaWavsXMujO9UhlvNdWQraXkXcI9B
1Cla6xCDGhvxe6yRxqWUELSoicLCUOptCd0u1/+gjaXMW9vvIcwKIK7LuB/Ru0LV2BMV04hWrHFQ
QkAitBzkfQva341EL48mzc5lToQgmxVH9XyruPx7J98P4N19xC7uK8tGj6aKbRy+6nLwJrVW3BmA
FUC0genYEt0/kmqt/D3K51dZGaynjjfO++1/2aiHtvpzVOag4YtRu+pXDX6NT8FvkaKTX2WL/nrT
jqmkMg+fDxd6FX+4DfEQBjY7Pih3ykycJRWRnW+yvNoBQtzkK9P1F+Fxxoo+YTxQShwK+ZBmfSr/
PIfpMx0msDqdT9FUzj/6HVOWbGML7XdzDok+H8H+nj87bs+Bkb1AyqoKzimbyIEoX8unDW+Fct/4
GVWCo4p7TW278lyGKlIqK25xVKXFlfsrUOcePHNajn46brk+SNo2Ae3JbP0Zo0CNs04oZwG0PV6J
7OGG8YvvIv0eVt958edeu/XZPj0cclN4AkjSbkz/uANyfPpBnaMWoaMajBu5PMcisOePsw217KCb
LEcYmdf3uL4w5rNJ3KXXkbk1WTJLb2DnhdqXzd0ovKKqsj/z5SG3p2BqR0WUthIIdFnPvrFsdrsk
2w+DkTmgIqTmdweA3KSvigdnz6fIJLUTOdI0cHRtPpBWa0F1mkCROztp//ZIdJtNPz6G3dLYuCXK
2IyfYF26J0mek1vkK6IGXNICBErEKthoPW88Ao0ZyozwLgYIxM+S8P92cI/E4VlhD32e8ZgjCzMJ
mR2MEoIHUf/WEId0oQCVPx1dmz+QLe42lCYoBwgaVaYoGBwZaxAWS1G4PAjpddh22OoJb/M6J2+9
Y/jmnif1bzKyQp7hCNqgkVXib02zFN3e78ntQZaVGPp52UgLafi9Zes3wKOU5g/VfVP4d985TxrB
8DgkUlmN0twm5MJH8FPvmFIJJWXGpoaVwIYvcP4lL8u0VTEBmVxIUtmA3vJpkEIiS6uc94tFfw3x
YOsgJNhadnLKySeXiaHLVeXch5SByUm8SAyQcdAg1FZYExeoXMf87Ovbp/BCOKeOndjSMQCaEZp6
W0g4bT/P8zEzhelKN0iivKMIzZVM6f7nMV5Anr4KiJDeBBHb/YWt2P9++/slLQK8K/y8NXezuh4G
YFJNXcSCf+4IIm+BukgQbV16xSVjtl7DmEIP1ygxgzQ0UUBpDuzg0z3oQeAHAfj9ORbRGIxZ2uzd
01PVSRnezffnNEvo54Z7STui8m6oQWOiesIUAl65+/1j1/4wtRpgiN53hwkGgM4by5IOgxwVmNWc
+iUMUdFjvo/ee+bNfkyu5pYeEJxTUf5Xheop5NWTpLsH54WNqft2KlHkAvmA/92nY2MgC7Z0oweX
c2ft6N85p0Ut34A+1Ud4c8uNAxItXNPd0NoiTm4inGmPBPnXBFMtdH1u7/RnQai8wq2gkfb+aOgO
3ts+cpTfI3cZPtrzM8TigLOsPaZgNWKodyJdY4Y1NWozX0wqqxyqP+kgY1sj3LxBMC1tdgqk6Rz6
VT7VwPQxdHdMgMwAEGuylmlbFgaN3pS2QK5h2njtkCuoAkbiEm830Mib+g1ByipNt5sLReOfzNMi
Z8NvfbvK8ZIGtGHrU9OQ8WR0GfdninAI3IV1ou1XLI9WBWAG25dlaJ3KAg6ImKAZSoPYKZ/hd8M0
r2Gmn2mSn/X3b71Orhg0T1lmbvjamTyhIel3XpE+v4/gUsrIiGTEgIJBZSJaKncXvMR48kbg14zC
j1P9v6uVmBskLhR6RVltKY40EXZ6LEuAmf9nAMmBtM0snz07oB+N0SZkbUnj1s7AeRTAPgTRNOMp
pIP0AwGhoau6p6J51fK8bV1JIc38VWAN/82PP+a0nd7NrJMycWo6IW4l7MY4ARDRUBeXITIRCFTc
t2qc6W0qWC57quDUnGagLetGpwK7e/TyuE0Uo9MENztu2PWnJoeUbo9f2BGfsE5rYhyZamuyhDkK
0vrHNH6moyzBnzSAT1fsXUO31wHn2NUlFDxA1zgHkTDtpVEYcdExUZ3N2/7GECarzK8dvUXRY7yw
3t7vgHn8egxyNjeHo1vRinYZqgoI8R690nrfrlvc/kEktyjmSqcGKScsCVeuS6y0YOLwjJJnbBp9
SeX10LQfVVQDNS7iabR7RNuLnarD1pAGxk/2MlAaeF3UDeldJKizpZ8G6pEKGcudldE0LZ1ABxTW
p8mjNwd4KCF3dRPB1R7KNhcP3B8flvqqBPtQxgLqb6uU+zCe40pze8fFeq5iOHIwVhLea8JiM9uy
FO/7B8/D+d/f8U2l1gRCKsFMjE3CkDQNbzqPQEBwNG2tVGInINibGplSo9bZQaLqv9gKYvLmBmnU
3wjPJtsTBmj8NNNT1LiLJcGSTkpgcaoQMfCT/Ut81pPTQ2fgIhttq8YqIiVpaQRtKi12cXgkWDod
lYoTMlEN3TAvrygQ00GS/YOaWkJo3LBnRo8YrID7Z3YCqIC5xsnVzPmir7YPavekJLIxtJAUtFht
sHR/CB2vCNBVdCe3OM9uNunIjaVeqt8SDmbTI8MKeV+msS1vhGnSaS8+9QTu4HhenKRa907UVqg2
SoV83QfjkSsG+qDG8Wh2c2atL7xn4MgAAi3ROyGSIlTheSNA8OTEHTwhwaEiMSd21sW2S9ONSXSi
Dp0LLdF4SbA1ZgugysNpGZ9rcP0plUkypKY7dWplgLuQihXvjHMVibddhV8rfqJDDexZ8kKIKNjM
kzOMRuA/r3FTvkDA7PeBidvSDiu9nSZLLQF1dOXZC//75a9HZv3entIaJpD1uO9dlm1vifFu6N5v
CfKMLsBVUQe15fP86s+bS9+xt45H3EF9YN6xlriG+niJ243OvT9Y54H58UwhTQWfd5FDN0nl/wjR
Vk0xtMT9Sy30+gpkeysGdE7IvPvxZfOtZKkXVeDsIep8x3Qm4MbwPuOYMlsCJxmcNI7dhmMWsi3L
pGMqiO/kZVXSrAEXfQEB6xcES8doPDTe5zxdityI/cmVimY5AmOWBJO2JdsKceX7v1BSRgEenXCI
cYj9YAJgTpobU2YdxiiNk3BoWNjLcEbHS4xtsfjtyYcj6rjZbHgFZkYItKglpVamXyYmZs/KUjQ2
0dIwLiUSLvtGF1Ay3c0EM4i9OlUSt68V6qtjFD71rFvXt772+kw4nzdEOAeAzvAwwnSvS9xAZpCr
+Xyrr3OF0y0oygUGqqkbeYdYEiYS2n+FgulTUVAW6odwrc+6Y1j0GPAzDIjQ9hMmh1f+2CKhT+Nx
RABWYHK/ys8Hokt15Ep6Ufe/Wq+iQbQgrSO37MC6r9k4e/nLUufZ0viAgs9THSXRT3ft8SKtejLa
tnegQJsnPxNAurNS5MtAGZpo7jSGnMR/HrskrCY2Makv/v2+1oCPsiRl7nE1X4LNKORl6bTY/WSy
4wFnZYJATXSVN7hhOMtYWEwrbAc1G4zsYWab4D9/tdEu9pXtnpA8XYgXdToStbqrmQ+C1pCHMcRY
zVokimgLZyIECMHRHCRxwa64YC3bvfjSVJTIj9wseLUuWAvLd/w/lA0J2+dFy60k9jp0nM1X8q82
aW+45DwPZw3XvtpD/UO34saPsvMdtFsAcX/JbJxyT4NSsvkUy4L8qIP45S8qiEMcET9uykfxesVY
4STsIbl+2vQaH4esE0yL7ZMCDeWlPvUAtb5PsfeUIlXSK7bIOTu0bE7DSq0BS8cMRoskfEpfvN0p
Ux8szl6Tsl8j3CTPMVgS9EHiGUs5eZspgL0jKRGt2qq6ADaxB+aHM1wCLeKU7Z/uXIw3GlDN74Cd
pPBFJNTWJ4m6jj/YPRq8nC//o5yXzH3iTm240V3ObTurLl2OhYuYHzsVsoU95RpMAEEz7oY/fdZn
gQk03tuOht0+gnTyIqH8wCwQ4TlIU17K9F3OpGMtxs27YnZC8z72t6APWXc3DsArWv2FJKE7OjAB
Y7mCojTW5GTKSj7otwjvSglmYbLvxnAa74WFxCiL9ubKocn0JE8QTDh/P6BWGgK8YeORcI1NMO63
TmXxEFb0uZcQ8AVZZWPM0U0uBzBkObfxQp9ag/x742XAXfAFW2rdFLmLIUxY+I1tfxV5E2vugl67
cW/3Evu1SgMC0B6VPig9kFlVcS+3R19MOA1CB/Psmf/EKYPaG0RyjtTiGo0l/17jC1B2aUPphCo2
04LnnHXBq0kfFegyi8CAb20R8akCBDqnpbM124YE7Xtj3xHG+WyQYT8gDREZYJJJRO5cAYBQdhwi
R29Itpll35AL0B8reJtRN9pgX38Xm/ZzczbnF/q4GNUItfM3Hb679qTIhqAlO0pie1Ud5ued3/Di
gCb/i0UZJ1zEy47D3wFA9UJcK+ZpdSZC4GskxQzmEc4UdVBl8MHgE54e9tv19BPQoKovmJDgBOvv
/ZekC44+VrWfU0TDqnbB2g9zThUGQ5PQ3rnXRwYjXRuGJwSYmbMGbZGT4e5+ccFe/41DWaAEE2E7
PdHzrY9VgmNx7rMFAB+rH66pw22kx3La4sTOlHJmX3egEN7Dd4331UUFiHKE0ChQx6dqEgDmLV5x
kjh9JA1QeisbY7H2j1YZYTYXmAr0yPEX8VJZOWJpaQsNlE+ADgOPG/g4frsWyXOxveYtupAHghK2
YkcQGxEv5WnK4kFghP4xLspcnxL1wdC52OhHcNiNK+R8ZoF+dA9e8f2VALmLSrjhZlGomq0x9rim
/wItMVDhLghh2UURIi/cm9c3AnR2QRrdHerM25v20GiAwgHyPpQXgQEd5vIMdMKzF3ZxqP4H+qDa
XltH0HHQnBkaDINVB/tJcX7qtBv6PY52UjBtNcOUNQw5RpWa+Rnmiey8Ifr5TVGtEsqKq+XMi3oL
vJKOwn6j/KGLZFKzBRtt7Lzgd1LXb1wafhihyuIFUeiwW8+tCR1rH4PW9KcpbwDER/wPXH0Jh8mn
NeCZqgo3ePUyhTFM/zF8x2PSBKdDbzxNRFjpOdoPdiEOZrwqqz8bSBRoYZcKtkHh3p1n7ocmt2X1
6pdhlxJH3b+rUtxCLG8ILtowjfY+Sh1BFFFGjpnDAX1eySuMzxPp5vbMi4x61IKrGnvu5RSs2tPF
3ytrso27hWVP8m6Z1FaNWyb3Uv45kWWZNLGnNqnYFl7DCmgDoXyo2gvT5I9vYOj3RscGWwhKxKXF
ekbcQliMqtskuLPki/QInim3lckHxgRULMgUUeNcnvXTKnyXaZ+KgbIQJ6w1/9nmvugaxKdLwr3I
fz7/wSyWcduG9FWSqk5q97zs8yU9qRd6y/vz5LhxT/UvzVw1JnN5pjfNnbP6MXreSjTyydPeo9PA
/XyoCH5znWPGym89lTxQIgiVG7XsmH1aVolcAEdV3/YuUCn2pxjB1+8AfkidgMuFnsK5ShGOdbas
oVPZt56ER+MUYf0MeDOMsmB1c5pUMEXJoqtWzCgaHM/hU92eH+9NvT9O8Ht1vyANHsfLedK1dUqT
BNq0j3mO32iUqfMrvyRrhC9oUQBXYlzG9DivX44915uDGp58soA1xIycxh9t8kYLFd9PCv/7LazO
cqNHlYykzXtGyP8uFyxytxDjva7SBhvLZnqdTWqUZ5dwh6I7sqRzibgDM/EMbwd9oHhCaVs6nKlP
hGruvsrOPmXQpW9VBjAEyMEQ1RgtP9Xw92AmmZ4pFYEhqJlsWH5Con5x48XEmQMBA0gHpOVn8X4V
vmL6jPOsVqh0sYKIfC7g9GxVyLC5cNfyRSaFVvOFd7/+euNrkzzIX+Jsc/O+edmK4eRo8bvbIyLN
jWMNJKusV50D8oWE8o0ldt4zNG7fn7oDWmiHEFHMrjQuO0iAgVakLrzCSBwS7VbelVe8fzjv1kec
2E5j/DE/lTH7Azuo3cTKoFBOidflb/edzvI72bWk+9o40jJ48gA1jN3hKkmNu1eJu7quhONYye1Q
wQSbJaWpN673bYmtBSTB2FjK0DYtNza8K2F36hLKOguY2Bp+3rPajnQ0sQadtgwm1aUmQKzCLeRV
2RcaslU3fkBo+H5ijK0hdBjwXLqiH0HaakbJHdp5eCOJQSoczoRMcIa1rC2Y+XcABq+chUYHpvz5
4SNbtcuU9jj1iT4kWRo7TAC7cg+TIrWTp6b0+fDM0OnJJRuvayrbGcY/liFq39eNIB4pgBRQE2Dj
/oLwjTwzwktETKO7lk4hGvwQ+YCw9MMBT/Sog3tC25YSxnDVIzM18Y0TIOddD7a8A54qy7n3mbIi
csjV2KdsNbk0rJbozIIkzhB8+LAkyMEy8hqvV2WKqIMDV9cEccqYJNH5LBwI+iySJ/iAOA9YtyTi
KlyIJWEHfNqwWQarSsYiGjxQZlMt6MUnL9a1XC3iicLrsOG4FhW9ruQA5xO7oGiG8HFeNegB23kz
fgs1PJKa+kV3rSg+hSacudTVaEhTuq6PgWVaXhIMz6G1aa+7W+txI65RTlLW0HaVChUlpS79/F9/
n2QwVxbLYhubg9Bkfv+sY41h0Gi/vdWkODNksE98/SPuPqb1ohy7XKrodHn/a22tch0ebObv+SvC
IMU4lwqMH0IlYi/xGQ0m2mCkDBaDynJSEpJA70SyFy08Og/P1JwDNR35dyBpuJrp/8agspR2yA/E
Mo3fOnKhaqAyd3QerwOEwr/z3vZmBSCY3f0GnltGHZtJ6xVsBzbDsVK/XKx1Dv4uXcMsPvfBq3Ew
KUvx2xnV6+wmh83e3KRSJ5luN8jCDsCmxsVO9sRrcuiyC1EW7ZLzJJq8bUma9OOG+Fm/qpMJQfVf
T5oWNcBqLLJj5bnlg3AdOaICza+JWOOJtA0hkezoxJ1A0GoLWq5wIgPLl2bvNAcZLubvqcrBIbMA
saqmTDIelosomKYs5Ph30jPowX8dVrW0bstRmaR2v7XOu2hfcMH60jcFJC4JaG10Wljl8Q7NEKZ1
TW2rn462sg8ceiq+WJy8cfXe4qA8pt0D/mGSprYrE5Pc0DsSddejpIav7n+XQuo1TR4hCF1DKuTA
j7UqodFr2BqcL7pes0voermjSfseqHFCCYqPj+TBOfwyT+xRluPXODpIQFO4UhCsO6lHHrVBDoKR
CiUDMrbjSCclOrv4+mvu3PEqFuZ9zRCz6mF0AOUC/JSB7gWWjZp1NkxsyW7T7zSr9wU+8f4pPur7
wCW5ZY61YDItC5NaD2IdWlsq+/pTrDqhwaFBp+fTTLAXMUga7n+Gso34jziAcjkpYtx/Rj87HknI
vZ4kIp2yLOwfVr5SdvyJHfyWZ4k9sYc9/LvB7ecBqWtiy8hbbMxfLi3U5pdNO2ywvbuDvHH1RkOo
RTzHH59KZorLoWj6ryGn06Qa55y9WfeUdsiSz1ubIXcext9NqXgA9hUAQ8VFzGW2hm9K7p4DT0QO
kOvN7I9dyULlMAzxenlPasMRWYfA7fjSMtbhaKkMDtkwjY9Cku84IJiTCQXZp6Lv6TvhnsgcRcb9
GI68wK4USn2i7HWd0wCQ+2kC/yibgQGjxKpQuHCg7e0t
`protect end_protected
