// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
cbMg5/3FY1spAqAjMBxnnfjiopba0rg6+02/eGZH8LhhqvEAzkFbBPnNY2HG2FX3XkE/weNIZHrx
5eQUk4Edn0n8wHuVouPzVBUwWLODBr3O1+59fAu/QZ0jFhrPNLP7ARqdR+aCYkauufHo80SEoOWU
tiW0sVWsOt5hanmVirnhZqjQrmcI1/3A9gao798dQqekRTvBq7h0F3AeLzHvHq++gj4EqUYxq+Sk
IOZiFTBGnGZra1BZmgY6t8HSXDiUXcc97PmtWI5UrPPX3lew7gRiFclX2CH1XmI5+yZuFPYldJr9
JLa4FntT9GTFND0lloRjAHSndDxaKSLWf0yGow==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
y9ChmHjsxE3qJR9arKSvbR2+QNGH9hIN6y9dnte1lwZ3Ax12YOR9F16MkNEohSEqDcWKWiejvot5
KtA7VTIKgVPeVNWevNfb0fGagTxJARMd4fP0TU/e8llGrY43kQGSRpcFFA8AtNg0NeahIcXN7yEl
/rYbbuWKXQc998LLTezA5l474lgpPDF3FSns7rJ1JlGH/BRq0QvAsahYM6C6+ZjysONdvevksM0e
vxzG6huP4YXgLamCOu4AQo63Z6YseSISGg1GxZN0P92bJlAhHG4rX+nv5kZM/x4l86l81nfZJ8dv
4eqC+V0NSZSfRZy3TSmSjwI6K9wVBc7jOQGisoQwe66qgUtLAH4C2ueb5Pk4TatTnrcJz6QAuXgq
h40mfvDe17LvNd51HQ2icqFachF3Icw4kq6T3RGTVqcvnucQpNiso65+os20CZ8AUQpwzaGJTjx7
V4Avb+JxBFZVKuqdnaHTVHwSpWTK/c+rYJxkvx5079YTUorhJMCjyCh1h7TLZlg/YoHJsHcOPhYm
Qp8KxDHYhCh+cmUAKFzDUbrKKoK904IVwKzIj/JNUmct1PuATCnxUvIaN6IieXw0wYaS1WtuGWrN
+Tt1Q48MfpJanUbDfaBi5e2o9ME2foC2tAdrBgweRihRF7O5mFus5QR1bsGr+mcsrKOCemMUltxz
P+h560gPNs2LojsSXxkYsVp4AUS0m95sGqDjUNZDOsgsawOPzXCDPwfEQLC1ptqHRL+qsapUAlRn
mLsPWNp9N5eub8WujTXaw2c8Dcv8mHjapK9ddapYGgFtKpUAzGYLvBXpup4LCBTq1y50xVxmxg+q
A9wtsJaOo83osVBI6YCBYVyFTgYSSm4BHGIIK12zJmGdza5xSehTFwp1gu0LkW5keqpJEe/5v8dk
5MiBZ+tiiAQyYYjWHSAO7lc/g7XjA4g5TdTqpx3HSBG5/OK4pSSko9cOKA4+WjOKXZitqlJ1q0lZ
NnUsEX8E1cZ8SJP/u0dKnk/Cu+sO0EABqTzrcjNhG/2vQdGGSBa3tyJhgzDqqJ41ru3ZW9NYbExB
kCIuJznufNDTSksVTJ1PZ/3MthweF8hVax6b+CCASlgghHqRGjMX5sy2uASQr4MlBY6tCpCoBqmo
MyKWtoUlPf68Tu7x0m2VViYbw4PdvzIjL9koC9sKIgjOch0j5dFi/aJ3wELkqm/UOUZwErocNUFb
enUA/ybHPg8v6GqjkayAEnfMa9G2JKUsmYOoXUfkJNb/p1mZOeXQfbD0sTNbkF5NCqQC0LqgPfv1
Be3RGMOQk56HQOSQMvXBcxq9VWWoNA6PSRbZb2wXmDWrvGGmw6F8myTW1TGZtV3RvQ2u4d3rYwVH
bTJmX6N9zZ8uhMzODk/kgjDFKlmUya2fidIalSvmpQMTsdOJqPzXmUgGF+VedgRpEs0qIfdNgAAu
igHDCoZuJ0hkPszlevNvYS5ObSJqDKfsLQ+i0UhD3Vk2RBMptkojnqH1eVsIoKZLJuy1tPmFfaHq
w2RwlciUjEu9Tn5XfXlqeRhVcDXtANwv5pRpIvtGOWDAbsFDdbQoYPeqURH6r1E/NEmuEVh0o5MX
igbL8aWxDPoVppY2Oo4tr+Jj34vXPgFsBOPeQCbls0qbLZtTifeP7xck36SD91nZ/Tka44dNZ72V
CajZNeU5nZUEcrNR2jn40Ym5+3dXmGRvk/dJteFVh5kY8j+k7fe9aDJih859mBhcDhagvKP7pWt3
5sQzL/AUEf6u9teuebzoFvsH7HFVR7nCTfCireT3OLMI4/DFyG+7g23XGblaaULl9cLc/+xTehhK
rvzLyXfuk+n3Vb0oZuYeWUEZ2YucsSzB50wMbqboyAGSTbkWsns8MIF4azVBZerx/YypmGVMWwIl
pYRns3/aA+s2BnbM17bjb/C4lNk8UzaZL65HyViesy4ffwS6BK5IOtaFxnoJenUMLApAavA4ZTpY
9sgn+MM2vCwHdn3aASmt0AYKpei/x9fBHCXioqoygXJ6zn4omGOJ+V59af5jz9dFe1b8Wxmkoxma
wduFIawDF3Y20x08fSS8+PXMrVX8vQAtw22q5NRv51a+uAMrCAroFxRlNaMujPrO3eSB9veBBTiZ
N1XTK+0ljPkD2BXUSwDS4wtDsJJP2QstMeCQJAlcxX923FR1z2l7S0Ktgrgw56oOljJrJGfre2G0
mEVG+ktpWKRb3Y8OjLsKsmzkB/xLWOfXV7Why7E1bTd6RpgYhctcu5x6iHbQfa1GORsTFDK7CAwC
5HkvWgfc7mqGHIBNDGE/4V2+0PrsTzDJ8gPEfPp6G4Kchzm9rC44ySEJ+3LazFGzA94AU+FDVaqn
qYwxZsODovmFgaZ+jLFmHcpSBOHUTCkiOqEzjGDNys6A+fRwcugqtq8p9wD+V6jzbkbi5Es/SjWX
iZDe0+wpVQlNh4dhS/6yBYwBSE7wU77RXDJdn7Y5YLMjWhiyBhCxrpqaGYW3LuvNTHDWZl3C39rK
Dk8sKclCeSty2b8NxYBohZHl960jdXdDqxXQwHh04OPPvRMFbgVvhAyamrhJ3FkCp9zEndIy2ygc
zAewqvEGnNpeHqtm62LDdbw7MaOWFQWA5tfbgotXU/PgIOo9WarJhm65AOgw3mTuwMLN5yc46CLC
j52JQeHAcWECQ4SC7wxP0uB6ENyBvouWN7aIpFdKGQfAKsJ6RDEXjH55OhNmdVd94W/o+eje/NI4
Inz06QibmN14tUJ1fVkUitfOS3mJwWXQNVfI7GPCUdGRfKizMxFMevgo0LA5kumsbWPeDgG8KCRO
lABDP/shTJGUU3lWRZB56mL9s0RVE5LN721tfdDJT0sPhq4TZdiehUjX3a0W4WE+rRgv70n6fGM0
7ESkFxg6CnAAuTAaoUoKYxKq2zIxJOiIhaI814MhE6bgGr50ZWr5OG33ewmrKbv98qGpd2ZMXiDu
TSB38maTpeV7XJTVmd0mg1S0OGYFX073ApPQmab/i9Ie2k6bTYf9nWZl4I2Y2BUdeYUJuAVsawW1
JwSNw/4UyJlrXzEYx5TONtF+c6fm2cam+eUPBIdANEuUYPwXrqdMIQMSSgOUwlyvretS39ezkOoT
KG3JPxfhamBnrE6s++11I9P1poAOlPEtrpfxpaaMO65bz2E2srFSfbOUAUvLrsnEFUHnx0mjxTks
E9rqIbNKusjj0rrr8i2JYj3MpVfgD7vRjex/rt7DzP9nKurmYeWyP/+0u7/TGd3dgg3tRDlySUCF
GQpwHF4K0IrOL1hFbRpTz6a8v5VuVLJMV7nSr5IaLSNcZwNAYJCrAwTkUOmEns7y2H+ZEzOwSq2q
VTADeLXXsnsQuIq2eNkd28yAWZqV9ub+IJrPR4inPHuEDFWUS7Ah1c9E7aIPq0e1vF38zoMnwR64
42x/SoV7yqL2v+cF9S9TirYMVG43wGOmEK+0BUpIygLiEd3Ae7alPBVXBvyfV9+ZBhNq4T21gGuE
0WFcbT7Npr9Jg5A9pw70Z/5oMnKlHXazS+5J3E12Sjvf7Xtcl5yLgv8AJr9KyGSbHgp3GL8fUp/Y
nbH1Qj38ue+g3SQrABrX9g9VgwI8HxYbZASFJghm3pNj2Er8ic5jdaIHOBZQs341vr7C7Qaj9AKO
CWXbxRftX8clQX4FAi7OC+WQMjKBrn09+A6nffu+FsV1CpG1DDS9eTjyQYuNezUG2rF1YBHHMjgr
+OQiaC2h7tyFStc2X5lUdWCEtW6qShoqcoUjFHwltZMaxZ/XPle+FZzXhhTlSNyojpSuEKtdwxDv
OiOnb9qAxfdZZj+UTjLi/w4xJC9dxaoQEg02GwUXvddCMdgQgB0od3H00ndXxbKXixfURI89COx6
2FNUR5twh2K+IZsAHV/vofbUO6ZEZXJYw2ACLJTEFz/CdBAA6m2uMgmzdI/yHFBWI2U+u7BuNBuA
A7HLAIT9231/JuVitWzLoBdmF3Efvwr/9b/EXtOUe6kw8nSBQQCvqnbeMPSyCCdkMBWjgmnSpeq9
4pNGv1Hi5D5AhwTI240Yx0KTq9pbomMtFeRL1+xcdfJCxmH2MAkhuL9jHZkDmyIml6HJzqSi75H+
i7gWvB5IXQDdmODb5KZKEuyKsMTEvAe4HjrnY3iujx/ycds5IuzNRmLnnrsATsjWz/8BYgIELvKr
ApoZzVZJlRniyirQx6p1H8c4hICgDu9+JVQN9GIR3Uqcwt2/F3Tt908hrryx/Q/3S1iKpmntJBQD
ayUy5uG8yL+kg4pnY+JOQ5eNaJ9CSc10HjVjXSpQvm5dVOpAds4TOzPBFtO3j3fc5eHGf849fKT+
3GnCtynknZV2tbuOx8g1ZfcnXb4veigWT0audLL2UGEwJcfu0UEvakAJVb6l6XGS7o4KU3tYQnCf
k1k0qLw9xszhQN/VUd+5NoVyG5aglyVsdI9gLQ/auwfuB3qM0X5Sn7ucdWYWvJdNB3Pk8d7OvL/D
geUTS4A5mzOR1/O9gOkpHammsEjLU5VCS6dbKUQx/Ha91WVO+YQs3BefgANLNKTntoUjRDUtfNBY
rFR1eWMd4VZHgqugROeSqFAu+XkIHasWw+hEbBVuhMZNCAI9A16LH4LQ3kYEJOpw2hgSDKmHn3uX
rjluM9osgbtXjnvb7pTCnAUpcItHNGW8s88/leW6UCzHoybpg1N5napIZ8olHYMKiWmmkmfUNhw6
dlcLhM0fm4xpTAu5rvyNKIbGb8Iz1gcuOV4IwQHjWtGkXKZaflXnWRJVRcV2uj6tAhlM3S2MerBr
UEQ77ShDsDU1FO78aHH00YnfuYS5AgOSHUfLJ0EY0WMhYO5JMJ7p1Mdn7bmUPqOkU2Dg/zKLMm1Y
oO4874/yo4yUbpX8x5+ZEaT4UtfYlkOzS15XJV6bMvP46m8EuQU22x4tmMcuxF2092aZA+GcIK06
CMsUgFCfVOGB5qCNNMk/MBEa6koeKIJmfHQu7rOOWFJ1YHRZFM+UuA7wnkhdVR8AV56PYVrURhFf
Co18tNpy+asdo6WRj/cpKeugWkLnQyvHA/4TC8JVeau3qq5yN9lLLdvuUO9hDZBD3nwkfpSOt55+
U3hwN91+siopDt0g7DXWD+WXvWZq93XdJitG02Mr5yo5SZrUa++lMR7EhOGp3L+RtfdNPPMv3d+U
UoIR0hY0Ze6s7D0UNuQyBm2HRcCbc55PuhKL7mf4GdO8L3qICr1UuHw7GtBhg5ZOMpZSxQ8d3rN3
K5iWQqw0ywbVTzsiOgsy7RGRL5Z4N+4QwYv6cLIXhlOvVSX3IbigBYLeYfPTKxUX72zEaarQohwf
tMNGIzOAGwzgHi4m23dvJbRynNmiGEqPYliktBFAsqCDfhV4kIi6LOj9Nmf/P5tlq50TwSMmc1V0
4DXIqA9msNZmk4LWQlG1pKfZnFPXLMsg4Cq9XZCRY+Xjsz0LCoPdYcEsRJktnKtFa8/As1OuAF4U
YfICbRWiX5yn5VT4ySp97IjgV6dKaSiakvvqiFc7OWtbI84xK7TnPoOCGyNsZ6s4PK665I9LI6oq
oTq8a+TyNO31dKBllyOTYBBPBdPqIYz2RM7xmhPpLSmFsVM7vwFXChWaXhSO0Rf4KztjRt/uhH/a
RDVeiajDdVt6aM9cKDFv8rie1FAzRdZKGAIz6UELZ8T6UQGtWROTpzU9EW8x4vTTLzA2FmWVt6V3
mdNC3QPwbzYYcc3J+pnBej9L0XR4kN55Oucd+GDAm4TX0axJBrMJ6eXHjTx16qz8RcXe/EXAK5Rm
l7ZUZTlWGchQqpjFOJ8N6d7ZddMsyNsEV2AE7d9QK5VbKz3V92WJleIhEFUKj+ucjUGYZVLLTgcX
N9PqQyWEtgR0ej1bQA3YBGsnJVIwLtqfb6En/WGj8v9moDads2jpyBH0IJkKL1oDjwiAVE8U7ly+
MybNLf56N5vajaoza6JRmn/XaYMTNOOlSerBpxV9re//zxl2MWNx6T03rQoaQ+bQFiV3kAXFecby
nAG6/XojTsfrpX+QCMoY4y3VZ/bgzHjw9ntg0duyKfPkRQonxhgqoDQ9mTZomNHaYI16J/yhGGdt
JQ2dgr+P7e0+3XGi78Sp7FMnEMruANBQoy8tfhAWm0YW4Oktc2snstreKcs3TkdEtPoqkBjhRIvV
SHSx0coZlAzwp8Rv0kJcQQ432yRzs8WScr/lBL/uuxzf5XCtn3Che0ki3zLAq2ZDZiKEoWlMJVwz
MFZIiKt/inS7mWQ/pEJLeTJcCdIS35I7X9kNQHVRfey2pr/NscXMrlKI7v85WMaJZYloVwHiRujT
u+GCxsKevvOEPXSh87utHLvYq5mPJJOgJTbt4pdWhGDUq/8s0A1RbrlO+5wTnYRbK3212ZSVr0mP
RQJ1LFjpr6sGFAa/b617igLB/CiiKUj9xKc1BHAwl3Nw2Go3CC0JBjkAk9i/n7Ue7ViblJfek5CM
7XJQ9CS1Z9nVoWlmwecY+ClS/3uFhl7gD0cmO8yslcdO7eXjwWhAId5uAb3gsR+Drk4vY71l2BS9
dPgDoQHl5VDuqUO15oV4RJa/uAaht327WUElqdoBQwNnJJsW61n+CsJjgn4xKLVMAOLaabyfAu0W
4Alv3220y+qgH3Ip8iVjSRdR6gWucCQvlRvdyC9W+7N36qzflSWrNA9WUuYk4xSxREe0+sUCsj8J
HSzn7gOSu9i/HxZgNxCKgmhL7d+T/ybg2NFILfva/IteoBAMTf/O2RbMZ2ixZcHVmrAyt7Lpaiq6
g6CwvB26954tXKRN1s9i723kBPqZ6Bf7+m57UAmV3lV7Q6zo7wP8ul0H8OxBsRKA3IZ8YLO00XFh
J//CxXzHcPKPq0fxHz/pAR4gq6BpnCJM5kgP814eZP3yEys/wk/3xixUhr/k+1107DPAIq61YqFB
7GJ2G4jfqL2ZCViPE/2+OdqhLLVG1pfboitk8e0q9jGjVHl5t+02fxOpxXujt8+4d16RP8em8i+E
paiXSUwg00Pi0Brb0IcGw7L6gUew8ratgE+JBYSp+qK+vjIdnVHX+NOB4qO5ayiYvaqry0axgQBF
RKSFS2VM2iCOODB1Ywkb2eDP2YQqFOrHcOGmbR+hcLrr1G7e8/i3TqLhUJuTJR472ayQOXv/s2F2
XPdJOKTD9uMMboFZH/yYnz/PJQUPvesZeY8UQ0EGuLvBbhKtbvqTH+xxg5TsOZDrLqQpiXrk7+U+
FHIkVz/ORD7DzT1Q9JmmLw3SUb9VWv8N/EVQQ8hnMepWABWGM1nxQK0eEj2KLi++ZYo587CRQWgW
nl6WmXFuAwuo8pCd96dGLXHCjUEgigvB/Q9Cp3salpoT1X2jhRKPNRfIZedOZFFEunF7QfyIIAMa
AzdaockBJPd+NaVcF+/wig37kAm8amAzZ8go3pwSkHOzkNba8pMHZ0RSSeOuID3708nIkyXbT1Iv
GZNh0C+2+4WF/54AhYKwel8o9bw+x0rxpGmf8lZe78fkH/psxGdzLBlFLrzRXaznG9GMratrovQo
fPd9kaDXPY2efGx2bc3C3hiRnUAjOe/obxsBk+Q01PRJ77pBEokCH9k4rVdnikACdNfCTYcrZOAD
wQrdSVl8qu/C+2dpYF4VdoLDAqFaWvkATkuuCRdtyKgX3Gi0rjzcj8indNJkl/snPAZS68Bnu53A
W7Rw6/6a7KAql+Tg3anKI9NWOdlDnkhj5Bv4epBZ/WLRo1Zzg//2D5r58tV6WpjVf+JApOClVHpO
VjpJDVSSocCzXZJ5KzdCddqdEGfb9ZwyLTZg3t6HN+kBs3kTivlR3/NwLy+O1wqVVnO2yqjjArh8
SDkExo/rkXlkJoixPDiharjfL8p2f1+0vjfOciuCeYhNvH/gKdTcePu+gWuPj4Y+D5qXJouLc8Xy
a35/1bNuJBdA04pvL3MHQNYQjDdyGH4CkYLnQ3tP13Hv9+LhYmhNb+/DlxuQbXcw7c6mJlWaU6LL
LiPW53Ga0sT0MmV0oGkQk46EcowpVNlxe7WOWq4StJGO1nqEJ2NKPC2xaRj1fyr1ZWdtA7D+6tFO
XzxXg01tZ0CgX3lYzZqkOHluYDGb07vAwZ3nt0tPoorxS93MzRYLnoDc9hJ8z7e9f76smQnU5bOI
sG9QtPuWV5DMDH7xQa9sXA7ZSFxmhD6FAbV2a1Ly9laRN5xHEoTvSgRFLqjrGmJX7YlXGlF1jIT3
jpb6UtQTQuV2OuQjwwJZ3RMO66b2SkCuREWtA18qV7yQ/HfnqwxygB2o/wix1GFhaR2U1BXuNCok
4awqR57efBCw9XDdVyxvACmH3cor9uAZBaI9bo11s0NuNQgzPBjD+XTjF85Wbl4gn5FQ+5MurVUN
yG0MsX0uh3D9m2Xb0pJhArHsDljr2/hmv4KMB/T/262gJ1i5FPwA5PF6eJM+obBKtJyjW5Io35u5
0FO0ldcTuzMLlhRX7o1Hj3rwMaUuuZW3uSmYs/7KYo9dkw376CH+vopM/Vwsehwom3k0AUoQ3Ogx
MCPTrWUYj5vO/F5D78vtqRO3TUCeJtfMvPgZcopSUds3IAMj+NgAfFmiCshQRR70A55UKwZqVK3u
aVAuBAqxal3yrmScHYfSu9kGrlFgfEsW6OADTWnj/GyWcQrSreyU2Yl0sCjiQIpl3cC23BoO81dH
DGr0Hb1XsKJV0pVHIvQ4e+1C3ar0vRqtI+ce5NmWZA3y6DbhiIAI+eCWvtxjCNjP9a9Yv0VlzMjj
vTegYFm8vn1gZ8Doba9Qnlco4/RlZwZK+HQyoXBOrpprxFGDR8g7NlgAFWX1BvBHil1w27E8et5w
aapd+/dpdEo5caNzoA4vnoctOe4vi/c2UBdBb6EetAqEKT/ml3qn47eDip72g/I7Bj4FmrFHo4r+
nCEdgOcXLg2QVdMhFdRZp/B93QG00lgVoLQx5tlLUg1eKoJXDIiT1Y+mA4kT4WLMgwToW/KKbILo
eTIpNdoXsW9obkLcMcOM8G3XMGjfHWjXoChdgiTGb0FiHPxAopGeeSIn1vYDAhpdjAXmKH0+4Dhh
1IjykHIT5m/5V77s0q+0R0lUj2sCZD8vNZPlgDHEhcJbETLK+I4Mp6KPZLGf8X0DfOl0UqbtVSLL
8MJVyDG5siE3ESjlunQ/q3MrYbMzx7Kuxb4yo6DTkfbShP1y0Ay+Gmnp8YqS3m6VdQO+7rAOn5JT
kcbDEhs5g0I2xiwBwaQFD8b4n/kyh5QM4Q++wzweNQyPbdQBZXkNrV44NPLPGNIn7zV++/7l8R3Q
DEObg2kOZf2w3f5RhtLB2K/mrzTmbUv1Fbur01R7qPAb/9if81J9oh05y63y59BZDEKy15HyQZUd
mTcIJTkeiRjFBpLjwybFqWKa9qFJZ4kA4GV+MmPdtI90hDQohFrNMT/tYY/0UNhHeY/UYRDR8Cvc
pf4BRddCDxpUauvPF4ho/YhV/CIp+l0PbiNE/ljudom5atAPmHg9Yekm34fkIjlBKV65EVDujuz9
6ucJJIY8jMz5QCJj5CEX4qyNeWdk2siJ9HB2u1wWic0alIWxR8cAvGqyb2Qh06598QPrj7yDyobj
a+3c4VGRb4qAS1Ta+Vj/0OMSk+m9EG2xIhdO6rWck5cUaKg1n37ZJmn9R4wY7XApCoDXpv+hvoHQ
4I8+LDBKcA5iRw7e/7EWqPs88xKO1mPSerdz3IqduNGckyNdwRvMISWLPwpgP1ON2MODVnlcsXcp
TR4Jv51c7klfDDCPSPf5YxKIaJKPECdfSUXpNBkq4A7gZVQGYN2JakBN7jTma5luKhxe9fatz5Gk
c/TlOCV6zLNeYejd7nuFMh5tQhGF9cescnteYZOCrOKgebOmLa8llI/+fhaarodgn/0H13v53UcX
EZpflh4j13lcmeztG1xsd0du89pfQBmAOG4tuEorwPqITYjDKJfpovBvYwFn79pH2+XhTb924M8O
1N/RllTSGNjYfJFfX5Ye8nD4O12Awn2uiDaRwCVFZBuXkNHTwsY8J+QtvmaMMmQ6D5P2+zIvDoZ5
iyGlvolRDEaCFefxuj4NqtOxzSiY2ydFaPPc8u0dN2DJHe97Lc4+1b9/VPbjUOasMlhCVRpN1D/E
pMgQGZXziUYXXkd3qtBsQIZyz3DeDUveLL585hQMQ8at94Lf83pWs+XK/R61TOnA3vJxMt3Ez16m
/BMT7AT9GcM80UaBqRSrvCnN+KZAdGw4ei3ShLwcLpDa+IeFVfFKSJxzLybcrDj/XhrNiWm4pLtx
nsOKqB4b1/el8xVoezy0Saqmb6rgJg4BSN3dJtfLfIbat9DwJ74yBVI8ILnAHFB/L6d4XY24SlIr
9Nmbo9f6Lw4pwLjXOaiZ9OJ60SX8OYVA5hLxlQ2ap0JcgOrwnGQra1kiemGF5QUBHV9351rPxeWd
gyznU+sIAhb78eXv9NYqLsrNabRUY+rG5WGqf1sByeI5tIPn9WhCDhHhX5IO6fWfVSh0zxzYOtRu
M4NPtvb8VyakWQqqb+9H+Bn5QltIZtpuckg9UOsoeQQT1JxJgfXXB+kAaLobSzXX3mV3n5z4DUqL
sVkkMkR/zQ8lPw6P6VXjqqJXQt2ynVcDfBG3AlnEJIhK+2aEDtFa5FJ+03uBeGZ/5PIbhThEdM8g
lds9Wyfr/H8yRyA1dXd1Y/NwGRG6YAc+uCWhg2C6kqQBVYvFOPvALGlUFQUu6xzW4jb0SNsyGmrY
MNo8vyT3GUtp8KtjQriYeT7e8sTs8ix+2gtE2uCKDql7TMlyXWXJnOxfycH/T5csi0IxhoC3c4C5
1Slp2VEs9P2HNLNYc7PbfC4lALKmCpO2PBgoK+uTEL12FZBVy8Q4aecZB30/yY7hZbDUPF20EQaF
P68iED2ZxM0aDrY6SwtVqKevb0DdvVCtH2vrGXDxrK+AvsSIT7XKE1HQfY5vCGHsztwjyft3GFyf
50woSLUmLLIawzRHDB4wfcpyD26091wfdyovWO+MFOhtJD9dmz2irYNIbxedE8FDEDN1zdrwemDa
mY43WT33BezLibM51XqGG09sGWwzUlxCLx6tsqsglZTkASxk+cCJG60B1IBH2IwWJe6VNog3xynT
DgpqKTgyqLuyumq/qohE1gicvfdDFoTCi9WaiAiM+mF2JVm5K1KETmgvdEMN1jBqvDZHF3d29LOW
Tra1uKKhSJwy/iN8678BhnBhJlbXZyZvG7vO7axTwipWgzpSR6ZsC7/3adOeTWVvOsQhj2XbPpfz
QezZW/rQ2VAtvUt15cdKg2YfJRB4l50rEHiEokGjHQt94PDCX37SvA1d2mgzjHjTAoHkBhDDaG8h
IuIpI5Crq1BuTuQYXcaDvvZsBMD7HqLBOXv6Km39KLvUHqGB5ArE7JPe5jG11aXGgrHvZylV1cIz
+J8VsDNS0mz2YCVU4a0D4lDv/mVVOwDmOkDXmagSdI8RsNuxMJ98egY+Eqnt1Lzes/G8jGzQNuqM
0my+qFeYl9+4ZoTr9AcDgv3pzz4ytu6YAJWEsTCt5Co1WlyqoJdjU4OJi23EAym2ZEuDbexmaHN+
KM0ZUry3urgEJElKovtPbBh0I8pbqFQrTHL18EoefpWj8fK7KIONFaVhj5gX+JdHVZCgbciZIpk1
AbKQF04zUf3AwburxsYbHZTHigALeuD/5KUsuH57Xaugqb9vT61g5BpCPUet7KQjTDxy8PN1XLQk
KOE/+QyMnH/0Kag/0I2RQgD4thL5ahjSR7e7lP6wrvrXTTdiW1fwAPQmR75Kq8QznnGUKzPBFfbM
fmo4sR+8K6JX/zPm5KinhVQ6Q5HGQYtI4/K1vF1nXmFtMgrXOCQrjiDICbgzYVECdmw49VSaJ4tN
aZ07maFAG7dlgqk9TeJCsuPOFwQQ2BICuK2ICzI5XJyR+Bo5TXg23YbiuFtkDD8nj3A5MZw5b4+W
PczR2HmQGkMuDWuZxOqCP+y6o2l14VdoSLVOkBxoN4AZbKSoFbmdgQxalfLlFXwrvVEjjLIVQfqc
x3WCOwPNn7Pj9UhNynlOawsXfcJGlsOlV+y1EOHHS3oxLX52lo3lm4Un2xkqp5Jxnl1BzjOtZI+R
9ZK1JHNYorombUCACPXQbyDbtgWrM+mi7STjUqCCCgrttpYllihlF0o/f8IabW5G6vA24xsXDKVo
OkOUGDf1h4n7/gpfnSlqGZxm79/Npqf4D+Mz+DhrZ8dkPliKCaRZ2o0JjdR8nqvn0oWU3AaG3MKX
SDGEhellzkkzfGCmKAFLEBGopC2j6cL7xWpfOZxUgRKrdeiPF1FjsNOC78bT4LfnweYRe250BsFs
g2N0aBypWdwIZQUPLkaJFT52lYo5BLvjLlU895Tvx7fAJx5flRQoM7p+R/hvtWylAfmhivXOAcrs
XT5XXyFjHq/XvK5zPr1sAJTCXFmPe5s+R7SJoEEwwwQ2iLoS+POMpO5vDLSWGz6R6JkHEENx/fH1
LLN6pk5MvChWBZby4dO562sjr1ynjm9DjUoFuSbZG/M3PTpE99dhdheZtQ3vGnkIcHQt0KI0lmi5
0d3/VapPsbPm5O1JvwO9RFlhvBerTXUnEvhWdJMsZ6GgiPwozMe7P3GIs0rWEs3X3DwZnvFwE0h/
xjVl4iUjl2dyLI69xZzIsRHn2qzOO0KdfDeU25inHTz+yrPogUZKp/1ADR2qjq1gKbZ9yvrydRKD
roHJZqiMJ8O1B2VfE6xBM4/h/DcTy/xto2BIM8Ml91RtRrYtXibFn1Z7RkiiqLU6Ab7ZFgkFpW7B
g5syEsHkvawOUI4+vmY+f5oJi5iA70XhoNbZiD2F4VwI4LKytpwNdltJdyh4yrX7KYuPPe+mZVTs
Ysty0H0rJyk/QW6T797ji4aCwBimDGiB9IfVLAMIXuDc0vRBkpnXkkf+BI/gM04hE+ye/BgtUjHX
PJnRYcPlD+6hX8OnotUjyJTqJv4+yzhIWb9Wj5cuV9jibnunncYrZUB8lbjtn2SYhYlY32p1MEWk
atHvrTi6VpOIIfC97PSsCUOogSWNzJPYL/h/vlK64ngfqnTaDlcOMWINqnLpyL+3UipnCX7CgUPC
5V3g9+DfJAYlLH0Yn71BUPAlihB5o4srvNxdnvc7Hz4HrJTC9Siljy+9obn87jvNcSEwRVfwYODz
F/UffWQRht93spYD6YWk+a0X9moojXhlVNZZeNMeZX57Sc20YD/9o/xLMewYuVEEXy6WVu9mBrv1
YGApjijOE/kdqZfNGrp0nO6c8E9aXIwemltGUJzYNAR/CjV1xqS5smK9FBxYtP8ygRTsBjia7gir
ht9Tabv5Gvf1tV4kNVmBKOsCyFYWmDN7d0groI3NqPMExQvxcXzG1Bfl6jnLYmWotJjb/TbEn8V5
1LdR52cfva6DwB5U2Ecx6NVleo4QRpuf09KSyibxF0xGUmy25WhYe/Q1YlfO4G8apLiGM3D9Ylie
TTbaj25YhFY76TzPr4hW3SoXiUXbgDHo2gPxw4As4B3uItT0Q43y+rUNoEF6RZjM9JEvtryttELL
TQKXfZhaFL1pvaSKIrDE9Hrq/zCq9dnBkunSvn7D41otN3vwbiiTStMaC/36HA2zMTXNs08PxXzk
a5yxSWwkU1DtXnUe1d2ViCv0FXa6uK5pzVKoEm//8QhuNAfnoKfCCt9qGtkcjqPYpaAbbvuIDqvX
ZDqbhR79p7nPNe4bFShgtvjr3gJVRm35czbhIoRA2CyxmCPh/i9rBm9CFLyYW7RDIRL8jVRrnJxF
sUfO87c7SqJwrdFuER0/EFklnLOm5pGGq9YvVeJzhoxuwHnWh3+JOAaL2l3+ItaJoLRbcjkoPv/9
l1rxP8SzWdWdCUedtJnp19eWwphQtmuI+2w+/ImtbXNblRgGTFApWLV3yrcgtb4rrf3UtsIrWhqp
VKgGddz/V149gvNgZQBBIyohDmpH+ra/2zRgssAA6LFHx+VVkSGU4VUq/4MRJ2s3fDRm4453+gL5
xJs8q04+k0jxpVCNmojLWcibluqntW7Ur+/+8p9TEo8mVW02dRhUnfv3vbluW4qKdpQACR2sRieY
bGCXbHZlNHQ8f1EjelKY8cA8Kw6/mZgeUlr/0/GI91fC4YbUdX2D3Tpkh8vML+IOcFN6fiApMlp6
X/yMIRj9lFj7SG5G8x0bO/NF/8YPJ5ezgCF8B1Lsp/CII0GKODEnc7aS/A6xUiaxFV+Q81q3DphK
Dq2xCQQAPpCPePwdijTx4aWvUtqriwA9O8bse2woxjnQjdJaO9eiJ2+ZEe7YcMa8N1Y6wepDm9Sp
FIk7x7098HnuiKQxls38+hVTETG2XQNqIui1mq8KDh6kwgWEBkljtHvwP95E8lDjS4ZI7UB+liQ7
NhrEgldIWeSKCJNPlAdeaTk6x8OSupO3qwaz7EZ4HnpGMO4XFDsrCL6ufVqiBjuy/uw6AivaSMKQ
D7NkfI7IvhqoJ4ZDUohguiO/w7oSSxmNGZE5MGkPjVw8KA3tKnGip9up9o6/lVEoTkQEnmrTW99I
5fcLZzeiFSR5YKvNSTRKQ28FRWze7UQTnNNPTyewokE+qbR0Hks9DihN8zfdG9Cmdl7SFXBz5QQK
wJzPjpjQHwJfQuWiI2xzESzJfxvwflE4fUeHEoTKcoSOT+NYLV6Vt5OgthhZ4RhlTjEV8FmY/22h
HC71GucD8OO/DNzfIG7YK1OPztBSJcMaR38OJeqTgvYm/yPuXmMk3Lw9FQLXL8fVCAlhtrCpBl0Z
jDjTNCr1mrVTQHChXDHl1OG8dh/5M0x7mosXsPV4jGnUDrmxmP+bYoZbqIf/J5CCIOcMfSVHBWiw
4vN5hGA=
`pragma protect end_protected
