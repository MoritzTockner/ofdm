-------------------------------------------------------------------------------
-- Title      : <title string>
-- Project    : 
-------------------------------------------------------------------------------
-- File       : rx_input-beh-a.vhd
-- Author     : 
-- Company    : 
-- Created    : 2021-12-13
-- Last update: 2021-12-13
-- Platform   : 
-- Standard   : VHDL'87
-------------------------------------------------------------------------------
-- Description: <cursor>
-------------------------------------------------------------------------------
-- Copyright (c) 2021 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2021-12-13  1.0      bauernfe	Created
-------------------------------------------------------------------------------





architecture beh of rx_input is

  -- signal sig1 : integer;
  -- signal sig2 : std_ulogic_vector(out2_o'range) ;

begin -- beh

  -- outreg: process( res, clk )
  -- begin
  --  if res=reset_active_c then
  --    out2_o <= (others => '0');
  --  elsif clk'event and clk='1' then
  --    out2_o <= sig2;
  --  end if;
  -- end process outreg;

end beh;  -- of rx_input
