-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qBddUAYg415c9odwV5nhUtEPxsqt/N1P8+IdIFPxlCils4jczRx1Ly2Wirhhw86bOa7rwAh4Z9Qb
isxHrXvvOODpAEHwsN+FBJr4Pw718T2GJx8wLn/x7ic1X0mbl9iJY6NUMM8/mBmIQW+wacCPKG/p
vqf+aq32VhnDper+ZAG8wVP4QghlqQMnNnFkGd2PuIkf84+x3iL2EISru6uhe+9npVVSNIs7KmTp
0XvMIUpYUHtZNClr1/LF8CmxyR7pAo9VrSQQDPceoqDwQ2ghyl1j8b6uVXXr0Q2c+CZ7/cTjbC1I
BpZ6xBJOEQAZIfki0fUJvSyTr34r3dcYy9ymYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
y/djSPvPUxMV2svCxz8kPm2brEcSUy5O/QJvXId1/QIQegwqHv17YssecOWGHkET70YWXwqJzpPp
1BAKXP6dEIHoQ7npQwmuuDUTYIP7yHpqvM7klCg1mq0guqSqV8eLg+rv4tUwR2gBnt8BeP36FmHm
n5XR2oWSDQ1UMdP+O6t4Lr3dyJXsOxfPzbdLcIKCWq+5V20MAucRQfqjxIIuxm3Jex/7vNdk15sw
qEz7OhWJHrr0AfrXcEx+mlYSe8tu/e1eO7zj0CNy5MeI8xlKCcQLeEJVSbjFWvIIW37ybfQgfoq3
LeGB4S+7TSriGlumYKEOM0ypDvspxtMbmZLI2+CwqS7ROAmQlZvVKesmstN6dyYXUpskTxYau4R/
s4+jXAEUlDo05TZcqE/zZeiBoJAw3K3ES657VLV4y8KE8g0w13yD/b58mIuGeFKArMjujXdUTZdT
eqg6LAuuSHDoQ5AmMvmFfVd7DcSHvFPugGvQGwauEFXrbCiOQ+OLoSK2wW7Z4KSt17/vzvHPWvyv
6GMfacbRpYq70zRMm20T8FbBIK46oNdI+E+ET4tBvbIbfdT09IuVmUILWx5FbVK++OtSVrjPMcD9
4AnSovL0zWTX7XtFOAxsMXCt5xmJP/kRdcF8fGWYMXumBszOfQ6Iev8THzfwHhTNNLQQO85Aq9q+
aSMDccmb/txObBfJQnisGOQaTowvEtvlU03yVtER/p7KdciNTZBQOw8Spff3JCZdz6h+G3RxD5Rm
IBn5u/iap3oV5mOAfPGYhOeZGH1vmIj+NrXSUbwmj51VyY5xJXtoufsRwyPr6RzLlDVbMg3tyUYZ
IOp0c3Q9eP6pNEwevEsM2Nv8tuXDhgt8dWLrtPCzzPZE65ORyMl+G8yQhgDWtsvT1nptoZjiQCTR
jKJr01qyOFaD5lyYOIbw6svJhqskdZ8sZx+GpTNVJaXfYghQF4Nzz+3d1uXf8/xWFVq2f4ooLgKa
hsfDXHrQct/sjZIY7w1c19LRyDiw2TB/ddzlgrLUdCMDZ6/yGcFLkF6nYOd48gcGyCn9PhwuR0Aj
RHROAwIkdQ/cikT4CvJMRDackZ2OyD5EAi1nqD22stI12RmVnQ/5UQp1AfwPWVBjXXdUpBesol+5
zBMls8+gimwuprlybHj0TTNdd0a6U/r6iz3ET/YD9UJs0HY0fESTw6BKuUPf/74bM33aCBnXYm1b
f4Vgtrz2J3ygfZCcs8x6+GAacOKdFYUvZgqH5n+kGFFXLhqMe4JZtWpwfoKaUgbjr73JPlQ1Sw53
1fM+SVe78SxbG/YDffkkzzOr+EjPyE3gUQfQMVeDRllsloD8sHYRVEpjW+XPUhzrkxxScJu/pMYG
/MJDR3dFUIleXqvcfbW/goUeHA2aiTIQMAHJ0s7MEb58b43+AVCkTCy/3BvBQyK3P+nQiJ7qnnPv
ZkBKiLLsYAAp8H5ql2ttIgCzh3jhONwNhtmWpYMOXg5uIXli2XPIvLHBX8K3h7lqpE0DAOGv12IP
4zSwIhA0YCRaCGnW7CjUc2JNq8MlizteTul/rLSipcrfQV7UaDFWWl0SrWRHzKAidxUJA83VyEa0
RzlO8lRtoxyfcruoYfTZ17LsygEYR3zgISBKvPqFS3wvBNIUGhLCHjfZoUrnU80whJ/4Vryb2YPa
Xh28nNlfkuczru6gc2SDUqp5C8uETTCmhAUu0nd4XXCD6T4HYyNONIF5+dp3qtsd2J1S7hAhXOPM
JAQdb/uJodrPMyPi22Jh5ci5rj+wCJndNpyp5+rhqLGlZ7qWhIFD6gqoUPDOD/tOTXD7/yb9hW7+
j2dWqLLJ3zq94Vp5AxRXmZuoVjp2Ezxi0ezCAxtKBtSyhZD2+QeHQtPrpzTM8vFSKo5PL6Rbjmic
QFwskIRfN4UtT6bq/A+1lcpfAwZKKX/GKLXCoJ5J+pi6Un5Agu+Bz6bJmKwZ+QqJxrTTLlsUNhwW
BSEp39SIUh1hqF/lJ/r38LdamQac3Ijb76KtacnaS5QNHv4h2/JP9/NDtLnVLZlybANn8J0iPmPE
B3rdlzcedHql9HnSMQYVBloPBuT9Nw4c7rfia8s4TvyEXMwQszQhZrn3s8W7Md6QOxvrJnBQDbNq
AgA80Mun5pP8ZDyjsqEKdm40TjtgSW8wGjN6nz1esGyVX9p09HYLYfYBwN0CuHcrxBkm5UCNG0/9
OMmtjlut688Efio4PhbL1/or+/sIuIYZN4/sUfFSG09lVsG7BeNKFC3LNtqZ0FbLonN71oeVu4bv
+EmOC7JUsL/orvGPJEt7F3pJpNe0yhQIIEhOCh8urTMOOiP2hUrpcRZx+52ZsnL/H6i69mICrvbG
9ngJwx18lqGFYpJf9wOF9l5wkmNIswojV6sX6JBlbb39u8+jFKFAFzGASGNWKxlouBdxoLIoye/h
gdTNxEO+UAkCYQUv9NKUXWvaCDC4JRXLJhgmZQyp6eaOc2haOq3nCrUCzInAHFhx2S8rDWYYWThJ
XIodQxluxn/AmWh7MKqtAoCjyw7MjTCjggUtkPANOqwMR9/fxeRsJM1hnzQhBl+nZDMTt0uEn+rk
q727S2YmOkpg40JI7hK5xWnnJtn5YWSHFWayuohDSCS73co4Q88tIbt1puqZabYViQ5TE2BauX+f
R/Z2+LWQxjdUEFPMijEho5d6rzlMpI97vUPMwQqtF1+p/A5gb28Kk3bJ5TZpf753gLjY3HK+v5Ds
ebz58EvHDJLUxPFzHuyNOlMM9INMNnMO2DFExHwCCx5rz8XcbuuJsopV4wsyx1HA/fXg+ymoZZ1U
rEQ81ZqTNqST0W+ZegMeJRjVmEqPDfnCDuRRRsYOKRDeaL6HIpHBqwRZvs5iAeWINuiT5XQXe8FX
l4ER7aLvXEo3wa8GqwpxSg5Y9VoHVwiCRFBlkHf0BITLsavRwvDvlEK22iinAt4goE/K4vvAhilm
4Aw2TGaZobSnm9fITPRoCa48Dc3c8woDIDzcGLYPGDRcH4UVN0mlcF++XIGMopD/lflPwm4GRGtr
Hkx7j97pxqrU6bCJHGDw9XI+djdMk1YV9RVi5j53BtFA8YSXppKsj7cpiVs7iKZMsr2Kpr9MCG6o
K+MyXtcnCM/i+vahQGGP4WKXnGVHgEspj9YKGKttFFWiuoG0mnyumOpcAkImYBTkHsSSUpErLYAE
JXEPq209JeaInOCBBFxTzsJaPRgrI50QqFnuT/6BWg6wfSqGlpznIJDLs/SEx1vtIxXZhIBs340u
Unj4OTOdrr21AAGHMXNI9rXc0pYBHTWGvQcFiXI4fIUSghp5TVY+HSe2dvBNbjHz2vZm1EnAg07w
qmntmJ9raR6XoOKsRhzzG14lEoP7PEs9XQEIH/gD85fQAUDWChr04RyOqWfu3b06ZYY5lqXdkrGK
sLvfqWgP5gPULQccfxcNkcMue0duTKYW3VXqBuXIHkRN9Mdy+1eBrv+RW/PhE4swK7mjYgQ/rKUD
T0y6QVQdUvl6KTaKSKgRzYNfaxdYBjYu5SEsQpFRvQc/NddQbGXMtHyZuC9YR/DLbwVg3HiR/+UU
r433q/zccJatAGgFlFwRZ2JHdU2UY/2UN3R0WmIYon3qntevhJfgXNOdcEZx6vKQD1OZdbuqHkng
NR0wded7L742hvZQfb15rsQWfl/H3nek0A6+dgTjzTzC3xOBxsufTIg9fEwfRa8JYfYenA0Rp9JK
Qid1xfQaWy8a0p81UTyWgtd1tQUBNRv+EHIBHkuV8kS1vK5TkWzCVO4SKc9bh8sbBFgTYqOOEQix
jDkdkGt30+Oc31gd/uAc4wL3svkJfm5gUZGEOX8kLFNBAgxZykzvbMMdhOau+0ixFuJqBoWJTuSp
C01MwzvCdKs68sdwA57rp2XNBgnEe3aSkQCtunFG95oZZROhv1XXWKuK4GqIto1mlwwdyctmer5H
CwA28Zpgi/GFqehOkkM8u91XvAgKCmRV2PHtii72YFU5cZ4vcAoFieiZpXQYUV70gjT2P9HUXUy7
bpQtichCTVzwd1BSyDfmR500mBNmWEx6rLMZiPsGD/RF1QI/AdL/pkF7SDR+yiNXY8LL+0X3MEx3
5mXw4a+ga8E4Mi8uBzVgtoFN+h3KYhk863J4Gyg6oeKE+2O4sk+I4K+1MAILUbo17ywsLrvj98rI
d9t53Jgopzhbr6G9JkfLYoI8E7KL8hja6eHC04BV+RCmL5C8ZUfwhsqhxlq+wkg9WLVFv8zYn4kD
1Pf719t8A3x1JMd2UQuM+VuJH6GuOfGwdd0iuHsGbvUElT3xad7j8jINbBN4ucZ5O7p0oWB6NcaS
KjP7e/+lA1N96ZFVkGTlQGWsBJ5KDIUem9G2ibIOFPsLLYbqKSwaF7Ool0VdRjEuqPpqrzkZxzY1
mm9fTh6OZQ0TyR6ORcsv4iAouW0XNUBxGJvbkAYqFM1OJjbWIMrj/1ZJjyzNRlDC9OZicr9VvLFZ
N9lRzesQs+fRxP9f+sABn37AMXd3yzzsoQLJOb2LEs8PDHVjSVnUGBTd/reSHW95jRtu+dXbAy8Q
uAXUvu7hyDait7SQWf3DmDfGV6/+7h5OzysZJCMxaX449asbyIe3dN2/E4H+zLTAlLAAAsRuhgf+
ewRbgqkTgUm4pP+aveKCi/I5HYhzEfvoyAU+8UK0E3RHaJrYJL00MOn7qm8A+3i4+9mOW986E5mB
o1bQsXhL2TibhEMvNbepwQ+v2x+bs0OlxhoQt5PmjiFRMhwP+Tb0prprflGFeIkUZqQ8ExYI3gQx
46eZJtKo2nq+SBroIFyjPuPCQPotLkX1rBsQs1u52JfMbQybvBCBuepLLdrwlF21ou+7f2dIUPpk
LTMpxGl3ee3BcmkasDmFsQFkrh07OlRS4YC1r5tRtvkVcGtuKThF+YT9m1CKcHBqLZI1OdTOJZCk
OmesKx2A3XuGOtiBXvAliJEFTMdxJxkhYp+zTP3eIAHqzJvc/MA4uU/Pl+8DQh7qJmtsIWvFCN3y
LdkvJk6Sl4BN3a10tbFA5kV3dXIlk7pILNnELfY6MdKd+ibp4AtYWZjI0GUWU1LREXwHOVO7wWNf
paxttLxdwBKzFY/d+NEdavRdy3NMMUWy4Hycb0qvK897GPQNqogBjE3lNpteuaJHp5ba2iUG1BsL
0dkzTwJx/EH47TB/mp8HZsa5MXbOCiW73TkvFTLNkyN4ctNvzIRUs88ErKNNNV9fDz9wEtXVE4+c
0uecNs9sHRSJGwbxkW6pZQiJAaKdy1vL5RKyvH+jCPhW+uuaUzCg/kAysfJhiyVIOq01YE31ZXEk
t5glF2fB3b4e3x7eJlXfjRJf1tCvHWp93NJMat9qrel6EeNSP0Dn5f/UbgND1EW3/VT52E0u0x6n
DTVeXlJSduHOy0+PwZCqX3RfvywBWBXHiPGZEs3FDgHhV1lxRGzGxLU3m6aISQGQ5qeDq5iusouW
0jXFHg07MSd1gQJJJJmUDNY7sNmXMMiMHH5cNsa5mViROeiTJqplzj26q9jf1OhQyk0U1Ygrr/oY
vTL2DpVM4hNTLKRrtyaxcN77d/7dXrkOO4wl2SVKvD0Wui43IPDece8BP7E8uoJt1yhE6VCD8IkF
ZHreBNtqMpv0r60mRWzx2m0g+NEmcBz6LRR0AehnzW6OvKd9jOCijJKRtb7M19HViWB2TJKb+2W2
FvpcvKJFBgSkayJUFEiMfH7SdeJOEWFuG2mfTGPHFslNUgcoAQwq9+aEJmHw9okYX9hmhgyUsPAL
YHIJUO3SsJdUlPeF6q8ITN0qhBSFWHbqp5peibYq/gf/opIycXrp4E6Q12+MHljQgByj5SWDzklm
AZLDH6rMRdBMuSME5chUYXnOYM1TnitfaB2o2Sij7vuySJ6mdAQGag21rYEHxnBxa3O5UOzC61Qt
6x/tpWY/VKF/VF/Iy/LuS/M0K9BmoALjq5ZYCLSpyuaFjsVA/rQw5k/WjqUEQk9YMr4uCfXdLtkU
j9gBEEO0P+5B8o+6LvA9P2uOFFlmAvqjMCkeWJTsBIJAnf8EhtKnE2OQLY7YbjHz3m/Ff2acnbIR
k49dNsooeUftAByTX6lMK/QiMZjCMiIxLdCrsLDRRfdZP1dlF3uSs2ca/VUTDXZoh4d0Iq2/IiuW
GaEIja7KlJ09S/tp9P/8DA8QaRafVUwHwm0jS4oJcCaIlRWCu+KHIi8mwgPxN7pDWFYxixqGX2Ri
YDYlDuuw9GfOXSrt7aUeuQlMXCLHBkN+8dEpIipRM7nONPM3GlU9Fy+zelIFgvdHhZvO8pdX9XmN
Tc90wyNB3Avd2YbBZDeGHeyS1lrUsX8rGGoGYmlXqi9kC/LCVVUiIPp+yo7CbUvndesqUJIJ0Rin
jDUByqtDpZE35sgvd0zALQD6K+sy5kkHQLi9Z3Kjs6bPAyRlI68XXnPASugNOdvavn2l/ftZLo6E
pfYXRT3o5n2yTZ/yBI1aD38HE4iUC+AN1eEi29Q5GhXhLylmbH5PyN1i0SMIDfLhj2YRLxciCZ1p
gftBxoKWa0T09fWJmKA0SIwgopMp/C45LG7/JgXKvlmK9sT6xXps0kqZbbKBVzGjHyDynjUpIsmf
wCetePDmsnVMOW56dcsowRvYwXV3hZtGFEiKTmBuHeAUDHIi3zBxhv/Er3LtaDj4GGony7PY6C0a
LXxC6Gy/UfjsYaOlxXcIo1uF+IO3bh38s/j4xE2Eqsh+KsxFzZV0l1PDrSXktebpLev4vvVCeCRk
IOmtSHXFeQIoAj6F4tiqGgKRl7kUSBW7oRvGvTSMTxxnfNpGrid72u6KXVQYzpUQvdOxEyjRBES3
nYK/76WiRVwjaxR70RYRF7BKwyRybZp2KELFCpwq/R6lKQ6kfiebVCLXlVEvRx8Y3zQsO+mny2RX
TB3UNcTwqKD0qsYyIjAfXsgZMysWIfWQI9XlIvSDrUgtRB7D8usUZ7c2qYWpKERsIHBJcOx3dFMf
+cnsNSfhbjIWPCVKxwXdPrNIylHLq19AAr18fMPKovVvjGSray2uH3ITRgz0iD04Y93oI7Ysi28z
9JAWbVHDtV7aZVFjVtmX67XHeoiCYzcE7Zl2qPH5eeI1oTjjPV/fVbiVBcyBJ7Io9ushUHpUj+9D
4zimvP0Zvj3ziEh50Hp6/rzRZlMOh5UP8Bzopc5jBA3SLPhaRTiPk8/kfR5vQI30hnfpuKlafSXp
InEybyhCR/Lbv6EkYJYjgdnl4WyNlPGMNhGRuwIGqUUiEXkjFedtk9T7QQzaDosjSHXdS5kyTbm8
E1FML0WoM3zPZc4z1PCx1eIWsgX0LulDWKeA1+fVDpw0E2o+ZTDbS6Cw3pFzdWbYKCE4kM5TFl3O
t9qa4JEyweeglcYsEHPr1EaTi7V8aehSvGqxLefUCNvKeo2I2xqFeLOlWT6fsQizRWeeRcQi6pTc
TVmd5jkUxIm2aCjH8jewkItW6Hn10V2IL+z3/P4mpS/1qofK0EdxzpjGcMtjXQHBaHM7GARmV3U4
iIs54rSeZU3uo9qzzQ+zWFRpIU7f8E+WS8UfWqcjGGUQigfW8MHhVb+Xpr1AyuzeGgg0Dr+YCaO6
Mg2vmxD/pjW1wVG3YA9wgxxd0Ycin9/Da5NMBbZ0N4xBEwPSN3/pRCUplHkYUJ+SYQ9zBNlugrtc
kVV+X/JaLh/nhxz5n2V1clpp2YUwOW4Ji+YGykgSMLVaLITSGBKl/A8GKR668eopaqqU+vQQuCav
dFZ5gLbPxaZPmsjoDWWuiz80oMOVid+ryyXwmFZqFU7RAk8zG2Jjscywq3WPCHn9ivPjK7odr2AP
K2hDR8ZqzqsWrvjQ0aq2r7bvC2M2qsTl2Z/qxK+GMMqCcaG5rzdZlWJiXa72A856sXC4nLfCrFzl
47JYlMcVSGWPyX9U+LPxxCG2nsKx9SuKAlesAtEGY+mtfxC1/I2HnaYE03dtOdNAwFBvDi4N9toL
sqrPDYiyv2IG8XyCyDVVUaV6NADL3Qcz3WRzq+6iSxv5fWjD/d6bMppw+ykuyKWewGHWHJ1vAgXD
vexG87Q7FB4exEar65m32yelpboVLKctp/pDuM+3zMk6XQLnDQ4veQTNWb1x3zLjDpnueyPaf6gw
IdbuhupC0aljia1j/I3l09GN5qG5usAzYCJ6QNMsAND3JpqR8De1bMhXzsVAhS+IstJfSTuhLVbx
mlJ4GsHFWGnjyvM8LcssMheZsYnYaMhg+FB6UUS9VA9/4BlSyLnQ7qQxVKxm9StQWFEr3uZ2Fq0d
ItIP7fSAJUQPoH8NOWC2TdKbwQkpSaRzr7Uk7m1NuNDzeyNT1fsmgiAuFa8cEj6CtPyySX2Qftf0
QxifNDK43kZ6fl3wBXQcVhDuRuPVwOONf0tWwbYJpd4IOUBMuoIdGPibseP3LDZmVVCGpMLSQOxm
3OicFjdEgr8MqATvZk4KSHzrVq/qJ++NwI+PIhLC4R2DGX6ucyASnKKnc5HZa13dgQHCc5Omv/0l
xw4mTjMhz/WbI8tu5mN01WF/8MZOMc/Vc8TV3LgVDflx1RAvZcG8+TvcvIdblJ7Rt56apDk6Ito8
1W1mdoA4ZGu/J2imIttEdZosI5e4PWjts48mGejX5Kg8rGb35T7MMgTtq6zSmr45jYsBXazcyVAX
W7TGT6yKr+eQn3BXVMpYvFx51RmKYXLYha8JSswOSPF+0o+y/Sv8LovdfQscTnPsYatc5c6E9BxA
BkpyvacMezjlYzoCeepl5QOnUfRklewhNG0FmVSS8IbC9cjPVFjGekqtlxAI1TzmcLqiFj6jPpDL
LZS86ttH5/NKOyPVUQJMN2ZmAZSpLxp363INyrZlL47Gtuum3f5d6alypD+deZwvPIy5J2VnTgpX
DWiA4EzmNV2sYMRHz77QWKv+Qh1Gv2dxw7PxuijlwjfMre/inr6ANEO80GdJVqFZGtbJWXv08jn7
JqP9emPfpMx2KaN63W+9driOTq8NzRLrqcd7YmJgKjLfH7XiI1D+gBeoR+U+qhPPHmIYPBigr4Ti
2IlBMY2kjX0NN2N0hicm3XwiD+vWJRKq7Afu6oD6HEQ1xQwlPaa4eO9aXXL0Bl7mIymGY9K9E8FN
b7XD6QExqiTRjkw1GjcIYBROmlitz0mY+uskHIua/4nMN7qeRrPVNuffY4QB3iw2Rvvag+6bwQ/H
xNmEsvyZf/fMrkb7XG0ZtWwmQWaHE0tESeLiLJSay6GaoOuH0h5wAbctkUzTMcLck1UEUNIXLaPr
orGyuR8xAXJH9rBq8MkRXRnbqpJ993sGPsd7VSB9Icvx3eimmTcEM0pJiHn4ZiOiS2sP/JTRgCGo
TtncCccIms8kJlxKRHaN5s5Hu03DD/LzAHfjlMKGHRmSYTmhTdTdxeChB9qotNHO6SskfaJFysLP
2PLLWJcY8O2mOGpE0L+SjSWAsDUJ21vVSCve7zKPnU9LPoSLNy3Ou6fTjJraB0eFyxrdHgAa88TR
JV3DIvq/krSZoebOvi//lHGZG43I3G+itiFSPO3FjFSc2LHtF0fsHG0FWVjF0pFpzMPqbZw1TYYn
SzytNyRn2Mqsva1z/Q9IhrcfNYftzzu2pbHzHEReEYH75PLszDrvV5K0MH5G91shuhUhH0q/Vupf
zTLPml/b0moN8WQAwnQAiLUH7e0tq74u3YVxM5IeHEwLY3PHroW/YWnyWmy6u8ffezJs3CiVfSw7
yCmmyZs7hWXDnJitAgJbNi/ruDzVmYp1A6eGizKyxop41zjE+vUe6X2dei5Foe8/zeWmj+1rRnX8
pEDhENkjDFYFivk7faSPRAgfpJD8+bZcDGaDf+vJ2tprpeNPdq0uPIQixGL8gGKgsfX+NCdyGywm
OmLuzLqo/Ostn9LJBJ/dpkle7O/csuAt7B0XEMEicHUmDHF3jl7X6Chj6d7pQ5PFEFUmnj8MOJND
GsxlNo1kWDXO8Whnj5gi1v3Xgw3Zt7tNaZ1hzsi3lUyaGOSSKJ//n/VS332ETl/SvO9xcLhlhVYB
KfIixWLFxuNk4XRdukLSmwhzN8mw3Lz+zEEB6TPxky+Ak3qxOCUWzfp9vu8JeXBaGD4374MsVl9w
EePn0wKZg//azC1aCVMAEoDZOqTXWW7prS83ElJGN2PLPoxYPphERHt1hFEv1yKCf94qycXMOjoF
AlTYkWMmMkZtMUznDwdNNo/AWmUpdXWwUyySJfTuERmKCkCbINsR3uNSLWwK0eBNOlobtsyBabkG
JMEXNKHdKfbDoezlwdJeHC2db6GpQKnf61mQ0sPT+HxG9EiP3z336Sj7cLAIj4vdgCqyYadz856g
RaNVd6JNPC7VLpwx4Kl2oKsxL8wM7FdadOgXFoUowMN3ui9evfD6Y42K37wv7DSXoeHxsuHDzcGm
iRn/aKWrBMZsnj2kVz8a8RuuofN7Zuq4Ci6s9hP2Su1bcOu7ephw5cmzQfZuQ75iDgQXx2wMPHCd
477r/R+aJRqZSPVCqsSnHcysQVk19pJwlxg3VXCIwuhOmPpJFKigeqcDU4/zs0fnZxAWHOssal7y
uzNCVHE6Jyt8d+qhh38S9BB+rlxGrc1o4MK4KxgT/FPGE+64OuuyzbgdpK+l5+uUDNtxiZYbDaGT
RjDHm5rR7rYfSjB7nqIKAybbFUWlrRCL3zpgiCzaWqUs2+tx2NpcKNf2yjpbSjsd+PFZi2L75zDK
0LI0pqLjRX0AkiMwRVFBMdclMdz+h8ah7ZJTlnzY7O29KU37p95Q/Rplz4KJEFh9hL1j7ztJELQQ
u+eTBSK95syRYCAXdVAcRPKk7EIK2Xe+FijZq5S2jIH5gevLJxUWODGMHjD+KaJNpr+Sdx4w3dFy
4wiLgpLTHGgg5NS+9t0pWzG07nZ2VqUV4yxvO7JocM0UqZX+waJxp6pt+1LOvPJ73TF2Udi/XR8t
7yco/XN2XDADiH0Nl0xO+4UNCk1E2ZZDHjr95DzvvjVtFYK2iJImcFvqFM1gudyX5OOC3DQQ/7g4
bmFC/36eqL7lZTLdoqpcHl6k+sJSEuMRRIvAXYJm4Rt70qhMTRY5yebMjzXvXdwtV5r5HQVqmbcf
UNLJ7ftsz0t2+7rLJBmtChXXilHIwdlMzi7bB/2xXZlwrJZk9eh3AQNMqXMXaLQpxeDsbD02h2Rq
ayA+HNJoQWTJsmS+gA/mQBP2Puql8asji+4w7f7Su0o4di3zN/woigKPhG0tzJhkRwnoGFZPNMLO
ocSHDqXe1pQBEStvQi/HvI6+KKgilmXLC8PBCkd2DQl2u/SmQtOO0lJMZoHAmSY6uOG4Che70P2S
dyN39+3yRx5xjwV+mVwn7SAv1ZVdEVy0s3A93MEopN65KXR/Sc1VhTUSjiRK5oujtzX5s5fexmWv
a2XzM5h5U7sav+ts8QuJbLm3eY0N9tfU7ykM8XsJPlpo96A2YE+vrDU8fnFD9bkMYh4qkkuKm+8/
7pQoUdp29nK1eMCGuQDM3dqq9ImlkjqPH3SkJPrmmdRh+yvfcRe5i940POE7LAnnePvseNtZqXpo
ZRwbMnDI3yAuc1J+421mDSapy7sSL7nkyZb+tVKVvJTUEHQabNp3CK9uqwwTJSocggVmUKylmQBn
DPL6qSPAU5uBZQjPLUp0EKKRn9Tek84jhgoy+2+NDzSCpOF2aWHGVYUL458Zj8pt8h49s7ujebKH
sJjHk/uQvcyKynQYAsaqIWhKiCYUB615TyjQpzQtVI8IhL2WbeiRRdULviNS1q/dyeVirUfgeDQL
s6Kt9BsMnXDj4VnWofi/ABZBdSRQW/GirnJkYt9WcqzKtb4rDQlYNKEFOdryywRqXd5KfmpbUiHm
XqZoleZrhSLG5mMJR1kB2WXuKu9WR7kS1WXB+b8w//uqnB47SuDCjhtpv9V9WCJEnkHzGp3czoga
esVC95l+wuOssjo/mxCNHVxFuriNtHd9io1LtkNvVl7z3Ukp/3LpHIILob93rk1qGEN03tF9Hime
Byeu0hTWL6luhugU87mIBZxC6h7uCt8XjhiW/aDY9wJW/KFFf84fVYYpbPHZD9kttX6JXHroGRwx
JmhtsO7GNCopFVlurtODMClWqwoCrQXZhvyzo8IB5mo0Ymz8wLM0VcSFWCgIEOHSABJ8bIeKHF0W
z5nppP3p0OacVw+O13WDosmyVxYgX44QzF8lkyJzAmtb0eMIaSzMuYOxtCrRzFZHUpZ/hGNWuOUw
beLJ5fhlnu3OSt5If4ABWUYMS5lhK+c2Edm8S6+MZWmTi3QcXRGGTRgoq47PktoszMyuftbwDikT
hXT4ntN80y73JjsNFyrfc+jRo+JH9NKrFZbyzTfODGZq+IIwoy+Ocn8okvlLoColjkoufd86lU6w
SO8dto6UdkTMvmKs8vNxz/duFBobPyY1HxOKNzrD3JJm3YGh6+h2jPvrBxs2ksjuU0TB2vUD70m6
EaF4mkkfcKuCnIDlX4AnrPgfNMnanoIR3iXnZhB6oWnJvRnly3sFHDoQCEN7q+Y1AK4UWFnKSUcY
btwc327zwhp16xHtJGrRQLsm+okyFmDcvbPDAsFm+JMcD/AIHTle9qgIfMEHQoSaMJKAHBP8riVJ
2zjzAjEYEPzR2J6F5eT8pFuL2Fc+2WEv8WIZhvPuKrocgsG9+nh03/7clgHPN5nB8FImv6g9juaW
23yFtcammZneB1Cm6A5euOpulAaDFICJbntKDTqIM7ZtjxlJFVOu1t+AhVsa7cEbWDA84WGrcvA9
UpJ8Tho6gspQb5Vnygu6r0sdbo9Hn9US693R+BO7Ffi4vXVZh2LUrdBMuIi+w1Ty1tFiETgT9kCe
tk+YjIbjkrhONxN4PjlQxakptbalf79iXi+ztsT0xoI2uNKbm9O374IQx8as63ijjR1c1HFhtEzG
aduTgbpjUWZh8C+Bwo5/b+NlvGVJ+TxuEvH6J2rE77P/B/BrSuhMyD8v2M/Ujji7m4KB/Ahdlz/b
PHMxTIcQ1vAj68GxkJ7Dyv0zHc3ZotK8O4Ixj/KaqTeYDJ0A9yF9eyIJi+Xz359picTaBC2SHjzv
Cxi8QAQJsiOsqZTf2OMQB7sw/P4QUSzI/SGmqsnWopWtXnh4Kv46whRrSQ3LY1rKxfiuDEociUgu
CzsH315pznAPl431E1h7/DYzpEtj3s8JwxpUW12DvgeGhY25aU3oe9c2oRVAKJ9iJ4IFOZ8A5k2O
C0byuwnWsAOUGQ8c+A/SKxagZLfajlFY1O0+U5NyTtFzRbnuFkjcZBxa2m+Tv3XhrapA78/4FQZM
u0NogDztbN52RgzgzZMilfroVFXcPlKNG7x2QKACs8U52UdhWrTrK6cKF7lHpYQGvpWMhloKjVGA
JAQig5Ml+GV1FgZZl8PADKJV1kkFt3+ctpGzutcPX0+koLXiS2opsPLNsER6aKKFfsxZxiHCEag2
K3fY8df0HLH3ISNX9M5o4PAT+28oZ3PWK7O2tjYgkHNQ7UfzIJfb86/lVPcmuvIPZdgjdBM7xeEt
zrca5heHiHTYnIrhoZqSofPkaiNAIxCs0VL3vn+t39YQYejd0qiihwOTMilOG4jmLvSMWHPXrQNY
KT9OrerU+IOLmiPFcyQ4PudSix0ECQLhsjXrZQgzSLyxVsMrmAR6AhKCwfDFwr8rPdQRnBgL+Fnx
csFms7JMiNubYn8HUJlbiEv1svyoCAOJhgbfnY/zQhgkpZ6dTOnKV0Np/AZDLVMR3PxuB7BVoZPl
G+tiv6XZ+ZlkpMhDQxqKSm4ydGoxU7hh6tjDHMtzchi73kFoMCH7zqU+MMPCyMpx+UbsIrkq74GK
xoCzl7uroOEDVt6N2aEfrWrlmMT304Xr10lILh9/uIuR15nIOb/o/EETbskAP+okADCiymZmHn+D
73hq+OVdtUF/Y+9CLgvRbixDxnb37r/fGb401t23jvE6bfYoyg7Tpn+4XoWXJZC7jAOZ9Jmv2o/A
ZKQVW0TZaUSKwT1ojWpFiRpj1WJ8cQs+sFqdRsnIGIlpj9Vc70bbPclm3zf3vj0D9IkuVVuPSXS3
NNcDj1RErbZkYnIK8EYPbULDL/tefU1jL1HPQ2ef167MU1mgxPvy4vpqXaD/DVs6DwN9//SbWL/F
G0Gmps0BjRWjRCAz6j9lVhTtUCamxV7ht0YgO6ZWgQQQsAsAcvg7HcbRlPmpoYaUzg+1kSHIqsXq
DOn4sZatDs+JxmjXz1kJ82f/rS09IsI04kzq3SKgsLxrprkPBUp4OOi2t2kaG5yBb7aZkBrD3yP0
oGgzz51+8npsipT5RXykIvI8FrbOI8Og+69aMHqAI4GbvZ2SMYgItKoWsmru4ewRYw+8U7QU5a7Z
YY5J6o9EodAz4HIySd+FskaS2IQZhyRJVmli2YnqvpNqPcrF0hJBW+20NvlL7HjjFsKle6cH+DNc
ME5jLIxRXEpwtvGzcJjL3AVyNHi4IdYPhppZw5Tasx0dWO6matWo4jKKzGeudtryu+X2tZhpVXVJ
Gq7LZnoyGzwISNylACnGKpHeATkYmP9cNPs2kMn1FcIeIHOCggiL2XcR8bSLj7RTJQARdJqUW16Q
6LDwYw8L0MvTbxrbI9H+AZTtVZZqFGkvUn5QR/NFFlFJYfJ/gke+ZR3+1BzZqYwQmlR2f7O5G+H9
bYnXP4YZmTzPwSx4rO6rQLDupy/Mm5uX+AFY4TZKDx/tW2pTsTL60iytiUtmgZOfePIe8/sVMywF
uUjoY4n4Cvj+TS03CStKexEon5+uZranKZ4Q9sH5+AsMxs+t8oLsTHa6rqDtPTJIKr+NoqzHb1kx
AMBbHYKJ/skvxOutgvuj7AllKyP1h8rNNE8397TkE9PwCaIhMgwHkkJkYWclNSmxaEp4WM/3G7XL
S+lh1RujvQfdBjTHPGqINDoPr395RlnNW+682HWnatQzkHXmHO/mWAx6qHN5XVR/B+eCD3HZ0wrK
CaDfC4DNAoM5cduZw9Ppv6HqoRRKoUXpLHxCDuQ5BlRcDwfOeABRGDJVl/xeYp89Uv+fouRIjz9p
w+/y05Sy3N6aTkUkOcroMOxKnCUJnMQ6H5QKIFxW0HD35fLt/zxVVJ0zypvJ43rG+amzaYTDJXPi
bkb1RmQhbF+RMqH6tx4342LScOPki0ei6LWz0+l6aGE7wDENbo4XN0sXWMPpv7UcmAPZIaF3Wuns
evuW6gk1cIId+zPJIZH1Qu1kHe5t6fGZf/yzNLRcDcNb4j4aXr4LNKk+Blz8cOa1IwsUE8D7KCnJ
pAkoV6nUiJg7I57VzyVH9nflHihQYXLtCu9xPa+9pyPjadUT2W0sQYAZrY6QjsPRyPsjmMQDvVlO
xlpqnKZE8dvKq3uNl/Og6LSrQOJCOMYzWquRizmpQpbQdb7859yP+L/ZUz6KPDIEKDIvjGypPDET
Oy9HmRIgtWNELHP6k9kA3U5squzvvC85ANy/8yowAiW+y5N5C0H8UP5+UMsNG0o23BT77lDUBaMg
K1zn2AMrJRSe30CqO3UHh+ERBoagtYDwMLkQwDBQpmIE879+o29aleylnqUTIcezgtrtzhOUBO8L
SB+CzVKA1oMbfHd5UnFYBrHsc6gbuxRSE4jNwHJrQVFvhz/7c0fkHlcR9G+IlWcWcrCZy8uwFw9r
go0U3hm1M04YmricO5ZIuLq9YWcveN+mIHzN1hLn9AMKUdGr+jhWMjaZ2PYCxYprDB4axP8lboNK
8CaIZU0mtW47sMs9s5seMweJVqLNpoo2Fepfjwf3oQxUMgloQ/BjLULGn04lrcEBPD2Q6E8EYMJQ
W+N3MKfP6A0eTyOiFAeE3PDPr346hPkvhXWLobLzEgjkfJhn9CL0R71fXAQ5SxfYi/IBwDJpZEFL
AhRLQLjBtSVpca9c2KVCj0LCFYMemNg9yZpcWtKDCQQp4zCMY+f1v18vFD9s6ZRlivXyDrpxP1m9
8EcRFy/QClZYtljNSsDwTar0ueqJ7OnOxZvHvcsqukJia0Mpd+0N3iRtlFxqQOO3pln7hhk+vdNX
dR92xjyJh4wNUAUolzTJ5U7p17Zi/bQto0TbJuTbIvu1KSLw6zB+ZhuKRTrmOwuPiGdA15drrTp5
jwHwpT50ybI31ZIcaFjXTFIlvXujDS6Rs7z5NjS4xgL6UTLz81jdJHw7G+F70vYp6U8twVMyBT+T
xTd9XMkMs/W1quuY5J0sN0dNk/+H7qeiu6B+PAUkhaIx9402SbisVVqgRNFVKqsUHh04t8z/aLNX
e2vglGS4H9rHg4PpI2WTV0CuGwJN9cXaNIfZpOUesHdCWhBHX17B3RTazBRPt3pkCoc4KgLIwuGN
kO/yOJ2zq9nWLy7/3lRiZfxBYbfds0U+Gp4kxrvbdzoRm3e5UO0q/poReDaVCtAFgzaCi5QUsasB
dGwNT8G4C9T2FkOWf4Eh58SoSt0FINHIbFnVY0VmYlOZRlwW/gNUXbUaIct0E5oZhqMXJo7BB2WH
RMqfTTpSiyq3+GK/qTUmdMPa0p7lrYul/GT9dqCZC6Wa4UrcFpsOtlX9LrI5hehVjeOf932HPVtm
lNURvq267/3bg1BOB32D42OgE8WFCStjMdy8j3i8cRiaX14WE3+canFo9WI6xdOFTr75WIdgY7IK
KocUY3SPb/LEKrQUjKX5Yo5f3+eduvLG8n1mSj4ew4MCC4uJ9PPKbQdaxEPwIf6AxeOCvHdq/6eN
3xYXpMVVpbK1r4vkpUAmmNowCO4TEV+3HGZ1uLb7invPszU6ny7niwVjwXHs/7lb9iAf/i2uCF97
q3plhJ06jJ7REoADjOB30i9WocXQy9jqMAllJlJT5EfoHfT48fMYz8ffRFaY4/AGKLbgAZ1wv+pq
MANEdXyJ9Otn7VP61QShjltA2uz8Jtxc5Z+/oRQBcBjfTm1U+CdyVWiEii/RDDjLW6c0R+9DSb4L
xyiBnfhdf+aWk75HwrbLPYy0keYIWpNigp9eoOH45CAfTgmwPkmyoaiOAUj++eg0J/Cm238xoMKq
SMcoFgPaYV9hBchP5PscN4lrNkncT/PTQSRcniXfcOOSKN897TLw2UZkrjvjUSvjaZHELOPdyVHl
Hk1RzpBlYBhWLj7qUrHigINjBlq/zXI26EIdpgml5COEFkEadty5Icr0g/PqB6ID6+foGefG6BUK
epK6YrVKVk1GCkSddUInJBn9BHJLB5LZVDeAoZP4r65TH2tCNpORzqcShIByTa3XykerTn9p6coq
11L8phBbAYV9tFcvPDpiecT+17UCz+kkJinCCt5L+C6w4Qigl2x4J2kKC57q8dyJAxCMWgYOKtq4
DokBWVtQrMwr7b2eCpaUnLyHKdwATYBRWRx4JteJLrEpHJdpQ23fSxIgiadDtVT5qeOdEVpbJv96
z01NFJ0FI0XMCM6Q2MY7lP9+/7vo+51WfvdGdLDWClWypHvfXe7o90Czj7CZSlety4zI9t+IvE9j
Vm5jakMbZTFYaty05RtZQC0VG6J0WXHvRHsYYDBTdbLNsBxRirqHy5TTY8u8VEfbgXl/2XYBhvvt
gqmQWIA9TtlUGw7AhodruT/4VQ3IIXmyFUjnOen4LTPEF5UBxtGybh+MVtP2F9KG+qD/kgtQp3oK
XDMMGbBnqHWEQsU81yZOqNPnG9LMJkAMDHEM6GNIHIZ9ByBNCd/pYKsBeoQ/UqJUx+VIvebSw3f1
UWhoeTcnbLxbLUMK5sRbTvDXGLRVDl+LoS/jQI+rSEn57tIK+voxi0fKTtOfBLMd3iIClfhBaTYS
pRdc3pM6K2wFJ8uKCsEqoChqjS5DUxhzU2TcWFFM2K9zIKMv4YDBRCdxSFREny5QBsgBqS/OiCLQ
VTwz4rxM2aQglNPGNLYA5YUlGpsnDYPATNO7G2tr5XGLlsylWEgfvAMBZ/l1
`protect end_protected
