-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Zl1qFRYOabNBEQ1OUERjiXut+825XFN/4sA6+v4M7b+ZVUVaktGFXcZD1kvetRdE/mwgbN3PIJHd
ibbOh/vv+k/uSiPx0jtjv6vQxTjIld6+L0R5dn/9h8/gmW4hq0COdT1xvQOOYg4HoqxYv2rcx8N+
2y5wfA2FpSkMv+qyOjLROh50y/4ftYngPbbNw8bcvjJifOTmenWGoY1Rku5Ou5g2uzsXJIRMOtPT
yykBqPZUb67rl53S/FkqBtvBcAXDIOmhitRyfPEsTVquVCZZTJHkwjdG8Jv1Yn9RaTFAy3MR7YEu
ggIFWwDlgPKfffq9TO93AQ/gw8e4uAE5iCqbpw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
n8EreKtPtt857JzROv+/J4ifxrrlfbd1Vuk1Ta3Lf1EozXRo5xPWM+GGRlgLSrSe58IcUxyIWSLV
iq9XNjTZh6oJ40lnQiCHGETNhqqu6xf8cPFwukrpfAcscm0z/dxKJs+6l3rXsUnD6BJ4mWJ+7fCx
iAyIEFIG4sC4uKVhjgrxkQNZBViIiUiI7L9i4MqDNQPry7WXoC9C1LI7qieWDw3wkf3yPVYGHB33
Ptg2FuT9iq0inUntagIKeLP3jhINdXkD2TIwv4t2Ysqc7aYB/1mh2BzJD0zBs09p+5HGF+zU2m5D
s7EeNAHbKIvvwxfMRJzUWob0+3a6ruOhrm48yag1iYHDIoAQ8+mzOMEluJ62Tp/jcMJIYTCCiXbc
Ad1j8Riqrel3cJIh3RkCoCuphJe9mLKUYWsaXR56EP50BxIoU9y3DLSZ4xGE5hdBFN3CmbpEVil/
I9UYQTxT6yCOFlfS+TAIYLc9oTs/juxUspr/f6M5UXq3gqqUEYaTtTnJSZnt6m03ctUUavUQgyd+
2nInUv5UmVWQ+WAT5d69wCHrwPrCzNoktsddENB+zub6REJg2ysbdpQ4Ibbm6F2oW2HHBifQWQPk
w8XVsNHNvUr45pXOYZcTbf/9KcsG65S2CN6NNnFChyXo4BoRCjDtpVabznIRWmdk0luOOK0BFauc
Q8rWXXFAaWjLXITPS1doFOtapiz59eu7SaQ9wZy18JBzdto8ieaA9tXVi9gwHs8eZXK2hmfmdJBD
/3xaxnyQsOE8yu0T6QxciUlt42bPiTtqggX/3qk7QnR/XTbF7M+u0bw0FKXgqIlHyvOd+kT7QsqU
pDaIdco9ikUJyrT/tqeEeVvoZO3bFRsPa5zKNzrp4UJinzxa6AhuCpNgfKqk8cpYLZXcbGtqNIGD
MVK/r4fN/ja/oAoQBuU+KYPP6quZxgRJpkSkECyn2igUfnFzAmcF0rmaTy4entfo6CZM/N2g8j2p
YJXFu1FUCn9OnHRITHc4QKqroPTDHwBDb27J9KP9ALWx5Gk5mtURGeVzL60yfMsAy34Prav5KB3/
8zrv5S/DOr41GmwOUJk14Dl9iF1ZOCnK51pI7B/9EykOxOM+cGt7QWNb8JITbSmr4HSgh4XC9rmo
2Fk5H8H4JwyXYrZxWX3yRB3NiKqBrwK16h0QAta0bzGWozx+jrAg7jelt6rXFWmvfRAaJ10m1O0N
PnOvMGaM2WpdjrCcnbOje79iAHR0SNbrVGlDnENk0FmrjtbGAlxMnH8zXGsBop9ZK3N94k0icci7
eewn3JyJMUp39pwoqzILkDhoazfNpU3X3rRTeDB5niGrxTfXEZuzNeisdqBOz8Bd8drqjk/WElDC
Pj508+tCjfkUVhb52wxCAM1h4T01cDHjoSwJpbAnkXLMSRS2V7N9HBfruz6tLWMyOpSg525hI+H2
6LRSb/J/otdaJa6lCIUmCm90wLRhHNCVBD2c78xBCZJVVoTodPLsLja//p7z/fX7UdBMIoFQyCOP
bP/aNxdDiaVm8z8MKqKy+o8GHpeaGVAHD6BUT9xcy7iv8w4kkrI0bk9rfuiDEBv0gvsJwItD/kjL
UR+n48GHCMZsfTnduqoyESRstF78YEAoWgVe2PnHw6rs2kjqkFzag8EHq3hVWd25jYbERfw8ZZ7N
xWLIM2P+29rKtFfqEcyjXtN/oB9BtWyxYJ7Ebi1JYjXDvYkemYkKYKylsbAqfqwtSVoaWrrc9t9I
xmmluNfI2s4tG10N70iiv+K6CYmTvIXfVJHTHtmlnYLGXP+e3x7SI2PgqT3xDTIl8jA2AyURXJKa
8oob9C8kQ0HKWV073/vFmZdh3/QVmrP4ntGwTRFh8GnUG3ft1h7IINZ0Ll8N+5T0u6z1JfHkMiNv
gXqmIYJ02KePLw5d7EIIs3rv23UZ3p90VY9I2aMTpj39jAbcWXSzscbsOzj4sPtP/ONBBu4t/mRD
2tDv8ZuovsAXdUBqdCU9SCZqZ2+BKEFalFq86E9HltHYTLTLWWmdOSSFa8jbOHIRshfTNOF4jCgo
ypYNmHr1eAtOSIxigFRyy92A6C9vJ0DTfqe8bHqlgT7AMw2oAsAQ9qn9LuZQ93RFLbcFDUxQPXLq
p2qIIcje6+HT4F1A0UC4q1my0kADCpCe15gJloslHCLxhJ18lYEZgNWiFva5qv8n3+lJyvSvMBLS
aaI/mZMTzwUIYC9uvrkV5dLOBLjDvs2mTp2mm/cFT/71vd3TJL1og4HnIQqQi13VhMhRuOEsqTPn
btRiFZ1HPjf+w3mgXJS8qsKL39DqEuyJqIYVuB8Kg97dBB945jtEZO0g2LZLBi94CGJ3795cQo0I
cltFLFbZOCCL65B1FkKfLSCnpml54DM36CLH8z9GBhlN6Fgz0u4DxGdXGw6AUNG1n4qOSe3OZSJv
mNRW6qLqDr4jn0I9m635b7oJom5MGQ7BbdmMHFXZYGNOCln/AEzywIp+3vw7FP/nRpmM6wCBeSbY
TbHVbQVp3/Ey8u8ivCUQLfZn/AQnO0LKctQioSvh5gFBBaJfYLvrWcwNa0waMuIz6gReQuhj4JgY
je6YmtT6tSPI0FYgt3ePLKd1ICjn0YAJfaJGCfvTnHOaQm4x7OMx93GZVNcWZR0iEz9maihDU/fp
esJ8V8mGZVYmENiDHhuITjQ/TpiXGEWJQkMLopztnCTMFIq77cDpEE4i4CS5dQwxc8brr6IWX/Yj
5D68d2BTasCq3TKFNCfQU/e2KSeE1e/J5n1C52Xywb+TEsHWJ3zClioNUspFK/yFQf55DjtvqM3u
XPRM0aMtfvc/TpuFw+l8VE1p4LFm6ROFI/VywLstyeXMpp756dMVkqOkKASpJ2nooEQW0rmqk7ng
LoHUnc9vVEOgmpp/ZG3SZew5uy5flWOjjSegY7MzZY3fiDGF8xwGovKEEJ0aPf85erQXnHeLyav7
j05FM6T/4pVsR462JLMZfVg3L/tI/+0ahY2K0AUeiFUVJwKnS7lJEod6O11CLrz2ljTpSvHg7NEX
0i8QPFTUwRssXNZyl5fq5IrX90kA4NoVhDPt7xwTq4qH99jZRxHZ3dImnlQpma6wkQt0OcwWjQ9Y
afdnUitnOAc92NP0CMJgnI6jI3bpSnbV5trzb3l1ZnWlrfwYC0yPEoIU7CzZkYtaU7qz1LG8Li1r
2LbciylBu6HymPMMvsJay9Rf1l7UxxbqmhJhOu9sos0UaIhY9AH1RUk3zSXbvss2yOMxa8+srTJj
UIEEAWp+1oHFoGd2Nq4aav0zAfcdLNI21JEedjuVvs9PqgBs80riws07SG8Hm5mx9abgFOOKEPto
l5Dwi7mIAJFHjbJFpt47nPP6X2azdQmrJ82g5H4e4YdKU1r7/iGGCNQX+2Rik9trbdMo8xh3jYiV
RWo6QDsCyXxvqbNFP71njfdlzy4q799HU1Xpm65juFnb9fv1vBEw7yzSAygse2YOLxXBRMWDa3hK
3UGs+Dm/Ax3fm9lKi9XISOuRfTABjKhGnP5+K4ynWsTJWxDVSLlmsk/hZN/a/7bLkklZe9Oxd+N2
W7Z+TQwwS+CCykUixKStD8rNRAvAKdXJzieejV5e9UhqnKRtqo7emNZTVx8xv3WOplDmEFgDIFxh
Baw7DI/f4DLngIx0veH/IeLdt2FuRllGMHaHbKOvhCetXkhvnB3MKfVIWvFOfxbc2aaSxGweZaBE
VHoibpJFi8hGD9nJyRbwD/dLsxP8PGF8PrsvYWRxvYJjVZS5UrQQO3KOYuKzXsuELXFcoc3RsIgV
euIVt1bzupYkyzMbiVteih22g1mnB9ZH85aFhE8d75e/c5WQx8dmGRNX+tID9ia0BNoO64jhq+1N
cBvKgOpFIvKW10NPbXvDTbFIOUVGDVmBKIFsi/ipD4Eb38E5peCRCDl+G181j4R+x3Azj0BPz7Y9
bFh9IpmqT+OwSXu7aYyUMKv6DcBoFX4f0reIzPWQwDjL8zVwCvofyHq+1aPmW6fScIvL28c+PnKl
wb8stFC21jUful6bzUCbaSeUApnja2sjhv/0kcdyKqDMRvnZiybIUykQSV5S2W1knoX+v1R7MEgP
VZKveU2aXsEwCUT6bfDm6/Ciqr1URcRKmepwieZ5Kpfkk+0GZnU/+R6Dx8yalb95G4CQGo5Gq5X7
WhI9i8jLNi6WvzRBYts85TPgLWPEn2EefF5rDe5IEopIGewR08D4+XdqKe2JY3V3OrcsL8sv+tpD
EaFKJiEJ4WeI0c9/1kzi5P5BhRdEahuYtLLQKStgrh1BpjvAl0qlaVSMUo2SLFKxOfg17wQnYbsL
loDbqCBCYghanGX7mFolP3dXMMwv0iBg+TsCrrLFayc2/1afz2k1prFxvIF6lbC+VnXaCXFiTMoY
+wSSDy6/E3J5WscwTqnfUNBpK9dUhgdniypF4rCp4DMydo8fepqtBcixnWjKByhqTOk4O/brRAb2
lDPC3p4NVXV8CgDoZ3JMLaIxTgY+7AVJ477TK/GFpptFwr4XQO9+L0p01HDu80ad2nt4pHpGDvh7
qHlCT1oy6YC0w2CTroNzM7Y8v8SNq4UYczVh7VFzSvoCVMoOGMfQ4Yp5QmiwnHiwA5jxw+2ei6og
Cu7l3dAiMjhTw25oA6AuhqzSufKyqxdojjBhCdeUIgMNevuBqk/IvYPicQKUvn+lYx88mFfo10If
D5QZCjcGuU+I9KtjQOPFKyud0jwIemVcpe01nO/qJvNIKukrw5/NjObuhyD82mFCFsXJeo2pjgGv
bmmUpcThbMbtTaS4qzmxrvp5TDtFrzUJNAg8EuBM91XEBfaFmH/u16a/6MWc+xxkkWofhUIpPp1L
2byTUlPp2o0xWxxu7bI1cVLQYMCVtjvPQh+gvqFnNFVkIKzgtKrgvYCBHZ5JzQmgnGWx9wUeSlWB
KToii+cBHfDSaOfY664ktupN7JeklL6ycoGtym/q7p3c66Gz8t/oBZGlB3Xbu+061BYj/fm/iubR
ITyVNH5tvQFFr3mImszvx8vbRqJ9B/u+IaKNwQNZKuQ60lg1KCeX8Khc0YzmyLw2SmKQmKAO3kpX
vn9Fq0ID6oQC0GJI+aqI/j9mVR3kITAI2w2mwSpYB0xjBYXqK8kAmerGycguVP3G3L9eOYUzHTb/
TctTlU8S8DFsBbbMq3S2UPqWWja3z2zu4l4VvCcGbSgGbcBpwWgZOesDcKG1ro4XKOODBsG2XqJJ
5Ul2BPcSFKxmCec7lKJANAj52U9zYaIhvRGoFijDVuQghSbJQodvk5iCzjlar/lmEL5HNBx/Sq00
EsBgO/3LQjM+DLndDwEU6pUazORXOlVuhkR1ix5RlleR4ohIPImApBvUSgUxzMjoFaIjC0kVRRP0
p9XdaSWgZq7IvXnButnkESXzQjR+dOTUBEjBleAHOpfElrZqguViTmAYeFZTk22rM4MEsNRUSqqf
+3h6pfI3zqiDwE/FRmRvT/op5pWjwncYwFtf8+miMPwlCw+AaHV69jd7O/ub7S4cJ50mOf8kqrOY
Qqpj020GZkn8sHFImWXQFtgpE6gg3XFOYkb7y2QUCs23Nn89p8fkD//K/SGcQd1yatZH1vsorzyT
uTXTZzj7vZd/40VBi07+lv045UFNDU2FpI/etEv/qmg1xO9U/mWnrt+V01X3qrgX5TXBdsbbkIYF
lKpjGINCqa5VTfgcY199kyIsgFpXYbMvsD8Yt4ubRZNhIMdo5XqqAxUmXKPAjZ7dbpcvW45ulCLz
f7SHKjslM0UR32h8nKiL4PjTcY4Rg3Dum49qzyCbfENWk6wfVIYmaNrVZYaB3KOQ2gTij7G2X6lc
ih0yF0B1nxULdavwpQX3iUf1AR+koLdn/cXvv/0We6O1qRyi+0ABBvsxzzKflUJtVxcjTYRia9YJ
jdDzDz873gGHYq12oUsynQy5JF2uRG78/arTzS9WI4wGQs8fc0zflZ442LIBICC+rgdN6HVB1fH4
hEV8cmU8YXHVDKyeh3NmI0uRgLycui8g//5G5C09SAImWsWZkKZqICCr4/7bV6tvo1+YrF0yCWRK
/lTcE2wuVPdYpIst1Hb4vYlbw5ta9lmMUCDOdnWLgPLZVcMG8Wh6oHtUmRhbLlPz2wUznZd8ztTh
Ira8Y1MnneodCWL8t8z9NEQKm5pQFvosdR8YS0F+wg/9/DapGfurSvGHQKGwonv8Ppopyp1WiygZ
jMATUkHe/HwnkGks0YCt5XYPWJvaKSW4EO3qSwTeb4yOF0ZoZsM61LhQ0A9858iDwK6lx90dMDW8
kTDSHTJtVI2r9NU6ioZ7wyjq1q+SjPsbqheHAUfROjIvKD2qePcn7FzBr+E/G5HQ3+LMM7V+wy+C
WOKJp+BWVsm+Vx3qO9/fPglKGBO/SABFn/ZNmC6/tF/UMfJ9potEdeKHGwSb8imDm5rSqHHTIbX9
dmL0VQxZiEt55IWUXtwE+Ox378psVSI3NH3F5jbLHB723lTTXrtdKiUVfrhHMpCZrQFYg3hCF+h7
hs8YGMY0cZvlJ6QY4EaHE5sxZo9WOvu/TkAeJOw4MAe3lej3w2jUnx2OM/9IvsBFnBKmW9LySgh6
dXFc0WDrXAhmH9eOBYoxIOh1JBJ0LW9iePm887tQIMKv7QzJqnAN6QjrNLDYFrxMQDTamqeES4lj
BjjnfDHeTTU4/mvWTwREVf+ZHabcww1Nen2qfQ7cmBfBFER/S/fnVa1AhVvWVWrEw2SBqgrurvBe
LXAtUJk9RnqWhJeFSIkS4To2zIGPTlBaZ4vintTmSpBP82VnDomXsuNbOOe6yRfKEc6z0Jj4UsAI
g+0gTb+DHu7RRiBFuAt34Gmf3opuOclvygeLWVcAczy48cj5wdbWEU9TDlMt17U/R41v8SN34FrX
LCQUue/flJ9fZ4Ul6flpxzpGhif+y6gxypo530kgXERdwXKQ0nlWrqXW0NavRiGEdXcVji/UHgPl
vi3EePGC5B6xrCV1MpnH6JOGmXieJUgF4tvzP1KagKfr2QnRC752nhkvUcsHYmw4shbKTWpsXGBR
UQe9fNdh40+ygydIgXedgEaekSLGEvWQ0P+vmXf8k7UljIqUG335rXqshlc69M36KVnLiDPQgW1i
9iZ0nhMbMveHFBwlG8VjnnJK4dA9/nDQiXi3AYy940cG+cORnVSPZfTYJUrsOFrq6SondXb3K9S2
J3fXVTSGqD3JMWEFVeqX9EC8OAbxd6gxvmyJ7rib8gtA9uQ08V9qTCYTUfpSRQPODfjCMWIaAG1d
0lu/u8TfwCVwnS4Bikjn6L3329xTmAvcZWR/AVhGosk/OTteVaAUMrGiB4B4zz+USN+1xqOJIa1c
a2Hu2oRG/YeM1FtVkFozUI5xm8XRusY3lhuf2mR07PFn8qSQQhE/BWqg7sz7WzQ4JmTO0wB54x2O
t4ogWF74wtwZEmK4M3s+RPD2X2CVruVyyNqrl8XruBpS8e+DKrvVKBgqAdkOmm1+0EmmMC/VC4Qo
mQwKKJgooOVYEYG2fn7eg5NMI4WnaMTqcke+AcM2Gc3VYG96t/I4c72PsmsbspU/kyYERkCJQM95
t7XjGMbF+EhTDXXYBD2Bp2+iJV5CA4hR0Q/zDdH+beklCrdCi+t+YE5fd3Y0CUwsyzmVuGGVu8HB
bt1s2x/QQB9NE9GYazg6NLPSdIwAo0axQ7jJGPbjV+HNhx/RZXYBU18CTsj53+XXrM2ra6mdZfj3
O2M6Cz4Gylf0g9aLbs5oHhNuBDwpfQFjz4Eh6B06sRdToCT2jEIX6zgnTHYNhKf7llfN5VHl+lQI
4nI363/Ak+l5rW9m1mp3TwFUU3PWDvkeTfBt5XTMbYyhAJXgVnmrIb4AKzvH4ADj3d7vyIEfBjJU
t2ZECU1Ndakek+H+6ZTYj2fEJJmTBVg7qTSsrexhHu47BcPahV6XmtrXAqKYsh0i59SYjEeNZC2v
D50YAlB9q2zxXo3k/9/94F+oa/5uqJqlS1Rl0EyKTrf/j5yy6+eBgn//hC6tjrlkd15qWiRRv4Uy
4Odz+adRe8O9d5jxDgFSOvgukvRhUkxC5gDuTpShJZxIhEIbtNyQsGOnf3zmv2qkmImkFDrEbjcq
4vXso/WY9FX+9GGo80dMqrVI0+GAk13grI8sbXi9qZ/GfPJs7WeDU3Wwp5S3gaoWlIuwQcM11MVf
2WJaVppGX4hjbYroVgYkuA2bxnIkEUPOCwq6x/7yCGwpa5G0ysfeuetbDpLp7WZrAHssPvAuPn4V
SAWaqCPkw5Vn1lSp5hHeIvROMTCnibmAVQXejr8gUUHNMQu/iUhMmpKk/dDwCTBnWvH+AcMJgeul
2cuy7JBaY2h+FqU0qISZLvLZf4pIBylfpDqmk6dsYojGWFkK/FUtxTXZYt7aXHrybK5sSjxGAgLY
BwEljrvrt1lykcbEUOJZnXqWAlNqlJinqJ52RSuLaw9nYnBYF+ZDwPkv9WL3yBO4Omfa5Z6QbV6U
azDrlJMj7SA3yCS8iWmqglok2Dtg8BOHYXPuEDWwJhEn7vPxjkuPjhbWOnXFCnl17YN+lrYeS/46
+FNaYPSsluVus4JyxRg1R6sSP/CTZoa1hzjSOh1lfKpgVEbikxiCwuwdjM8fKW3seKiAxyVnGYRo
KRYDELNxUHX4eXqSTlMdqtn41kDaOHABtSeMKubeg6L3brQGGSOYIDm3eH7OeNTWcaa2GNfAgbJA
l91VEb6QarniYfscLRAw3k/QNA+6aYeseQuZomg820NtnQcgxgnXVditnQwOB4CkEZIeUcLCFvMI
SKvvwg3DDxvYApT8yZqchk8cTJVTeyXGEk3f9OIbXpET+ZNEi8E6xTja5gwtKmGqhDj6Fxr0kBaR
bUraPiNrRlk50SFH0qvTZjeOr3Rtyi2WXqs4odgDCqrYryymcbishHwOArpsroJX0hwLR569eWOG
+EhAfhPGj5W4gePHWACX5uMkK6r1TohrWvenXeS29A019ikkaKBIDx8hd7h6PPR0d7uCT9bBT/M1
dE1QLumKAE7WMb50QmKYEvejhY1A03aAwt2vIv8JWOpAYx91lTbserfawlN37UfIpckFhxMtm5gr
wsNOAaZX5EZ71pGdPSpfDQSdVfhlcC0X+s5LVMrcmDO0/Ihc604wqyW5mnSWKQuXvUYSyl7XLN0q
9ze4KdBx5B8TiPE23v0XPkp4IgAyWLvyq2fUlLaak8hibL6PL29T4c1zEY4RFDI6Yoe/xndwCtTN
WHTKsvOTWDwtz+ET/8ynmrmR0bILB677RU6nt59rycQ64qNwOgB+NESLtLXVc0fFrNB646+0OVZI
mFeW9yVeAmKEhoxOK74oQ3/rtd0r9e1gvMY/RjLFGIFuu4qVmYIoLv2ziEUobiLKG4LdkBzux1ce
G3Y2NW/2bX4SLang4ZuTDaPT+zOLNf3BiNUPM9a80ldjivxR4rbj+O7g4IRYfyBszW6B5JYJeboP
VkQ1jF3CqEGTB2FUfEj7eh1ZS79lm35268StutxDMB7dleuVHKQwpptsbvcfqhwl8+9FI40LjfKx
m4j2S1XN6eWSX0/2yv5nfaKfRg1A8q/BLn71UQu7YJfRXpaLC1j2WPZ4pEhcOUQwDDIFix2B9gDb
bbzgblY0e8LCDLBKetLDrZwK1gMl/CaiHRKfe6h9et/H4RZQvybjpjc65rGZR2sx9MhIvrZUMrML
8509nUAl/0GCc/r/yBu17iHVJuXuX+JL8wAzgFCuM2/dxNnqlE1ck3SKpDAWhVc46CNHL17A1F1E
iqXcjatdx75N0YIKJlToO2UwqRas6mbPa9sWNGIL0DNEb8Il8eGwgSdPT43lFViOKn/4sa/9pk87
GfsXmBskDTOLDNR1fZAPKIQ+379A6m7hachnzitI2Cp1/h7g7NyRX+NgBUaj2Xtju+GmShTUl9oL
Y6jNfv8CkhhC2+D8j7HBqw8UhJCTJhUPAf7f8ZOmPAgLSzF2Tzg9p3mPtBqxoypFwJK1elmavWy6
6JAew1S2bvWZC9xCJhpxWQsZUC/It0UZBAldtdcJ8NJNXmHwdwoAeJz+wVvVbmt+8iRUpP/IXD5X
Kz8lpWFVzVZnmAarFdWBCNZm3daxPFsaMAc/ReIgwDXLej6Bue30GtTQidNb5JecfaUl1a+UIL2f
TuqGu7E9rO6zwBzxBJNI1ZqY1VLffANl+N/tq33s28c7RZxUhheFMLYux1sX4YdV6YfeufieM5bT
DeeMnuB0kGNgUySkaCTDsnvFM12zkldnpvIJgCt16e/Mg2sGga5FshvNC2ElpXB8QTHCwcDyEtEk
byDb6hyuQO/NvTj/7Pvb7mRdosLLqwgyaFqe6+994+Yjkdf5IsAi1XZtjp2yDaX2JvuTHB4CNz0Q
8xlLLbtqcMvPC3UTelNLDf128bcYSFmy4fXES23Q+qWQNalFG6Y2ia2cALLvtlF8iezDNsgP37pJ
dqjC1f3cVJHxM6YLSyYze4tAOvGqKpe0jfPtemcXfHuPaBAVDAzJyBNX5zdpLpI8AEwrv4aGGLoN
34tu1q/a2UXLvmcJGB6KoEgXFcJk6uBVzHxiRbIwmZ04qY3hhMTpWh6MMJEYcXpiDlE/4BgQd2eK
L2HcXgcxzp9m7J0jDzXDQuIP6rh6N7yYU+K/EadMM0tKKSonGcn5yOMICEkpBeRrO6TKQLux9gq1
Fwvy4w/zWNx28W8JQDSGl+ppBVE/cFt3XfJumArzQs6NyuqDkYH6KoxOY34//o55zvEjTX+fN3oa
638UQNEzyfJNIntN4wdt3uCq5/6A5wUchMlYX1YcLQi/oyH3gYTizU81iVZwP10B1EwdbcU58ihR
IzmUQjFR+Spa/obqZLz2a2FYqSUlR1phQ0ArvROBlHZsZ3N9zec4LllMpTNVVIEqVb1jjQt13GUc
DO8o9FN29Kkc6KtefbZzy3Z6+R8a6QXGARAOhRfPZeMDdp5QETsq3JbO2t4fdRYfCqq6vu3A1w5C
2uBuCLszuCU1HjblZ3SiEvwGav8bM39LgCO1JKmLMZg39Z4AeAtt5R+eA3VX4XDhjPERv2mOQw0T
YCbi5o6mfGJc8ouoJC/pjV8jAxsKVUFMMyLHJb+V209hyWwXsEHup634ezo74wigvBbVeFRpK+W4
vpHsyvXE0mpH6YeXFAK4oZ2yLjUrDB0txnwMlE7xtOEAGr4qXUlxP2xAw1rJbzglgLNprvW4KpNM
cTWuEK/7YA0C4irXPN7tulzQNtBELgUs80fuzoOK6WhX+RaPqKK6404z23MhZukE0Ev83mWMZ4jK
Cv+vwJ0fcgOO7WcE463IyM7Vw4dWcUeB4A3eUdex6bH7nMf8K63yuDlCPS4swUWsIIwpoUh5iS+a
0tJTaV43JCjv8i9msQTcwZYxpVhcvApnBo+Ohj1hseIGVDgikQhPPWETFmLcGzW2RuU5PP2csP95
q/PdxPS4XmCm+ec8Z/IG67Woq2qjNVq8W8/FLD8CU5ejoA5BrC1G1HM55xfQMwaJDqMge3Ridwmn
DPA4D9wAaIhUPE1CkaVfrpSUi3sUpN7cMHZ5lH7wA/p3ZwNKBeLbBAg65PYa/x3oe/9FBUsGJBCX
6QNMHtU34GgpgX7k8X97e2vj5uAORwo7muSZ4axco2kTDC8ICQJ502ttD24TZ5/PekmIPt7jxvxK
ZmVvT/2uKM5qp7WJz7Ndkn1hBm7Ae9Fbv1LPdrH8ya1TsyJBeHH8kxbPhx173diAB207awAbgyMn
r+I5K8Za+VAsfvBA/t2/QaMZySWwJRikZ+01YOrrbIO7fDzxy4FCipZc21NyhsJuheJBxnHQ7KW1
vvugTfGt2tuz3MhVL3fFsSrqzvEGthY+sgsEzk+7YEuxqDnUVJW4acDPBF4V+7B0DxpYPEspqSPt
qMLTEMtCKnzU4FBe45p/s1SjwaUIaToH05rDrLWCHk68VdH091wV8FQIZ74adThDW2iFm/Wriq3A
mO4BkEkvKtZkecGCsmyXEZR0kiqDM2DlOBcoyEXSJp6Y7LKLABF5BdwDK8nSnQ9qr+Oh2kVENdgj
xrUZhtZXLESmdEX0ZTfN3LvzV04nP/2mv/pZHyUwanlqy3gF6USjbcHYuK38yh2Ar8km0vhuW02N
iLBsCJp6J/Zhkt3HhBCS1Rvux0ncRgR6JH18DX+URvuyXxeYMvW4MvZhUsu8tu8upiYkFULDJQA4
1xjMHpyTGliw9kPr/Of6FnkDXkEaixribLN6GdNMIPn/8BQNYKkXscExaaPsxPgLcYcWb+rlL9YP
5/SiS4mhZH3PiEWvbzC9DFojfiV+gO2LX4N1ECxQAh6HvjzKqC3u05vgAbDNCZKJwRcp/34E369v
kNeckDTH2ZnULlUrZmemd+Drxj7nNMXbPOEXTLXzRJeanFd4bSc05jnfL+bWE41mKp2exwu9eVOY
NX5FUntcaw0UvXoCilzUP//aDSmt1XiOyCrIn63BauQhPo64chNxyXzxDFskkoErCK5PPM93Fc5m
VtSe3LRn+n5w/fJu1VIKmNlUMHlXRi/xVMMvuml2WdVdcs1myyorKAt5m1QkdwlGXkULL1QQi3v4
4Qx2J6idNcyAH2dX0OK8KBDi0VjHzKA6BxbgQM7uS+iged7oflbYqMJ1aKd9W1MlKBqlkjpo/U5r
D2coipG5SxFpoNoIOPNVyp25RDlwQpbnyqfcQUX3Vdgn2f36ls9WRGfuJl3O0jfguny1PS03q3ch
8gNn2MA2yKEvzfPIyiqW62Jey/gGPX4tY97+bVfDWPqi2Uov7y+PEVsg1hP2eu4kC4OBqhgHYhea
nlSdp+aTII+yWrY6NUJUR5LKJLhISqDy9gJeraV9hHw5JLVAIo5LsJCzZtjEYjkUGL/ZqnXp64D/
eAGMftoIS6/UZJN/YdDCXef6Rg3eBYimjt1Olv8y7uqWVtHMmoKFzhmcII+OJo2dBbZ8g1I5JU3n
CLSQ5FZQ/1YjdQlrLSiNFRIJ0dXa39fyIfrwzVufsCtv/ekQG40dmFMCpF6nyi/jGxN8xaLHU5F0
k+qBFEvR0ZtMMiDqy+rcRReO5Ichlv9nc0j94hE+wwrv8756vEXzxVYKT1BOpQV8dSqMMcVqqW+v
xArrCA1oCM/3dPvDQ+gmSUTea7ixup6x4AUFXkqzVOlT5DDr/eYCzWVNGegB68qC3F4JZNUlPBwy
k5KI5ms5RHLAe7TeDDkXzt7eguTW4DjiGr7CjXwPMPPOh/TsYBs8iDJV5QD43sXoniPc+hQ82C1O
pBFmzOgYI6tn3QRKvf0YAClC2E9LP9/FfyUpeCTi4D7nTrDIBxPeeT+hd40KPLtRLTBx5h0nyqUJ
XF+9ise9Z9+15ZpzLqnl2x4yuoKrOvYra2wjgRGoMlY+8uXwOB3Uk+uZCm3zBdrhanl/GXm0mmkF
F6R/HHHlyum2Ry5mfn81WOJXhiN9AEm3IIs+u6lpTmIwPREMbvLV61izBbyYuPug/QiyACstjqjd
dDc5hH6vEdSpkTPAXaFWsVXNMP4Q5dHaZphL5VRI07osrFv47MZPQ9l+irM4AMkvuRjNPnzjKDQU
PhrAtuGa0Ktsx6fW2x3cv36VtaxuCOakHOTAjmF18+CodvOEIQtBoueicRbYI44tsFHiuG4=
`protect end_protected
