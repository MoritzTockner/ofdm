-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aGtbUBAm8/4+cWCtogN6ZjMfzomV7b8luzL9ssYsUaN2cWBsSY1oITh3XcOGP82mEjNlMHpwiTg4
I/9djXkY+qVc24PwtDJ51CE6dMgL52Xl9l5jhB2mRpXK4xF7iL191ILZsWyNP2/n3QOWXLan8TYG
2KQ3GuJT7Sftj48k5F/vfwB64OX49XbgVqtxczD/qqnKv8H+AL0rsTkAGahalPbqUJcPAk9+G88q
K8j+0OWPuK1spMSOXEun47EU4oaW+c7jvlIlOyms/Cn2YtPyGOehRYy1QIDp2Mrijdu6Hx9u7mTi
ULLF6KZQRhD1LR8vmusPDvdw171udyI4Do0zSw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
9/Otm4xC+kqLoGTv+1dECqGcdNqJDU4TL2eSmuM92UnbtDC8AfjVEZXDQ2KLXycipk6oSicB/d0T
CXQd8jcHezR03CCsm344EZD5XEWkpaG1WeNIozQqA/OKiqS4m+6AR3qorfFydYc3XejlWbTHrK1q
gQHQSxf5+nvlBV5yL/7oRpmS631z8w8JtiL3wHklQvW2/syCDGojneOLdh8Kg9vxjz1ir4TCr8st
gG/3J1/t9CJ+txd3IwXMLYOEArYRKLL8PFSrcTd/koqsdoS2r6LLms1oDlPcteY5RZ6H2q9ZkrSv
LgP/KGJJ4goRwQULbyxPwzcBKstXvLIbwS2Q74gMA0aNgdam8tLHW2Gzc+qTvxEtF97SQd5qAAb5
+qQDPhxaatQ++mnWgIXO3u/7MXBa/0UZEvZQ1LhJtZubQ8CtQDqyUB5YEgn3Q5uoSmhy++AT/jbw
5yp4IqcRvxYqNxtdZpM3s3mmTOkIf9V7WMcyVjTlZYVkDS+6yphhwdefR9W3JxAUVXAEtCxGWCqN
FIW02bIBASPMUeT0iz0jU5db6wXxmhtHlaoKNnNXKi98mfg75l+oCq4jVthtbYdegxxB2KaCZIw4
15DsTDCUnWXZxk+TQqebCmDNJZb8I9PSBkvmNbc2B6/oEqdXi2viqsgNWyEcESqtETeLX0h/YyV0
/cht2S63C2sh3ov4n2duXMWIZLPdLJkL2QdVC7j/qspcTbOY1r2hmWMEwOZmfbzhVaUaVPTowmwK
nKyiooY1+FqY2lxlqvDYWccLEOIMjjcolb7QCFnGe1SjaGaiRxHSgMVbOrbvR01ZhZkvYTbjlbf5
cxeRSDlgg3W9xhXtS5Ji4ZRLfRC77rnpwW623M3Ni6DhKCF5/Hqt/uqHSLmincrEozVEGS+3K+RZ
VBO0H42NKHIP0h69J/7BE3Z9lJHMI/3wpIzCV1mmSp+0xo7YDhg44Cq3+UhEmqHgr9RIJHESy6Ug
dftPOmwUZdU9hQNtPEj6zC5fJulofaL7jhiDpQsbEuKRdHTXLUS6516TL4pnAgt6Emp3dg3ysaiy
+TCyMrXnG7xDGi7YsqX6JTiI5jnhJ9occE9GMIqSrpmasqkqOigzXaOUUWpmLIAbj4GJSPs1Bpjp
4spUNPBvS4JanmLwtuzTBhnMIarpHLyHl6h4fuFt+Hm0VSf76RMnfpvlNtC0+Jg5Hv0M1W/WyDsI
UAagH35fYSLdqZhhWGmW8//uX59yzTGjVIC9jt1vbXkhqDz0SPNsqREGUTayKj2/fXAkL5Jt0Vhk
Um0lMU5NW/ubqONSg8Mvp+DXl0OSGVqH6ZwJFv47qLvoxQCMZVpwErNbglNAtd4n1nMK5SjiICk/
oNxyxlYUzIleQjOGG33ajwD8juZq4DENjwjMVBE392wR6mmNEpiwN2zq2SXemtP/CVNhRH4Ql4ue
30/2ZJHSybijotDZqRssoa0JOFz+88Y1jtPAgfMjWJy9Z36RQPGWMxKI0pMhkkMSGH162/5fzZlC
b6rXiEMv5nQeRpqtGGPjJ4J5jvI0gZF4LhF1+N4iYGI4uHfuhW0qH8FvLXdXLiEyrP6rjTs0ejnO
myAZLJiG0XRtPNU7OS8+Vg3v/yuEmst0bzYdiH10USrVaHN2Lzf0G6y6nlFlRIcLWzuta0LjoAd2
TjZXhSNfh7IWFGh0rUDl63i8EiHlaBA6ibozuF9OAF8p7Umr1M4ESuFEXAqujY+bVvRTuW7ekcB+
qPU6v0rlUrdqglZPy+itbhJQCq8nYwZ8oRYzjhvcn/r0WI6ObPaPlpUfTIvMesCU28TVayWIvl8T
w08xflWTgX7TfhKbbzrcSijCX5TABtmswb5z3XR9f16M6F/zOo8aujT2i1vPkeCBu9mMp982xlXV
ZuswDKIU55MZvukUbU8uk0EbCPi9Gs+P1+K5CKPBsHFeC1BteEiQCO/S0jozRCSU5MPgrcMmMZeW
wp8mzpFtEEEqaEzamsjxr3D+U3TOaz+ohe0OUPpUUSVtCIqx5N4lGmuQjNyjigIqtM+IOEid0gIV
+O/4o0YrbyRZhWBApslDjyXsiMcYzWL/L0r+VQPIAoxahk+aCFJFwZUW/GUOkxTWCYGPqAwQXMVV
75MBMs7TEVnvrqYAd49qxRQcyjjl1cnxdJ4mBPCz6exUU5mFe1ckxI4tJwcNCovn8hPPag1LCNsK
DbmnvWUOCLFOAMHMMB2IJas5niXz3QoTqBTonC6mupCh6GNa4sVsuyTsCacE9WZBMvUvSz91pnW7
5TA5moqPSYMDfrA3aix7al21Atdu/BbqAOftFiU0YhqollUPYWW0IhX4s5eZ8S/b18Uyx/qq+33o
UXdiLc6dY1ZDIKoVUwFIwWpb9w40+0o2c5zZ2qPo6DyJFHa2jytIhkqfclwHY/S+2pk9drubnnMR
K/N9i+0vMc5LkbxgnhlY0TLswnIvbJBBxsHKFH+rrTrA5HizgS0LK2L+HF0EUXRDwfIdey+/O8pY
HJwT1B10IReo8y9Pb1PdoVEgA8jzrpHDh+FLjKDQeBIlLUGtpezkyRHMtZzlmU0KdL+y1IE0gui7
HDYcE3AdhdnpWvYYpaJzJLcWLVuzfNRsnCuuzE0T9LpbGY9aHM12sR7oKTviPKEnU0hUsvcQaIpn
Wq+EFZzEmrg7BEBPnYy1woZzpd11QxCZ9mKfUJYigAznHKHU8s4ny1xGfKy6iArUxdFiZ3haaIdl
zA6Lqg06ZwRvsQS/z1RfBGBHbitnPeTYj9xYm1XDrPDqSadq0zAptt3nI+1iFW/65FQUxh5kGCC0
Md5MntVriE602Owt8auWoByK01GlfGHANq9KfxIs9AoQv1EsDKqmQD4XgeMUeBImagufagW+S2od
IA2e6kdf96bYh7XxiNiTI/Gp3fY6QtKDj6bY/kPGJFkVWcjJ/NLbmFFRx4cvMIylc1+mNRGizBoA
WxZEz9k6+817Ly0dAhP3sMeAK+YG+9Apj+IDHdT60XJNTAHkSdg4I1/lG3czRdNJ2VKmzbBplPJ/
v/qQclyiIQRkSKu386tx4wkB4qvunGMF4dkvnVR9+ANYERRygsqEIligVUcUlhxLIgtdOCUZtGYl
5+Rrl4OPxtb1XIj/CcQST0gAQfjTFuOr2kNNVtmEI17ua/ZGhijy2UfkgoQaSQPG9anZpha6tcUM
XDfd1OY8bG0Tz8wpluls907OitYIClFDdhZqzhNTD64IcSN8FaiS9tifZd5F9q7KQzu8qoEWLfRT
8ALevAsNhhc4QtcQy7F9hCc9uL7H3z0mFhTdLW7ZyOfp5S0/dKlB9gtmeiF4VFVOns3zVJHRRG9V
PHwJMNj62octwq9xWWgMKhi2Ejplfw/NDtIvXkYSeccY9XGhaBi//nY2kfsW8NAryfiKc+pTNrV5
pdFE8Xzu4mkcJN74poJx5B37iZFmi7VPz0rh+q7vo+chnMiLNwaBjTKv8RRGSp+J7TalBVfyj5fh
ZbJvWzJLTg/HdkiM0DfaxLAzgUT8LFjhJ2+PbDZmXsO/m0o6frEHAxCRt/zy6vg1v1SWOtWc34cI
DgGyDabspjmCcdrLQukDd76lXzl8yIidllYVYdY7N3wIU5sWkX+1YSiRTrjELat4ZTeqjLj5AmIG
lNgXyekDYGtaT1B6MRmv6b2wmL0UumZgbF1TRPfLrJO6xIZgWtxJCX10mnVjlwXC6NPwUnB4ZeOA
ULcobfg8UmI6eUzB8FGSWfV5Xv8GWXFvsO6vejo7Vcua7dT9zRBtBHkALcM9Q9qcanzUjTbjCnqQ
YKUrpR49sZU7By2YYH3ob7V/mPapbSgC4jciw/oU6IF1JQCePObDhLDRhOJIrCFDRmH9CYg9s27L
t58DppqMQzgx3bCw2uXVDchMNbMPO38vEkeY5bWmaSOC6CUHVRH5Jaahe1p21uX8ZPx0flnovnmk
kmKuBMpNDRAFpmtrlXTsPQ0DaPxZ1J8qHxcayHa37lnSdoINGrjwAQWNxLgcoNdV6ZSe3mpSbyrf
YdVMbHeMG/NMll35VkEnk+v+z/hu/F+TWeUySiR1tqlgdkGD3tIUIcETXEG9QE7ldGoGtUap/yz8
zeghEkUGc6SgE9+opVBVZ07eY+i7PxUwtZYllDinhdrNNx7t7fCD8eLepwgwRpqqS7yYi+3sBcEm
yk0XsNpsfxNQCyELzokcDmBA1i9629n5nFEFk7IkZ5kwXvl+6u8gz++4bOuCbk9m2lPu6GiuFe+m
3v1bb/8IutHSQNE12zUWnzJiz5XWWLy+nZJ1ec6nYRdpcUtT9MYwLLjyShVff289VjGeBWKUreYi
eiO+OZ4qxKBkyd40YzlyhjNpXONlMFd7wYTVwLI11W9hSQ/iYSfWWy7n2+3WOVfa6hoT+lmgJJo+
Zzc0o394edej1CVWIP0x6CH3JklgVC8hd2H/MVjMHC9B07H+SdQjMLHR2R/ZFmHhjZVknD3a3Qvx
bEmLIwtM69Y43G4tfGscV3RWJCXXqn5TcqgsFnuWHxg/5hkTWY7hEMtV7PD/Ipcf3Zn9xsqKe29T
iSB1bjrU3NP2YTSFdcx31qNCqOOWFs4BxmfcDUv/3QxCun9/8ekU6k5g6qpnHiJZFFwFOEDvnxdV
hR2sqTrqEgxiUJNX1POoXn8/R0UQfxKetXXQ2TEBxhS1oC9zC1you/WMs4QKNlx35Xu8wpr8hoS1
3r1j4QvPw0xgqGZcjUhh+o1D520XXNr6v09hL/soQ74imZDxH49J2bLHEo0MdOmKMhqP/y9/NPrK
cdJkXR3l7dXxzxgF1xk8aEmQbTm9bemMpczWsCtkgVOPp0RiPjMeUqoQvQm0RTfl65QHRtoDzXeH
n2I3gl9uE2RWK4pxZJui7axlt51q21LNAgZe4lRp7bvcJuoE0X9CSoMpX1UKeUXlhLnKT26ZIJPS
v2dG60JGdPuMAKIS0A1w6LDZvzL8AHYUNQPuYIj2MHiNXLTBZ+pbwjzl7emFMhTgJNbW0gIav2FP
ESAc9MmGFiRPLODGE2DLlIt1sBv6GmCXAGfmxFOFMvEI7umE68lMMrQjINSGapQ5yci3VS6Ojw5s
9RsgYgZuSV3nowbIqz4LGFmXtEhj1Z1DSlbuN8B9GwkG2zjrGzRltmDKjfYpz4qyc5sSJ5y2p1pd
X5nrht/Go8PQeBn2A7Dy+93zm+2SksFAYfkKt50YUVFJPDEtt6iPUrA7Os1UjNvMa9QI292gtxfx
WcRCCobIWU7u6l6kfYhP5AfN/65SoEsM5qNOZ8lBMGFN3n3GPffnkzyjugE9TzIGNQAdTBVEnw0J
JYlORknMntOS4sRTAIfsIudF2gUu5amBYQ5TZZEffp+sP5Xbp9SGuKBqvi6RBW4xhA40gfYb2BOQ
ShljbrhvQWcrY7VLjT9uiymz26QQHKpjsLjQg3a9cfeDEAYmKC2NUxL2kFnXcADNuQ3HrkgNGzKE
HH1PB/bLQs8MovsnbwbAG+bDtMHgIb5KW5yyLdooRvZJX8G0kJUdoWaimMNxuRnZPEXoceDWwVUX
x6+njRvH41ejF6exwoxyomIsV00EvglAfheg1kNGX6gs9qly6fLHEnaX/EWkERrIdKxqCXDrcTdT
t7BA837u/qXoi28QY2m0ohe8rVhTnm2zKzPjUmQ6WWhktIzr37OKwNpp2yNyrn2A8TyXIR56oQJZ
NiawEruNKeQmDOqVVEjh2upPF/Y5vBCeJ0+V4a6aPMO8+1rOdSB0rGKhD7oPQzK5cdvmk+yfJpoM
wZ9HwG2LB3OCz7BGZQZ0g37e51qP89hvO3mjV9h6T5acrpgsf8BSKN0MVeR92uH+E/eu+q7tzDa2
aDuDKUU4o5FeO4pmrSN9FESW/PQ25S1o66GN4YPRkPlijjdJzxg78eszHvEBd+rc6aQB9XBG2Gnj
awZgYS9c8t3QSirDbGT5psh7Drz3A+lFm2lT2+QyHI7gsc7AhTP3EuCbXv14I9n2QtMMuawuQ5kw
hQFxbx5xlcLR119HMFU9vIRycnhGuGgD8IYIIwKQOj7kzsWwCtazZvg7CComlNC/8l4H6XmBsevB
6Q+MdKkRjf6o3PH6S/3cL34GA/oHEkn6LuCzrJ1oYPfymd99SW0dPwtdeEwXcGopIko6w5TPI+kW
2Q1rPqFZrPVLiYLOaOCUSGqUzHPUZex8t+QmgIf9qrHoZFYPBh1xLDldFFnRnOqJhSdCQiIi77JT
vYE9XFjA+F+NjBL08jMp8PZk/x+rgWcfaTr0AEI5BTWXH4SfO1O7mbkzuT/SGZJFMFaj717U+p3a
q6kMYLEwfiqv445+iEaI1CMqdR2rgI38mFcH/aqamlakAccg5+54U5h36ttniOC6rEEkVBzGB6Pg
E5+EZL91Xq6JiWk94fPEXQLav1sViBu6Kz1Qrxfw7EeaYaY6QDHhmOfCyAVypCbKXkbymwn4xMdv
xJJJroj8Ih4fXm35oNH8j26KzHCmwyVZmQvihAG4wfRcqCSWhGJ8Wh8oXS3PCZYAwy+9aWXtC5cR
4vrF+d8bli5KX1xH2C46QD2xMsbwgNVNy53UkehPElZ2Ed49tFVM9ZcH9GrT42Ibf3ltWgAXhByG
on/tFB/mMnrnuPFNqMeAKGnHZ20PZOKtu9yajSNrxvOB9K7E3ojbbKUVcr8IUtxhRAlRDJ0uKH9c
Av0RyFjetnqcRLq11X/1A/fW7yEM5oeNYTZfmArpYE3HqDs5jAs+Rj0Xof0AFriMuPzoC/PfJGs/
/iSGk6q0IqNTEquABTCcFNYtbB8xkErmJP/lyyNxfmDASdm7Y9Q30dou74teT5iyGWQxbKS29xTD
O59hEUbg89wRk1degsn5dn8AZ2w86zi21QCPxZCiZs7C/p9KcS7uB5E48/6Tq9Xhjzo913XiapC2
eL4Rep3+f32wU201GqYlSb1JJFlcY4UOf5E0pQ2QoM9pX9cN92g2ZE4G4NHe/QxBKG+RdEQXCdTm
oLapNXVCZ7oMe4sCTWHQ9mRE1vuF7ugL8gCaJ5bqIPDiCbbpy+wIebT4pA0aO8GHaEx8jjVpbGVe
LBhIEpfn1WLM0GTWNgL1ZSfxydTIT8PSAnwC1V0fLzFY64rYUBmXSZmz9E7RTlrQzug2qKvzNKKt
O6l9KEaTrViMzlyroqD5GfgWz6arTjJG/OQOKRhwmWY5KLhVhcU5ZEvXHkDyb27TCweA4XSqGQpr
efNATPDyaWN3kQO1kkAuq5YICNbaBLcM03ykPR1KaIG6IDTGiwZ2d91i7blCp57O6SH9fK5jctmX
CIr26balFGrMfdGKYfHcx+dKlxFotHikH4YFwK3g3jbXaNsrmbgySio5H8iEgmU5erC/KEFBVHVQ
xwex2fXwUsE4yOeN6rBDVdNpBm/DAqUhTnoxUeEr0WzWH3HvbLb/fE9y2CmbYxtAh24uMewMLdaX
NFN6bcg46qQIkxEP3bCqcWymCUmDKH/Q9p2V8r0Ddq+UqxXurcdEBNNVlC7bFUeBfgyg7mXJtgI4
DMwVI4COTi6HIjG8c7WK1U123yPMTTY1xgzs0jrVBALkOO3UwwaVpRLtRI9YGCMYJ79Oc6h1y9jW
Tamp16pn67B1d4aNKW+hZGJtdVkoRSsjEPJDuGmzRuohAuDj33tHoJBaR+ZDehJDPTXrsnzJrNZZ
SYRcD0Vym5UPsO/x8asbgQo2m4+k3bkhDfnkLRxei0SXjUaQQpaTgPZLPuMro1XZDGw/YESnMwVB
J1ryTUhSH/hbkUGqOwohpsboDeJz1qL5mXXAvaIlhnarRxPXX9piB/2SlpN0WfCKpqhq5ZkHLR0l
7UbiQMeIdT679OHrlffPMmwW29fICSnbSHSdWJHnlP8Z10qkydSWBZ7fl1xbM/0zz/mhTus9OSjE
QxKz9phFlZ+XZXVGRVVrvERAm6fFO33u2o/YVm+js3sNZVtwmWmYdrTFCS7h4L4zPxDNGywvUckQ
i10yqaF0GXdR2tuOfrxFthxo3kI3udp6uX161HG6QC3tkSqfDgjjU0Rp3YiIrbiucL/a59yWDRPC
w3mJ0cwxlaj4dWl/1LKItDFlRZb4Hj//BswbFCL0Td5tf8ArDG1v05scZcAJ/7qlMG7qpYxHM+k1
EZD9f60vl0IB86TiMPeFkt865Pu5LePlVJsivsdMQefZG8/JZ4cQ8H1R6nxgxfMtbq3ulmvnvBD/
XuS0+YFSOuKyr7vkB+bFTMKGSIpcqU8NFL5WQAM8KjhtdkDK1Hzp6JMoIdS9IM194Zee3pGK2X4v
3/rO3TB+0/PNb3hox/7WZ19FJ0/8Vrq2RcsVY6yZVtPRctYSAUchyTtbeTaYU+bYmiluW5UVQdWE
Q+1cbyoRNMNgD02qbiXR1eK/5TIfvMGBaxAlOKTPAP3pKigKBNXLUrjRifzZwH4lYVnUWn3tIp65
V0vavEVkIiIMwms6fmd2jfAhUzf6g7XFMq+TOyg7MvrZa8gZFYCKkNEi6U4SB5iH03nbdIpLscBI
0e6WP+MajwrOx9Ua3Mk8MiIsSGf2KSopq3a7NzqH4nVINBS1xj7tCdxV8PMpdo8BfZmUz4UZOGBs
J+nVOMP90NTRhdeeEF+83pp4T5ai/jZXQMjx/4W6xMCRFmRxM0wDcNuuZ048HLJ75sTCUjh7jCmL
lRk4UgfjV7plW7onwajTPQshkdnynrrM6PcU+53oYziUsfq9LYkH/NFK6lTC4nR3Z+li6BdA6JPU
QdEEXw5Df3UDv14847dhREXAhIgxTx8y1Pv+jRg5/c4z/VKm+n9nDmJ5NGvh96mSdtxJ/H1MUqKv
zYZaYeKoBNhISdrxH+clD5BXBmMmlEtmnfqeQsvrBLeNssnmnTrre9xEEHtuuiUzpJPoVFl55XyP
T5WL2M5gz+UOYoxYEIZF92LdAZgT8JtZWNiiOT2Fwwek7wyjBFrnYn3FnpiIAJQBX3VwtjNFrjIR
O38z7AEy2aOY7+p4d6s6s+Oz3Yeo5jFUHgTr7SqStmW81nJ2u7u8IJoFjBhYRFc7K1XBHqhxRD4b
K9Zlmc3eWE4mZ1/5N8HlFR5w6we+5An9q5u32jV5ADjyRFSOa1e11N1vlsLmTiqhgCN6xB8ik6/L
LQ1BxGh3rFH4N7LBIjaK2+mOdy6WExHUbdrgg70wg0fzmJOtVlNhdy2Dy/BWLsoVmDoKMWwij/gb
edO6Zvj4skOLZ5TruroT9j6HZCtGp3k73tsO5oBpAulaaN/T+8YPB5eL3b9LB2tzaOMWbl3B2C43
3ykC8ZhnCEJSCWEVqU4hWffOFte/J1IvjTNhs/sKPFEMtAyfh4pQfFCu1eQKgbWGdqo88WFk9fng
lxDrE/fJrcYoTeDkhXojyBauHXTKSAXvPFXiuS3KzJ10/e0k5yc+XCeFQrIkpDIp+hq9viN++i8i
o/JmuV28MRZ4RDl9Jgku+HGEjpJZNIZ7WLSg7uL2ZqiTbEZZ6KRFOrAAsNW9uHtcYJhTTdAlyDR7
3+Kntu39Da04pBssoVvVndjLWEJG4m61lW2XGBg463QYH3UYfe9/GhFJ1M4jBs/NBEuMz5IRmMen
/2X8E0H3kNUvlLaPzMHaSGuw6JGX+t6SMd3z6WpYwVDnQEZPCP5JJ9y/nrQEEjXdtWSELWCb1N/b
joSJjJ0Ibo3FxlarlpksAIMjqNxcqArgziA0uSR84TZJ42GlAh9wZELCeq+Pf5OkGKek6REF4MY3
k8YDxCaC3xGTKUFOCvGQVutVr05h3jzBYRmKSDTrfCo++TNhliKqq+jqRr2E67JfVTrJzC++ZEnp
mZKe4uDIFkKGC6N0uwx3TgphsYplwTf2RBk1+n2LKebMwpF05eZwFg8uuCPsiD8BFcbcRSpfrfrd
FjZCXAjzyXQGqmQ5JB9gfsJskUkIZ5kejcFZF7DHzN/tPnJTCJlDX70+fHAv9WLFTUG0ome0uo/7
fytvI3qr0adCm+fiOktxVRP/yABocpBX7ADykvlKOnt5F0LZb/OcgVfbUuzuJgAfLaDWKJKki2i8
rOZduUig8xkCUkHffn+h2KBu6to6z76g4oB+JDjUnNXfi/D5DcTPwNnLQgA3R3EfJvLjgY+4C4aY
I0HTbMGA15mf86z27sr/Q6pPetFcmv+81wU81qcqrtDYk+GMk/+4ZyRLwmw2hDGHPBeWvbn1KO3K
pOZFyW0oXjMvPqw5hPjKt3j7FsoMV97IzLJT5ODTEs6sVhGwPlQWUjEYiXG8kLzuk7G+xnw9mhr4
4dSt6ohgZTDhnCFFjGRBdV48zB6C38VjpoLKIkXw5pWXznH67dAA0BNeFtaqnmw7iPh2azS02U98
mLlrjMOUODNE7jyitVMmEp4lyjAM/zpeUrEHQuY9R1qzRZCn/w+/4e4daApwWs/NF2B9C4IJzQfT
I6xSpJ4uBJeyV3EUC4bmpqMZxJQfkaOzZmI/T+kewm2cRIYLZsNQrKbT1xvBaYjg0WzR/TbAbkdm
J/1ljzhMrNNuQySo+jIOucvFTRHhX/AcWcMCxviVSrOzhiYq1v8jO7tK7Ai90g0dfDYp+w2wL/BL
7mq4Tqt3mJaNaRkveeDwIBgQHBA6G7jCYAZu66Biw1NR773RpD9yqsE1MN9O1Xo0lLW/qheeuvcY
H6BWJqcHu+f2qREYBpqdQzbU97X3apeVlERpUzHuMTe0jbv4SMuEda6Js8O1/iCi6Urv4nN188gb
a3ThqPOiy4eb2uAn2NacJik9tXyOlHDPxE6kO8wgYP1qTGoDeimgRnoAredT0ToUKoXrQzw0Ydkl
IK8NfjeYA4VoqYYExD3a7xEn46q9wg2DxvIxjHFVRs7YDoknU/8JiaT6lOSlJfQQRdgeVeelqWXa
kbBei9aI6JVhFWVIIY424beXvctkB0WhZXL7tVavVDsn54tiXTuX2W6KgyKNPurSWNkCXCplxKW+
3957bpQeZO2qCvaeIyzCajF03nMUBC7t4pgUNASrO07cp08y55DEfMmt4ny5AlLPN3U3Lwfe8vuf
E3GjywDlIM0IOgdqPrA7LhAnQpNmHkr8X7I7Po+ff596VDnCbOSbVN2YRKRu9W8n0hCWxPAfVhHd
/nBU23/y5ZYnC0aAdkAgcPUt5oC5XPCqlepRkO2S5uRggm8fFGnwGKYdodm4SmWDJvKkwtb+eVpP
ZF48Ve4PT9whBuX/OiOqZ2oXjHMC60EtSHg84uX+xUt4IFmUmfTbN5u1AtLiUPldSrLQKDy6H5x3
k6Bes5SIngHdOjQxaT75s9T36ciVXPIPqF+4oE/GlyvE7N/BQeoAA7Xpr35h1Tl9Clp/HkIlyVRU
VVqzCPBtS6WkEjnPdnt+2zJWYdmmD47CRegtFLokX3H1AmhZU8J0NTOBk9sf7uU17ulpY2eYQJio
JdYVEKXajxw0kv0NwmqDkY3FYrB4qx3Yrgz9odiDZKj1UW2Y2zSf6kcEJaC/nmBj66GXh74TWfhc
C8NIoBvBsXRNY7JXllkhvChqg+TFyHEMqg4F92G8GXAX8a9MdRq9pWh1JUeELF/PIQ8ohBQMKwaH
Dx8+fkjUPjq8mIZPLXs9okkDMR/7/6OHNevYNP8mr4Ue5UQvNUuC/oj5hCXpRuMKwh5M0alJ3I94
iKqUfSJkF3Th4UB4hEjNmjentxDeATs8ajvgc5P/ZYBelSkMhicclIPiIG6UzCrnEnMa2oC+V6nH
pAkoOfkulNKwy0L8n0h+8SHwcxHAQRAKgkRb4VczeF6MdFzI5TizCbCXK9ZfU1L/VpEXlinVDQjT
0+8z5VBqGdvokk+E03ugCRPSZVKX3OwUzi0NozmyOwpRsDqPfVcVatgmckiRSaR+jtsZWSf+KExC
Xg67pdqMV4QpBadepNkUpOAw9OnpKeWPogLS6G+w85T2R+3nSTmR4ZuEAZQ5zyIP0lQJ8oyRpcFJ
XAhaQjcA4pwlo3TIeukybZPuqeKBjeiIlKae5iOlON2lLZP9jQ5TLim/Z2I8dL9/P7VPRioKLitN
THecGxOgXJnu63ao176q+W84sDvWtcp+Cde3jmgPfjK9X5db009ydWDw4+VNtpGjP3s7FzkAO+oY
1EpPJezCoXuXK9+sWaqO7qxznfFl2kAORjOmitaPRugybFPERonimAFrQqmkHZJGOCpYWd/mDVvD
1p6r/vQ5g18+0NpCKZjRSCDJA/MY+R+Ryh0UAfkmmx2K0wihjNB3JiuzkDeY3Bzmz7qGwTzNiJlD
FwvP1Up6aNPv4mvHKjuBP5JEJybO4chk53FddIoSUTAC50t1vhI19CUrWhbLKA2/OEMPlP8m9gPC
migsgFX6trvAxRdfT5aQKgBWrgSg0EHf0vP08jntD7lpqPiA6bqYVaoSeWAUbwYLEQkzAFRy9lGz
+uoxlunLdeF9Z8YydmiU/mXLZD4YDzpWstD05Axq1UJzyfqH7LU14U10X2Z+pGH20hHNbUbDsiDO
9+rlhtidYw5jMGm63HaWb1LnzVWwkBU406Q8psATF1wn2i6x6+KYiHL2LgcqWDLc23O767/AzIX1
HpcTY1yqZtfV1RJUmhaB5u8WFntn/i0XSprC0cXmejFeUqnEuCXKuZLI4NW2OlpZbhzC+d+LEOfW
b1HKh2Z4yhDI6mTX1r0AlehZE3GuiyMH/0FSoRVrTM9EQVbXSOldWm14VZL9995/peUjuyc7OUnN
czKctRsLg/0ktUKMV79eHbAYrLyGZUgHD/tVz6abbR6ZhTPi4QxCpjWcD+QTO+xuuHEmX1gXbOOI
DTJbVpNtMbVw4zwW1CFMNT2Y6ZMlQp7e3iJoGO5helGQnrWUnjo9e/CM+hoSMfn2E5l7SdY8vsXm
ffoOuVfkoqM1/OmfemQaw5ggZ1zoj1XFqVYO3qAvp01Qc7RoU1XRaU3yHi3wN9iBq9khB7FgWZsT
tdIxbilGm7OTbe6bAgQvvd6owVofvtY7Ng2WBf/6fGYdtH/dYmmE+ei73yANMHb2ZH4a14ixil+W
KMNEnH5PUELXpGlR5ZCzW7TVJCV9ZbMz6reIDc5iz6sD5Bnx4GXETeOFQZ4dulWpqpg4PQcKYjjl
vVed+B6mbYj2BSypOTDEuIA6gwOBd471tAKFj0lw8mOZoMuxi7UUEOPru76G3HeXqg//dLHOMTgP
5oH+vRe93Md+kx7taAK8gJ8ukMHicSsKwAUefaqw/15rqh4jw8kWKqH1SUHPpSaKNlueIRw7HpoG
/kdsBy795OeYNYSB3SljT4r0DYAkRW4rEHlLxr1/IHbSywy0ljJVIWO6Y5OwGp0U+XgPzLMi4p36
VHERKsdFT06oE2uScPtnN+THn/FSCelEPocZ6v1GQQ8PjUdvSjzUoiKMcTitWbScGyKbI084ed2/
bACLaHg+h+jZXtAiEj2SrHNN/0OP25lHCDolKY7bHmFcoZdrO67J9JmBCdNeWArJ12dKznz8EBBu
SxlIS5NO4g3sRiMvqcOKsnNJdKKtSp+OKLS4ZmaELoYsS2hU3ym4m4coAjhRgj2NOk4WrQI9Y1nD
8HXauz89Q6M4TkeDR0zi5OFO5HPsNBVjI7ApehAZvaHBHfxNjOxPbEHC2C9LVvfuJ7YW+0VMTbCT
C78vSlg2rY4OqL8hWf6/Rj2u5ReJnvZIX4CtF0TPZiUZHueuYhHX47DQUtD/rMm+bSHQ7bvWMP3j
07c0n7xDp9EB0xtt+M28ut7wvzHiaMYmIV4Po8BdW4Q4TfIWGqRBZNOhLR5dYhZ61e8M4/EzYv0H
PxO0WTbrbK3LFZtVKZa0V9O/Bi1QDl+0A9X1L5I/WR6ENI1+4cE+arMgriQxbQOQtYyVwwsIyii+
Pjm7YFA8fDT4vZEOQoVogQmwRmIwj2ldC7mxwwO6Q5RjXbDKAsi8LyI+mn4cqehJcen1fyj+HGoR
TzhM8nk16u0bMrn1Wnl1i27b1L3G4gD/o8vRlOKnDLvscMFqV0xpPAJ2uEvTV46PB5gk3y3zO6Rv
yYSP2EC+DayRvPgNtdADtZo33qVQqmXx7+OBGRrQP3u0Accl++YFirpX/3fXtzZkgBOWhvVCrR2W
JNcGTQZr1NkmrPGe1cSgz97QDoQdTGYH4GW/MQXpNlKtHce5+GQKJC6fg6g4zcrb3bqMf3+xLd3u
tVD/kiAA+J+FMnRXnXjWcpALnwd17u/e9LvvdEiFUglL6YHaSXupVvPoUlq8EJ2IwBhWfOw9e52P
Rrv9fX+eritFnbziXGCHz0lfh6ZqqVdpa3uzhh0zfzXBWgT6FHfiKooLNdwQtd6vnYPLYIF4TMb5
TZ4kzE+Z+GjAzZ+kW3PVxXyOxKnYXYL2y3U/7ZQJyUtU0ed1LzcPMeu2tUrv1DbYMl/IjM8qTtqg
yCyRXoGsFeHZh4Uqv1WwtDQing7xHk+8PGZ8/+baI2IVrDFxWmNbfglc0mMl2vdKpBbGM65QY6YX
aRf0+CPabjydV9nWnvIAuNR4hbhU9MEfpY7BDu9YQ6ckLArv5LHcb7uofbbncm1onTU++hBAC6O+
jV494AIY/O+FzQVzxGYfDsznAfzZ51P5R7IHTYjrnOr0m58QwGF43PH/Nbk+BaHZW6AoP9mwOWyv
FV8/sZH4hYoskF4YJyUXUU7rjV55SEzpUFj3WPn069qe7v5JnPwa18ajVVwQwLxapQKqsixtmNj4
lj6JTguDEE6avWvmBwhbpOoD+qAC7a4Qw+X9BzzFs1Qquz6tjlDNF7YLgUM6nZ3TJku7BzZ9DXoB
ttrieeIiiDNzVNn7rm5/Md3DqEzdQSUsK2uH3KEKa9NXdEvzY7icp0XYilihn17Qhf9KvF3Zu6wI
cAni6eKzCLDRKg9/Kd4gVXwW1vEtE8XgashcKShzzd0xg0LYYyTQt1siNTPE/+aJEpD3u2bAlK3U
cKSQUwwZS2TQQ0bXzrnwZhOn/xlE2jCEQdVtT926jfOJvXbyV5PF8N3DTxO0Y9Gl5BFwlsjOY7Ea
0VZE4umphhRZcN1LxnYGn7XePBv1sVeFZ/PcbstjywRiN9A9KLA1hesnuwtTQh+yfIcIrl7iZT2a
wCUGuxNWoD7DqVnh32+4C3wAwRMrv2CbCdar9lx27f86ed8hi8JPvEoAyFPn+xmd9z0o3FlNKBdX
pt831kjaiTa7DFYX2hac7w+LSC11g0er+5MCptwsOnHeoG4QKLlORRe9PDCJOFEW9dih9RVJoJbC
VVZ0sp4cU3EdDN5NcN2P2rrtU0Dd8zfeobaYstSL1RyUkWQZZq3wd6DtF4zNjmDZVyweA2/C2kPP
3DhxE4JSeufoZdP7NmXRO+PxYMTb3CSCYx+u6kp5HVPSjmvRyRvtIzVdWXa06QzAXIapvgqc+P4j
m0OCRI4ttX4vKi8P1cLgyQYlNvARGZlyqDgOiaKkqcNW7VpGni74khHiOCB7YqBD7GL7eT59R+rT
g3102B940X6+uVKZAEeewuBYHMYAGUNLILuBzW9SaG0DSXphvApH3Unz5/edxRO8mVZ4fq2A04P2
H/lMUhfOGyg2c3ZOq2XpnGnYTisQ+vQ9ZcNzqySbyMtpbMfAlBFnarTs9MHwTQRMoaWi7AmkAckJ
MjucGyZja0ULUO30MsUCZWK8hibnysg9ZSXCbBINLRZDiLjwgmzLe59sE2GkrjKXDomqf6fILWFq
2/unBXjK3/yNMfKprUdUpbuhyXnZ9deAPn8R5k+gADqz9u3iOVmLOkSpzT4eW97nkG++Yrt+FLVd
tQjh9V+FZ4U3FBaLtyu1xmnF7Jnp0qveCJ3nzdIpB+2343iw/E4GTJ6i3YvdowZXDmmDBN+AD9zL
24S8VSXGeTNNejVJp+RESP63oSdxVUPIWoXzGAhVb+4pXLHwR6VhcM/H47dtIK2fxxAH8MdQiDhS
vcCDT8oLMbe5QVXkXlEAKRxtHMeAx6MeGtNZOBPHIN5r+ssd6xXxNIFycCCuQKFiVelh3LzbHRJC
rimUsEuyEA9wWgQVIRljxtGP1vp+ZstjnDFsyKxZCXOda4GZzjvII7JYOp8QYAjMxgI9iw7xoJxT
WYmcbEHKDpa8/aHlmLthvVO9t+mh0LbUrTw0RQV8kw/7AS4YVh6FNUXEh8qhveyrTH6QetdXWIIX
4SFCvrKPE+KLu1YK7Iw+zH2dWEWk5HsuDeSv05yVbWaAJ8e6SjB7oWeeGLGeTyyHsecS/tS0Svbh
eE3fczgzh97/xIfV7bWe0GCpdGZKrsGgZMx53ioX7jdgFBqZul2BqDTd22+HJAYE90rZqa5WI0+H
cVOkz3xS7QPAKUN9o1Z/vVa0kl+x9JSg1oaH1XGk8oXqWQhBks1DpWtmKbAwk3gLgi0CwuJusNjW
Q1OckLK2GmtVZEPljDF0KmfkkpHAYUBAUS+NtFMmFRztwRIrcjXtvsTw1Hj0M0mLQfaHd8kDM/A5
Y3ZiBGrebSlhwmazNpIyD/e7YDXThslhCALuiNH3NSdj9BJuD+k9dWOUuo23+SuZ0yr6v6BbG5Pr
VE8yjODn6bihMQn1TIDNEBx0fX/MTqZbLDLtkObrkRwml9YrHBg2URGDjFbS/pMfo8N5NxeaZhnH
nP3dcLwZ2O1X/V5qskHz3GGrNBX6QspQlx/uGyo4TQciYwl1uo977FPmlP6lOXYeKmqQAch6llJG
0dzj/Ug4Mfz+hc6S42LFuWf/lnU01/zbNbi+cvlU2xqRcq+XLuXFEIEQ5C2HIZSnJelpMFyiQ7bB
SFIY4/NaH3+7jbQFVDwqN0E1NhXYZp6IH8iEWHYmKdvW7dhVVLFf5Alpf4FImNXkn7wM/8YctX52
9+JKqSxrX6XuUs14Ni9ITuo4t3OOzkjObo3/JD6uYuYltf7XKmQ2rX80k6/jYp5pAb+Eyd+6pM5j
cAdrT3UoeijBZ6eNDqjKIdyWwnPb+S0oHcNf4C9WLjG1q/pX/lWIdeUngKHUSJ47onYoSC3jT7yV
JDTqIQgncRLU0dtlkiAO/SAvNOgszch2iObZUmKCorV0BHQy0JsF4T97Duy75RT5QElq+7OJ4WlG
ngY1ufOFvMM4SQROzNdnSICg1+KVTJ19FmZUMRUtAf75xIGxZ5Cx03Np4ZyD6hvYVX0tp8g3XHCf
gYntg89G1bjVK+tcjKLiUD3LuR932osvF6qgq18xiAouHZTWdqj/byJsaWNaGATG0Dqh/lasbRuU
dWGKyGcouSpFReLZ0uufsZShEd5lyxTm4Yi00C/QuvMHKGYuVgDMJqhYStpS6rAiQqzdSgAxWx2a
DEvnPtwjclFlM+kza527rsVSExJ0WAbeoBpgAMfMuoc41yaxLD9wOFycsQ6jhFVCEdgzJvdgZZMi
Jy0Xx9S7L2jCq4o4C7I+KBPXTFlyBl+i9FJUttC9ZHMNT7JE1LrNcIA5opnqBXu/c55EfKWKbgm/
ITBy6zLHGSsEmuK8MSNqW6a/4lCEGYErGRFNwWxt0pVxgc16+eJ0CktEe6rNVCumRTaRl4WyyJrb
ta0LqPenDuGE4lR9x+e83AAKo+wcOUh+GqsVHo/JGXjIN86f6Y7qOQZWaQElsoOiz/CK9ZV08vWq
qs3OOXoSsKMeWA78a2LyyH0xvvUN8rEMm2BzVBhHhvNrvmEI1GaEe9aHw3Ls0C0uXHY0YBMUqwoa
hUyzesqcuTqNHBj2Meu64LR+k1s6KQtyWDAgCqQklDkd8tanEkXM2CL5AGAY4RNHqBj6JK6ZbJ9G
mdAbdbLzea8sePqDcQbYFT3SfUmvQ1reyRNKWhFh1hBE43RbdQmq+msr5/445wL652Q2Z/VT2VYD
jXEs97im2mYfSvuW4KSGHWJNABLXfpFltUvLznfwtb6iWxowS0hOr3qE5m0i7VbOVi2bB0FlwTMR
c/MpG58mFCtssxo8Ix6Wrw1dTry4zmU6IzpYyEAk5luFztYJ+00DLRgJpg1SpC8XsoArjgga3FeK
E34sCAsskB+Q1FPteezHLpUjJxBIPNMPO9K0vqDM2f56AVFqtw7ypFCM62hYjtWVhtFtxPn4Pgf0
CIFLyt5B1kDH1RYGWEOYDXBFydHrKZuB0DiJinH1PbbQMNFHHqG3azkpcthdew3iNh9/iL9QUsm1
QhhSMkB0GEOAWGnF4Jv2rWq0SbYk5AJSpLBVl9Tb/A9VCAfTpWX6Ya27Y26pJAHBi3ZVJqOVeRSO
cIut67XIC86c2SU4Y50PZGAy/9IpewUXF2mI+ZK5hwTC8qEQF4YkaNMC21Rkvj9AYm0ns4lJhtM/
vqr8vMhcFroSdNUHusb5Kdjr90WP2hQs6TLirxseK1P4ocIHENSAMt9xl9k/73iWayd3XuYkedLV
FLIBC2yluS1TYy6nODXKYdM6YzsxZowma6WLbr3LEunpTO7+x4s5OPxWrVkr3HiTtO9Op/PWMvjm
F04Q+csGJealLm4ZVPGOTG9NjzChwNJwp7qBBJXQuwN7mtJb25rSBh69iMN35ZOED6l2XaVr3Q85
nRGRAqltMW3yVVlt8AE+EFsgx4JyqyQHvMxGYjIuCbylXALoR9YuBTIoIYOZwgvIJHpOGaAB/Yu4
XqQVLBC8MtjBhzyYe9u0oE8OI6dvr2i+HVgO+6Ti817Z+LuAlulnNAy2jP0tspdT0f7/AdpD30Yw
sEK4H80kP8JiPWt2k1a2eUc28jBNtW8GtOluO/AW8kk39z31/NuFj52AQKvfLmS2zM5oSDmS/QH1
IEx9iMORzh3vOma1Ugo77YLxsv3OYikgGw8vLYxpicyAeDqN87d6gnTxsi9YyU9WgB+zBGcwwnVm
2wZ2G7qSxMfaAjPZJ1avPmx+K4xoWdKbPTkC1nc5Edgqf6hbrm68QJBlE7RAG8+r83N2LHZbC7QW
NZMlISAh9k1BAQQu7+uCguyYt2jhVZRdh7BYCSbX23QGIAAJlcZF0/VqwUiNU1efy3jfDo0NSMWD
43Wl1nuqHcNY79Ls9TICJpqqK2r0nqONVJh3d6+XKNhqdA1/lu/fSEJ1F9C92vlaeY3TbMlup4LX
S/nZjt+dguJz1ZkokMrg/c6XeD0NkkzIR17ISDbQs+g52YitzuDGR3uRsV3SH2yr6LvfGWAv4Nn7
9FrmS21SSmBL/KiYxmQYYIke1o1fucznH/cZRlfcCxLu4LX44fnGyRGjLxPdjJBA0gzYrjdS0Z0Z
UwBEdrqNYMH8telShO9I5agZeoZBMnQ2SXLrXFlkHy/KaBrjfhMbEM0DMX24XXmom1S+TZCDp4PR
EPZlgt1jImRuXU5taOsNwEtNLNz9Nlhl/bgvdSFIPlifHlxGBa5pKKLiVB2HhdUA+eYQmdoksVJS
taDHEDn2mi3qC5LeRqqqEnTSAuIJDgmpEkp1/u0ghb8DHVOk3Cx4/9ue3Pu88BdQbkDvYF474aUU
vn4PwwOleh0hgC2X+FgLhhQjfUec9Pb9evsR6UeA9ZiTI8yH/Wo6pouildgVRVXB5aJtLlC/gnvK
U1/nW/qOQr92LKHaPkDMKtekIDKorX7UU7Ma4jKzMjO2QqPXe6QI0B/rpNfPCpPwomWsZrmksvUI
a3cHKIziGofx0h2U3HjX9Rvb2Y2v9xZrGFu7rfDIeSCqARcXf7Ta5ftd9x0SQqoTIUtPJmKlA9k+
+2yqhxFSEQn1rZgfp4mghkHWF2+OSoUojezjHqv7xBh9xjeSt30WTA2L4CFcnPt6HWxnSls8oNhD
p9W+nENDDlJ+erETxo1/UZxLCzj4nb/2zsn5qWhiiibB1JqtnjVtwAQhw0JOEE2prj/I3LuUb3Op
jv13NzAEcIdnhmDPPF2WE7SZiDHU10uI77pTkfikv3aqX3n3Xbx6dZYIcsIKxsKvPy6s9Qo1eHAv
oDIJ4Mr/84nA67Rb66+QK44315GtIwEXZj8wTnheldown9rYUucVJkZFxnK4qS3b17bG1czesXrl
daZmTuRkL2GqRoakEb4eE/+ZNr+fV2BMK7gxxpNXwuzTSYtqQ99gXePj5+bRDBRDh27nJEZlDKLW
pfJE2Fp4xvYNZdai9w9paelrPTgsZ/riaFUxjDaVcMbHI+37a1MgVHevOpGodK5ljywPtNQZNIxt
lbCuDaIDOaQ5Rc8L5m/BReLeJ6sBw7F51YKJ7nHFt27k1NI0VMui+clQjIIsoSoN6wP8FOlrLG/L
uNTAh2mDbpL71dwqs1MIR0Znd4OXvVz28zhIVGGkCF3+ddgr7RwExntZiKalKdq1vsyMqeNVXn8Z
4PeXKuSre5kODfc219LmY0yKRByy72lpFt71ea9OJER4XjGl84MxSOcdmoKRBh0usa/HqhD3jCa5
sup7OgNXH7437LE4eOP/B6yHYWjyfj+Mauc7KYOSfNQMdaFR2oxpVefQqAwVDCpeNza1GDFIuLt6
/cTCnWfG8wfyBd2y4U4e/INW9npocBiwZMzVhX0nCizHIKO8ev14TD5i+vx8rl1TKMel+zgxBIVb
VUUMignwr3N2I0i/1gVFH/xpukAvMo3wQa7aeNAsDd4Awsq2NaRxWu6N4MnGwua72GnbyICNCcWU
47rsN856lYI825qS2PU7mj6ZuaRD5PHvTNKV1jHr2De6T7nmJ/wYZeto+ZPViUJJHv/H8QU0PcUy
HtXF4s1POupPtueiyYP0KokxgX/91aHIpJz3c379aWfGmCDPspxUZXc2sX53poTUsvvfIlx3Cd7j
GK5PB4vYcptJD1j6EeU281gvJhJyMtirZKEclxDnnsjDqGVgLo5j7dPQcH+WzOzquekfHSVXZUp4
D4YxzPr5XcxxwQ2Xoxz2FOe25aRWSEYQVPVNYDfnIN3xlTBih9QjOUzo0PbfuwDZoNUyuAUgpVsE
n/zDqGFaptGo7sgK6tAlF0q2Ed5J6vsg3NcZx8us1sUIK2pZGfyDvD7ikk4jqHWi2ajYAdbaOKUh
wunLOoIcsYxvcpXrYtRGsp/WU+MXlsntvOk6aipAh0Nko62QXYwGpN99MadspeY64xnCJ0uRlb7w
A2puwJMNuYaHVDPts9pTP7inzEkW1bipixsIYJfIowB0ISooabPADN6+pdNpaKP1P3uY4Yu56Yy0
qxck0qgSNVuoToEH1i87jpMIX9/dZwdEGiqUd9GrQ2KOShQBIeIGUKTQ28IgCwysSyw0h9Hu7zjC
Qj4wdOK6IlKzc4qAbbZnYP55KbMLolLHeJOBc+hTnfAvwOAxUkA++dmTfQKmM3qxGOjmUDrT/kBZ
crLkoYX96IpJQScuetdq+ZeaXBCub7tENlyGUaKWQfMGuRPCxDV0J1HtVph1wYwYVtXzfgtogTFT
M0F1A3QcPPiWM922E77iWnVfL+8Qxyr9GPflIO54o/GgjJJ/QaeR/0DYCqVnHJtofKDSCvl0//Rz
jXkRzigOnRKdD8uh97qu+tUZJjIgaY05LkVvpFewjA8nCmJ7ok7CzM4XkvQjV6Od/Pa9hODMXxv8
cUAA0VKuqt5/PpYQG3Yq1/oGw7RKHhCTAwlRr8acuUqNMDxJYUrRdPn7J4Bh9GcsnL6zlhiH5NAs
lSZEuUmJCT31qwlvB9/6jt/x+5Bq34QiMF2ArFkQ2QNQScOBnTWEb5z4S1e1ADeTUsEQR+NFv2xb
LSkGlpNgUn1NUv9Cmc1eiAtU12NRdUyLKmSxhvFgmaPB+M83vi04OYKGfhvJPAm2VMdW6T9VIGM7
FXUIRCWIV5jGejMzU2HaZ0Fk/FkBAF8KZgZdcrWQVEcc+2owmYknwU3Fr2ScBbNypXvNFTO2jyBJ
lyPcHbUQ5X/zGY2RzilvpCfl1IDEZDV3a3AfXrc3UDQmKrcG8kX49NZk/mdBi9FnlehdZAQT1Wma
/B60Y3lCZDyDsuVA08yv37T+Pyy0fPiIAulnfQqvwGMhQfc/FKQonZip5GvzBveTo/ToXDZ3uBO/
hHK5wbKa0Gi0Gny8kwbNb6HU/CBDtLZL8vYua+D0dbtmH2eRTmXkqXUPhm7vGBMvipiFuVnqY2aW
aGa62qepnzAfU0+KrC/2DFsieaBzbIQGiEv8IKy9aPOGwV4qXIcBppiuZGDPq+KsVg3I5GIhA6Ls
ATBDaaNuU4GWzThfadDwDhG3d/4+PdOU4bD7P4BxiwCanKV0YG6yhQWKW1p8WtZC+qWAArZPYIGO
VQ2+YNU0fhuCSHcCQERC9woxJyXlCfVhyg26MjrtrSnD/asHJ4uIgcpZRTr+LtslgdSrzFNQzB/H
TyWWiWbQkove+EdAvblv+H3WusrVG9j6vlLf5AFXbbQld5lyACwdeVgSFvbXGGmsSL0f9zVkcV1u
tYFo1qoavGEZf43C6LfGSBw/SesCSNlxxuY4athePuh+mUFlvH1y58M1v5fcd3S1svtHQr11AaPN
whJxncqz4+w5ZJr0K1GJqc9YfAu/9X/Gjd5ByP/7AWYCxmfgLMYA88R5P1uSffJXR2Jx7xb3LDcZ
KZmqJTh8dYH/GgUgdONcRcMRJ8D8kZGY0IVePZS7nq7JNZVAwYWFDPpbuOgM2ViuWPE+EqlOlbQ8
q4lTmX8v1n66nJ0Fa+MSwFYwZVrO8ymIGFRXJqjmYtkPKd+uDYqsuTZlwEsuR/lZnHsVvTQ/Eucp
Iv6e1mKyPidFja2z0D1XFg3vCsJlxnFNn4J+8e5f/Oo5Xbz0JqS0/RG9lSr4OxevuDzNUFcSlT61
AbnmhK9hsG7kxCLPDZQq6VlY5IGwJ+FeVOliw6YTIUm3XsMG+JpvolJO6b+ZV7Sr0AWML5ay/7Ev
eRR0JgFW9cndIiouZM8eccsK8LvFksz2U5CQCk5UIHfDIqSf8en1uVrBlYFLGc2SM/4Xv4M0KRLU
l6eliSVQEwqT8ZB0nYoHba3AWPqChpzXbSrKmzDzECoxEAT6F/aOcb0x1z5vNphpLBM+JvcMdI9f
HipPqw4LZ/eYpFLSDHsil/sXYmZw7PfIDiPtMj58kFtc0iVsvBrXyx5B3sOpCDqxlT9T0qCp/41B
RjNXt/SNacKtUhM7Q5p84C5G5MrJPJAWTxo4RBfvZ93mU90ioFS8ymWeSQ3iSJ1/2P9y+HCDlrJT
8YEOy7j5r5DG7mvG2zsh9ufsAs6MwAakJtcNfbDNQwNQDfg8mcmsAgMEVOdem8bMpgHrn50GtQRD
uuAaAhMyZw7sNnGcvUB0A3Z/GK40lY/iguhy+RoHc0m7+y4dWUvF8oRIwkABmJYUpqHmrjVYGTBG
KMuOB+YjCLphAVakxoCMN++zzBC47UWWaerZYIPY40jqZRGRL8fX0J337O6Sjn+MnZYGb8HQTIcd
OHOykk+0EBp4SQZ7vdFCc2vfTbtnnXiZr5dOLEmiIoNgsP5czuPZWUdMoKAwcFXyVXibiU43BewQ
V8JWjSBBqkcjQYNUpBZ7bTjDck9WhcKk/pw4SIFWpBQbcF0SR9YyAU9q5m8RwPD/CkHZl+jjYC/I
iMLIrcfT4gfAQY0RvhKuAfAlOzy9KhNokO1R+ytF9nbGYACMxW8XZNrqVYsjVA4KwscIiKnIUv5L
44I/NiXrWTXMB1vy2abZY4zZ1t3YyjpegUTvW+z2ifKD33H6QXytiRWUXbMkeVqdsnhXadd9AzPE
PorcM2hujiB95n8XIoPDCD4SzG6S08uZQZ+HFEgV9XoZ/nDE/2qbF8Wbtuog7daJGNDCub9EuIna
qKQJjX0JqJlH3R/h06SGV/PDzs2QhKMVe5iGSymxx3/FXzyxKEUrFR3kxXOV7k6ACJykH6rC8w1W
BdNXucwscYjn9VcPvTF5hahfdLQlZHlGGkSTZVplTxSPHaofQlcyj4N5vHekVo04Qzkx3P6EAa3L
mOIBtsFKzyU3n2pNGuVwjTxEomzEQFtCHY8ydGdVUNUQFj/PC2nAixeo3sg0Mcm0fUgaF5LpWu4a
IQVCIRMsGkfHRWcCO284zgAZoi9Oe3/krdF1/AqDPC1bzGIdl9o3Ng7iQCLxhGd8FXmJClvNfcHm
XTDVevqkPhR5M7NYlmNrel4MxzY5iJCFc8Q6iuYI61m8FHtujxGlTraTd9TUMyhW/L2GsotRoBBv
xD9zJwQhiJeKArNSacqFyk0e7Ift4ODzUY3+tTSPtzLQY6rCbEl1FH5wOIG7egaPRWfFz2lDUS3Q
f1tkzvsqr+8HgEK1m6NzNEhUq3k2uA3jo9pUuzDKLYq2V2RCqBEo+kPJTe7y1+uRWtuslgv+noTw
sS9/PuTVFm3Fzu/2cs4nshJCSJN6XAkXPDtQgS8bPUooGSM3QyOWZnaYlUm6iy1dzdA9VnjxGcgB
6Sf19ZRyAfI1okk7uxwZhZuEx5hWK0B+c1E4MJwPXfxK2cLHYsOOGjaElOqVrzbxEl2A5fiwJQeY
HWVGESI7PxYbXMMpZwtq4mM5P4Rcbcl7398ZCczIhoX9+8mSJBt/rF20JtP4BvnOxuvFkhQQo2OB
gf3XPDytFTOErEUBVa26OwiqOehq0HQhriZ1nFG0eqAeBOo8V65G4iKpQZ73A1ROERdA6b/j6MPi
FUETKuJcOfUVjkqhwvPbu3weaCmFYXo/VOBVX6+u9U/BwkJMmA9Bsjg1faibjrC2+kJbgtb+TbUY
bmDQo9m2yrniKhECYyStbFjQa5lCuvFABTChPil2j0VIV0KjfKrfMbMzV9h1/4Cz5ROWpiu6+7Pc
+R4E1fcpebtDY5qlFs8NBlnJF2Zyw74OoX8rzgmm1SYWl8Lj/0Dykk6wkj1ldWQhPQeljbSMpy7h
UZYnF9FuwQ+32Lmpnh9Edx49/nAsx0//BKdkYjGMOvnr/2xKvGbGlYKN9shp/mTywMdlO+V46bVn
+m1pJAE7kmWUeDo7RUrv/Q8saSF2quSLMQfNbfPlWO9YI7AB1yHkA0CS9stPaelB/cUg+2eqjGUT
M7YfJ4jiNlEkjUxG/jPVtyBnuRiBxJXrNEbZ88Nd7M/LS+x3zYGH7emcKFbD+G54/hj+6UkszWYI
ti/KG7/gRRW9QjOwCIM5U/dj3sAWdLMJUhQcT7PJ6Ze20THLZR99CqZk7uCgnFLVtD8DgtGp+GYR
GqBJ9gRXF6oCkuR+2frMfqf87n5+PRhxi7KWDGoAIjFUGqvAZtZfySMktvbTPedvEZxlaNkLCj8L
sZz6YD6DJQ/RBGs73clDrterhj+HEe/4ylK3tGn53zJOqwB8eiPDhI10lbx3xMHDPb9KFPrEqdhp
oo71Na2RjweIvrsglJ8j1SStPDFsULxBSxlbrXCJwlzdyaA1M4Bh5vYxLs1Lrz96WJ+qVUfvLFe0
AgG56OCC+N6ojEqEk05rlKjXXEnfZob25RmWCsHLexnI5BDmbZEx/kxF4Rfv7nCwMeMRQP1+sXO1
hdyH4ac8s5GK6cZ5Z5QZqBz1t/UhBxuG5o5Cj303KGaaPindZlQc62Euv7hJp2eWW0lIAHZWabvS
mu03GQ+XFdHiVGKnBo3U6666hD5JFWNi5mxCi4Rvr7Ifp3y5CYcFR7G/95KZResO1GJ4qbImMIsK
37xrSxMgjHcoyrYdU8KzEbrnSElcWkmeCdO/1MPfqhM2PGGrpXL2udq7ty93UmpFtGa1JcjbeGUy
HXT9wAD4+5n2gVyeGMeDqk1EVSzb8HeH28CWgdyUuFgD6D/kMKBhhyjBKt0O/mKnmtlNfMfcAJS6
GZFI2+0/y78T4gXGmoUzrWIPJ23E3O5mL5TOfLpPAO7zcuhElG9OJMjRp66EPWJkDZdEh4F5hHAD
GfygYh9v8LHlXy37WRYyX2FKTn2LH20eBstUxOzfBls58bkqG+nJZDsWx4eKJIpDgOPqnJyc1SRp
RbDlrfrHlRIgJcM55DnNkLeo1FMocIvd/aMMBMALREVMvFzD2s0F2kyoiOYKihX/1IMelTyKTaTG
Z4ioyQkferCl1Q5YWCiPuBs9n8h6dblid3PFruHTeH3RyJO5L4ZNqh8IbUQD4fEX1Ir1r9HduUZB
PHYF01OZZLS+VYz6invdHK8RQbuj+O5VobsWoaBl5lFoI88aviG7E59YMIoyKhI6wnRJ7GMvSVNK
V99HCZvliwKGd6vaN7ZgjoRo4BCVUdeBfYz37l68nWPay9v/zb+S3JqfKLPdKfPuA6ptGFvvM9Ds
rKeZBwYmss97x70YSfzCFcPZULVvggqki5UTwKNb6zWSXW4lJPuJI4vIE+a2sjsGudrCVMwe4QwN
n3IZrzhVmB4ozBn+vWeoisObzred+JG3rpzaKZ808CxFR2+cSygUdyX+uNG7LcgqkuffxSkXujLE
N/2dfeM4pDyNO1vFIEnSmFCt+Sx9+37LV1/kO52psy2zoAQEWmYVMa3lOGTN+OD2SL/CDBQb4Dos
3FY+iVzjbkxnuJepKCh/M6fRSmThekVnYAvusXkjmrpjrhqKdm2f9o4s2XGL9e2qa7HoV8PEkWxn
h366DGVIZkwT1ZVtbv4xOs9sHkuWHxhBXjcBRg5QGUk9fFZiH0yDZ3Zia5QeFZtqR7sF1LvJx5vg
q9+IW29UmiAvnwIZHxnJPsAXWXu1W80qqhPmFdIZTkD3gOde+6e350LHfeiHTkK6lPa1YdrBGZk5
U43fPJPbVjZ+dw6wE7V+T7LqTLnsTUzfdI1TwxTJoSc/RcFbMHFkAF9CkPkFZPdwlSKX2AdF/Vd4
Toy0Bk7Dph/gO1IlCbIWWDrjH1sKvrmCx3LtjQYNmmH4Q8VbzHJwnhJWx5aVKuTc2lsEGa42j0pF
tXxz1RalwW/dz/eRYDNlT8i+o39bTSCwTiv3wP28CPNpdhHWTpzmEg3H2r5WE1P6g3mzZMTzzXl8
yRZ/AAiv+T6rlAJ95j3X1lnluoGCKngNtdvqgIfgE3IVNyho+lV34k+Py/Ogx9dupXdQe1mE7lGB
WiG3uygvABDS8XxzaS9OqVDIJCqUiu3Tiz+egKVArVWpGCwLqhJEDUchA0HmBE3mn3LPZNronTby
yG4g1WE9Ral6Ia7uNcS2jD5MYRfF6p2JQStm2KcQ0l3YJV5tJzhVuytBesr0WzHSVPJtUa2wvjNH
4iRveyyeB8l3eNc+1kjM4VC91Ff83zOoOMJmGlskc58cNbXMwKUjKfBTOt1DdDtsFp5/RlfVvIsK
2LiK5RwQ27WaDwGXFqRckkUhE6h/NhpAMCVr6WDb2ZN61UjmEh2/xbkYZkn+ql3pXHHOIxmHSjwi
sc9bnrE407gooyZkjtXYaFygc+rm6qGM4jSayrBfJN8dfy2Xt6aIUQlzGIms3lZ0GN+Z6ST9Qdfg
BW5JAs/7ShG+q96FEJrlZ/8S3lcOR6sBIB04oBsS1brBua2bADupfHWvpJWafh69lc+XTnVFkmto
RBXOCKMpO8FcxyjckonnFmu2BcSiGBaqMwMIET4wBnJ8iTIsfdfh15AcCv+GmFIj3Eoy7cSfhGR6
DS8a2BnnGoDsGXziIaMgdHLvQWdOe/F9fxOOq1WYh3UgQCYQ5WAUSHLNspkgKlxBrid5cjOqvjV7
lFUi5ch0SF4DNehlHh/0kd1HM9OGMWA3YoTy9QxDvEtm8MvVZMIeIwnq+I9efYKHbasN7sN1UWEr
I5FoH4Jf02f8CyqVjwfIm8mUYJSSdIuBJIbY3en5Uiar5EqkOHjaDYydZpaPH0TrLQdAfyavvoPx
Ju6Pe+NkaxOMsMWqY+sTHKe3O4ikqrMmjVSqjmZ6TDsrh8hjBW4wyaSVD7ccHE5DWRqBunEPLlOP
DDt/TURyHkx+hsrishFGbgkgOxZ0dInDxq8lRbApBI+KwgvSc0wjPamvwsIArwlfywH+lmrOAjZz
hxf2K517mIdbVTsdjt5EafvJptJV4w7IBoC9zNi1ARNJ9+PGbs11ZSjU3sxR2mqi5XFV1SH63Oen
E2+fsfos7S8H6fTlXQoLbohmOyh3NSv/bMvkUP9w12g8+RIXNZmuBxxybJ1YJ316dUwpuNJFOQeJ
/ZFUYnLw7HfFowe17H/wHMZnAjOfGWFj3+UioldrZycz7vhhB+hKFidTzKwznFG80VeIe+HiIVFV
YoAH1sX41aNSkCcqTyOwZYCUI9kCoRU6aHyVKCVtSowWjgXQuXEkmWYOxjy3faPvjn4RX6vIu/ZB
7WIbPD4AMlfOOaDNoZezpG9+PEpLOj5w+J8IBDSkaDAG1T6dvp+5HcB5NIRWGvX47SVY+sV5M0p4
n5SJ9VxLOp64ZCX721qrFUfQEuiJg2AvT0dGL28hNcS4AyagBiUfYipEmYiW87U+VhE33+oa7zcv
Fgz5ljXjDbgGq9N88U4oXMG7p1q4Crb/v9Tnq1DNZdBxxt4LZUtY4ufF4pPES6lJXrjY0tDpFA/W
L3A07v2rv2DZ3JRRmG1yy9Q31uTYKjk+7isZMohCQclOIHiuSPOGYmHUOwbD9OXknmZAb40lBD+E
8eab38Uxv7hreDBDLn3XhR9+JvPcPjpcN2dV6vWx/6hB+b2zeKvkKYszcsTvE0cH8JCuRG0pss4g
1orduEsUtunvLHJE6L5l3/1VUUMEbh66XyRTozcxdASyePq2VAtJlr/Ia+sqkoX5jZuR4A0wI0Ed
9VQgQflBh0/9EsLAFggqTztHs0ov8ex6OmCIIhlpwwV70gVF6e3jP/Y7PniPetXWmvlk8y4USKc+
8evk4m37T5cR7q0hluhxQ3KXeUEiJ1ECqsxjIPxVeEkHbWGTQfcrVXQOFbTgwBI6Onv8LoPYI1Qi
7U61RUya/LZ3gqQv4yXvlJZtqGscyJrJrxkSeRdtfPqk7EA36d9/yPuOAa8htUzQvY8z1dlI+pzT
sbHyNtXMhzFHUQKsg2QjrmyP+x3NbIA79gTh+6dmeFALfBHMueBnayExbf1VmifylGn7wSf2mDFI
UxLVloJRQr99N+tVxn7w2ciIPvykspjRkHG8/QP2mrmrFGbFqxifBlGdjpC/Y23lzf8v/2z3/Nwn
LHLX1fwEXajEn0JtioN2fP7yN9d/oM4JmHGB1Rl4bX1qksqdNOpgMVfgC8MXNS/0WCT+qzrQEDpw
q9LKkjj2wCYoVq59P9bM/VydRjA0Bn2ham4PVCvm+prXtafXOfmgKKtCcUIC+YqL2MOOOlJtbVfO
xjTG4+FIzFdkQQdTHvIn0Ah94XPQEZtBRofW9yO0Ezww/Iw4M1bMLCqr6VIAeiQWfI3/tQqQ0UA7
fAGnkBnJjQpPNCVKBwELbb3dx2GxlUJrY8Y9GLgOwQyXPyLuc+HRXK/L1N18R5ua2PD8zZBblzkt
SImDR74mqARAZy3Vw2qcXszpnYx5aoCqvgb3LD1DO4PG7ykmz8dcA5KSDq8J/+Rvh91Lg1XpDYeh
hwCNjhwRwoOFt3ExKiYc6cJL/ep6TiauZzbnpqCdT/lxkXZQ/eH++C79Xe3ngGr4rjhabwYwZ7jE
/p6NEMkGFXBjy2VeFjgISrVU6lUrfBpDKaWxTyoDI2ZNCZg87C0ZyAiV5vTeBIKri1BG5e0Bz3R1
jsU/scEdHHLRdhRW/zKNAE9AeAwySwWBt4wLmKs2GHPzWe1yT3SdosAWc5sgbOwLj5ecOGxijY4I
VuiPD61HGWKkrcVKzt151rFRF+dtmQ42Ib0vX7eg6S5Yq2ZJqZXADtg5DnBXj2W9YrlB9RxtkyQr
NX9TYIEo/RaMmw6uLTBKzDRlZ73a3RvCEMMwqZOnnFQAOgnjnTh3KIx3Q8iud7YErMCQ2Or7c5KX
wo8YvCZv/SP5kyEFFun9D5AZvzIIN9dLe2oi6vpJp7B3Q8iMFOKi9eZ6veXdwWV2D0KZNmsJ5cn6
0/xO49G+704P501bavmOLAw8oq0nXbd0P80zSuwtd97MgbbAVZWqoE4BVukBed3ohDt44xD9M98t
Lef3JMpS33jHO0vRC2Zl47hUHTGLFiwSsQzNmGVojQKO/3L/gCe318LKvy/TdlTKgk3kYUHWJqQm
1zn2R1yi1hYp0EUjVnca3+BXlxRRUja1w0SfnJgsL4X0yErC6G+wDlW5cVTLWWeH/6+emR0FhOAZ
/3rsiOlXFtNX/7U12Vmek4/aTJvhYbfNhaLPdM1It25+BMCpuCA8KNMT6M5swXfwiUY2tKvpf3dw
lQh9ZjEbsVqVHqrK3GznyjueHAur8ct7qU1J1dOc95OjtZP4CHxCFiBnL4NZKFOhN4QALFPI0a+n
GYHuVzyQjb2hdhi/0ZusbQOCttMvNsjCtSGmt2hfD5eP51oGl6n9YPA+hsF0TEh/RgHwG4LXCUFr
FPmzRHdFBhY2mQ/s9nSLO3oSwiXL2DZ/Yj6IhosMrDVQv8uYcZdzVRTqS+prnlKapzfbPNIXIpLW
CLMty7iXTTKE77HxL3j7bfayW6DvzmXqMARr5tY7zOoOgvWv9meb62PMjTQbDsue2/PzihBnDOE7
QNDIJ3C3BFyIFO8wHGnDfyeAyopLMW36CxLTd2dH5J4C3rHGAexQO68bsyyxNsRA3LJlqZ82lp+c
KgyxWh/Qp5mR8+F/Btu6hco8hPl638OM6o8hUtj7U+R+clzQDwUWuWNDxiRUYqmrjYoTYmyhxYU3
om5d8ceU3PtoyEWLtSaP4g4ZFujoPgbCHD7RZvLxyvfidUtUu/J3CLiuBbRsYM54058FwyjwAY/l
OQ6RE7mwR0H3k0UYGGCtQat+hzRCzQUWUz6vIDtcR4NjLcPfHnYdCLfnQermrqDevBlS0XYxByza
+fd+UGl301S+hOW8hDmfzQJNS7UGN2G34JGEllCyw5EdPFFPZyggYqIR4NGbmsRuFlPSbKDL5M+n
RIQojIZANFTIjLo1VhlIXqm/ypklyXPQzsGgvIaWpbvQkWJWRm2lv//9HJfZCIfapnei9/vSWH4v
ZT+qdaVGUYFYu6XAlGk0xUvp8hLy+JhjfODk8GjKTQJi3a3g8QoYuw/Wcrz581UA6JkdofMG1Rlc
+oJOes4IxVMPtyCcp3EmdikoHAZtScWPX85VM39KYucq3ILHc5EBrnUXY37PulG7Jqofp4s4S5ck
WSaXPDbhqqmsEwvuAFRnkqVtWraxVKndDXCgCYn1mKPow9xTN2SixKnec9feLXNIj1oPAWJNrsl+
lNYQn0gl53g4RNuOXa2j4oZfyhSh+R/2al8fKaHKxXdiYinkU5NtpPE7UAwn/Eu5kM1NYfD4UcPp
X3CKmwBpsu5sLO6k66F0Lh+6ZEOcW0UJnWx3TY3VlQSSOYCviBMsm9XItmEDbmKh1ZhAq1L17djI
EEEH8gQOqZYL6w/11fL7zt7PxnrmDDPKbrzYlRjHi4BZTSSaoMuqh0NBt7xiFldscJc/Ls0opM6u
mG2Oa4Xta/BAOiiLtg8GqJrlTklBqvZGSYFQ2i7sQWnQ42OfobS624Xmbs69vP8qfaU1NjSO0kLU
/l8iUV+NejtLzE4Ife+z60dvPBbmarWZF9UJVy4paPYisZykKjpFekXqwFlQ7LAohl3T8NcWNX4W
iYmcpjG24KmwMKedSHjn/WMq+VEYXnl0rEfAmaJAxQADMussdBi71fr8JMOZZ7GBvmaMyk6YpA78
epvX7+XG+/gr/w8IiMFivTMnybm3baPOhy8kubihkTUwRzB/zKs5+/pE/D+YdZNmbqorQgZHwLsU
JQxgo6B8UFaL8TVOGb8zwm8uoA/Ov3FaQoCziVtK0OBdA3j7ESXvyBJNcBMJBSuw4lYRB7of4UTl
bGLF4f0+XAJOf9iBN5/CXLZmpZA7/ncifj4DC7YWGDydPLapbIGCWFJDyBaLDhtx3+C0dLtcTgRo
Z1rKZsX70Qm1rtbIrksDuZBlE8/lljjrIYjvsgJcLCbZ1TSpuOiQs0sDjvqfGR2jh5HnAWsBCLFS
6DqzRb2FUXhUXu++ACUihmvoZzZ13iO2rEn8ClLb6rXHKEdh5WyQbDPkm41tQoowp/1WOXL1sVD1
epVS0PIsMmUoptg5QoQdj3+S1Cc+3C/fysvwkmID4Mf86ehVKX7NGnk+PFCO/0/yCstv+TIjitSh
P4NKquMgs5j2FiHve+sgQLVfJAWF95wiDrTQ+ILRv1bmTACTrqn4toeevrTp2hSXbqRh0D08RB2m
okZnEMF7Dk0SBy9y4UggtbbTb6xeDgq25+Ul8tsZkaY+F/94tUm5oEn/JXOBHCA1jwDCh+6MOSR6
BcsSZrL11Fw60GgX+YTmgFTG6kt7HHmCJJmN2Eyq3cPLWJFYG5YO3nFdHOsIYEC2KVJzSmFMzUdd
21bsuMe8YUTxAcvHjfs6/PT0W6rgCNCL5AIaZJu2PJM1rmcWHusAGNowReMj/SQQGlFeFAhuhf42
UFMRB8E9xoMDEMET29vkBTEbNUsFhg5WYGII1ED0zboX1ewXj5Ix+vY6RZJu8ChdOrMSk7/nyxcl
W9H4rzMCb5yQAaxjeSJ827dfw7USiuNdGzdUq4LoeofCeCiBU/cp9lz1xRXNQoFR+7FP/uxpuB19
nmsqfk6cnz383LktSirWZvjSk9HreEHXTipj5/rQBht09Kj5Cbl3VLBXIh70GxDIzCGmT0zjl4XR
Wia5ThouydKoOrRy1qxHYR8DO7Hww42YF6XLZPDF4OxdTcS6s0gzUwQuD5kd+bXptnmZicJnbonI
urTc6OgiMa4dQFWwDuX0lUiABb4M33KPQ2bo9SzF7QY15QWRTj7X16/ZzOXHnwihPoiprM7j/AE6
tJoluhPeNlWSkhMk2Xj/rhwpdVCeTgVIbG15/bvcQQr/rvrw9tfT0/mmdeugGyTK4HbW4VEXojQP
lOLfxAvYRRumD7UjCmE/lA1gTLK2Efbt8AqMKvVmpufQyUpeN6w7aHVclehK2XYx9ivMWbbgKhz9
C70bTAERpEUBg8xEeStXPoDKhGTomZ+9GbAL0q/B9USjlweMmaxYw/i53NcWBRTkt8r49sYs5tvz
njJrnDeatrOSV3hw5WRHUkxmej/FTWiKnD0C3CaB+zke5HvYrlrkd5g2TjTLzQk4dMXDvatq8lAU
Wqh7QdAHyVC541jCX6Rn/QgKuv1jRsPwIH9/72OY+gb7+GVZjMSziEBbV8q811fDc5dvfAHXaDJ8
ic8Jzrkr6px+wkf9XCQYNPpUwbWdVs0jQFT5AoUn+qHYMREFPrq/glZAJ6nqED10kAY2t6rHRT/O
b9PkK+WGOHwKg0xBzGLqqeaz824rpPpCydCTXFa8U8g0YcUhRUTAxjCt5pGueCDNxjYQECLqnaDn
yPAYtq0oZMH/wg785LCdqJYyjiupI4O6LKPGsNp/ULKbWu06feD/or3LXd2LqEJBS1XGLB10OBj+
XkbkUi2ckI9926rFbiBrGnXSw/bq5o2SMqwOhwNLu6XHoNkHBcZGYKzqHtw2Y7naVj6Ea7xvSYbR
vRdMUYrTb0ajH5K8n1bMwat8GSMgcA0IRv0lze0aOiNZK9uAcXc7Pk5DLbgKZup5hrJhxsx+L9Ld
FNyVL+NGA69ZL0PMMbBF/eBP0s3R1Mua3VcbJ5ZN/RhzgtwCh6PK7b2RlgvhVbJYs+eD6CCHJl5p
x76IigXqYmwpsWlNuueiZKYvsWutGNJc/MReSGUTSoivNqZ4PoxcUEotJRHEaYJL06kQ6z6HoLhh
er1K10B2QEtmPLbcWX8ENm8OuD9gw9Rsl9VbMzLenEY0EBF0XzG5KIGa9/knOlcxt0H2DYUbd9MN
T9VGp759aZefLjSVR6qwOJAmE0ADD3/fM5NwYudoDo7cfnpntcgxREocSmDdO5gDxXv3wSsLZSYy
oCNPvFalusqcQSVZYGkvintw4vJn5zinoTG8nLO+TGmO7E39p2kYw1Hcz2LmK7ft8wdH+eDj6ojh
RIfIWk5Dpph/aNt5NzvnAjvu2x/gRyKj5dmaak0X2NJMvIYK6JCepzhcsSa3muC5aVm68HB3CIDR
i72trD/tW+SxcL9Jxfi5QYSb+LRC0OF1o67I+lofinNZYSVtGeNh4zOiSYdrBJwDBAcbEttLB2+O
XXmQQeTX+0dPWcqZ9woU8E8uRrP4JZb0ymPW2sI6vjLv7UeCfTKn42OF7ilmn9T770Cj/gOnCr+2
exQfPEW+ctdZ0S0r5NpSMjdG2QXoQQqz4S3chgpFPPDcjQWPy1E5MQ+DUr/OZPsTAcrr83vikW7f
9LzlkEwUEF2Fa7oooJXUIxPNmxLZCn/H5k8FGwls8TlM1MlvU+zpeBZCnP20d8UyHFsw/qP56LV2
0g7r9s2Noeg7qfveF4zm6EGDPSR7sb+kp1Coq2wqSBjodFzuOjH/xr99DCukeMmDvv+5UaN2RqLX
Owxmc6XJeqSTV0uJA7C/9fjrS6ksy5KbxEadYV5pQxLlymo9RFczJiq0w7cmsrDXlNdoc84VIe48
a+tZtcTVm3D+QhhcnhGybkVOHSh1FezNBIo/4BLiqDYNDMiHMzu/VaOeRt8amNTqiA513M4UNsEP
egwUGo47pL/tQ738oQc8PGTH9JP7Rca2GKmm2GcUju6mP9w6cc2gV8++XoPp3dwx2ZUnAOtFOU6O
D1yYbmTZKkFsnGQK6U0vXw09UDwi+P13y2WFbKxMEpOuGlmm/fITdJtbevJkRoUjQcaCEk/fyPwb
OrX4gH1ASj93rrR+y4Q80NXgs9QvvkDXsuVC2+9/bFRS/aVI2+sIdIDm+I+CRIr5JzNvGoYMn0OX
quBr4JqX134Iefz1btVn+zm7Nk0TMhD3XpPUF3scFzdzmSx77Ukjx3z+sHEjUUXVoUu/ZsslE+f3
GdCms/P4a/VatKmZhQ2JpGrDdTNRtLzmrEirVpNT8spwzd1y06zF3EY0yjJCfeTUcPRvyVmNwvv8
Q5MaThQ/0OpJR0Hc8EdMK7iuoI19WuZSgG6gqHJALI4X/kaE5VKACuQLSah3oin4XvVq9hhzUS9f
jfPcnHqAci4FZrUwgnZEbQ8Ix56NvNcCHtEgCcFzrSCmIwONvBAdDgbbiQlEmPsSR5Y9f6q9Duqr
OhHqBS2+IEmml0LAZ6owsukgj5K54i472oc3SW3YG9nXtNovLkEMhF4B7CRRXYAuIP7lI0RiiiG1
2w9WaJUZe1oUdaQXpGuebwhZVyAvrvIpiCI87g9Br12tIDeqBydmiPAHr8IjZZz660of1KuMSPFZ
vY981lWKn8NXe8dsvnrxYTDT3S03b+heSeysGXVOWSyRY43CX0k5jTCUYLaZuGJSXosFUJ9vvJ/Q
EQcCLst/6oTDDxHWbNiEr280578Q2fxGA3eY4CQs1j8E063TlNvm4aOdAP9KyacXoVs8nVbU+OSe
cN9krt6uGO01f00An4M6lVNFRwWTHySihL6XLFijrP7DSZxj+QRVDgpzdSxqSXkz1vDcVSZtnMCb
ZgEzhYwZNA/jJVKCm+E167NTwXUh8jtDfIDn64xPb3aeKWerJFWJ2oT8PoesDzqzEwLTPeTtM5JM
3PWvqyFErHtx3qLBlCEwjiAJktVaVlHhDQXvMVi/htHvG/RhvY0xox3pzDrHK3koqrIej/vR+YPm
N2QkRFK1329wXRWggQZ6Miq7d4kVsbx6f8RaCB7LApiIX74XQgZP/I8sGDH8gCWN7TDorLErYKEJ
svY7Du6abIocvZs2pjXtzbHKVcagvWwQjRmgbLc0tY2Ja4mJDlZxpMOsHSAqrgHRfM6Ie/qOxAo7
RXSTxAm9UsPfPbeAYftJfvBKLPS4wEypL9W6ZkHRrMekck5rNmL84kppcFciZhFffEQSOjeTBHRU
+1Oicpe3LDj/jQ4WIQ6BjeCMPwPRLe/z5zK2nTfZNKQvCbEnQz+guWfI99K56pNoi/IjHvtvHpge
8QyBeaBcn+o9NiQOXZSdak9Mo66NZKgqx9V7ytSNzG29CJfRkL/UJMszqVVW257AR9kpKDmbrYKp
VuKRTNlR55CAPlJW+YRVwb4AdmCkop4SaNIqx7TAgn8ZNkzCk2W1PhcfIExVCe52DAiV3ZVad0KR
x9l8oM8MjpERXE2/8QdXBXvEMuWk+7l1fFTtDc5sGI1m21FzXzuhDoxXQJaeGcRKhycJzenOeO52
ohGDNsFgMe+Bg1KSnbICgKfHz5SjGw+wGQHb8IZ87g5GQz6GaoK84UxWHTFN4XgOcnqq7faivn7N
Ry71l8Irs4pxFM9+/4XGUb9LvL3FENRdRQ27adzenyz3X5WwRdaXZtgCmTOcPycAmm7piu6barNH
00Rm+cFeKZr7I/R+Ed6d/wxwBVCGcRLEL/gbrKm+lEzBKqcdvzHjyhzPM4al+JWZY1g60tD/gfAt
gJgwllUUBwEbv06vA6wsrbe7feD0qfvrRcxlfBRGH8fpSYG4EdW9tk8qreHGbX1fddWoE6d48LD6
G5Jp25C1drPdKnJdy0Gpv5akOWyZQeSrKczPF2B4kOZ6t+M0Q+mFlmI5fGqeBHEA+UNER2gmQK0t
PoC0ojmtg7rm80/YSc5eaQbVMpoQt4BL9VcZxhMv4otvLokeLEIr5qsd7QYHVVOooX7RwhlJKby+
dfwJeRBj4osn84J+izMFFt3r+nbCoK5drbIdP8oAJ3j6LU82lU8KqVVhArrocwwiIKqhzrq8e/WS
SbgnICaSzklAw69kcCY9XWRS8Vtfle4AFgo7VCbe9pWZtTEftFu99DnQIc0mjIAfSGF9SbabJ4N2
r5oaar5Z/vd+UVGYFLqIlWgt+SuTHu4vtZ0vn4oKKkYZn+Re1ypYpv29yyXoqDeWniZvK2a6Uy3E
YnaoxIdw3K91HOWc4Cagw9D5imWVCgkbqorVJ8tWvY19DB9ihMTWEJ8rm9OM0323g4iHbD4j7qvh
nHqKNt0i3BMbwQH7pRM5VXwx1RowL0hic2L93cDgZ2dfIeVxQ65M9bydMX4GW3HAqvWItxdylTJa
x4en/95o4fIOYYsv7gZ3bH55nHuc8f0CL7YApa++WIms8JLY7xjudg24RVzmAZP1aqxJklRT96mq
Og7ZrOJtnG0RZzHylJdCP4vHnSPtGJ4uzujEkdYGxRt+wrsmMJTNGsescTaIhjal+a/dgke60AKr
V290HICFxJE+ioQxIbEH6XEhTyjpoqDFvf2xwkByuUMzimymx1MJXCwDTo/zOThT6jJGHs6Ss3DX
J42KpbnqPd7Tm+oAbXHJouPUOQjgbVtC7sCUDri97IslP16/5WMM+e9gndcIW9olHbEY65R+GCBH
BwG/s2DSNvYHF0IHGZwBlAPHHvM0avIdYzb/upen1LEX3ZMMw2vuGCkdt1F5cM4RuxqlJX0NkHGQ
RYN2hHZQI38KrB5w7N42nKIZujOfa/pSkkVszgq+sqalYqhpoW63OSNyH/mXCHawZNywzx18FQHN
3KsdtTtVeFh1o0toLlAou5ncpwFBq1X8XLYjQnWBPccinTQEyDJusk+Xwm/h9Wa7zd4vJEgxsUB4
9Ry4sT3iUuA2+KtapKpSHsbK2Q/IUFjDW4ySD/aB1lXQteup8DjX9kDeW1UpuiAoOkXEIxNhNRj0
JCFkmKUN5ta6E1BMyt3XMEC00bW9U5ybH1nHFV4oLdUUN1FAfyl/YGPGGFlTVhQ5KDsP/2C+xstX
egRVrdwSvB82gd+lfHZRq/JnG+6yOOaN5dzM+unMYvFEmCde4Ppg7mpKC5r/eD54njTw6AGTc7tz
E+mQ21fNvQUD5b4t6iZxN/9usGquxTd40qdXXh/DIPNQcoxjlxQaMGOajg1XKWNs/XFe8To6iXon
64/67WeT5/v+njakRzs5aCxGe65ZsarVXaYly1CMxTonN9Wn5CHXGqDsv9IalmfIcxeIKzP49+1D
ojdxZRn9RvQNEYFjd/gogugGhzAmJxqFCUjx8fJpEzUL3psUw2EKG/SmdH9T5JOsPOf54CMS5QZA
CXKmU+3JxE1CAUXM0s2U6IgZV2RbWlzuPtPw8j5cmdJY4CBDLOM/oo3EtAeZDQNxwDR1XKpyv1Nr
kvnCVLRBnDmwcYROOWT3Bl4dIKtUc+/xi2VCe6uM5/+s5JkLiQbA9Fjg8g50XT+qowQX9H+qLYyP
XHUT/ugun1MdtusbBPYG2ocpoIZx5vvAKsZ67yuuz2xy5+usIkgIEK9ovpTmx+x20LiW+AGu1VYi
EQc19s2SAVCkPsg2Ad4ap/ZhhaexxYwBQQZyE13JsG3+vExoE2Zcej24LDCkP8dJFv2iVDM8CbiS
i9L+FTjLrxQEbbfNyNotmcmY8w7lCfOuH36IsdB7+N39jyD7iVw+TQsUqtNJQyWfynVyA+VzsRsQ
XY737TU59Nj977Fn5gOwvu+ZapxOfM9VEw4yh6LFtjsjoqyf8l6bSf8KtEpyKZuFR/WLb0stMHu8
zafa3KcpLlLkoHBJQ2kRrmtM7xP5rHJmLye5SM2OMhLhVD18qKvJZw1+hjqEpiKEZU0JfaCxnnAo
In4jhIokw5Y=
`protect end_protected
