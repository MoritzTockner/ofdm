-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i/6guCxaflbTsUnF/XKHIoRGtE20YUvorlG81PRFwkKmDVun+A/d3uxibcqatoAvsz4/nL7uw433
VqqlCxsk0In2jylMCymL/HS5M6M+SniR801loBBPvSuf8bq7h3oLlLD+2EUYqk32cvIXGUcy7w0E
H1xeo5KPUlux6sHBavTqu+ocamlnFtppt/ewc83d3h1gJD4RoiUmBByUAApm5jACqwQMuXIgQIIY
EgrY0q4OZFweyAHq6KepBQoWy/1bmNOyOzC8BugrvMf7KR8UljAnP6efFBBg7/yfpEJmJFqppvyi
yivYSo7R8R166uMAot/BwOyWwpHqi1CZ5JaC1g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
BYlpSMDhS6CVowC1PvyBc06Yv27aphlT4Ml+KrOQE+nOKchRO01ew8xrAWKpB1x7DCoSV9l85xoG
jwQUBle8JoNeKQlCkonK6Na84qUNp+Wt0L72WVsdrFSyobNqOqZlDZJrZGgYDcd4o6Wck2Q/3UtD
tDFRJvrZoircK+oZhPI3v9RdkRGppWnVZINRHeVp9uthbfI39iDYgg99S9t6ZxyLy2LbYD9hSbtd
PzjuhNUVbvk9GbdHKxoiyKE0r/XiVrCh0rnT/VHjAg47zvOowu7y/+LhOhIZgrUhD8YEHt454qOT
UiA9KwmoICAn9Atcj7X15ETdBO3fxEeUgcosLviFzCdUJX/h1UYq0YLhsjyXuA7WI9s/AHkZSOQF
8see58u3rpzTISckJT1O7UZBBm85FbgtSwY7XWky+m2FB7H/CC5Sn3lFmy48CRTcWReXlO+ugG6A
IsaKut5EgXVla0ePWkcmehrp2sQfv/MltNhWjymVuIY9rNieMFE1Ju4CBvs2mbXiZE5HmLunJClz
bjluBd2uuUtotfDO/UhyqjYignjWzcLL74E+C2brj3xMVYSTs2FA2u9xycSZllotnYSaQdfevjBW
0wkL6FOFSHABy3OlKHTgQCw85cj4JYyViQfqMIZGwayRLN5hiD/KUapos8v4jnxV97Md89koiL3j
TIKUcyQuCOz4gNedBZPiGWnXK1nlMgGFFCGP60axGU4QULaXvuCU2vVh1Yzh44ITalz/4u7xZO/g
sx8O2htC6AxRd2mjuHmbj9w0QQdnqDIrlRpBlxysOBYEAX8n0ZnNP/rphSScHkxDP9/KXVKUNTBE
2y+YKc1nsAybvPV8YpJvY1EP3D8Ny+UdW+BRQ4ttqpCCiZ653tTSVjBtA8VD2T/0zrekbbGZ5PAn
PrwYG3k07BwgK6MKzyGbtfytxV4yrODVhngRaftGRuhAoD0c5Yip/xqUiz31M5MdALpyvgK6nCMo
u+K2IBzqusgCJoXjWKO2WyAdLS6obliaKXyU0yLNqeuh9RuUwmP/tUNPk5F4mULmHERS+s7UEL4g
p25znFQsgLHaZOf9M4E0hKViAnKp2l1pG01i8OrH18oMw9men3Whfu3fnftcW8qoNbtfuHOmWwAb
8Kyq+ewVsCx5sycaSmqJAVDiuIBt+a7mt2rl1s545+MGrSS9uYXPUGk4X7ReldrnGgO9gkBPBVkg
u1MK8Tx3WqPTQ7o0e252W9w6SFshoGvk9zOtmPv87s1GaqjpXeZeUyhJvaoGMHJuBaRUVa5+5Qke
dwBiwtw5tF8iWlJw0vBY4OjQnRDeZjaOPbgBOHWaqz5P3PkHUuvXWAy+59YcONzv9kqsdRZgu2+X
XOENlD9gRWb5CrNZEx9uiAv4qUGHnKUoIkTijD7wFc22YaG0kfsZt7/prCwE0DK01Th849hhNTCq
wHaBQVbvsTsLcAg/RRnDrZY/ABg+cenbR4sAXd3C748aETjoQh/4LZjACoKvBWdMtgB9gbxnfoWF
W7jlkrR5BdsHNiMmkSJMoXZMSdy/x8Ws1C1A6Lr+eTWLrIXLFQHvQc9r3WUi+DXQsdayA/BevHg/
nUTcl4rPoI6oy+k0U1g+B/b1lopbdNNIcxkp4Sj514IKIWDC+X0TnJoX9v7h+snk+/ecYSmkTu46
Hk9HkK5H4Y+sTynudi8KaOZ5JANMRk4r5mHLcTAcH8giVP87ms9/BMgKff//Cq/t1HBYkFsXEc4W
t0cdd3b8vu9yGblSxu2qoYPZPqKb7HU2XtzVBGxlgf6Mz8wvoSUA1fnO32G17c9XHNdNKKBxltIf
qQPiGqPdhkPhXQ2GAZnWJYaXrPtsR95RIatarhFKxuCxvdNFzdG9TG7ugnbvXzMCgFp+bSLPN0SN
IIo3xk/YSsL9PrsO2j/ZATKCp5fyT2iqdGkvqyj6gb2Op+eXldJKFJWo83ckoG1cmEv/C2DXwy0/
ArSwrEDZexhE1jwO3aZ3bI43yWD4q4uk8deaSqrNWMIvNS9/Z5VoKeoE82YBHUauIprQuX8waJXz
MRycKLB7E6nZRvz692iLEBG3cmIoQ74ZAa5Rog8zBjSKE1grMmtgAEIiqhjw4gyVJv7Xwu7KbG++
Co6wH6543cTX4I4xF2MyxAKl+Np8NExKcAKCsMCap+yKhEpFTTsYM1miKFzYS8GqewHg/GrfZC3E
6sxVfLqL8wh2AS+3VwQRBA57NWehkPTibeQ8L0ZosokTeMu5rfaDvuxQtaRx0DAqItZlYmw7eBGR
Yd4Yh3WU1P9rbmWXLfhRqriIzC0+S3CE3edL5zH9zcusOZvwAbyf53lkmof8tKS15NEFX+qzk281
Uq3BkvpO8M3ChuadAkwpIDNciyhVqKGHBQyV1zXXE3vVxJ0lT66uFww5gpb8oOtY4c0ziAoVu6hU
yfwLwkBhdFrHLh3rp37pLY+8vt2SLMT7DFcbvF0bFDil/84utmKWgmihH7ag+0O76fSN/fdOOlxU
Hc+VBH+xUDIVECEFpll97mT1wGyqtDz5Cnn0scarwYAZhUzm4uN7e7/EAMBupZIf7CWc7U9sfEp2
0ZHhFp49dePl7nfaCn3Qeqdt4nStbUnuagvjx7TEyFlflGJUAHIJp1H/hPZwO0wU0XfB3miXUtvC
5Z/WMA8tgt6nndrp8ueufBGVRfFRtQO6dCg5GCsOSFqPrVrnz2kt84z1GCkh1JhTfw7kNf2Da9Eu
0vutQIGUC9XvjXLj7gmGmKDRix70mCnQp+8Iw1fnWA6vQVp9Ip55lU8DZV9BYeYh1NHczvwBNW1C
COVgHq8VR3Bdz8fRVD+stKlp0+nXvjzvAcNnypK7YrLmTlTVqmEoD3ZkYOsjv6uZyGKPbfhZ2Jaa
3FENAjgmsZYGk5/ak9YvvDc4kzZWuKPhMSUNoAoF2hnCfb+oSYUSsGMOspSj8v7o92xor7uuZEdM
JPU/UZJTIu2sJgHB2Ps5p7m0CIQrU0MFBvpOpgslraLIE1cUwNSyc6M3JTN0IQXHuYyJaANfINn/
QHfJAQwl1ZSMb47XcL79uawmo1zyplin9nYv+HL4hsYo5+/Z8yPkQoz6iTfTLQOcDBcQ5C7sT45J
aoeWgef2TyIORKb8O5xqN2d88ouP6VgYxlQKnn8uapDrYpVxmdZxXhtSjtsampdcJSyyXgrBX/cr
giDKYP58gz1ao4TGAqCxJBIl1j0zC2nd1TwYlD3JUwCAcnNKd/AZcx+IoBhQ/r7L0KhYrxRt8Oue
EGompJnvVez7Kbdo+mXYVRoDoE05DFHObhEy6v7bUzxNhZj//eSkYhB/7ZjzYz5hf0kgCkDxqOWM
pYZWbbI2jqMP/ilxHjgIJatGgYYkkOQipQe8Y7UuKfrfETmygT3sNc0qn48OneBuGz/ncalL1uMg
rFjsH9kHBavTvSH+xS6roDqW9QwiEMhVbY4PbjjsNN3lZ9HNT8OGo5AOXljRII63Q5N81q5Bn/KH
Drxksocx68cDBTzomeG9/YkHlHMk6KiHnXEz+KWSjqiJOyFrdbpT9iQK8Kvpr3Agl4wrKveAPn8O
qN7ZLfttT6O9S1+L8+AUlhhf9Bh8OaDqgZ5cFw7bZKlI7/9LSn6NEILa+GCkjcGvB5TPj5bgrP5Z
wLC3FUba2T46lO94S5hqFB3vNmlyyrkcoPcmMKXFdSt76Dckd5MDhpo+YCffosjad6lKfCe9dQSX
m7j9ct5IY9poscsoXtfUMuxgsEUsvGgLIlqMy5uOlVBYZ01N/XOYoHDounBpz1bg9Zsu0A52tkIi
NC/KqYkRHO7bP9YJeEqSscyjGbhnM2WbxkyxYuKYxkTbKiKCZ3SZ8Ua4SPJbLhqFp8lB4gWsLc7M
bSNtBOdmnfPN5Pe9mO1iBz1KHha3ZkAnB41i9Rd4ALC3rLG6wl8KfJbSBM01pvcws1BgdV3kVv+c
qGNvTuweb2H0kXH4JMIBWNx1zluB/kS4vE+V8MGwAD9yo1YYudOA7oMf+K8iALH/plL8bR7RB5zS
E7etmr6WNysKUvVKLU/EMgu6in3L38hqgiEuEDT05rPW9VeNk2OvdzG5w5fuNtK00ZD+E3T9z1qK
47/FDte9YRf4uZur7Iy1YxznJ9+eENuwAn6ZUpBMnj37KP7DwhBgW1MvC6lfeESYOmtej1/t4e4B
QV0VeeGAzhwwDlFTuzXdSYH3nZ9GITjEbn6deEjFUFEZpekih6DoYfoh3WOOVk/VNX5zxnUF6ufn
d61LH76jZmi+1D2bGZlh/pHHgEWQR+f6MkTt1EPWzern2LR6PrF4UbRlAurUfhx4b5P8lfeA5qj7
JTF0Y6hO2QR0t4FjCtb5p7+1jgG1zICoCtFZ4xLoS5VlrJGhbZzHcCsDCR3FRG7WAFd88Hi5zM74
eZ6kzV679QZGhNfQgKUOHdkDF0ODjZslkEqdyXqBnla5lw7SK0ZKhtI5ccPPK/mfaRkXOssvdgHF
57YL6OmFURdO6ja1LBWxVm2fm7POuTr5434tNYflcmIr2Riw4Y1QLRPVf6qNeFh9Mgv+nfr7w05A
Rnu59SZ+O3i7IrB7CsLpxdZ2RQYUS+wAsGUZE6MwPvNzoRUusaXyGcEJ/TgxR6qYs43z3CFsz7xP
7e7jpLknB6pLjzlwad8Q24xBaaV1MYBGg/j3Cen9MLD0NSH4M1KZqKiJbc6bGP38ltyxR7I8pFUz
USanC6ZmS1WBxvnutA3ob2lb5FApZQ+0aMQ1PzwgqTIZyA/+qyLWAwVxUy5ONmDKsQZj+AnmjK6F
Z8FhnqTItvINxNN573p8+e26WLm2w2Zrpf8RFXfSwXFks2enGmxsRRh4oJDh1cw5sX3kMtfY00VI
YbI42F1hWPwRt1YDXJBZQ0OEmke9YeZdutJtFSGT+mUdUGWtsLtGdphimks54qtHXOv6UGJ7lQXX
MvJrjjCAogU7Md5i6eVv/RSiV0OeCe/wdaINfNe3MxKSPP30PYIWh/wW8i85zWGCcE1qZdhNgOpe
iXBpjrzhF7H2lMjdfbQ2YctbZ6ryNMvJgG+56P9cJaqT9TJ6E6orVbRxFGhGAENxoRVj7W11Js0r
P3shqZsE1E7cKJ/boIVlINxDRpnB+NOh60C54iDpvdTkmgJ2YiC44UWc8EKk+sEy+1bTVv7C97K5
p+B5JqAbKThJiLsHKuBeU72mBrImL+opxzsF7BcaZxsYn2yh41epkG20107xZqVMnZWdexaVvsQQ
KhHFs/LJNz+uozvKsJp8YaA63rMoqhrfqXarMHZklrjkjHm5jlo+Lft1bWoUk/aGOSIZYZpUjlsY
bZHK0/TYYImsw/IKnZXCpf1TYegUiylNhqwirlmElvFamwgAfuXHXp/a2JF+RT4r86nu9SwfFS6u
Qcl/hnK4JUsuLOGg7UXfW8G/7tzW6hRimsdBqNXNpMnA7yDD5UMG9tX1uypjIW07jrJRzH/5o6dV
+pNHm0G4Som0TQEpvDvPYP8KDvI/2CO1lCYzsoklF7tcQEJSyIuNCoUNHTQn2kNNKrAps0jPazRE
kJZUfQuV83EOL8+Gf9Q0UFUDaAtWBLSy73uWI/brXY4V+ZLgg6w7JZXz7Kmey/jDM1NAMk7+OliH
gm57otTXswL9zWdvkxXRuYIovRPa8rLpQuJF2ELLDxWTvXTsFmNHGIg2LWj/2x10Vooan/p6Uizb
zbDi/6Hf/hzrgqRCeVNdm1X6DsdwiwP1QWgFd2UM5s/jFPDbk0Voody5u/TDnEMS13GBndO3FX/A
JKJV+Vo+P1Mjdj5u7FIOFVCKeUtTAS8CVkmyWzj0qUYQt9gOI0/8P3G8Ph6OKQVxVUVq9snXbBav
Z6oKJPaQ1ZdO/QuuOgSabPXpHgDX3L/cmKea2YvzJGUw/XEIKlMDvKwp9smL2rLOQX7/nPUYIppH
h6jjjBUifBIZKLnvKN+G1MNkiLSi37tgfJ4bEA/nZ22VH84D535rD4Bd+meCGvrOJB8KOGOqR2b6
0Wau8EgVe/pAXUsY8bI8YFiRFA1wpY2f3ql7M5pO6NTMkgA8NxldVLFVvts4s3n+VVWi4V4aE09W
kufLoTo1f2jN5qt+dKORDXw7xvcanN9h3stWDrhcbLFCwAssdxHN/l08rb0PvRA3emWoFlh0bILx
WzVYCq6AHKUlGT32SamQmUD8Lk7FVmAww3heZ53NQVai53QWNYD9haTs+ylLHxGKeEb8X0X1aXrC
KuTJGDNYwOaOUed75K2JkfLdMnz+AqR2G3msd4M8+QAuRfvu/qVKbmtQLh/ILQYKjScn4eA884Cy
Um3xags2NIrCXuowXX/pGLBpjSh6CNg20cf/kyJBwpnD04721Y/ODPa8P4dzV/nA2oHfQEvTaUfd
wOP1UWLi+atj/6dYpOMz6iw4Kee+Xro/1/a6qx73UJ9PZOB7hGAo/7N455A3DdU4ejaefk84QTZy
8C9r9XuOqUJNdZkK8Ih5F1s+AjYWzbocsOrXZd1WyydVehGeqJs+g9+ufx3Cs+n2sBoevnFOMcWn
XTZcqWvlc1wdPWPyKZfYpQXl87PrX9cmhtVCCDsNP7kTdiwf/rJfdbrfDwZVl8Ycb02sFpR2uYSa
0lPoG4BV+g1FN67eofcZgqdG/ExJWgTIlODy2Xas7hsJ3rkIcjFYmosFfGAZmHYsz/p3YRzJl9x3
ODSkmgq0wemg0H5D4qv/Oxx4YQqMb8vEZsV6ave4UaDSEzqoAUjtj0OkNtSvDfdOgT6REINzpKzN
w6FMWo3hoWIQ3s07S7a4i/sMT0ZTSH6ZezXGkFm0+eIJUDlN0/9gKxnHma8E993hYw2jsVnL2ePw
9lZ1q5Wn2kytzEFhcf1o6j4E0HCD37UdaRjR+P3EGZNP4PzcpeNYlvs/uhD0jnIqB43dlO6vaZhy
1lNYV3cmwjlnFarmqbPDXeWkdxDQCZLkVrXY+AR/3LlaToBs5dy4VhrRftDVTBeZRpxvMEwADxLq
FSz6F2IpAn84CI4sF0V4OCyP1cUivTdr38OjGvwGh8hu1jbtU6hjSYvznG/6ShATe5IFU/GWYJoS
9pjrygIy4vbnSsVi3qGm2UjPpOLptw/Hicz9RaIPHhokPUZokGBjlHIIDKke7Gz2nRV65m///r+5
O7uZFDBOkcMHpbMbpgl72Gqyf0mvP1dIDZX68XKJKdKoa9I1nSE8X45R5URq6hnL5KyfQC80s8Jz
4X4lZ1ba1m9Y6wcOaAOrZ895g1D0jVzZQ2kSXyypvwQ0/DeXHc9TMgA2E1CV8J8XwO2xMqAgd7vP
eVy/m1dc9gr6PMo168RjLWz0wRXjaedVLZ+cj7r0WSe/eraLH7RutgvOLAmHnZxfAvwAE70P0ptI
VDujTqvnN74GZw/wQfeOhiyo/oOAPD9rZoS9UUd5obAf7FQHokN8TwLFcQPHV+JhqwxNNGKXx83Y
jVzem2ZO2ljH3JUETxTluZ8lUc/U9bcqEu6Fo4nGFZn7PeCvlUbDAZlU8s51SD+XN7yXVhxNgtox
NMYHUYJoGsmmbDlfabGLMKK6rnfo/n3PYCbVZ7SNrOyrGM+oXNVqouBvC2JmLAOxXicBjfc3Psdq
lGzKD4gSv/R9UCYVHJUMNAwkQguie3wZcW90ha+1ZmNllOAq6kit35h5ItzrclZZTM2n8k1Uaucc
Y2H+ZHaoqLxnFOC+wdNjUPjrccPuRIqGioP9G5KLyAvfOVsmWsILJladtvZhKGgIuXDL9kJEe8bV
KyfNIb7MjK7Yarq+gregXupdUcmUEaU9FfC3q5mm7jqS0w2tkN7zdz0+Ipga8unXeyez0suHaw5c
vTz0EGKAtgcKj4tqUYxx1bwVciK0kkwq9z7Qlg4XSFjPmg/Tv9L97iIT8HSJN3qyVT42Bdh9cZOg
wy5tcsXuZy5nIjebbVM6RErJBdg9DCmoN9vpLamLNP7wEHFc/4z6p/iYHSx+e2qUqPv2KJRVmhsW
311OjYwjfJafpgKcOm3lfOtfYnqx4E/Bu+LUUi5UC13zzCnTGomZqre/8O/bDoJn3D7+yWK2An3x
XHjy/7QstweDLUbv6CS7fAhqQr37mAwWAYyePpfQcasv/nff+w55+jNqsxsr/DIFMGjkPUUIlUJf
0SPrQB65PbqdB1aHRrUpeyfiuCbl+CXrMmrILTzRUNKpmWFu8ouivrRdfjiGEf74sqVPXUK046f4
URBA1qNmdh0dEgDBlNgI+7kpDLWz4S0McuMsSST2PECnhmoN612jAyClVmcRVIvzpLGYdGh0xUjt
4KecQbf4/Rok0OIzlqwe8JvG6eoqHIqFqYIi51bOTpeYZuXDuQFbCfneIa0YQ4dBgvLazrcNtpc/
xPXcAs5DmDmyvrKih323E3L4BWeuL9Xy9BF1NzX9R4KwV4VPHz/1/zug4kfhaiBYSSngan8VqWGC
nKiDOCx9gWsDOGU1YSRsFuJTndGyNDtfuIC6tLyf7PUp2lwBZ5i2gsDOEWwPpDY/l9NF5nKS/0GW
WuTGbEj/27ewu/MjEA2xrtK1Jg6ExkGhnaUtLIN9qM16vPZjyTGoBIKLYZMuyKhL+yn1UWQUL2GF
Dfbd3cU9JDvJgruFeBIK8CMOiNSFiN8uxalsVjzU98EeRNCVyu0YuiBU8K1jP/xZDI97RBN+onvA
Sz2sUjf4dDzWYip3wN+GegOXlw9nDuLYzNeQAUMRI+4+CWxmKlcOrZt4waWj1OuZPo/d9xhuKIB6
Yi1SgGcVmDjxT0lofVPpmWxvy7cc9ciVYyEetbVAblMwNuzjQgZl7TgxAfnuHJ7S6rzEzE7kE+sb
x2sjx+ciDN4T3oLUsUleZIX+jDEWOwTSWp/qc85HsAJ0zQmkls086O82v1PYE4DXFlSxlcwlVbJ0
51GWZni6oiG2uaX/E9kJLZIda6ww4er8B4h6armSaIbn/SjyqLjSC5CyfC2qL7pFz+EVVZxpw8hf
eSov5J64ETvIByWb4KxmY0ttv2lO3sNwBFs06JMjppQl6B76tcRhSahdSGFhRt8kgyN7F7W9HT8Y
WuC45Uty3hs56PgdXg78UUzEO+UEY8e4i8i40qCKl2yxfWNo2WEpjrXRgLOQJ1ujRspZ4zVdjCj9
2GYkoQdouE0uJy1pjUT8Ow1NWNVb51zwn6WdlH4ukbzOcFLDULzRj9OFopT/moXcJGLKmXXtHgbE
TG8nObtFAC5ucfggGuQ0gw9Hi1L1wzbMYV4Ov5CEzTQ4156wkaYM6bSJg1iEH1XrUwLM6+ac34Yp
FDrnkPdEr5c3HMDY0fFMxcUX3WcFljtR76HgWqfOHEaQAcOVWm66VI94OL70UQv/MMuabVnq/sqv
RIER/xI0AV/y64zrAy9mqBQA/QJCwtU4HmjmPYJYeCyKXlZDBDwfM7Ye7m1/tFuALCsTwjgeNNHH
XlqUn7KzI7cuRFwHpPj+mgZ4VSLTlBbJf27lZM1ADl/z7Sg4XghfmybXbT09TMwuIlZYFB00X+Y6
tfsnr276qtZ4UPnFA5a6Z66TF5FPo2DsOwL3rPlkqjZF92Ksfn+CUMNPzr/zxHN1ubKgObnEedfy
NM6ddZYZKKFzrsqOvBD5ixUM1IPQ6BcmcPg57OSOc9K/fs1zswwSvN/cva18A+yfBL2v43pVMVZl
KhgYg83RryenOXyk+uLTCcR5giH5Qi+fS3s7KBFU2kN097Ij8zgac8h0viZWr7N9+8skxWa1pyxu
lEQiM1FnjH0MXB2/8RhCzJIwRrAygxFzxObmqYZ9lG/AdjKKfP2nvXapgFKuU/tzkbTQ+8H6aWm8
iA5b7fCUKGgeprDdTYIZ32Gau1RTLydF/F9s3z0GRybolBQXRDW8zOXd6WhmyoLBxXEXlIWTTDWA
LSvlVw4gqMShRDC4jYP9qbjI84gnpJuoNGMIj7MPVd7YtingAU0ZzNSuI0HQIF61vVnMjBAUnd+P
40bVxo25SEowl9V9mz0dZRU8yi08tDgvXnsT3OLAKr834wLgxlMFeiFwpjd7i8Pc6LMvrpsGXjj4
wQdYGO4ADwRrDYYnBGOK8GqWx/oXWLAvT5JDvja+1httAGcdcoGQsEaqk/OaNF5EoNt+F38Zqmh4
kFjgeZr05qSRyv71kEDH+dIVyxQ6g+2kKZhPTnGCEamI4jewSSueVPx95DnC2u9W5rLgWqnj2M+P
9909aQzDzPaYy3rfb9zqLtB0zI6MEHAFTntZ8aPo2kGSmpjqYP4w5qskYhIgtsSFRevNqR2od2B8
5uyBv7RBSBNy5reEimKnMGFlgu0aWfdt8/sSJwmfDoo4wZ3j6ZBZdn2HMmNSYAor4rhLuDxtSH+c
qj8axK2JIOe1KZGsciTi8d6rzzeKLK9LF0V2TrqoF/sh8Bcqa4rSr9iBlVGunxeMSTMT+UC7Lcxe
Cgro3/3D20VNAN4Wv/5VGXdVfi7h21r5n3ZHPCI2auTqGCnsUkQiHL5DIAfP1K2kCfL3Nqwy+LKK
+FZTrt63kCpkKFeDH0KNXq5xD3BzzunbL3XJmXz95xEfoZLtrSYqKfOdr6Wue03Eqa0Oob1lP3ve
YNn0w/oMuFSjg/5YNhv78OxeK5uieRxsvyx7Dpw8Cknsaqvu9CJsK0A9Pkz3T4A3+A/MqHwh72oW
NqCvjsXouam9zw0sUbVWq1i4S2wZKzp7rlKh8jRGUoxBtvjbBwWxvvHQCnW9Z+htvLHyIoIawP71
MdkVxpliNMUB7sra0Fnbm4stFmoKl/2gHwqWUV14kwnuCUz5uaRl6UTZrBe+X4sQlVnJABRV9Vud
b+9lOt3fEEdMwEQjGuXJvqZ7ryrV3r5I7RuFoF4mFLu2JPW8ZmrF14jX68WVCKSSYEtN/pgeypm9
uuQCFrDi5XAvulTPnXVtE+ZFTY6jFYRJTqG9KmNQEZ/UQ+z2JmvCYy5TxRtxH69OpSXyZLlKXIFW
huSJKWMuYweVuqtCbF+YGyr/bbXR1WmhaiMcgUmhKBSbuQzpX5RuNv3O643E2XwVvwxKxUr4VQ5/
VhW4ErVekqgku+uJf4XhDAzvDDq6K/sr+u4mJFfFSs2FameuoKgfa+aJlarmHonAYLcFf5eqpNvD
UUTuVamPAqcoxIPMf5EHS7DvlYDyh0ikezY5P8bRw/eDiuZe169ZHjHx9xhXIdMM+a4RLpqwBDv5
SRF/QROFuga5Mz9iRu3FzFMfklSsYTxdlRPKE92x5s8L5PqiYlZCHTK50z5hHV2cLSYSIrVgljqe
WeAKNS4GVnP4VtP2UVrgFGltlMrME2iKZ6xK86+fncXYsoZYB9yzAvo4uOuL8QXIM3SwCbhvixgY
pn9CmOGisAT1aNBj2tj4Fpvs8L2DKKfK9OydAig5Hdrj1fHcznPHKbgrzrxnP+ee9Jp/iaWuYFht
YdlDOKIyFCLr8fVGB7kiu3OMZA9PPsm5XmpkvsuKqJUIudA2UAMYrQeziS/QxmK3NdbnCnu0hvno
VDj7euLXVWUL2x0kg21RPFiR1LZ7TBPfpOtiedSFzzMZwS5fOZEPJaiNkcwqp8W6bdbWvDGBNBiN
4WeFIig2VHqwgbPGggfZe+gEsnWMAoXFeWB/vYftD5OSUURtcfQMWj/hYNBU/FOvvlo1mpCbj0WF
HPoqlfdP08NhLy8rVsxkzyhAInmG3+F/PYkuni7wvgaCpFmySGXJ6kE/+BKwCLyQUBCdlU0Dyj2Q
H2He24hWhvONtu+lBL6Aedexuv2UjFu9F2E6/EPkLjZZsNfDp56NGrTU0qxQglhDrbsSZGgp2UQm
R0D5jzv5z5au0H39CCXa7yh2jJs0gyZbgBc8yOS6WamjlYpL2t1r7ad4pSTU/JO4U3HsGr2Ar73R
+WiwRiUwvZfwb2MXflaoc/cGX2xhi7HhlVs2OVaybkwbiiSLZgobJF3NMJU3yaTOUOVm9VCzefFL
/4JLHMeXDku4iVHaoIoca9RTLas4KUx3qZPBUucTaoRTFPhG8q5Rm71mV+z2CVzZpEwxgoKg+iEW
bbGO94WwDOpwhd6DHvznmUGyUvvYeTG7oBUpZX1/yP7/QMguonYaxq7mJDtHLDmuemB2VHlh4XAJ
7LLCxzrj4jgPMPF26LSEq08ykILPR+9t+fj3VuRuSPbmXSzCoLDkVPsFyj+04sJhOlXw7SNDfYrQ
ct9Vvm8QUKPl2ACig3YavCc1WU6QT6VBnVcV9de0/3UI/mOOix+/Ls+oO0nWjTB1JiJAIwt5/BWj
47EjTfnDVMeiM20HNIMFosItQTOd/OCtawDLSUa8Ess64QV43c29LqzV4pLE9BDd67MZpOWO9Aa5
5WF4Wy1qETSutcuhI9FseM35QhHPWjBnQfoDWNUrPrNOmyvheHFW7OEGzznsO8fquueqG4FrICvF
p/+frvAuaMJutR4KRHsfRQFbk4JRbs5QY7F2+hmZEp6LzKZ33WE6IiE7RR6IzwtMswMkv2OJGqri
gWAHRinQg3CK1frkDKAlbaGd4a7gr4sk8yvXmzaoJ/SQZDtP/Ao1EJ0tW/HrZX9GXOhkoY+h/XKo
kY5UX0MPvL6SP+mOh0p6vmUz9OWkVFEhYcpbLaGDV6CbdBZj6ae9NoyW2D0tJ1NV4Tm37DbnjSWt
aSlAfxlSGSA6eNFlH3if8CLb7OH5/NXwiMgrQJnKKJ9dLlhx09a/HRUSP4Z6NUf6xIZw4TgUqRmd
eOav+TUCtrh5ODEwypTsAv6HVY49ozbc/KGcJ3uTKD/JXgwQBMoWhn3Y4yA8/g7MVg+QSHjn8kyd
xemNjmWE0anG2rfpoRrWz5E39343K6hbqRxijDaZiAWYp6fueaDR2iKQslrlKfYUtnpLy4WCFvTd
DX9cf+uQHmgSH6ryIaq5IOuiE+YGhBctAeklvroI/CYh7VW+OsZBnGLCU03MzFDTuXJPoSM2x6QM
eOR8H2Wm/A3jkp+zLbC4VyRW3u/HGAraauEYbtuYuOlEljkKw86Csg0PJHDG8/wYYSQxcoio7eCf
P3+5cYKGaX2aXlnMVK1h8QhuX0Tg17tlizhHWCwoIJ0/dGELEatgEyZ3Hjns+CIyFV3uZrv94Rf+
YUkiRxrUPYh4axNWMNF89naxVuDZFPoaroaboH8oHOVqcQVHDMdO706W8S8NiZDR0d+V8vQ5s4dG
lwfJAUBdNh7C9ZG8w8cXFboq96YkDzfh7fEgAg3/j+jfuSBPkVwTntD7xxMZO61EUeIRHkDAQSjb
bLMn5PQzJq7y0HiSq+xTC658jfHOy7GF5vWK8fly+8770q2Uf/tgy04fN1iV6qMyNH7rzmb2uIFU
/jzCxeFnrCHynNmD27f673qDq34rrEneHosMVEWApCKkf4GegN4f/j+8Wq4nvhIHUHXiLNbSQoSS
ZkleBSF8Un8FT7tNfq//rffwymSeKMfGi8sqDLpB42Svy003Hu4CpeB+dySV8pPuyuTixPLblqwD
iV3RsrOem4HxrK6gNL+goNLfHHTJWOH0nnEi9vMUxqyGSTRQdqUXCS+izCE7o8sMUZLH4S5HTj04
9fJJS8Pt2s3jObigtks5a94SXSpU4o+ZCaGslDaoduFXutFqrHpm2dWwD1P8p5zmQjYaB4FdsmAQ
3umhntEf9q9nes8vxRw9HPQ0B+fKPsypjwNTwY2qxPVTRl+r52gFv86MXi8tBjGmnis1zDpQkdhG
FdaorUY+ynlYkCQNZOzvuBFKX55s5eNBBnnA0Lmf6rrj4Fsq8Hp/6pj14r4L7Si4ujY2MDbukq7S
/K//I2nO8DOqyQlQDANvkzM5dlDqQNUD3aKOS2R1YAax+JnLT83kRMjGR4sx67TF+FjpDJ+UUjZB
PkMxzW4QOs2CT3FlMVc/eLK5cQdqV92gNQIKQ2r24bxgH7dtlLz4t6jf7ObSvpIbs4qzKn1Qqi6C
HcRSHCxSNmga1fiuUSbfEqSkQKuvyKlQHDHC9DdWwbJaGKG32GzMqDt/pHHnWbGzRRU4LKEsxf+3
fnu/JUT2/G5RltySVz9PA3ocZmVqtMQIDjYr1GzScbVkFmw++Lje1OEnOZXxxIjoJclw01IhLq+H
FGFvXjIZjxKF+udkh/fYqSZeX7N5wAkRGLK0qWgObnHpTrZ848grqX2CMmC+byVtL1nd16juSQCS
MCzL0DtthzgdjA8rlomSL+HNQIMcSuLFp3f161jsylYRfEQhLs0ougH3udrqXgrtlGv6U0tXAXHv
7rNQMfnuADAslZIW1Ij8IYfiJpQ5KRawZnZfAeo0SFg+xf7dechOo60kuuSP7Jif1KGPgVJqWhxL
uz3ZgcEthVQb1Nfnj/nlf17FEmRdkG1m0tvrv2BIV59fVUYtVUlpmEujciv+XkYFx8/xN0deEsYu
orY/NBIZGcAJPL1yOJv2ucRUAMmOzs7bk0T/Pue9AQce5P4senPPH/3viWs9VwpyTQFkS0ZEzvwv
J5URhwN2HmO/lthwX1mRAUL+ISED3tTZ51Tl6uju3/bYpsUHkD3vntk3n6DgtsDQxLIKrdcZO7yA
CL9TXoAyZduHlH39+WD40+Wa0xCs2eskaygjjpd4jBb8E1gce4EJxODylLwfFulUim1qWe6z4wAQ
7OzseqYIO7mOxKsuKZsLMUZe5Sd4FWtwQ+kx6tF1Ll2ocgy4xQzHCjYpdEDo0TVvBK95AdIDfUPD
e7cYi7bpNPlZWxCRJeU2DxffncAa2vp484pn+UfX7gi1DqF69w37VsAYfMfkMLnLG+bTLF3obBW2
VHD8lLsMfII5KCGo5EcNaMPn3e1qUbtBZSqhHDoqUPMolbEp48pZNYugyIWcZ8kfI64v54X8TDuA
YEBHZcjPtKzhB1Dk+7ixdudjhP3VMNIaaQL2KNkv/b48TnKTZpZc1SiZ0qJkiMKQfqWTwvole1cv
d/XJb4WonkcRnf77O7ronLUVeRkIMu4+VzxwCYsQ9SQJiCv5Xowdq+nENER72q4Tqf+QzyzBrHh6
MQXIG2e3Yly0Muy7oqHcyOssYRl5hKR8C1gBPZdNXQ0s5U+KcuTooOG6ygdN/m5DbMs9zpmuU5M5
w6sGeDQJ5pbtL2z794kMCib0vMtGc/6CAtpZgu/ejl32x7iMLvk5uomnmr97FQH8UAg1eBuTscGK
DI2jcxDmpmX60WDxhbu8gavcH5FqNjm4sCRf4NU+MPhkq3WjYpDdAQ3AJZjSxBqdKDffd3iGXfeN
3fHw93dPujLFaLexPwF3Yr9GQ6uPc4yCdc5dS/EtMEJBmOGQ7vOZEYsgRTvgtCsfcw83iykfcLIV
TRxtI9yz+a0h1d9AttwawtBQIDUvSFDHyyMCSMYn2H4CgEbVJZtBEbdpm0k5PD6Zye8HxyfU8IIw
BD33QSBoH2DvHs+FAVZKQ42ByiKPkDjcEwaagNG6GpSxGRVbD6QlQc68vHA/Zy66ZGv/bGSAJSPT
FVTtRImPwIlkewrcIFVOwLAw7L/yVitavh0KhAYInY5jA1JQy6wFyOGqa/WcAE6kiMMe0YlZGPL/
KVUZOel6uZfsyoILAASzIMndTVZiOU8qaWGcjeZl+xE2Nu6/vTX+Uyir+77JBR8c2HIhCrTRDTsq
FYcZ91XqZzsf6j5s1LslBzQPnZMXELY1BCu5Va4Q4dfKF0bKDRo2BlVJ7XlzsSEdUp2y7dhp6j1P
FfmK4PYNJjjviaWOT0SMKlatrHWLJ8bHM3y35ow5Kac7/3YVXhShVxCSDJtFgfPeZEn3dK+Fv4yf
xCjKaHCH8UPuvBVEGAdIq7QoDPylTdN/RYBjYIcbzuLcMcWewk6rEM6yzV0s5lWfZoXTe3wSL8yb
1C37cFnrcFk+4ry3MIr2/6fl0kb5QUrK+OKdmFnr9Qz9UOyQBBIVTC6Qh3onqr5chmbHnbiHyB/4
xqe/yOsTly5WlYin21PfPOjmL9EccfWO+QG+KPUPBPUsVnWXIj5M5tUPyV56lRmg6+VRcu9I15QZ
dWRIqW6bf4HnJxh4zJHmMXJvfyC3XLh1MkiB1RspE0YPl2LaLHpQ43I/W7CNNCzrDK3zQUhsnfA3
yROVlMM6bsqXpTv0CLNePDDXIXMx6fFJ8aQB6SekmdzN20O8uK/OZSdbRabdaocvq3Uw69i9tOgi
WMSZii2MeyMfoJef0BsYtVgfJayWMkslbHWOZvwi2ztojxK+OmnYcw4gr/41P/oFi9TrQ7eDwVob
Ky7VTsx6+Nq648+UmC9l7pIZPE8eUKoPqjEnEjoxUhgftAtWt3WiK2FuHRdqz2To4Mdad/4oM7k2
NMvrxzcE32Nhrb/MOcuefzQ59hGqMmlQFYOQNhU4sW9q9cII9NvG0UimBHLGaLvYzpN9wzQLBl28
r6/SWnDBClRM7icBBIyIlgjWAspS69OfrhiUy+hkaTViFjXXKOwhV89iA7le59biBY8DYIPskFf3
or0Mq0hiLtRplCxfqUUX0+Ae+JASCl2vXUQMb0Nv8sQQBLs79tJTIu+hPpVjxZGRo96M0bd2ypJr
6mV4whFpHHOATStmKCx7Zg7sYgxaTXF0PMnpQGnNnetk5E3Gro7tbicT6MsmelYIgfSwmCg2IGs+
z/LMSMuKBMQ2nI6CxI+/zQfIZYeRsdpAetHoQr1LIf2O/zb8qHhq4X+k+0QGbxqV1cj286IaCxiD
u5zp+t3yo3g3UAy0Hy6qBWJcPMMbwafCkvpn/8vra898qoS9tMdUP/MMdQ0QpN3/asesZrhMgBWv
KjoCnfiuw4fMA0hU083XwNLt9Sy4/tJIknLWmY49eSqrqGGjHLxaYxIulW9d2Iocu56kTPajb0ht
VSvLiKL8EVZzlJH8D6+MXGA1q4Z99LODT82xNu8nIKT7vmaIQhSlmKnSWSxkRHEahTvT5V53Ggju
YO/IKuZYWTMrrOz6ancz3Jz2Y1hWL6ihiy0nucb45lvsSDiXsuTAaVZBxuOOedJkePTpjbEcoObs
FUnjICw+S2g/Zq+R95TsYajlCEPyj2zadQAHD7gZu4EJk/+uXivvm9lwZtqbQtoxOxtPmxEuosBw
nzN5P0d/wU5E095igkUDgEmjZM0fugaOX6nHHLDYh2OObOGzlDrNw5NcLuwmy2yezwoB3azR60ra
IV0MsY5Asd2DRIbCKkXl+1KjoCJN88oqCksD8gYTx2xMn9RR6TbkJlFOIuaV+7VpCjNPno86Bx0y
Am+Xx/VzVtBp2LlUcvJBPABaRRPqAM4KPOsKtEnfQr76lHBatrq5YUCxisLMSZuCKDf4fYfbu7/t
ZjisE9a+V7povRiZd8IXsh+ob315lulMHbcYLleTVg0ZzWj2ooR98EA4dHt+7lHa8sPa4eNHg9hV
FgBOHMYrQ6oMfofPKMDCZKUlhrnKrNNRV7z2Ps7Qpin5Q6rnnOqmyV6v0zfpizMnZxIIFOGM+9ev
wC8TA9PDc0MpQk0mbruLhp3Zg/2Ac2ZY+BFNF8jBzYmpjeUPH8TB/V0+01B3O7UKqvfw4kIIhD1E
FcBSAwV29nG8Of6Pc279fU3/tFwJVT4QxcZS6UB8RtKowi8XWs5PbRI+zL/6sBeierUzczvqMxK3
JaI+7rknnzp4ERm4Af7CeowQGEowUL1id/+7at5rhZDTXoSZIpYvvhiRqqypqyDe6Xa7W6GxavZ1
5TVCnM8FTWIg5af9dl7Ts7gM35tlpcEuSPN5l/0JWOgGf5kPjr/07LSF/6XcRo0bnnF+U12kK/WS
l20RJg5bkXX0RM0f6hvCFqf+kTVLa5mefG59N+YavTqz1JF+lO4DtQQw9Nt6oDInvri4gaSRD6yu
beW27zwSH9Z7ob0cLhj56uChxl2UwlvwTOE3YAvPfYw7CUol7L43VnlDolEoNwNuI2snU/z47zaj
LvSkLifw7tMiUP1rJIhBrKnOxrNGuIhYO2jUbM7rOnYAxV+0a3JLUAPWx/q+AEn7zEVIVSq72eZt
vxsR51/HqF8CJSa9gGoF2j4nQpie+BEZG9OHShMiEIttlE5dCBMY/nRL++Gu+7F5Yl+0RA9ShVxu
JusVKbDPteg76RRld4CLxmeFr157e5yxgVRQy04p3Dc2Nj0InaKqiY20DNa7uKX73t4Fm0AuUsPu
7Zv7VhLT+ozQyyb6oe1fIi6YO6mO4ue5SjgH91SshpjlqFcl+X+XTcUqOIntZbpf7EzUm4e/nzux
P7fFZnLsmTNfgmB5UvqslZCy7/QZ2lYG2kiooGIofKH0BuZHvditCPGMDsp71ydQ8xssa4HmKRo2
2+mi+sE4/9eqliOPcrlHhcWP3wJhtkm3jPPJP84UML8CE/lMzFyZB48nTFkFcq/jClxu62M7kh5p
1WChZSbU7SQQl1c/aZc6pipc9NJLMtekaLXANvm2Vd9uFB9Ta2paV7fiA5ds+IPh23ilKkiY8mXD
4hsOxi1cTTUpxdW8dQU1Hfe9J1/NFR5BMuPkhHUEFdfyGqcaaFGhpqtaB49QPRERC81mdmHE6ozo
e5rsNn2OS8F+9eb2j2jr56IcPyxPh4tWNJFdjKImPiS+LzBTayHpIiy8FM9jOTEYUfJJFjtxNsxX
aGPPgxp+Au+rvruqM7RrrW5R97dqZ9+/HFTp4EQbjwzhz+yzFxwi8KeAOu2HfQ5K8W4s1/CdB4kP
QquglLe1M/Hm1TaS4X2LH5u7K8/PGN0wZiZZ0c3+92aAUgEt9fwnhHZLnbAqeu0LiE7TFVh195j8
QwOjkB81onhHaUwispDKR14P0tmZ8WbHMTDogcMA1DLL/3NMuTDjv+UXMe/hYCL+ET8bjk/rbAPb
WrQDRiM0SyIqqHS+JOAMFPQh1PqgK24IpzB9z+3iAktbw6PZNs9fZ3N6VQVlU/vtOY9Lc4x8j/uN
ZTaN/yh7lfsz3ycQj0VueHKgIfkystBazOCZqmdksi3LUNdwOPRQDkEJLLtA/VAuDkSwo0hhr0TU
OtQskQ/GTu68kNMP1vPurydL4WWcvgqdIb94CHYSjZJYDShcnc7bezOXjnsTCzC33sNUwrypm6Bf
tdlvMCtkKpTsbOLaWS1/pCSWqYEaA9mzVCiSsl9eohoZpovQmg5UOP3ot/qC3gQu6XTWr9Y82GHL
00pXf+xOpESFsraQ0ISK1O4Uc08NvwxEZkwEwiPagHzRC9gFdzcer+4UGIJrxT10YOPn8YYhPFfa
AYRcjJT07nttRnGgtH3OkvR9FRKHv9E4o1LBagmyxR00C6qAlFS4lWz1ZEAQJgP7spSUVBfNT5jT
JnV2+h7FJq7stMX9iavPohMkH6v1nbfmXP3By83w0txZ0W4jHRhWs3siC+GejYUK33Wahk3IwXsG
qqYTpfVGCj7BBlVzR4y5kZDXyFkivrZz0910BTWDmLfp/OfOMMnAxd+kAZivCIATkyWBP16vMQa+
W7F10piSs2qCc2EHgOYXUL6ECCLpyFPrvbaz4Euja7XhEXlEAqL6q9mfFSOeUxhOc4CecG/uGyIo
Kvbp+bdDFf7wzIj5h8swzILBVR8a37zsJC7hvvsiItfxEZnnxvt6miiDHjYEiQRriX/vd0+094YR
Q8qg9z/MfJJenjFcq2xLVfmqJM3PNylFkcvEqYkh2yIC7PsBTvEwL7eNU65NdKncjVVWAllBeFTa
KYHx4+DDNf9YpMNgzQbOAr3QcYBL91jdj8rzwCWCa8+ADAUo3Pbh7j7i8Ru63fY9gA95fyLIf/Wg
U5b/hYzjOKOaJvhWfdabP4E5UNHdGJR8i9LKS33AjYcKMKvlE8KcppLX7FQqIMiU2UyfXu/Gy5Gu
tQSY8AtddHg5QvI9mBJhBhehOJsKC9oxVOzp2fw9O5DNcxVUfIxTAKQRrIr3k4Ncum7xPuOJiach
nxunOnmBGiB6Q022dSAKXlKAZJrokmrObTQlwU3pnF1HUDF8yG8p1CHdfAYsnWYWkQPGFTb/sPdU
qqiD7p/iNe4yEwHDXD8HXET2ZWb5YmbzVscAeAb//epwKfxzIaZxCBOM0vH1IfS8P2RK7TqpLv2h
e1g+ppcd8HlZZpbIkbtzMkynNnv6Xf8DBHJS0mYR9HyeYAOBQqwXogVZxTilwpRJzH3FOwR4bP3R
u60IxmlGDgnaMqYovCYnTPbCnF0p9G2h8+E3XqzYTNUPVjTWP21NsiWz8KGxcGSZ6EJRVQGWFP7d
b1hH/kBejIPcMfZcJuenKQNEVp/eWEYb8QCV92HoLOZjxo2C+wDU1kdRZQMmYMFYhRByfjPtV+w6
q1z74vElga8qkF6Icox+/SC+eQxTH6Qu1nBEqBFxJglWHGDzS2vNj+NWigQTj4YXBUnOAKqGRJTF
h0OpvH9kueCa3wiXpDoqmZKX+T/lAj2GEAjmLqKDs9iuotx14ZW8eclHeeHKblpDs9lX2A0Pgxt/
8XXD6TAIAKZ/pPH9S9W+JITdgoYcEECZwJppVJ6DG22aaBAbsuvhYQFEW3+FPdtxJCirDYbueFQT
NefcJuiLeYJgPg80/QgetzMWrlPN+u6xaZWO9Q6lCTqEiFc/H2pI9hxWeFiCxgd1a5VTTGmhs9M9
kvFyXrXCsMdaoxJDaWGOYGRMbpzKZlsWPO0Z+U1dAelQ9nEMrtfN8AJdyhduQ/OekdccVRP/v9nv
d6MI5YDKXbEG7GssuGzzX8jN7c1ieqALzuy+nlEPqxS9kUXyro6Mi7jK4T0pBdQ/x2dWqp8vRCQB
TkaEayexLE9odk+hxQhIiRS8JmnzYxsJAmDK6wpMLYxP8pcQKMUjMMHmfzLIpIpc1vr2X1Z6ZWwE
37txHJbZ91vS5kiaUc2BKkOaptX3bqCOxThEG0aFc8eXGNXAs5jzVuBziZIJ21KUTY1AcDUkQBpG
aD7Kz+Uir21FVOEZG77osUYu1Qc1nhoZmmiQLT+HIZ8Y85VZI38ex0T6pzaIkYq0zC7VfliJ5S0u
Xdv8kr+N0KIjP1uEtpt2XDVnVTqyb3912bBa+ZL/4cgQlJNjwy23YZWpS4G6/S0dNnLm33pwuQYl
3nqZGWr4guQLlxd4v+u6xab3Kg+n3ds0VBUyW86mJPTuxkpx/PS+vSe39XhOYHLXMPGRccZFLAlQ
ecDyY/DBUx9vHTvaqbG15Pfw2Q4XJuZlc8ZxhdNq0Bm0KqRrZn93RrioVg13RmHFs0NAxItj5K3u
fZ2Q88jdmmXcryMXcD/s6u6mCqf37nAWZWFjY9mdQ0aj/hA/vypiMkc3JC+OOZX4KveYmSrXINIL
KU+UgiwDWrOYflFfUNpa++moUbDBALxzd9QYD+7RlDKfYKHTE6PM/jAfM6b8rhXLq5CgcPecCg04
ZnpFyZS64oqQdx58TPLbvxA4eoYjhOlWWj84jr5HLQo9whfl7j8ZyXCQLoM8Xt3D3ilk1KWvo6lU
usWaBeOWBsEw4VWUOlydjfOWQBQqaOECHv4s+d43CS7zKQI1akRK56CfmVhPxrM9Wlxmh7mNW3qY
qH1IR+jiWKNeQbDZYca9jZj/F3px2qLfz5WdmjSyosHhix+C+WSejpqRTJFlLg1kNZECq2z14AwT
5eHrO80yXSx9gI2+LNJny6X4DdTQVCrRmtEKJQK0SFXEEdLxPVnRaAxqvTYBTzJrGwzg8YFFXafH
GgrfnW5V68SUpSvpnPlRJDJ3V2uXzyQHhOtF1+TFtVQ9APBLB4/H190g4l+sKKASfOlX1Zb3oVtv
gxAem94r4SRJZKsousYp2b+19qusa6fMWnyt1gBRJn4Wuvo+96HUqtaFDtcAs1L182eaqWKWwOJJ
ZQLfoW7r7HtyE/VsbK6mlyP4apt183GLC5HgKEZBW2QAdxKZLuYoF6V+D1kBeGwbCGWgDqCehsBc
0zHglVoYSikndXHNtTNV+eIwhQ/Zro3iTVKUySLYzumPpUWqYg/ph5jpnTEYPHr8sMtbCmTi8oyn
Dw3KKTrSCghQLuCEnoAP1X2FbUwoVDASqrnCZNlmKwMoBEKkiozEuuxM9VDKYr4QwKJCsnKj0QTP
F1ccJ5aPTIJsLKzBrCsIYe9mbosOyWi6O0pBDYXFeEohF0nBhT9wbEbXgv/We6o48M2Jm/JyKDr1
lmLS6eVtI8kzr30PD3IcIGJl/VgoTce3r0N3VcmUh13ovTl6FEVIwOFM2KnM3ZUHI/N/9dYNM54d
LaoZu0ewP6lNyFxlTEncxvbrqpPqWlA/7L3r/C32IUjfs/+JLTVf4s6O5/nQ3CSLWoLNlzmqU0Zw
Uk1tbgBN+FLklTcqMdLwOxxKPx7e7sXUgJbFHkoGmujhZKHKHfq0IeHqwEeeBaA0fMXr1JI9IuDV
yXg7C4KThz1Q4LVrcyIY/LuiMjzVAv0IKeKYnPfnq4kozfOnoMucTxhlL0cDcBFZkGYvAJ38UU6A
pRQqe4CLqWDkHhvhvsS2fcfn/uw/hSyN2vfwpVnEIXkJH2zY1PHhMHBQF0SmHowHT/k5p+5NLj/F
/nm8ieCiLFiC6aL8OveOFZnRAntKMkpef+vvrhDcIolAHWbg9W5UuvOknWFnejfw4vFJLDjBXXOl
zSnMCIYMqMBbYGTkrpxWMEWn56PwSV/DeQ7svdikSM707qO7aYaMgtF7fEMqvF6BfBDSDPbF1/hG
8cRHFBNNCxDiqHp1yFgTRTiLdrPmA9tN8aJfrUnECKeUS/KEb/9TkCzQaIP7nkny2PzbYVVPFxTz
Xlhsmpsd3GAPfs6Funlos3c10Nr3gz/LOq9jIIxJGSN3voWZOG+h/inrupywRDm6ZtzKKcQ3Md1L
sCNflkX8mK8b0Slrq2If127X/ZtAHNF6FkMWKefbZFriTnP6YiDMSwHHBguDUc/ZRFcJBFGMZMwp
q1GljvMnxl+5jhwOmxfWFLxcor4+YRb2ryxIZjvhv6skOG/EjOE24MMX0ElNhoLJ2l22r2NwbuHy
Pf9KGelj8LAOZJ3fJ6OwWws3VODUU62SY7DUuISHgPcmU736ajohSMO2Knkg7CgeP/z17Oa91ZWk
rN6j1s5B2fcWaPYrGiWzlBILE//1FgQ9/b+cz00+FpcVM+kObVSs+awe9iGZbh7sTfHnJPg6H2K7
ds+cGcQ9PyqDZjlH7wu2+mP4trsbDa6KqBak/K8RMo1p6uXQyhjC7WwdbPM1AQV8Zd1fCf4mKf8H
nPZKPjfKqiyd+2WZ5KzueIp/pwIxk+eR1Gx9iw3GgGLV+KPSbmSCWt0vBVYLTLDRWGnXvBDdHm/h
RveQuW/jktkRI7BxN0CA4eWcmxjpgkK1LLF90aaziZGtqBYxpKnE68S3eih3uO9Sj+vXgnKzHPtI
fHNj5+GFY7XIoURE04WT3w4Q0x4hsTDReNqqAozXoJ5gPA+t7MwL2h8Hx5IfODCQNd2VZi3mE6Wa
8y23EgSXenU9EXa7d9fT9E43ZeQjOLxzhV7ffjnRm+xlr0bw7h8EC+CB1uJIpBN4xQB+kpBshqQL
jWAXy+E1bA0dQaB7qAtTSaxEcpS/qhybspz8wA330bztVc2SvB/GUhDrl6ri6N6z8Qi/nAAAGvuL
Hbh6dz28Kz+5dqg8Axx9KZvOVwnFjIf6p1Hq5IjxK3CEumxGOz+fWLS6iMyUX6RaTTCtNBu/IqXc
Wfl2p6V6OyUkdeFRSNHN+dOxM+lJW/osjflOYJjDAybJiXmzzE9v+W6YU0xXiT6BEOKxLMRovnuE
VTHSK+soy61q7ErUYLuAM2PR4MJkIWGxKmeHvjldaF+NutcoPfRWEiCqrxBrCuvxh7WZAFp/lwWn
diLtmXrhdcl/D+t4gupRZ+S7o0gBR+mabdd+DE57Ix9ko7FZAPaZRJJ3CI4ZlxhJELAmTBbj80P/
Sn30G8UGOI+n6TGmh1XJWVj9/O34z83wXAjp/LwCeP8v8XuZxly7unFMWMFueVDlDx/6yWbrJVrE
DYTHYPZwpbXGaqdPwPWJfNbEq+jBG+030RW0mGPMPUIp0oPwr3AON3wwqCMSnz33RhUAOlSTvWhr
YRYgerHtn2iBjZEKO5oH8zLDCqgbtLYqpSj9e4V2RoOqNVyN5Y56yXxi6yeE3L5npoTBQ4iY2dP1
hGMKBo+Yz9Kh8a3ksnotzsDbZ7505YdvKfYJDafDB2u12VX+x44YTcAu5kMd+fiU8bQYF3t9cWig
BIKdEDtnXwS/YAKbTXRlujN3+H90QzYXCi+FUmDKatIcFwGecBUoYV1ji5NfuuYMPOf3Wy324bXC
ivBxHggPbyz15KMjdnebpNp+reUtb+wgzKounHVwp3FBw1Zi0nBwNV3JTYAr+lRzRKdQtuv2scHg
n5tQYuQktSY0oA1HIl0+pYK92Imz1UsUlIe6B19BIoMG7tezQS/uBns+vPPP33Gl9s0nmVBfEua/
dHEuhmUZCzc0hHTuXie1RCffU++e/mm9fyc9cnLZ7PQXq23tBkxiWj65IRV7FoFrqqqU3KOE91Is
h22JYu3vZwWaRAQmXXkgXJiM5/SDBUWG0OJrOZ5Gtgxps7vGiy35zzO94GU2lEiUe9GcaIrNG9fR
/TVuIpyVRoq4w1aEFMlaVjQbJtT89UE1mq1GwmyaTnl3gmVkWXvaCNwHqdiv9CZVeZSYQP5pA5fs
/iWKqTiZJTfvhuUv/ZZF6JD/rUPDUy11rFeBw1Z2vlKkdq5lrNR5pTeWvfkf3ldtG+qHh7UftzjR
TNGy4kgQxejvfLkWAkv3VsTUcyY75bMxxaoKmEsXtsLSMaNAmmsNTKUJZvkZB3xTThJBO2RXKuWN
2kykVp5GE1FfIgD6g2yPIictGAyM9lTyiDMvlk9cYHkAs5QbuBHKYAvPUbL+7YJ/K3vdOPfrhL8f
oylZNzYpOvPUW74EA7a54tYX8fTnqrxOnFMoC1I+hlD7TN7RMvNR3Hc0O9ude6lAuyRfeijFKlAB
OnyMydt2chyNsibz4eaHcgZBOxh33of9CoGOVfeIH2oVy7E3Oyg67Xol0ANudHdJmnWp0K8J4/bZ
JwQKcCQ/tVvkQVuV3cta/3skDjQT1Soo8mgGtqzvQFsGzp2DFiArUdHszTq9lInTyLaQsz15BfCt
XldhcdL4RFcj+am+w89cDsqqAeMel5WHsyWK9PJTclQ/o+vfkULSZr8yBefR2E2/SUn5NBo7u1iZ
oEkLOn2yIzFEkIa3YxcmCs6A0MZ+CGJFMWa2dsibKLcjuHyXLOyQ/BSAXk7MopEffX/9hMInLBQ7
w2eTy8O6r2BPP2PUv0xxtF1bp7hg7yRb78310cJlL9eM1IFrnos82T+HaxGcojCZa5hnNvPd0Ft9
L7OIRPHPbLnAo+D4CkESyvRLryYLYiXjm8qo4dyYna6C5/NdR4asJFJ+85ZyEZvSjOY+b317dsCs
f5Q+QxOJpZLjkgoDQXtdv11W3h45JGX3OCrxxr0CFKHDnjeS3Tt9sr0XItmItsRQun7kPojKPSRI
Ip8uiIR0b076t8pTsGNNw5/Cndo2T5XwbvR7Yz0OU9gx2lsJIoZ5u0raQyFaVtJ2X4hEaKB71m9V
9hupJ5X/qcEGDtciyiLqZ6fQZORtsJg9x0K7JXzm5MgIY7nJ9G32kcTdfXNAuf3wr6xWXwx5XbeT
ncnDiBiW7AeOg8LP7a3Mai5aOnUBv/VAp1gLMy30q1vMObaw/HxmHXzwUoUrOf5Q3dtrRP65ZnZf
F+kEMLvn3+yb6KrOn6sdLlO2/no/+4aiMs2DolM7CIt2IErA2PWXN4RJ09GaHAANcS8NCnq+OvTl
OUNeqsEojG/sQLdCqh5Hyw3l7vZbM+B67/XahR88aJWNuflxuER1ay0xKp4hG35++JAUmM2ZtfYv
65OL7ksiBkYBc+mQZLdQd++b0GT/ADimRtYt5P383TOwVCJ3R79CPlfoTjKeluDX7qgJvA6goWvR
NHcU2ch6s5mjZ/QJfhww5+XDmtnFGIVZq/bicUfRhp+CAPB9QPtMU1dfsDBm0B5YNSWkaJwRXv1l
XXQbM2P4oCjHVj1nZEFoi16oJ87OQXFBscoDAyhm+57ZC5DxqSvtl+ZPxb/1AyaGQe1ZhfHy31sa
YpUCMsDnRYQvB0tbYSyMdKNc8pzZhl2fCmE/mXle3g6oJWe2EK3Wj4TkOGrbG/SMnacESIgmEwCN
q4IEaKCiWH10TN4nDTZPUMHZESeAEa9UXw/6GdUJpyr8o+mjpGx6RglvgClYGihoCHsklHKfnZx5
7mrR0SHsgYDyMMMu0iA+OdSihfltuOaRvk6HY4rVrOdFlzO4OH4MtQxGs7a47yVYlgZDJesq/Usx
XezdtqZmUoyyrM66SDzAL0FlM+gOP1frvZwC2tEUUOlWYyUdYcQpdxJ5Jzqb7t7wQ4t6kBbUEr+o
CQGTtcGAsf3xw9Da1mIoJbu41g8WJpE+0BDHGl1MTRM7RKU8cgYgEY9VZVyGPlFHVIR7uIjk4/Dr
II4lcK7dN7iyLyzPA174R2tf6fommVsb66YfjC8DPpPPYulxLvAlt5sBg6uo4e1UtYTZpIBn1zhI
EPpvN+Abu0V9lCWYXnpdi4N11FHmamLPTXFMmqV6OXEZbg8whDYn2XLBPPqbVrv/Anu8bjU3zdYX
14XflutUcLB0G+Pnl5iyQaaflkeMLoTQNyGpeL25sEOkrSDcyS7yKHY2AudXCAju0ncaPtEFGU+2
3dhQXffLdTbVjFV8RPmcWDX2V9+qrvJ/8Dbr9MWSleU+qMQcZ0UjB2kSiiO37Gkfkd7Msr/QzMtT
MJI2/YPs1kj+Y86+B9ThxYztYU173y9unD1BBWO5LCCg6Obow0vmUTEFz1TIU8hqIKKAynQFkRie
AZYAdA6qe9lDrsVDVOMbGSmMwjfoGseKTceYs+EcmR3LZQ3xxATgZAp5dlZWteYIVgozZ97vfRiR
QKCQG4aOTRivdhtiuzxdlTTmr63jjfRJJSxCK5N9Vz++sfeFT1keI8VMnReRdCh4XrvhYjSv/kRn
rj8QSPatehrdS+Zl1+AqxIZJwhXnCHX5jeV2Eoju7j+/3Cz/vTC/CU8Yhs7TdUKGH8XJBayzLlSZ
vqY25xveBAvm1F1oQOfcosvF58gdiHYf6Sr+7afLihIFZXBgzWnGv1IqH3ISnjjpoujg7+VDQHeV
Wwc3nqgtPu5euCXRiDh4HWptQXkYWzjvYwcGbqMhlbLYnXalEGEHApEnUr+efGTISMqyAhCyubLT
WoeE4eh5hCt+yr1TxJjfXH6WYv4CuVcIO32OgBpBrMkpXBWF9r+QsUo0MwTolla86Se6kDVlDd8A
y1FU2aCerK4Io+fpxvBLXkao9ncIhzktyijKTp/4fGQEGuQFxms5IEujf+t/g7VP+KvRlLTyu/FT
O3TlpFN7vi6h4MbZy5//D5kL9jfgDLxC9/EVmV6A3J2QXzlLBnAWy4stcM26gnqFjYL1tKG3bHjk
PulhICzbYYstH8aKzzya0aKSlA/OAr0BrmVHlso061yJUb02O+b1iUXeMYYDHpBv5UxhrmK9Q88o
RvGhlWcyuEvxyzIDURERGruowSM3hAhGp5IbYZsFcQvjPLPQHspGnlWGrlhGirWZ/3nZnMkGINqZ
1dgk2Fp1nW1qztEHPNoofEukDaUHXY8mG6JlKs+E7v9O23vw3Y6cFWN5InPfUtA0do9fwb7bhCO0
2TeNtDVz//FZaqxBf/cWqYW+6rbSs72XUTJ6MYxnjAJ3fZe3y+ib/ryo7+/TOjS3DdeMqOeCm0XG
hOautTshArr9sa1c1+ESwveeMF0gpbT0OR1VqLHbeM9H3O8EFeMHmHVQKctTeGIJmbvU3V64QQni
ik7dmZHeGQCYIlxalUbK/K++pe8Ht5dZR3SDKatgJ0xEW2ZhaYYEx6cH1hQUJGbUe5w9Fke9VWZI
gx0hrVOGDIkf85JiLMnFCrmckyYKnMWUizfrKrKZdAcF7ho6L4EU/x7AxqjrLSRfIrTWg6k86Fh3
HEOfCVaq2B+elWmBJDom75yZ8fPbVcg8FeZUmKQOC41YKQrskh/YoeET0yYCrav/fpurxv2XYtJ7
7MHrOIRX9P3ZkYF88MTTl5tDUrJh4L9mFYb9VJLN2h0BntC2xrwzMBxjDFDnrdIom+oDyfIkrBEz
mIRjYAMwd6iRXYO6ieMWywV2hpdQKwb9zUfw/vT1xr4osrKq4S+G23Esz1s6XLubYQ1piYOBIBdH
gRb004DMdriI7xObYbU9TnOy1gYC9Dt4IcQ9GLfZodT+cmqDnW6psOZrqNkq0kyKczd+i3bHpB55
W0i+tM4E/GJXNacEM2yPH+unmStqN1adgirwhlP7uft9+9/K1Ow+NSdq5o6gxW/1+jN/GrhXAVGl
iQ5OeNS6XvLkb7xtlBg+n1rzQLV7NKooEeSzuJ4LlYhPLrFR2ZLrqCNtTuyMYBzEgEKS6+25z/8U
RyYQa1E5c0y8PXwp2B2/gnCShFnU6OT0JSdMhfNjbFLRUraLkuOjPy0+FtWzPFhzeW7jzLL2n9Kv
b8GGR3MVTEJeKWIREP1sSp8LpoQEv4euJLzEr6lTSNV5LNlRuY9LoZfeVcoWe17yTKI89L3JDgm1
BuJM/Xql+1muzP3dazevwAYti2tQ4D7WSjty9jwKbRQGZRvve+hBMPGoh3QCsx3XjLLg7cnGjsgJ
bDiWHV11pBYCn0Au89VwM4xhA8MmF5g4MNKq1HMF7M3x4cVmApLliKuWL/JszHH6tkeFhi6rUf4+
UOjmANfYq+o0XWEwgLTO8CMIJtp/FryvhDPvTXyoA3k081D9NWjKMM4q8i2Eko491pDbo+GT2sVF
/ajR4G95IN3zcSqnA50/Yf5VbjfgHaaILokO4Xm6t68xC5lS/+C7icvByR8sljFoHNC1AJLGOPn4
ObZ8xAFIxqpY4g8N1qy6gMCfKOZvuZfVv8KaoJL/jkunn/oZuhp/qV5p7bwyUJprOmxrxV7NXKHe
U4dQDnMhxeIjJGjhGg41lDrovlMiOK+u0UHdEUnxpzmG0PGkzrZzh5YPPVUbKEXAIYvzyOky+Xyg
mB0zm8ttTvqUpCW57CeweiHwUd3rWm6AI5Pjnri6iHF2Cjiq8EoiUsf+atJtO2dP+1fdZ42+ckmS
oD9engOzENeGkt0GXn6pkHhhHW3L1BWdN69mX21FrTgpOrh62XMydEsLXZnxj2Mfci5ndyYsmfiG
VsxKUjYPvoSE5o/AZq3mS3GmoQ3xFDiigBO7oX46eXVeUvXvyTfppxbpIzUJi4bEROF45j0IA9Fv
PL2+GI1ENRmyzEnufQaSNushOmGi7kXSdAGoGTpbtfZqDToNMt8evx0JmAahuIsClz+xLBaa7hfP
wvuUQrTOkEf/DG2aa9H1sr3kkys+0nYzV4axVNAAhxJA9nctGEoZRLnRLiLNHMrxFpxGzNgcPLMJ
Rmw9zKH0wyobiwPyOnNh6vdWLon5D4HXQ3HRLdYZuw1rGS1u+KosiGLHzfDeIaXX6Ye8wfORh+/d
xdW+FTuwcYc1rppubU6XYSFw7zx7gOhY1l214iRZFy4xZf8OM7Mlepj5CJMWXZDZIBaKqafmsSVd
nqph9ZmJiPl9RCXHuKvlT6Z6opZdUazPU8Ohg0MitudSgI8cOysS9EY1pk0eo5tILYYxVeane7gA
x7LhQ6Nzy6j2hCmh6DvcAHrsj5jG1sSCVfPWTR8c3Ci6ikZkBK6bXkASjAm49Vodbk5suTfpqCJq
Q3GTaGubSacl3jh4D38HYb12PsFMSri5ky83phvuus9N+9v1jinDdS89zzGlGRUJJTVv7QakK2UX
Cd584TzZzjlJ9OQRDpFhu7msoZ8VxyIqxIa6VBErYpgZt93onrGqF5g2D45WG2q84n4SB0rWjZpx
rS+RNQLfqNboBr0glmZGebfXRCR7CiMB3KBGW+WgRAn+8nn5f1Ml7VgniCHZf96YsaBRhVozjnLj
YvmP4j4FaC/3wH1qj0sZ4nPchlprgt6Pfz7miLrpl/Bt149IRrCYZi2BVOy8o1Ao/+kNkjxMlWjl
ZQFOrcFb/VBvWlaCvzZ7qQ7iJbpKxgFyx/UohuUKF7aatcPrUj8aP26yTfDMbnglzCxtqRlARPIG
UebavmDFK0Hug/6lrUq7A3esc8vSConOcHfWmaqCq/iU9cEJtHd5ylLWuDnL1vy4VQ0uQ6oz7NYU
3lTRMDaNIiTVyJSSvUKYbdS+HaapzRnSmfIOxj5j3yyRvuZYOYIIg27sqZcUXXun4MftwPObWDEN
iXXl0NM1GKKUw28+X/u4UtO0gg85DEW0kLeSNbnzaNAtH5B6e+mVjyHbiV8kqXr9hiNH2ledjxzr
ORZt27KvSC5ZntX9DRIRSs3z+VKp//4YukuOiT5TZXyNi3tuBNAl00n3Kdvzf7DmWGkF2S3dcrrF
eIPwbyCu1BerLBMOhIcdBgobnNm8W+SNwo5q6axNiZ40qumkewYyfKuYwvcEObxUEw+t/MHsi60U
AkN68wQQlsirnUnb1kERjldjc67egYWZul45nADpRfsC+o66aaYAqBGyKMzqI8BYjo7SW35/QrTP
0YFQcS/EA8OXxmt59izGVrlXTcigk5aRoTIQnG7BNmsMv/MNRsi1rIj6e0snQwAPLQMoqW/zheiq
cnEyiKMqV85lMaOjSaJQih/MxI554qPlkxyPaE5HfdMv0bidChUeltnCw3JSe33l+woG5JbfyOfY
iv13jYVyGz8voRAE/B3EygRVurThVeqkwaeDj3zaLFPLubSrWupNpuPiAFNoBz1V3i18drJFrJXd
EJ/6GPnM31CvcFz8JVkgzTy1o/QNhRtiZ6ybxoR9yUMQXQSIco8+3jSeoo0/gKwblLBYPpualUIL
QY+U3pHojX82t6JDwESEfhnTS6fJTtg2umkBT/qz8RcXE9qsUxPrOTq5fj8qRVoZa/5f9OoAsIui
WSS7hA4KyAryjcLeyIzMzZUMHEwNyU7DU9Jogk43I+FSr3gok3mk5BfgBOcy1rfA1qNUaDi+FmVD
TpOSJ5BMRJpbGp3UhAqlNXNh5gqPhhM46xtSfio18TKeIs8IsI5Vdh9HcsKP4i8ypWlC8/ltOR54
MWmVcXpAsfz+vz3CgR4F7WuialWI3Nj3Yie/kr06OFUb6TIu780EyUW0Knd3cckQezSwICB/DUbo
lXCaL0J3Qy+Why3A+bRwBsqajwSdyR00CNlAvdE9V5jI895ZlSB0/eeXDidIwcJnegHvLGMzMN21
zyk/xi1Jwac4JEQLxNY65u1RQLE+JyLP9VqZMee6WpRd2ddhCL+DA5RCBTfaqKmpD2G1GPrK0uzc
A0fzC+uw70BFI0dD1WgySyl1gsHosgNyjG4VRX7YW1w9XTZFk4r451zJsImIyQl55qblGshhloMR
554x1zmaNwlrpFLLaWwVPGPsQtbpTnmzE5vgnt2y3kqntB/9ZM8pebaUPOcIGDMw9PRm/bBTaRgi
57S5d1zVd6zqeqL1yhtG2iGWvAMYf+c4q9JjwmZaV4ovbUmxxwtQxFr4w91sJhbMI7H7+tZYg51E
9G6hD7fzkKnR+WVSAZiTSV0rQTMZM9NLF4omvPXy7+HsRmWEKg3EZ+GAX/R3Fkth/smw6EGX9fWc
t20o33iMxGUENs/VpzzLpZdQIHj4Pi7K2J4x5WYMx1SVptLiXpGpXrVM9Y+i/kAv+/e6gTgz5vpK
1l5+chy3M2B7R41aoLdTJ8Cie2ad1tDW/bNVGjgyuv+JcRbHCehBaXEiyVwk2SHHmBzMm2a24wGU
UojDgpjuFFjqRab8V8JFvnjcA/s9uDsB7PWgO5LH/9ngWHmWb2D6kBe8ZJURKSDVtAHzUAT34gvO
iM4tjPMDMuh/iwAwqzgWDlZ1ZHJ6YlS9RuveUlYz8asK20mXMeHG6ebMV6EJqNsrHFUb+qU9TS5y
Tny1H5cENP5jQfVZnIRcH2oEIfS8Oc9XImdVuhT7y9k73uP441r3JQBewya8ZWUiHNrbUVoI5YvG
rTaAlevrZdAQd7MZBGAPBOflq0nYl2NTeYjF+rCKpyshmXGoGwP0FQhK/UJjLUyvSUUqVVXcf9X9
dYexq1f8ApMMz4B/4b+6G09EsB/qHre8VBEd//rvpvG6RjTLJMD/lxZO111SmM8vpOeQKTPFK4Ml
GkhgMewkktnkxOvXp/+jNtrZoT8u/HEOnOJafnsFrRM8/FJ9aopqnsPjbhyGWCKv3MXsQkZrsCWD
I/cQmaPC/PNo5tUC5oFaGmrNfYrk0xtmZXpTjP+apb4brxn7o2DjLO+U1hjFH8vCJxNTG1qTrc/3
Hi5rbvc8NNqmTO53IECa9JQ9EfoJR+rfsNa1qQr8xiejFdr6rpOqzMGVJWyK+2PlnOZFJHnvFmKO
24LS1yIdYW0Y3j6ZtzXh1FGBV8PiUSiE8XbJN6Nw+/b9380XqrY530Rz/JyAVnu61UzTHRDLFgqg
LopEaDCG+k2EOXH1bCPMlXS6Y132CBtkOVu7jrVSYiL3uH94Z48oHzLO/R2ZFt3073c2W9QgIpJQ
S4ZetE9BXNweXMo8lR0Nzw+AYS8thRubWlNHQJtqINUyP6r0l+dMuJQS/WZzVQHvwxhVWTxBm0sL
1am9DKavD2VHaPjz6IZ5e2Zq7ykdWeT+94MhV4lfDzR8FY//j7nXwX09r6jq1BnfZirlVIZqjhzR
pvK3kwneSX6IicTo6V2JGr00/6YmLu3kinpN3CMQyIXkKvm4LW4dtzpKA2VtVyAwawN4J836Esl0
wFH1Vqyxpa27zUDH8YWz9tPAgrBOJbM3qkQ79Yqg04yfXewJP9Dsr3JvP1FoCuLFATwkx7Mp6DE7
2oHsoAy9SVg8vRruCVXy/9YhKgQpZr7muHVU7fAY1COFfplxldhWHsg4bgsdKPWJYoPwY5dcCCiY
wMOU6GcFN61MN20qHPL/V1jkF3x2K5obDqS3tGFFC8dpPdH/eXRp9gjQZf1FmPCw+sHgBk+fUFzU
vGPwttaZFRTsT6R3bZRKRfISuT4/EQQZY8dBZhOdRjFRwCXlGgM+2Q3zQGvAD1Dx7SPrW2ReEkC4
W7AFfwl3quan9Cn6eQ22/R+2f470oUBzFF5Y+lcJwuzX0CM+OyFRbdMEu9vEnkLsTwB8rE9SWNp8
3WmISOy3+X3lOcHtlPWbYS3tUk0bpSWKzfdsLt3c52IsgykrQZ9lsxNI30v4zzgJeAW4/vcOh0og
ySFKuuOkDbjPZLp6PMCdpeJGB0xxPL8G455ugM7iyKgsPHd5/VbKzqlvA5Y6walRQF18IlnFsqao
cdQQvkRVnsMC6zjMUCPs9FM/AUHfzgEuiYH0b3FEd/hezfcyMDVcQrV8okCwHktx3AHtMYEYBEgv
MjitLByQvHTdyGaxkhvamOMT4keYYVRwz/iEwU54GC19x4MAq7MpnTr9yas/d4J7iDbr2/4G6Kyg
30/SkldVoC5H87YW/g//1R8kYG0VHOLh/oCvh/wlxdIRG4Bbz1R9tTM1/FTJXPgvO89iWO0doshg
FiUakrlzZH0C6rNrVPjPyvcYrsM6Hcyef6oaICe2xpHhnOFTj6WNIe0bBdFYJ2ZJx8ugYHAcyttx
Lue7XxMtTPD5s5qUI6iqpghMKvu+ZlAh4RkEm0ZiIsDDc7pp/UrtucrnKFCX+27KOCH5qBmhguUN
WpKo4FJngFmXjs2OcujMk+NLtVvmijyjE8cWh/BRRw563QEjprHXXJjJTiTc+1GUvk6r1t18Bl+E
Ew0C3cTTBLtefsf2uuD1ancJLuePYnFLZrfEeYqA+Pz7mMPqoypiJtSvTZsT+F4KLTrY/RQeHiT3
mMd5SsJloN2AwuoUkpreGCCzpfGxR3t21qQ0H4iZ24ZNH+scLvq4yrx/Bu4XF8lvB8wllzg5Yctw
ej+q4ZOk6B25OJTRjwKbBLNPpboCoLfI+9540U4Df2SdSv9/OWbQOGX55C8yiEadENWIQRgjgR5M
F8CcSlGqBELPKVeRS2ml32DCGhhSCwJgNuC5KbxyvnSLyt4L6MsidTqKQGyBUDdNvgnN/crxVlVo
yJO02jzz3OZ3HJMxXXCRmNU59rsNYqUh37boMC3vW8cmkFh+O1s/ZaSUEInOg23AsLmTsmKuWewO
JVRWLO1r15P38hgf1nrI35SB/bc9j8HiV0K18g4MiQxWEAhzP4Zkqx1GKsXgp++OycQDhgyYFdnz
EqHrcZRAXdrFN9Sc2OhQkqg443aDPlSYYCCWlz0vPvALZ1nSJY6/f/tny5HBlF2q02taG4GLQSIN
YZaMW06L9IRbUNh6or7Kqw918vFgmnBPuPb98v/V9c86eEJ7eGX1KcqnZvy41VQYZrutVxHz1pWB
KLEfdbl9OpSG1w4WpyyGtwolZzGrGvfTXf5yM3mPucfFFkeIgT3hRffShmYUQK/epw5wi17HOuN1
zrbEtxYAfYLgH64KjOKQXp4Oez24L35086lkdvh2Pd7VU8kiQ3snVyR4uXK01+ISHLV7n5ahuN/d
XUXKR6y0MM4HMzjC/Z8ZIug9mX2ClN+WgLdzvVg69OLF5R6Gfh3NZyTMgqj6UlaJnrvT6GflVHop
YJhvvMCyLZqjd7rYCY8FQeKvoMH4QDEkGXCnlKA60xuiy1++idrAQZ4i6w/WSlyM6DO4Qcj7r3JQ
jFeGSfjJ6Qv2afihHqK/9l8rGti0SdQxUD3JJyY5VdQywFNm/vpDx2TsXUuaDATYJRHByp2UrDZN
ijQx9Xqm2VXKTQpQ0PbdCuDrgXrZJLukjYLy9oLan7Sluyu3oANJAq7diECkarSLt1kEGW+VRWDK
0uQ1Hg+tl0npWgorCeSzVgPXQgrIlrpxn3tebFNvJk+c5kJ1GmCxlJHQZUaI53C5x7uPB/2q80Cd
gCM21BarfUTND/nyopW/7n7mT/ix1QEG7rl9ENq/QJyhpKzDBCtZdSHd0wZ8zwehFxELZfOr8LHG
gxuRBXOg7wFrV3H9TgCWFXK4Na15l//f+z2P1kNswaV4zwchUl+FB/t1wNP3goCXSpjWHZqGkz7C
2H/E1ruorf+HI9746HpoxI/bN0VoIPN+syPajKzFVJ7s9lpSk5J2asIMRgpZ4NSvXk+NkBd+0ChW
CZARDXZgUUy4d6O1o7Gde2oGNJsK0uIBvI0HBc3CNicseDxDZlJM1IlmOOBMX42G/L078yK4ycx8
EkT5xyhXRVQjQImktTcbz6Z9Nuj8S4KtxLuftRgYD9sbNAnswAV2jgR5CelHrf7sx+IueRovunnt
fECBt4wSgIZ6nQiR+RzeOo9vzuTyeKQhv0UDAjDz4jFL90HndbpuzLWIZ9AofOfW2T0B25rHnJHu
EKp2Q2H229izpa66d//aH3zNv6SdZ+RtxPmwfly5xri8Lwm3g/3CZnieoHx7HKXkwUG6mmgaFjmK
56aDa1CZZoLIn2MJcnT0k0QboWsLoDDNkjBU0mcW7Z5viwNb23713S80yRJ2qv6mCjqamlH+ZL9G
wS1yzBF7qXouiTsUGUB0YLIDY21X3WnBIbL03n4xlhbT10vt/B6sW4F36c4vD4gao2HUKyHZYFax
/aPrVaug+lvZE1EK4TeNACJxRTWGvIjGpmycwhE8ODwNocIcIl38sSA6oEWFvWxriGGWzmndDUjx
SiFFOVM62uukHHtDMGjSTclWffO4UuD9BfvoWsEXQrXLhhH8WHch4Oz7/D010/UD0grydDB6qOvq
Dzx+g2g3z2FzQ2Ac7wSMNxqiWQjUI1bL0pVpLPW1vF+SzW9rag8BzQye9xcfsEtg26oZmVYYmOum
ni/7RWbU1hzZHfgQGB9eDxg6LNAFxKsRks8di15rv0Aytu8ZysDEZevJfxWbg3wCXhHNt5v5/D8N
fZJ8/v9zH4rkN940oxGg78oai9hiIuOTO/A5g9gQmJCtxRLpf0sw6JSsQw/qYEqYMl001KvY6Z7C
qR23hb/bhha+2MQURr9KF2IYUqqrq1gmpxJnLlv+hhBXFBc19KNPFvPYqe7LTEyIa6uZgwX8FpA8
Q3nBGYrl4bwFolbbaO83kFz8PojcXzUjXvznkaW12Mux3lOFoWy5breO67R3qBuSrLucSLcgQ+na
pgsJy33QRfQzyfCCDu4arBB02vAF85BwT7nqX0xfo6x5xp2dsGl29IX2BJfr3t6O3XXCfcUzsdZx
JJoGvdcT9lAfwpzEv1Sr27FqxuSer/UHvRnolXmSKrlKXphivJs/m+AzuMXduWT57iBiApfG8uAO
dcFZ0fP/lJdfO6EmV+yE760TkxgP+sb6AghhBQzDOBq2j0EB7I/LzocbxrILcvxmgXS72OP7mC5x
DtQpBCsXkT++5PWqFPRG/Dn6H5hJZ1La4KcrULkXFEhuOBk5IJszLHicPFkgrCmyBOHs3AZbVjCa
50W8UA766R/oOn9zp2lhu5XmNXZ8e0apve5zYoOeLVo1Ae7l5IqgYDy9AKhar0IXlecXY/cdy/V/
rXsGOw5+ud/xc+UeCKFk6DTsPpG2PzrKcIWyqMyBLVjpcJHH4ACa2QMzxtd/GNaPm6GWydMwGz9B
VDgtGyw4kaQTJ8tNLQzNM8Ux5qZn80RJ4eARWde+f+wJrThBvTro5bg9WMD3lI5RTUZtgbxfQJ7J
vzeio4a2scFttBRVEDeMW43/Q4zsvMn7wIt9J7Zs6cI/co7xFTYfMJu+o/2qi9QdtfJZBj6utivC
7SjZCiCLh71ZXh4rTd/wvSP08GbdiHA/E+oGoC3AsLphvccc710OT/3dykkn1elPT4tr2u5q3fLe
ZFUYOF9vQSfqYYhYE445XcIwQ/R+EkOlN3DDWWSejMCbwNN/t/OBTZUll0E51794yWr8aBUK4scC
Taxis/kT21jKWslJ9w/8Zhl0zIrKa8Nu+ma2/dyKUuSjMsbUGnEfnlx3bZ5ci8fnhduRfWjA161j
PAFyw3xrVbSkXJTZvB3MYbgHkbJghBKUIxdWU7f+hqyitHPKNyqPvSqUGSCskVLNHnNTUVVBKX2V
2DvRZiXKQnLFE+C1BorMzjXEs7Njf+CR/Q0FmPntBVhx5kyErpY8BvHSuyAl9+Y1JJfsdC2LSzzf
qLruSk42wfEFa7j3hoiZ8HAsQ165IhNQZ+pNpTLuIEHshkcS6ZTl2/wSQdQrNKnK28Mh+Zc+zi8+
hj+VZfdMzqJVyrFjzbOhyOTiYScAHGYOnNXpKazB7PQqDLeeQrp71SHYBqNfv1hLe0gPXVKuA83T
Wh3COC5XMTOoWy872cKRyO0rZHfea6Wq3dxt0+cfReJAnZsp7jqpkyVF+wcqBnVkyc2pM5jU6w5U
15Hz3Xo1uU22HaAF5It6d7CFrPITeyoxqBQePh6mo5/JxkieiqHs7zA2NywKq1XCcHIZrjsgWBt8
KjjooU38G3G107YptLtcwO0pua9XWE/BgV3kRhgsXJlpSwJXJeK8UoM++jDxxD3NV8oWGqQI93GM
+8pHtZOsPXO12Tmphr05gpqt673CyzKRtNuIlvyj7WyuMDRhuWIipqbOQNCjcES9FxT8wBizVSDq
xwrEhIh5OMqYnv4BfOFNC4pNq3jHvIl/0gXMkEcV5tfMTRTki1GbG9d/pBFLXCyQyB05cL79QVMB
46TgB07ZaigJeVyckl77ybWV635t+71A/ggNRbTKLD0dJ96mrpL2qfp1MoEciZmz14c8tbcpVPzO
N0ez2nVRfIUiZjkfOes3au+36KBSYc7ih1NHkBU9z3YBAGsdNbufWyReKf/ZzWVAMfrjQfazNF6U
WhpBTwBVQNtjsARPGlkuNIedbqc/DF61ieinfEFci4pqHDb0aJuAbPqT5KLOBO6ZK5QyMPAjTdRd
9Fs7/zaShLU20MrSnMLMIH56+yPFcULCLbNVKxuX4glR/GA4jqiUTv6BZBzesqT9WvYjifkRqf09
F6hcjh1yv1QXuCwbGZn11oWxfwfBz4c1+YYaJIBuXHGrjfW1pC14QczC+kN06tUbK36CBJXLj+y+
pNMMMtDU/c0M8Z/zbT4oHCRCPHBHEjQJYUyDwhzZHlxRUfSTX60brXFIw47EYIMmfvgnWnD/a6CA
Ip9ujwVvAm5+wNjWSPz/vmYmhCgOjDeLgP22Fa2VmZdoVNcOEQwNZcAi6Q+NlZJAu+0O6LozCKZw
j5X1E46Oktoqy/d5hNfdm7ZCW6juZzmUw+loqFe1BHKlvTwRHsQixhxJVF8wn8LrkYh3oupYUmR2
lmZWTMePUjEZM6j65X0dIScGzvIISNvBi9+psEXYX2NUsE23+O0O+v1LI99G9hCatsCBET1SHO4B
o9nBUNGbWycEkjaADDpRssLECx7e/N/nUx2lT2IyMfPuMtwTbOe8KBntljmD4ZpBtAf5z2vlNX75
mc9QvkITlHwq1lNbykLbJnY7KuESM3wXth/UhGuEN6ZAqDMvqwKnEMDViMx7RdL9u7T+GLLVhSpZ
xgUrkggpFy70+8cWrZQF++tS4mEQryndoy8gtyGjl8JWVWIL95k93ZiGxLpKF1wUYFaE0nBsNhuH
iJWcoIb+oVcedhzJv3cDLQNfxmivgRrKl84D3dlTIz6pwycO7FrEP7o4OXCirinqGfLahXkNClfH
61nb/q/XueTbu6t2vSdujQLYP4RaYYrTM3P+fnS37ZcpP4JDspP4I/apO5MOsYft2derOVUtD2nY
L6uYgV5eM2OcNIngkIYdSLqu/cVBC/JLb9+d+Xum/hOzJjIfLybf7YwxgSVzaIQaiEWqi0Qpo+W3
hw3nnGIqeRyqgLZxIG5cRc+4r3oWicleIldxcVMq5LRED0ZALhsupRBgk2IDklumRCqtZxYZJmSe
nPhEJ2DFQPi0vi7+QyaS7b2cgQg+7CehzuiZjGZEwXW3nbtXJQ2syY396W8b1IhE72bOzjw9odFb
cEiD2XhL32Ht0Qo3X4xGD0z0cqsUT+2bp3/w1OI4KVRH8R4Sgj6qwlogTXqK0AfN21XU+tz8W9TL
IrsuE0TtYZDEua3TdjBMBBXv1zNV9Mfydn6Xisl9hPwckBC9Djwz3d8vxrYPyrrH0JLgU983emkL
dNrAExeQVV0c6a7VL9sQbvR2lpyf/2EHujQdn1QkUmUyr+Mfck5Oj3AqBKHU2BiSrXeRGD9kM7JN
8IqEQ03h2hykaDv+55vOYE5PbnnO0+8JfTE7XcMrPcjWN4FFB06pd9X3RGBTjBxj+2736V5jsmBs
PrYi+mlJsoRFNFMuzQ6s2NAbA4JOSV1KnH4V1OcJSlFjOipMAN2AeTRD7duFdb6qikxwtIwlJbTE
PoV6tWtmosKeJ3HVTe4lfWXPU4VWKlsbs/lcNBtgNOZ3uLMfGlaD4NHnY3qS8q3d1NkO57rjr/sx
1/a9yUZ1DEuguMKKeLJplngXObQEGoALC0tmCNAb/LakUnA9RBEqrGA4dRQvi/KJOE64vozi1fmg
4zoYYXKKoS1W4E6J1etc6BH8df+zz+b6eWDf6UXOphSwhCmD9nBYQs+nV4cB9UGTUrBM84IL4+HL
kytiVR8IUTzDjPvhc41R29B1MmRx984PtkLLt2hSanU6YNJCzEXvfssXcHnZbRw6TfAx1UGmNLyp
Np+ca5gXI4lJ+Ed5LZ86DX7Nry7h5QDDfdI8xTs+MOTDisd0txhgvGDq+QabJF3mWmsmyRdAZ1pH
P0bLXGyVaR4IJj4fgeCn4H8IEA1vOtfYwa2iA+aQ8lmLtuV4IVSE/QjyMWUl5XyRegPe1JmfiF6Z
IE0T+djItI/2vrwdQC/Sx9avsDnv5YcfUrR/CkH638vI9e8JHcStxMWiR5zl9lOqlNq0FAd5AIDv
KomUpYwYRJxqBh2MOqa8CDNp6SYacdxXAC3oES3VqNXIaS9Hrhq+ffxAIME6BFPmzIW+YFNex9mX
O1Nghvu2WMGBJ/Ie7opeYWIxflnK7a4jwi4ePiR6+l6MHRp08znY/e9GQJGYwLlCeMcrZfrYQhcc
3/NvleLNrBhabhcD7c81Tc0De4VYiU/rPEMBmGEiHgEL2aY2KAv7gQ8d8SaRVRVrWq1PvzV8VDMX
Za7hD72nude4INYhlxTHudugGLnrSyctXCGNUv8Mzt9Dgj+7dF6Vx62IEyugqe8Av7KkHaw81O+0
Sx3ez0imAfQXvJ/JHiKfTHTIWe/vpxGRgh2e/Iz9U1Y+S7xR1pEGQqmk8TgbER8uG8FXG10r6s80
4IpqNpxrSsLpQpCvRvGpaSBk95JDxdEDdWFPtcJop//QAVmaidMFmY6S73bDvKb2rNnbRYk8jWlZ
xT46huOZwSjVo4XKVcKZh3piCKVAl9QDiD2XDx3oR2P6M7kx8UDyYl3C61v9C4WGUkivhVzkjP3R
OaQ/UUZW3cugC068LyQvh8qKAlrcY9d5XVERj9QQtA9hEH7Bl8UuCtCsJ60OiksdH0kjpkidPjYB
02hdUiUMrqRGqZQt7VQvtvmBhLdSNnokLt1N593cG1YQrIULEvrYDfWn/Y3WWZeAD7t/hbNfqZhf
G1mNDOBhbwzQXwGUKYoiv2I/41w10en6reQDjgs3uwOHUUM7eXhfxkE8UTq3btE1I12LeJREd3JV
h9PX5lxWxyYnsAx/aSPm2lIJZtG+Vbls8kBG04tg9o2ZiQzjDkr4HauiyRPY5aZ48c4ODeI5yoix
oY1bwQLyqR+NmL7gb/prcT3DDjWID43cr0OZLmnWNs1gDPLJ9C9eO905ho3jJzyo/0pPUaFWOISX
kOTUWfBS2+C8AMwVd5/fFRS1qd0OvStW3632mlFrAW11J8lyHEqdX0hat9aEfCRVXukqRLwj76ac
f+2CWwolHYGE7lYLflUJPRREl5Bfx2XV71hGqPqplpIqfMpTjHal7UwTEQ+047jvz5NLUZexJ7sf
JZkmEJMbVS2jOmFAVw8tUOYB/ug4SGoEu/Ru3wPJy2p6aKTfdCBYMQZ7gAKuDJW+qv4xmXTQnj8L
LaCGALjVN0GcNa+GEu3CyPypUfkXdqUSxxBZ1auomtHq1da0IdkELNkmFTQO4HrQ5lki+9/2UDty
62RTuXN6dhNkJmfxQGjgPU6Tjo3jVc4xbMhbJCRYDO5chO2Kb6rqBeDSEAQvDTkZaKoE8clCvJ+o
qFKJlj/7xv3bItFMyVJog+TBwh6Y9lfXULsRvF9X8DgSqit62DdBnNIQzGHjl09MDtPpRioWUHW2
MuTaOjuEiva2sgRTTRTOwLjp4LbA9Ache1if+3dOgUa9X4yNFshTwVv/lVbXjYh5uupoIivg8xuZ
YrzThO6fB4BdCuS9LPEjhbcIr9/tuMO+Y9Zk9g1jOK/36kn04Iu+zYm1aY1qh+qr1NbIeO6waYxS
6t/Rtm7wW1nW/qV704cFqPX4uzfVob9x0ow2pfa+J36Rai/skq4+0oIG/Mia/GcGeWRe8HLu3xM0
sh3+AI5fmSiv226tp6S4TZweAw/MS7MO92O8ufwcXFZ7uNh2ZLU7iSmxKqNkcij1gNuIJMLWzbC+
17TOGEQXDmYcaqrvD4KFlwlfaq1YJPNMB8g/TptESQe4JhgTUhWMWTZ+Yhk64jQq2R8Cw5tafEaE
gNNsFQIPtqOw/9PTlnOYCxlMsaSBG0Qu9SqWGFL50S9KaNlLWeuysFxu5P7nJAELYhhoFuXEf6dy
D3iQIf8Xz++9HSeV1mY5PysI88UYS71YY56+vHofemElXKtxM31tns0bhMpw6pinBEmPG1hUDpoE
qlIIFgxK+DgJxSbGMweZqtLKob3gOaEaIxfpDRXWC/Ysqyn+yiMCyAoqE0QI99NnKftZIH8joSEd
yOVrVrwp5Soo0CrFb86Aej4vdpxfZosf3fDBtnnTdcJjX+uBI4XNnDpJcLCWyQ6xK2amPpubnUte
nj2+5zYQKevK7+d78OMM4cmXjtSYe/Mbrgjg34DkAIH9LQMx4rGOftKylc68JifX0iMvZPlBqv6L
ZffUCg3w8xWiO0rqwZ9tz1e1zciGZSGmr25j9mdxSYE8C70dSWnWdKeI4rSe+S1ziSJqgy8EqzRN
CF+caclMfMUdugiKpXDZBYA/nhOKoWe3jlJ1MGflsJ8J24jSrm9RbH57bsm+yo26qMhYlir4N9Vn
IgROXpDrsUBoSID8S5qJhYo+ZvBImE7caS2gLp/Q6+cCk3T1QnlhUV2dKHN4sEAD3jUynkjAhO93
POqT4h53KoRH8gDN4mBFw0bYPQabZtnQXOGM2gEt1w4Txpbl0DRJ3PJHDvrwqPkUwybkxhru0EvE
8CbiVF/6CEAfse9kX1AWavBe9Pz/JsGVtkV1TiFzj3dRqc9KT5fBKL6SbzbCmnzwdTnpF1s5rEvp
zQSS8yPIhGCoRNGCMK/EI2/9BJonsZmwlkdHjOq4C5+vzMTOg8Cgr+Fp5pzHyWiV6V+y2Y2WBX6g
LEdMMellTPrEWsvCJtTc3DxxR8KTcJZyfyv4bPms0rWINqGNaVpHq4+coz3gPuSV3zP83pKfjP93
YQ5TKOFiZAL674LxLLcxTMsFPoFz/eHWRVAqkt0LDQP8aJckbqNiGB3fPj+RyX6KWvieLKUMQpTf
EIGaz7QtXVnjmIb5skPshGiA29aiv669qZtt2hJmHjOH9VTpSsLXEowTmZOUMl9nTl0fQubL1QyV
pjyUd1uTVngFUbz3GSEySONJhNSJoZxe4wmjV+0a7S5bl8ajOibeyNikqg846fj/xiU0jZzttmoa
kM8p4k1fO3/HFUBCe9dv7dGNv/AWKb7EPU0va4a11A6caFB4MU9wsvngf4ZgfU1qINp5vIDRuyhv
zXVGlas4Ym+ahFoHGKH0ZSPUnMvkcRUiDJMC1yxBKLQXJnqDVrFxjdZWeZwdA7oDQkb+htOYrDiP
NOS9oRbSQsZZcBEIWwPtZtbnePBIJuPFxUraiO4yIlINQz2jRyIdw/GMFT2x8TjV3QyNAnD060kl
B9DIfYr9m6OTKGG6fK6V2K5NrLWDnHqAbdiQ1ZihMisdPzzBji4sTKWoUaNfLic8zNr4/U5DbFQz
/kPTnERWszrit9lO81gMcFpWFH64LZBJDYq1M1Nyit8BK2RWrH75s3EXapvvT5j2bnneIZ/8C0j7
yA/K7lJMQitKkXjCdpXuNqyOnk8ZwPbuKbYgHfjn1m6wRKYawHqOUE2IzbJgKlXPJSFcpNlP2Avp
xHoU262GpdM09/rV6yiq39akyflScZtq3WEFpTLA88sP2kt5athf9WDHQCbtDwIdi0iYPZZrEpbu
1/l7BWI0eeCxR2AcAAful3/HjIkqrcOJeZLnsQvj/aWN1EMPhIQ+3+EATfgsnqWvdOHmSxuXY3sX
gnaOYuR22rvsJSpKHz+mVPGnE1vEteXs8OVVFQZ+4c6wiAVmqZXlCclbZJejReh7KhsH9/DMoBQg
AfJ4no3xvDNaXIvRtL9Q0lf6/A1+1+MoHk6HiyQ72yhmXdRlyrgnzhu0HL329aKcmixC55Et8cpM
we2JWIYjMgMUBMw/J4Zc8rdEmootPz3wgVYxvTeilrRfLrtfyOPyUAYTATdluY3NGtiQ3+rGS8+V
mNY4CqiGMbwpHtnie1sr+OpDeO3tmVbTmIwTU7QpP8hMocvvCQ4IEhYT1Xrrh0xOM3pLlP0jo48Q
QPEn3eurpyVQgP6hglvvWzUOPSciMM74H9Eoz3U3ugF5aYebfQaPcbFcB1oUBIICNXeCJtb2jz1v
eXdQhuUZng/0ChHmjyRR8vX9f0kRYc54s4nZg6d1Jn44oKQlNY69u04e4kCR2XGBSlfxylKmptbJ
DHqSygtRd581SGzF2ojE0lDhrr20cUHAg0MRWuN9z98E6wu2Z1Ha4jgGZLUAKIDP+SWP/hPH45k7
+TlY7vgh0po2/1eRSza73lIbwkpIZJiT4MhtM4HLDLjOmSl0INR7q599zztnWVDSqivChl+BrqEu
Xk/Ec/CLhCTaTKeE0QYyNRo9Ep0JyR9J0OjE6XUzOljJ7ivfqlO52u1Gkj0v34Q+Ye0nPFiMiiaP
ciYr8StAMlC8y1HuNfpX67EaBRqhuvUMkMFm9TDZb4EJcL9Ypc1YFtfTq4WgUCrCuuX6TjmdE1SZ
h4Ber/jhBdYr5oMShLlM5tctvZ7VDUFT5SPUwmLyrAYp9Wt+MGI7Cax5MyUcPHPVlA/6KNQuioB8
zm+wggUCk4XmfV0z2O02AtZ2iR7HixYhgAnzjJDDJaExBCbVIh1I/sFYjnBx2/akxoHYX7t29skp
AF9sFw4/AscKdUB8QL9/mQJ1iy89KCWSPOnOKdPvxjnASBUKos+QY2msEfGoKUHmzGgCcs/Sv26X
EfGERtPsTyEhZSrrFwO8vi1tjXxhNZuZ6utneIslayXvB0aceKVMC299E/edUcQwao374YnLjOeL
wv20k9ge3iK2wjkSG2nMNrkRQyjk1/eRoQPM9hfADMlno4PxmdZ0aYi34uZiAvY9VKJhaT3eSO2S
z2nSlbRamuHccHMH/2O0Z1vL5ORwvHWa5Wx5p62BiHq0+V6HD0XgbtEH3u6EBPU2yiFnS8R8Bkla
gdtHv8tyjUFDFcVd8RcA1IAXb32yrmzm1v1oKgId+yMeZeVvM6Cm1sgU/traWvn0QJXQxvJ/P4uz
S92NAK03jejPDxJISVvU0l5yLIRJf4ZM5sak6kVMuhwOlint3OdtLXUVWbdJUTueWBdbwSrEM6qe
VaBA5hpg0TEN/mpuxKML7DvgCLYx4ySzY+yiOzYfokyIiiFVLww06f+BGE/57FyEdQhZ9Hs6t/xf
C6QtGPuuwpT1SICVQHBaZp4MK/uq6Vqp67eTut6VCP8/q6JcB3FTDbYpcdALlJ39XyKVDhmOc7bM
VgLMmDC55yWpwB5tr3YATjSCqR8eHhlDDONMnyvPnVlpHw7Wp/9D7gQrb7oYLTiPzOWaD1Ln0OmH
X8xU5pvR8Xqf3jXtt03JvihIMqpywKlrSRuALlVUusGDeKB6oGyzaArjsA0EOpAO61IrbB4Dx5X+
4kf1lCDZGPdFLSzbWxLC/fl69xfVRuaR3tqthOAOyzD3yyujyfrWueh6teiAI32RG6W0W48PAthl
rc1A4uqHBX7LkMOQr2etTAMo0Hdssa9Nos1NfHVJum+LNvayxs4FsQfWLa4KOxW6WwzxdcF92rrO
eZzbBBYBqN2BO/LkR8KwOu+WoN+jVWsxpCUC6uzOaHuF3EpbFzj5IFfR2YEKW02+RaW/8a26gzTD
Rwnp8Ut2OqcfA+F8Y37N4NoOOmwU3X4simcupWhEhCI+obT2ab0xJRAHht4MuRZ5GxK+OlF01FVn
GpD+2JArU+ulLFZoTyGzhEwOAXpE83yLzxmecMds1ROMUpT6BPB590CaXAp21Pl8atlzx1YhFkN6
nGBYiBzmB96SyhSQ4a8sx0ovio+c6dKePsgUWJ/mKd0Ltx6dhp7dcziyar+wgxgENMf+dNcb77o5
+PD8w3KSNOt0LaxvxtSDtEtfInHy/Ettk5AUptMLEzEgpQSvH8LGVLZEeX8EMnQvIFt+pFW99uDu
kZJmWzxT0RpUkN3NXy7COTaSnWS9fDVXdsJq3ICmoz03hLzVBmGQ7zinE3XEzIWnlGvFHeVPXqFR
re3VYQqC9O1/i+Nln7hAtDoq/0eQj+o6BDAF9yBAIP+lr6Q2P7zSmIsbnhe5yaDeLZmGZU4WNoya
501C8txkwVA0lAmjP/fd7jKJ3vsCS+FUPptuJMq/bccpzCLtiX52gGF/eZhI/7OPhqfGq66hv4Ut
P5xM1Fa19KQGUn8JSCo//3ofh4fG17Mp+5SopIo3sqny7mvkk8ClaSXZQd3vEaH+aSZWNilrErik
14DVaBMKe8FMYiJ3wZGkcVkcwYIDNxA2O+0ON3Fy4elYRLV3ZB9gJdo4sMCKtkP3BJe03pS/l6OX
ig9RJNPusJANh5cuxaIBsptk/QsGBmcbzVy4k4/Q+hajaihSk1D41TmfIud5eUMuECu3YPHxxwF3
7W/H9FvaFcySUbSCd3dZekVaW+iieDIox9k/7dv4HgDkikuGUQcHd4qbr3X0FpjVd/ONDa+McUiO
aiU7kRajJ6lrl4gVvAh/is0R58f/Q2WDzkGnqDJjnvBmBzofUe3IR9Vrn/dtAF1g+b4rQPj+FCZl
Qiarrg8zJ0cJuu+6EjUtnnDpdp3RGQYkLAFW+t4Hmu8gJ+mWM/Xuutwp6k1hY7thRzcALqjIZoak
PTgQhHqBN7UmyJjbx25l85NN7p9ymvwGoCaHStNoLYcXKmIRiCbqvOKKK8MF7ZHvrF6CxN6K7e1E
litpKEJ2wXaH7NMBqi2WB77ueAGHhFgreR0h7NzVHTmDMbZgZV5URZqbvdJlNU2L+JK8BFtNnhzr
PowjURqkcx7EsavPU/FcXWJimBw2iBfI1sxTcjVbilqvoc4F6kn1WLXUyY6TSiQ4IgHHMENYRFZI
ytC1dVZ+C9jQZ0I7uJWT2zBLCBMyh3jALMGjcUHDp0lZDnUjEslezd+mwq1rrEERRpAfuQdMRUZj
Jm6HpQgGXvoy0SyTeFAT41wioOmw3Y5CstWGhkaU/aQtqjGQj1gFd4af/GRY/zpeLsubUWBXOAHC
0+rp2BBnF3WnGHOBF78I9LdJEfkMCQ8JA5Cilva94aSB2JUpNCYn4rtZYTbw9XnCQ9Hydaa9CFLp
z/9rU02cpYufhVVhJU7i4n7jiV8zZcgU1x7GM2c0Z5DjFkneXp69fxY/Vzp3pgHQO6HfFw45/2qn
yuYodXrRvDETnnMmTT296cnFcPfiQgL2g0uMg3MkQNSWdbHwdzSTUTIMvO+EiW68JYW67zrnPsdQ
lKzB4DQlxi8L3Jqwq3oJXSyY+GXCBe1HS7M5TDilB/59wnWvzCj9qOgwfdqepxmFzi/xxRS/OLNo
T93rVmcti9r+TvLOq96PaWTpTGYoFDCLqXNHoro9LP6IzK3MvYbXzgM1kO1xGQKNxYDydj6aBBDh
vjZVWsEqwgYv+nnOa2XDfgnKEI+N8ExzGqbPKW2i7CNti9wRpY+yY4JlPGYCSzikmtANDbinql/Y
U0H75kUat0rsO+1upLaDOhFoUBeWxF/8IcFkeMiQZg318I56APgMMB4oKR20KvP4FxwdBpU2uZQk
fC7B29yBPNZUywBeksmbZ/+RuCnxUPp98TxIxd/rqbLq2fhGKBEwCpjX28PWw+0/srXDUxxLXbKh
2U25onKNY/Sih3rJ+48AMh/+sE6wDb3DFBpCkFdcg8pnvVT/JSooFXBvFTCdl4cklCB9jfzzcBR9
Vj7dgvUfv5h++y9QGD4LgZe9JYNrxHZbyT5KMzCLpfaUMHAM96kYTJkModHtfUr+YnlMF+AAncOh
MiOB1iuCh5GqnUnRVlVnJFSCOoN50EYHeDFW//bk/o+wNFt4wD6uAVyMPIr8YWe4IfCAVCmkVwMS
tY0fvjpau9jOmjJKfrImv0RvHJUvXBlnXdy2blGupzwV7jCd02p+IgZge/G0NmfsuxJ6hmt0YfVn
dfXNofBFaVYs+vGGo6gemd0fGm00X+uZA+bJY5XNItH/1qITmjLgmf8dFfYFJbk6QzshAiuCrhZj
8mfX1mBZO4UHJMgMVvTf9N1EuNH842scOxz/ccPalmehCEZNNL+lVzVeWYa0hMZ0iP5ghCwhMAEb
pgpSGBYYLMZI1SUqg4u/ZL5a1jJ5qV6QlBqlePgHjxSdjuxA6myK8AWsK623PvlTjgvZBcsCx0/8
ocOOKioQY03ePVpwuVt2s9xKqxL3Yci+hcPmqAJ1xjMcKavzxmVEQ0vRrWy3FJPs1q5WNQ7TO1dm
jiRUZIh3s41eOYXEkO8OsSf6kUGLjb00XY+rJHnur8YC24p8qZdPbxdKhIXorARlYIpg6qbmUb8D
oxIw6+jQQyj60aGhorlRl+KZzjurgN9o7Jd9JhlJZK2DKBZB0mV6pNEYyR5Mur5rcoY3ili5VDq1
JzbLFS+zKlL/BQo5LW/9NZR8+ukKPGH2Qd2uOx484SZgco07mhMvpjmgA/ebpAyXI86QtOsFXEEi
bGjDuUMw+sajzX2xEy2K5/939Iu81POeLdpsSSEarl9lf4Y41d0eEcWmdJBUyc5C3n09s47iJdaF
i1sz4v7Oc9LqSznt5anqABBaWwmmBQN1J5/J0H4y/fb/imn99SSEgOLoe5/g2M72oJfFQu+tLSPV
XK7sp+zYshrFXFQUZFdQ901JhHnn+6ZZ+YAY0coUJXoQKmkS6i9OzGNRbHqbFPcmqFcliP+Pc8+J
QPc16sc0flkSf0Br1Xj0fCkp0TgFwB6PGzRdcskz+iFu/D4hv2jU44QLEmtRuLeYuvRRG9LaL1+t
/sznkfdxZ0fKa7Vb4PONszQyo0h+YCMxUU+NrLa7a+QV1UaLaYzC55lq4ywBbUWDZDcBqr54g4i8
46MYFnAqAp2CYRPvKS3m3Bj2tKdom/gIgsaKtGs8mUPO39k4mg0MwOQrteu2pzcAPyIE/xA+ka12
Pi/qmnkV/pLgkJDvXIb2ZSLjlFOD5RpLRTu4pOxfrRTlAPzIdvBhQBd9D8SWfpEyvocJCKJMUcPu
Bx40yhu2BXH3lPUDBX6tj4RSPBvModRoMg5iCeFpBzZO9zyuQ/Qds64J5w4EfJ1bM06Y4radgkoj
08Ml3bWp9TbA2wDspGWt9LHggnYjUiG5nUJTujCBUF9GhgZ/V2rw2BiUYoEhipgvAhX9048Liz2t
wHAZKd9tJYqw6hQpzZeXBh4WzSTysgdZMOBAx84cnInIsMowomNQAMXKAbFfX8kTk8U0n0nY2Jnq
IpS7wfatXlnOxY+VtCEw+IejAok+bwLh0kmafu3v3QdCiJ1Gileu7MXuNV0ti7FWkc74PxjVBnLp
BEqrxw55AWgNgPwB4YzmrzyLFfZw6FO3/ySlRScTBvHGVClPK6l6Sg1vhs7OxSW+Sqp2rOR0d6Va
ocU2ry5xBKAi6vtDLxcF6B9MHoiyUQkFmCYktShOEY7HQOv9VXvBC82gLLS4o1pYkfSLKbVTRLox
rWJAbQrpZMHZWnDf2nbFd3d4syiFdumwthxLHldVLz3/7MBRZbNmdGHymb/Bzr7KVB4/8ACjOfuu
DxmUkEMK5+LftQ9uJQ76P0kpKedAv70560bV0ZEFpAbXNPGKyUgJ/tQ7mBF0HIfj4AgTX/Ium/oe
7+YQs3EeBJZKvXg2H482CIkelPTvrspnzDO2/+fZoM8vkSc16X3vMaXwcpjcIA8EP2VB/OUhinPg
nq19+tnlmoQdgNtSAWxE7PZr4Dw/Ew/cpKwogQQyuhvPwrl2KxoQryaLgJoYOxtIUdB5qr++yY36
lLQjZ5LO2dT5UE49AO3AborrpFXR6yIeXRp6OKwsCk9XMf/ad+XeVufifSA66YURLxcZWBq9xXdU
UXht7uCrpyhCOtdfczF4wZ3nY7aQ/WlGt+yl3ST+5mxh6cDmXMCJ/l7kjkoB7TkJ6nj68Q+U16L+
02Gz4ozvvSbecsbBhhskIy26S+dU14zPUZETCYgxqChGepcUI417AS+Vrp7uPt4j8cxoJ9CZPUTE
iqJSSwFVWdHw34lyTy+tJ0KOpknJNX/6dWF5k4KhSlOPU9/ThcCNAtSiqJ5PA4V61a0e8JxHXc1h
8NftE4Zb9naJqKS/8chdTsQsEE8JUT/YLZ4XTOJJh+YkjCbUSBdqOxvcat+KYP3rSzultG6ryaZd
QjcaOeOI9nVgJnfKHfW3EV0WGVfK658nhqkonMM77bgUfueNTtdIt4JWTSScIMmj+BgJGUhg7/yc
nbsJ2ONsm/HBYful2cwlWZgPevNZjafD8ICGeUMaEXrYK/7qYV6aRUOWOIIlEqAu0Z8K/ZO3vrKx
8ywX73/crrPCCy1Cq1IVY3S0fAt6awuhbZ92N/ZNBmr3nGxZbMJoAVIX3qQWSAEf9PkSDMQhV1ZA
S3ZUGSb/I3xFB5GrMbeR2WcA0ovkHH3vB4ie5xagb+oy2yMUnHwlyu7DIazOBnqB+90/k3UA+PkE
XBtggpQm9Seh1QyQW4LboO0dWrafTpKwW3i7eM+kewJWoZ2V3l0WFSCAnKBPFk+70Q5zowJbcczb
W4uo03dg0smTXL4GM6/+7kYnsG2CFr7Shc/ow+aeOqbiYT8jq15LwOVvvqGGq3fdsWniEy1kuSd7
jBiDz45cpo5Hp+n2HwJLybXv5Cb/FXBdArmjwMStYGKn9Ws6Td5gbVBvZL8+hd07m7mENhq6p+dy
tjlEkp5ZoVMadjgftdtEztCzOS13+P3P5IrjokKp40+GGgjelbWaIVo8adRXHe+XyaQo1j3H9R7l
6wWuw1kNvy+FDu7sIgvdHoiIuHTQQQWGPpJD2DAsXFbd92RiWTKbXXE5mDhy3FQlk/zK/1Bu9GKR
4B/Yoxybc5+5R9fM7widlvB8F3fK2e2ua2lUZVPatPAT3Hu4ZLOcm9C+PEIgp7dkNmyZ0pqH0ib6
bncEO4gGWRrSBzZAcJpmdofQ8vc5EgNfLmGFgJ3UF2VqhN1ZKuT78uaJo2YqndWXBccigPcRqiuM
J2P9Tu4uROFTbBKJpgPGHvWq6z+fbC3rOv2zDmvkQOoR0UWJ7W8oxrU7Q5ggvz/mbszI7uQsPi1v
WSfEHBfqBhT3QX/+Sd5tYTbPlk+zmzhaqG2GsZK/IKGXZG483i7jcsuAmo/6tnmIvFxZ2uuYiVM4
PftS/hPnaCJlAVylQkkaKw+TDoZQLHZ0H4klWgz7rrfRzjjCmJf80mwYcss+ztI8ML8tpXHYHmay
0xzqdT8Gi6i04m6equsmkhwd3S/6+7fCCQ0JOoxROEeAhPlZhN0sK2TPwl4cNHDhHRQ0zQiRQNat
nWdiBlo6yRgEMfptlZBRG1+KZkH8+FCR9/8HHHUdVTUbGwsLyEVCNti2YPrXCdwWDd1bm+AzufLE
sta+agD1l7RYylxg/Hc8y17n5FJTz0CozG15fe5nuUjpP5evSdXCWV7DY2Q5oWL53DemSRHnhclV
pUBoK965irMXEXnf4WF4xpkT0YIaf13/C7DBEvk5mG2yVifSRQJhbPCKkZHWtbtiH2Yq8g2G1bIs
pTwhCWBNYgUhsHhxt4IdKJAHZBtq4nnUWxNaDGyd2Oehi/aC6jgBdO59XdKl5uDjVhmQYrQeKo1O
HXg3nv5UFwqwXeYP/zyMh9zjqX/1KHZtePPCs4CyuhI8j3/n2cCD86lzBLIbEAIN0LMGnyibgSrV
Uxp/rNyLpPpset0Aq4XO/cvXAqzBKjYenlONUmz12jf7iuUo4IlZdjQK5PSK7RyIE94/mLWpz2Oi
3ViwhwsBhY72TWwzYXDZ2wxUxJyPigLeQi3uYCkxqP4xV5uG11vPn4PKELRNz4oLDiHHNHy2FVF9
9jN88+0EBtz4SeSIx24Z0+lPwPTDs4tSQkxC2Vbh5vMjMue7ifFWGnpcW2q9dAxEPul0+Wfxin0n
d18uBPWFw/KL/c9DqrYxNUi5cK77acwBvFul6Ffk0+Scs/kUvqxI1LynOHMGqzrg34xlalk3FN3B
vFq2pXAqK+L2A0HPMvv3ygW3FLW9bMI/wtaqpbq2Y8v/h8XHBaSH2wbVhAlBHQ7LMi/bap409ITE
Z4r2VqpVu+D8ivG92oTfOeO37tlZPypbRxrJUumy/ywu801VKMtCAUfmdSgYW6JwFAtz+rhzPzIh
TFGh3qTiXCKXJo/UB5O+WJPnSLbETmEZ7rSxe4MQ38hQ+EouX5vI7cIUeZ8nm1CnX69wHy00mOFc
AHw2RUUiinOGqQTRT3Zp7sixyrpXqTwH83gjSgBhoOxoXXG5maRqVVJGPT/qzd0SJAgjhjwArMJe
bQbMOzwvYwYNoq+rVHS2/stidr5vMRXM6A8w/U2pQOghCe4BKS4rtlaYZK0tJwGUsBMREiX9WaN1
PMPL7I7+mTW4ddiW0GfAUw+f0aq2So709aP7yuv0Q71HAnFEevUhAyquBz1Zc1I9/Hgc8m3xxAd2
lfVDEOjW7K0zYxRqifzbn01LLHEwWrnfP7k5kQ9DxWYP/C3JDenGXNKDyYb+5Bq4jRdjeBHvxW5t
M1itas951IEhsBPEoMEiVSle+6nLMN0ZdpZFzZeq5dU8HkBjxoKNg1mzpjXF+zYycuGgqYARlSKs
401WN/k2PlX2ni97qD1AsiOnzVANaE5oYvk1vTSVKZh8bPJWAb+asJ7lyQnUnV/M/4aRS2bgG5mx
Ia4lLHlWPOvQn6yNddszN/B3oUdmbh8EXNm2riQ2mOFPFvu6qKNbA95H033QW3j1d1uiVY2hmB0B
uMaWPmCZ4qGcObdLwJgo28/+Gbo3UeqSPjgGJRHcS9IYMcOvT+H2DKRp4F9WG9Y6ZZKQ/wcQwFce
Ukj9qjMyFvcFJLtwht8CCIrOM0Y5CQ1Qf64Di+LKFMdol4ii5LOfmSU24sVVWZ4NYGcGf4YcXdts
YokBdikGB7VXY/TJpMgy+YmzhjUxl73f51SCgAVQf2dnh8E63II4d2nHRtfAwLnqNktxGRk7IgRt
eEKqq+uY/rT5oh0oDezot6Z87CaG1LLGlBdlDyu7U0X/W419kJ+5zY+tPctQc4bGDeAPFzwLndRH
RlqQqHbp6Qy0PcSPvgFz+ZMHCkaaYXWi9urqJ3j+2kzickddp5JyjfXu6m+hVOhCCxe/N/h5sfHL
HHkjinfD+6RlRyo7fUaP00A8r70LqOrKC12r7U/6sX0lHjHBtD45rS1c9tRvrBL66HH70shrTSG9
5KEJYAax13YJEtO3C7i7n6nsWrZrLinqfM4zgryjz8VUgmXIoMUxG92oYp+NNUDaiFsaTgouP8Ew
c5Ep9gfxe2cywtwhGOj377NYH0+tC1EbkEetbqiNDO7m7+1W3zgJ4B/g/wU//CaqAYaHFBqy4L4D
ODq22EQo4PbIlcaEzTv8OlsyDxUsZnkRA1fQm5Ob+zirBRNqCBmrhBP4gSN7ig0oNLtC3JOqJm15
iLwGD1Gw0CBMeNSoJx/W0x5viGGhRTa5oATlYWwvbfohG5Q7BFS6EpoHN+PoHqAoS5ys3z0T2Xw1
WLepJyeAPNVT13j42kEk4J4OIK3RrN/8wR1U9F/vXij9Dpqh8y8jWLNHI1+R7TSmfOocWb/nHH3P
PuixEeouIg5jUILy8tycAkjXMjgE5sjIYAg+rYn4DlJUX96M+IFQDIzg0QDl3YRl5FSkBNgHnFZl
gQthekNVP6ilqd/LHLfM0tgIUNBrpXscV6WcThax9l6UQUP4tXNNO80TQQnnPe2k0pMjiLPyjJ6Z
6apkWWEMTcaG9ghXPkD9lqNKLKSCLLC073OenIqZxKdBrZ4V6hVUoy+fW1dSTkIihwqlHNGSGj+T
pC/IjAKdNQpxt2jPxsLmF2/wRetJVuHK3OB33Mvz/OWpg5vro425YrTA5upothI36MFHUKgbAz82
zZ0i+3rLQL2d3t1g5v088yTjGNY+qmno/81w6ep/vdamqxvBdy+Fsy88OjjDxL+pN4J7nHUakB/l
bJWQZKqeXdBIO1246uriHGNtALtmh83NHHMmnumMBTTh47yzVYJ6hNF2YbXm+8tZ41UTAiruEt0P
bGijrxUXps7tFLZWY83++dq+++G0HarhtZb1VE8JwrO7IN7e+G+v+A25/oHUmtkVJrVVhzNZkLVa
aBPGbQkbbNhlPKtATrvGpOQi/OYk3U4x2HaKaF1F7FZpbUBNfHU++4hQrSvR7RcekXerw08pKOa/
ZLGaM21rucUfhlp3CRNzmdsN8Q0QQ7NlKR5zUuY4x3DsK7uuefPB/aTqpDWldKLOt9fVb6SdW+f5
efg+C1MRCSMDeLSMYejdru5cOaXwdsdJBRhNW6NIzG0MUjQaU2/V+6Jul/xVWir/NvD6/B5Zudpn
79uqQhcPIecQOHiOVw+X/bOUnlPKHHM3goXZ1vIPolm4+tkXZS7xx3XCWYXygeRs9yY5IYHBugaP
wKplwXUOlH0KbZIF78N2NCGWn+Qlyo1fsGdSnYmDssdzFaqYs07q10zWK4/LtUvc7BkLIr+/cPuO
vAQjRHzRIDawqdR54BAiDO2SVzttvwgN1c39S7a/KOFNuDJvz6YSQJCwdP/XO6JrH8FimpRTpXJR
L4X8BuHlVwudtn9Wl3KU0tH0+SdOcASbsWSGjeb+BbE20Ay37xiVRdXQN6VA4wi8WpAIn6tzhXSS
7E607G6Kyhz94Ut5/TIGpsEGp0euC6AwSwGT0DLr5e/aQwCC7FrIpGWQoKWXMXGSV2KYg6clBg3d
Wzf7nMJI5wv+75KHCA1uQEk4W4OcEPH5zTwOWZwzlVgVESLVtm9vQKy7Uj8PXppi0i2yYzoDUPeK
osxCIZTUttYPdqdCl3f+v3/N/vMD1gbzbvTfyCqLpePhjc/Wda/gyAp6FArp7jHE7vFUkoCdfJlx
1fqjxVPiztZbOIVogTgw6Gvunwp8h/Iy70lUN2AII1OsyL3CDFIRA4vEkKOEMKC/tL+zknOLa6IB
42lzcbIJmARgxxq9yHS8RHmbCvOaph7u9ZialU9SGFYqb4ZRl6Al/5E18y51sMlWNqITrlIqRlh5
AbyR+XCIXw3duAng9PoMYAffYrMsq2BbGxwU5uzvcmAQN7jUZSeP2Oc7Ug29YAL+vQXxX3j3HcKI
oSV8u/u0suRQMp1jpxG9N3L/UUVVxQ+mGT3w5YN9+9rmOEQ3Q+1XC0lLL2O0iUXvEZp1Lgzh1v5K
vWoFgwFpuFxUaZw44DbwYIpYy1UMj7VcZWCBkNWvg1qdmY1saAcM7hTFxAmxLHBlg71+f34ImAoc
KF3VdsRoZB1+kAO3z67NDKseAWF6MKgUKZxL9jnwV/wfqx3wVzKJ7iAcYNe8/aJf3FUALywB7Kk5
czEyKISwE0nEge9E7u+SPI1cUWhHNuO9aR8kiutnTW82AvLHu46O19QyNB0g3xb1HpJIVI8kfhjz
kb3774QYzbM8Uhj2XmCOM+yJZYmBSfKfSwhoxetXsZhkxkyFBJQT+z+Fl0NTyKRdf+gQVvAuM8dX
W4Z65HudAdnpO2OlKHYLYW2IMr/BPzSure3qPSaiMl5lH7Wt2Q7ojJQapBlSQ5ukCuNXb/4QpTt/
DCXBoQd1kCZ3rY5eudAAVi8cdIWCg8gFKZfEVtM+kg1z0R944i5+TGyciVZ9kvFpuVnjL8Vb4/Ee
wrL2nGAJi2xLzk7Azw0L2B6CYZrjDoVGr+uY9ReT878gsTWo8iUvaX8cODqXlwqSL61MVxMW3tDl
f/ihoDLMfkv4ajCr1u+PYog0JsSBb6qHcfpjJOcL0ScrGoMJZUzHdvJ+jVfW9lAcnnrdbfbxuQq3
Z6KuaL49Mi4NC8QZKQMhJJ09PhnRWIMo7MAcQHfA8GHQBAgD6LlbH+uZ+ABWfBL7MF2Gp+8PcLQb
OfSjn2ihe7qTcz8Yu9zMdeyYyXLaSTFVSffggPFWPkdFvek092JMdegxZlxBHpSHk/xg2ZlbC7Um
YvFd4HX+/SVZRrhkOd6gEwFaBXNYUM8aJt8BCU8sGZlA2HMWXd74N2pdN6LNvRtHPieKel6rDLY3
h/yjvFfg9lftQuPmwe12WfWjtxoZbsGj7J6ttOS5DtSvgASWWKSFPs3DReDrwklmCym64RXwVxzv
aD5a8dTEaeV9K413yLe9tXJRP6+baTEC5piJbQ8NcctM6W7knAbD2I5Kp4/xJkGFgK9UI4OnY2fA
Ajtths/+ew3GqZXRdMjx0//FE4JlbdEfT+mixDWKSsw8uvV2ucincnN8resBzL3yqYCWGXM9wOS9
lDPMml9p6UzX79sPoMsPrLcH0t8EkS9OUwEXRlBSU/HiJqVc8MDy+xILQYGgWVSLddaEd/IgoHcd
qw0222UJrgx5aNly+PZpRWWIYXSwS8mF5dywf+r8kDbx+Bn4+WcqHiwizAvuZYq9q+SIhopfRsfF
sg2gujFBpAcw7c0VFpvOXHngnbahF2bHCgD7Dca0RhP2e7zsLokZDMnjMzJZVEHcFXr72j4IfNjb
ZiVqARc6h2VZnWiYDS0kParvRIOwdhCMF7qDxGvk/YYZ9YUKybPa8+wOx4RwcBIyVqgNBeaauD6z
sDoHuNlir8o1QXuHIjJY5MnCBStJNvC96pI0La6MinxpsaRJjyMf+D4AT+u7M8cMzoHZJjKnTRJI
cLynLOMET/p8ACNmFjibjw7+Opw2+XERQJms8JPh+xloyKVTuRRgr/sgRGMPJVMA8uJlJgu20RYX
XiJKA3YX8Brx5XEmfcLs4wKaf87ccg37nGqVVUO+3d69r8bbO68ZiZTqNoWkxBwhBUMcw2rNr5PL
yQVe2gpEWqUuirXG6gUUIJH2rZP1bGuV+4qgSdGGDmzeg2AbcPSZQmJ32qzoFxCZFm30kNSZzrlx
09GZiGq7cAwibbiFe1NMY3EAbKg4AncYYf7R+VpLDlsxd1TTjPC9D06xy3tsEW5i7+SBDgxwy3cn
oJd4yxSpOdt3GDM07rLml/FNk2UqMDRpJDZrKAd67eS/nqoBL1RgnsAHclazFyWxDFCQXOz3RXop
YyzYIUjQeuEgkVxYXDrWipye9VwH43o643Y+vIIZ5xcT2C80BCW9kJqkEZI8Vj0GuwdLjVQ2i+Yz
UpwmBaTTR2AS0pcvt7xzupTKEN84/ytNIVxp8chJp4egLKEiI7uw8xdoylqF+uCJiS70sUykjsog
GHYtvxigviD4P/aE0jj2UcyXZdRPfQ8ZMtLZRnnx3TKbxrwgKIJyV3neXBe8GU30OLkwUxYsvtgD
4DHskVEwhbjlyOe3VN7aedFuHE3Lzg/V2D0TV/0GfB21jOx8NEIw0exXyl7K3m61Qn84TKTBXT/A
CesS8IkvpKi8iImTMmYhl22W0Hd6I1EHt023h5wI9YiOW4KCNOSJgz2oRhhliocGwYpBLlT7Xw4t
1NSh6RZB5Cd4T79cTeL6njfkOz/f+VghiQZbJmstUqwDPdYCMyxhmH4eLVyWvQHtXW+dgFUGYGQ8
0lQWBSEyEnYSzRf3F19tbscKNfgHwldAvK5AvzJ7hP9gcG/Qf5wzoHqlNtZI7hKKAULyMc1CpANc
Bfw1WtiNUMUpxwmsYD/kPyX3aLOgCx1laKBkVrQdGr3773xkpxelrxOaGsYbFKXWKOkixzDZeKRR
0y08CREfcGILdRU8pOEWiX15By5mOOei5zKAc2fOYbcqSyHz22q/jhNh0pk04eIsTsbM+DO6a7Ee
haCmliB7QTM+hl5A9tRHac7j1XQKs735T7hr/qFpa9kAHZZLe9/AJF+yeWPBwiPcpXG90ScO1iEa
aaes5J1W9yaTRyJqAM7RGBCzKXXwDZXu8zTYgwHGtEWB99K6WprETxuONWCWQKrPJggh/xet03P/
gq3TrMjniUnaJJBgWKMyNgtkMna3rQAugBPeV1DmqNPF9Bi3eY3v5BdSBOR1uDNchs0u/QIRIUJU
YxgrR7+Tyvip4gG79f6pnFEAA3qEtnqdmw/RllAbldPwGAP8B8xw+YSC7sACNsHV69wyo5yyOe/5
tT8NiW/Ig4pf4jwpuBiP9QrnSpHNRshTVoQn1ZqgAgnYuSzm95mO9nGgohYs4xPK2lPGqJZX7n33
Gbcj8oSaPxY+StvGA5k3Nk/1nxih3sSnl9OBRixkV8SQFeUuJGJsnW94y9CHGj/S7hnpwjEpOPOn
0dB2eJPdWtEN6nyKxbDmNyyJ1ueg2uCcYViVU3Ur0rc4Om7oH7fC3g52D/DJeZVYgeijb1UgfYFL
1KvimSED1smg1l7SLa7yMyLfJcz07w9Xv4sc8feCSjRMrHNbvwrD2wWgHJyuj0dAcPlhccO5gA7m
NV0uSpyUrYSKPrQTNp0Nv3CczpGGwmCd0NIyEE9iuom+6tmvRM22YyfUtd3CJ75ow6/6rvf4LC8P
RKkNn6D7MLHKw4keETK5AeA6+LVGI4M3kirm77AuyyeSSq/WdU4R8VvnuzlWeT/Lo2f/lXaLLQCm
5490IvYjxKtDGjmM4o8HLXyywIunLA/aYjGl69OXmVfEz95y6CAoVjqNHRnGYisodurnvXhO5rcW
iBhq+F68JFYu5RkmWxRRu3OAe0N9FQah+zMd40UACgf6gi9qnQEsOMrRVYv7/iERPVQ2SWOd26D9
GX0xnF4EvkWGW6Ox4s9uqRKBxpC3qhaSmQxT46BNfIRg7JDQ0k65XM42TJv2HnYBrpXBf3FsA7Ys
aF03DD1zmI2nqL8qoks/dFk7rmwlAUBrWrrDcFjKNpxDN4mntWRQ4pvW+p7rbOuSvu7o+pz6B5Zh
Idp8BWNQalE9jnnmwRVcAYua+9Mq2dvVyBJI/fYWKd0Xj13vj5QrkhD0Bm9qG9htPoOBcm0ThSA8
gLMvzHQy4Oja/fUAEZ2MjuMLKNOZQeZxxLsgVskiqeeECIQ4sr33fkyhJP4QXUh72zyFMcmi4QIj
ym9ZgDNEuOD9+yjvkOSkWWFBBtO1Wmnaf4XFLZfKt2wjM/j9tg07nVgx59FIkNx49tLc8+769NBm
n/79NN/Mcdg2aoSPv9HV/9joQUmB89cB1oXIYTxnCIeZxJnBbO6d+QpGhSgOGnNGK22CtXWJ99l3
PPWvJZUiCp50OJ1tYxnqegWk1ftQRdvKclbH71kVw9n6FGDlbcOqcvpP5Lo0s1haT/NNZ68Qs+25
8jsEHdPJ1FCmzHAgoDktCQEhJsJcyB4+EkDe0kWQO0+WiMaIof/KdUdXyUoMsyrVluPX75X96Klz
j4D4VtSqqanWSOEhWr8OlDGg7NK9Z+mXWDhvNocAb/f590YbUncM9PTUo91oLztlsk8r331ubTUS
SRpk2v+nQ4bC1SqTeybUTwN5Jjb3Z37LoZxTaB0KEGsxWrzthsdBm5Tra1+NGbNSpQqZpRDL9EEI
F/CbdpGP+fnNghN1XGZw0px0C54vtduiSCzH9wdZ0AO3FPKOZgNeMiAYpRmEuIi8+fjp8kpakJAZ
z+uPG0nLJof71pEoGD9WFhkjgrS/3zygsbcdFuIay0WSbIDQMlngMU1GjngI/6qEyhkUoXRwr44X
cdyc4Uo5VbGE+9v8dKJcVtUnRMWgYd0PmntdJEDIzl1PWelCLQOLxsOpFNKJep1+1NCm2ojgs8jp
/ws6EDaVPdFLEGg6RDQ/CSfQy3d5yhMRBC9aQANX6j+X2s671ckQtgzTlz11z2sI7wOXW0pfm+0i
T3tB3fuNl4g0yOSUdXqp5zcEdaTY3H+H8eTzUhthaYpJDTIKfB9ETHYcJ59OjJAfZkfDwvTVsub5
dufCaTq9FK7AS76bJEQyaa2dMVIyhn4VLu+7DP4s8fwMhu7/nuorwdvx60d1zt1G2EHIJmG97d5o
XydUJcLSZcafiK3CdHr88vCvyNziQrBaFDcYRq++ccUkea/IE6AGw5B3ApIQpt8QYko6bHIqo5o0
uGFvHb6VxHSvCCHp+Ic3Q+QiQnqhYCKSDtoMhVM+jjHqmU0IlTlpDUarpM+3K17MmarKqMKkF8gF
PRAPpR/u8MZuFscLZszrwk82PKEFy31UGZACkaqGN4VACpn10Fldy82jSynBgAEae41E1zylzja4
e5SC4ixQ503R41kct1VayTwuFwxb+uFaag/NkOfsMdIRjJOaPkBvhLw4IZx+c8Rka31+vwUmoqWp
6aiDBs7Y/0gXVe5fDwgZlPmJ/+WwxNgkvkY1vMJbpx8DKDtMKH/SgJwGQEZ1OjlYA6Ml2aBU8irI
0sTcFfCLNRkhvlyFkjk3zcukUi+/joTMM6cCgzLUKQHBHfDhiSzVojV0ckSmbI9g1hGDaYrqautn
/OABN+1gjt1uhlsgL3qfS5bBssXkjcnSvap/I8e7i4RgI1XWXoMJDzS3qphOW0ekXRW3QhRwqty/
Lo47MpyNkGQJG4siIJtsRhPEkaQvAAin5p36f+nIcePFXfBSJSm2BVB7PkovMX51rzHRFU1v+aul
/i0eEsgKBlVOmpKUoNE1lfiZ5FTi99W379WjJmrgmxeE29Y+f3xTgTRIl2WtD8+71SUztDuK+TEO
sic/G70dOE20tYZsUOY4YVAN+iB4gthYW1jaaI0OzN/N00VvQ2QxKtDMM+1hYrf6zQs9uhi/qhYw
kJlyDgK+gfOirKwhq7YhgWKnZg4M0NLT8YyHOLRKu5zufhfRq/cR6LFUxpKmulULq8gtyV0A85u/
VlHdPpiwM4llUUaQ0JQEdNvMAgbeetwsR1lXHrVaucJpNugbvXG9MmwyGAugGfcSAvAtvzIeN7oV
yPW4L0QdkdNZWrtFdXKdBUuqaBS5G+17wT3pGOI2zSD7kqvrXASWXOrQHrQRYCyMcthxOG4d+Hfd
SwfarnnF2GjbBFOxboB0lseouQjssCP+YBGgWJbl3v/lxRrTntLORVwEzy7tjEIMD9kSNWJ/xna3
jAI7RzpDvGEaRarc6kTvpS5yF2PCDTgMt80DB7P4JFpT74kScSEx6ZOjfVOvOQuC7rtpsqsUlVG4
9q5Tu0Y9kJICNn/X1Z8TnMhsicr+bddvGnonesl7UjPmhmPknlBxs/jnqBjnGMn+RS0jMUaWtXYQ
kim2C4wIvYvgjbsslW6lMiWwrU6C6dPWEIwBDLYHiybybEOPT6d0IsEBHWbQH7H6356dPQlOHE3/
2TlkbVkvcuxU6vQuuiGsp4WPb25OQKuROiF5tmJLWTQk9jus34/GuS3gFFEPL4D7Fc0K6cu88k6z
oZ1g9RJIkXqQeX/Drm1CiaGgqSoW0iFJ3YncSJlc+pXRy+tapDG44E5VwwHZ+rRo/zReuug72WCw
ylGNBeSnAz+KSmHlz8qTIDjsB0wBOoux4crh27oZGuD7ixxHLFaqfUrx2ugLzMsMNesSDwlJeYwB
bcgqZgYAzqwMoMQ4Gmh+EFHJZsyX/BqPmt7erXN0TsIiuBkXRNfFAZgx6XTdgxXFp2EWHkj9jceB
A1uBP/9YIl2fSPvp3HAPwAM50s8Ho4W/+vBzKDfDKYmKzSRepxCXDlTYR8Eml4cQvGS4TCYGTPrF
6a3kA33IueY9fYfT3MttXU55sFO7iVkDoCmpD7WX57FJCfEPWQ8Eeb+upLDM2eZ5m09nP5CoZnQR
aTgPXure2wW7pnLgI4t8OIRa3+z82tYrH5/28gKeWt42/nLhtvVd2AdKdSQU7PhmUKXUq/bGidfc
Jzk+gXj1zYPi22RDKky2kwvQZ+6uABKTwKb5jzmXKZ6ywxLEeYCUHCRWtJ+/FOEuob//5Kpm+OJ2
VVAnogLqXOIU+av4hAaRHDjOeO02njxfdMCioy+nQjuvukSD9IQ+Jkec/vkU6/Fefht2nuC6CDKj
AzdXODNqI9Vp2GoJQEzlkXMrR8kLr2wQ3KUwdD/qrNfHyjh5cSLx+8hFyOpo3ZE28nx2P8SYoi7k
jSyAc8Vep6vq4LLb3lFeZknIzNAOnAHt+ucnNTB/izjNa4iY8wL+tY+bm2byShVv4Pi+rsHezFqg
PLK9RVt/NF8BfcUHr23KoeHOLe9heDHWEzhu7MYVxKThB5g0tMhpYVdgH5+7+jb2Vwtd46Nb2ReQ
R2emj4TIFb7vsPQb0220BSF4InkWOgULp56EvbiEajN+u7sDAu3rnz8aKWhcVJU+Qgn9KTHE+Js0
0QXnRWX+KIdBDgZSpr8LvMOe6xQMvycj0zuQUgfFPya61t7zFTFCeRVbYGvqZKrFyPDIFx6YO2hN
+GLDEcEF74oPcY3oAkSyZ4DoK5X204+/ca8dPRbdTzxCiMX+xZoAOPlATbzKwrBBWc4spHv4vu1B
I1n1wDBCEcWmnCgflkKdQYHKqfH0VKrRftZxvv382JZaiadwRB/vOocGojYx1u8XXO4PNl+/anuP
a1DWZkfX5ln/a/OoyeP6vcEXBhelPlRKJYOUtiDr1qyyXDBPqBO8tBK5pRXzZKotPvyf4m3aCIbz
oOcJrP0yrt6hYVmmmTsr9DEHSXQ8i0WOW5+P+lMnVCQnb81KgHoWQ5915IUM0CEaFAAbMnMo9aj2
6Xvmvzzo8P3Czl7SOiRSA6iztKWTSWoqpDVfTZzFyuXHRNOXpRerBl5V3vQvkS3OexSU76SSk2ZD
YjDyp7N7KUcFtpdK5cVmIHmr1tOuP/mz3SwQv17PWBqkeD5eAn2sQQjK2rvsl8ZiB5URbBNZqi50
s8IQK2Oree+9Vs1i5TfOsRjUJp3onxCjqlYDTLDlSzDUTAezVepsGeRovohPe6/NUbRzf05pU5Fe
1uGYc8+G31nj2VNNl4qtbar2lLSE0nHJ76F300GcLLzoqnqBPN10yl88umXofFxZDYmqGJXx/R6L
BK1yV6xXKbJiTgYIS4g6Ik+tuLZGJQoylaNRwEJJJ5DtjPgF0HpSNt+2NTsal/HpMghnCQF+FgPw
CtimsP1kA/wrM0PtSPYrc37bXZj3KusZd3NwFm+JPf4uQ4aPZB00XpSPe/sedlTNpcRJxsdR5fk9
ma5PXl/Rof1gCB2azT9IUD2UlcTPcFGSP4MUCXtyZ9ZI/xfzEr+/SqvQ9lTtx8oCkjhNdPgfPnLD
r95MWjXugu8zn/0bTNPn0t4zwAjpQJBJvDUHUFwt7/q1Qcopwku9o07ah6wWh8nfZqARbzQzRGyl
IIDJaUXu6BD8eKXYWEKQr++ULLtL48/FHqnYJ02F6HdwnfNhzNY/EXVYiXgfu6hdpkWdBXxgZcCv
NYwLDBlJxzntvBwEk/F3asM29iLto2CeQ3/jIgc/8TllLa7IbVhBWTxP4+DySNMHH+xwQAAN/2c7
BuVERm6+scGm8ty4GSVVXBGAl/75ly3OxsxvYS68MLq74QrX/gG4yaCWfMptU13xIP4khMLa2/TK
EA2niucAF2Ny/9HCQv2iMAAMrUyL5x8EB8ItmYTZIBz+D2VDqTTvPtAC7VFxeGJffFhbid6BbG8Q
TiBczTSOlRynS48MJHQfItwSvzy0JPRkauNRJ+FINnQiaMOf1RnZgzGGlWR5Asco5+QP6OB0xO2Z
eN6VyHr6nmqq3JMt/mGObCbF/Pp9F9wUEdadQpDoMKlbFUxTDgQdbES132ph54b9XIKJC3b3Ym12
LHOTb14Jt1DJuBeNLeQn77RVL9NZhs2Oet6gMeD1f0rZh8RakWm2csavBfnYtNXh4QuU/epDLw7F
NiHcTlnIvJt+BukIglA5nfDNG3cL3yzRkErVpWy3ShZnr30STwVLWp/rvMVPFAlOPNs1AQbYGK+j
no0NYs3O2LV489DrmwDFbmdDVEbmmkYxUdLbXgHH0kGSUk4f6rFBQmiwN6eS3qQC8Oayhw47el5k
KhUvHUVp08Wxyreat4gyQl2BLroRelXsfCR/EuhKGJ/8+F9DhdukRAc4N8JTo9cXbFyvbgnAAS3O
Ed7wzn6JqMHG82J5qpf2pWofDyN94LMYsH7Yun85RgreSJi/DtMkBjG5+5YSc1sM2bTdCV6z8AHG
h49J0KeUQKAsGyx4hsWKzsl+iJaZMdcKCNF9rUNAUY0s3qy8WGWSIKURK2dC8rVicbqgN0zevhBd
liJi+H+N987XQLFCLuLIRe2kw3VmXlNOKu5Uoe9S2UPO2VuMurxj7Q/LpgtAXbEnAZ/QS7pG6HzB
4ijKS3/r+C68LG0Z/PYTN9PGIXkgYb3ZZG7x/5luwzimZuLQUrCOjvSp+THdwQZvaR3X47vnX8gb
OuH+91jhUFzWmQDSFMK68oz7kGT7F8+ldAm8XYZfDTF24h04dum1Jbi6vrZGUQ/O0w0QYT13OQsV
e33GqrUDyD/Yu/yFjEbgnYonwWHyg0ZmOIhaZSBEZHCKhE4NOPLY4a9vtDMl1iUIluo1bPXCOilP
mZEtaGeTLi5feZ0bcGeHi0Ig7gdbXx9ypd9jul59A+SRd2TjzQurCv+UHMm+Y5iG52WhwHG38azy
+B7j2bwHm0he+n/0JzOu9kUt+/OMjzsUBxArk40CAkeWXumpuQqcx9jgPoMLFXONO6NKRkwxDVI7
J7scJ2XZrIEDX3LmquUEcWUlVJcgCg1gy3HF0LwKal5CQAcbugv6qLPXsrHG5VrCzaVT914MH49q
BunUjLGX1yuGqAvZwCXUme8rZZ3zFPVRHPFEQDT9cpbtHBj8f8B7pvgTMR+Va3yWwtRZZBSBNr1I
jHxd1JMUVkhlkLEiH6egxX4CkmPyX7Do+o9Pca7V19cjHtk0DGwLuDagtvGoD6/q3Oq16ar1pSxL
Kpxn3+c5ivjNZmn9e6Giks+mPiFS6ykUB1dSnASLbZ5DGuw7V2I7h3T6lZXzVMOg6I+kt0szWOUg
MzeE9KO1yhwSUotMdkkOoN3vm7AH2guFdnzWslt8hbvx/n8k0o7b8zIaOUWMbTRJXLonqlxUBs0j
4Qrw49UTHXS4/qhI/IHxceVnhhaO1Pb/JZcYVehbvuzu1o5ffBfiUh3V2XjXR719PJh4ZDZMH7W+
IdoxHrnrXlzeJDCDRKUrtlzqQK7uadrKasmMD2qnjyXDQG3B6PA9uq9jzi4StHcIPlalKGlnqq7F
lZ2JaecHNVTRAYNkRiWRKzlTKkSxvdzuNlDwqOGVjGObIXnE9L2roRuuNIFJdzcNDHc/j/IKozL+
8M4Et6kN0P8FEYU8pooZeShAyO/QaMCftbnml9RUkntn1AZcfyqxRaRnoYOgA8tFMz+rBMlFmb9u
h26+ZArmzMoBpje9/xMJ298vntcwXVb6ZDTP8u05wkwZHH5Q+PriSivJtDuQC1Yqlqgq7/W86jEE
dJPHbeRMnCM1D2Y2WmAp+QTuL2JhKHwWsBZ6R5DZtr5CqCyVvkD0Va/9+ZwvFLLPLUN8r+Niw89p
4fPyDNBBoh6XD+CyR5KxX7trdFG9CUcr82m7NMJ7faAaPOwGq4sYVR0p/7HOqRk0RH4IrKHVU9zT
gB8h2QaPdhmjpd4IwnxbYUPQorg/HAApALekag8zVCVSgg1jeJwR7KUUZpO0XylKQavyMCW5OaWm
5sh/FXTFwSdVlr/kJacuvn4Gx0E/A8G1stwJVgSPDXCsh7IUhY2hdUpRm/mTde7HcDGTd/W0k4w6
Cza+QR1fHUt1iBV5WNGFsyT5ddXJ8E8mK9rm80VUhgKRADT9XaA/j/GWEgsMrmEPCv9fB4ShWV/n
4c3+y0URkQnDvq5wtMt/sI5BEYr7v63j8F+P2wwmWvUkEke540YqsWtvBimA5WGWVToDYRcUmuNS
NsCWS/RF53Ucrl9ncRjMm/QzRyNiLYAuYqF6swIDqW2dmjgMKMaWH671lRPFZ84iH+vj4pnLIRIP
/l60+9CLOgHEKLWOrT3g3ri/blgT/eNQADXwjVpAqds6a6UGF+b2O6X3SOmPkzJ2qKQ1a97nsI8i
ipOrqvHJLYdSHSbWZxRY98FJwPkWUAyCoC0/Pozxb4y1JnyM+npwcFyzg0DdbohRW30pLfzXVsHV
cQbuVITHI5lFRbHarSkQi6qzDhiD4vdR4+531xHyGoq1Diny83R8OBL8SSJoxPZHEAyPqVUwYmZW
qv9tXylF+zuez4/wgY2De4+vBetvxrmc4Ym2lDjSMqhGQ9C3/8Gm/6RIKhs9R8otl1vE0QFLJVrq
3GfSjXZSwHCHwcb6nRExdUDxWHn2jSKIa6q9dV8ZFWSBLA9j7m3Ifz2I2dGzDqq9642/MFTGIpiR
phtcFfQGK8s0rmpM5PKfgXgwgqmgnYSCdHU2IQa9x6wxwX/FpobAqpc9AKCG4NXeR240aFvvu+0/
qziWxGUeE9itkR3aEAX1dbDftN/q7AoIBBiFW5aiTRygU+NutslmXmzzsrA6athk9fArYxs+03x4
pVWOX8ETB7w9YtgfGi2hLk+N+xNNnVRSmWdNu7KOE+TY7BE7HXndHBiNzrmoXwoWCdvVDUybUQq4
WcQ8IsASrkW82ZyBoMpL8hbcr6OKUAW2ANn1dcdI3hSlIBAeq/eOHp911v+POlhm99C8NFYDTmLC
u78M8xwlSyjcZV0+59+cuWj2NQezymx/hdbtGyLtQkd94la78InDTS/dN80/tvR351tSC9OvP2OD
GuU2m+269qJZMri05FH3iHfX9FZxLJgwfHJ2l3Zbk0SKN5KcX4izmdjCalsaYO+0gXcTVZRK8P1G
1iesb0UNvd1sk0a91x0+qNB8K3NKE9QCBJawJjwGsXrYqi4PkojGvIa2GGeMjH5/l+MN5FcxsTUS
ZlkK4UnUi5ESfZnyPLejyZNUO6wEvCuqJBiJo3bzNOEdVRA/MDoXMjlH/JQCA9NxwfZVZeIhy0ie
SUOlHO3G02wP5mMaUd2YthGho7MY8T61a7NYLammC9ViFDnuGCm7XbukKOlwMFnUFFf9x2LJ+TLo
Ub1QdlDRp1tHntr7q+TexdZ0jy/9QPqbaB+fYpk75bQyld7U9DDSe86iYCOujUF3UP6y3WaqpH/H
3YUD2G5p4+nULa0su4TphqfqRxsfzewcj8NV6+4nHTd245nUaJNI/a0ZpkC/v3gSCWfiqLOjj0CP
0SSRgGjArCZl8C2ZU73GIpOij05QCZlh8pqirHkz6kDwX+erpqYtFH9gl3y65puL+xvH7MSmBPBX
MUEmB2qpuzRDUwTu0RPjJSyZnai+g7VqSlLSEIr/SDYtRqVQl5Lk9eouOlwAE0qHrHh+mo0YUtSn
COdtsXB6d84j0ikItrlyGbmn1RZTmHNWdan/Cyh+npmbHV4CI6kB2bNf2yDebr1bpT/FlXvBK9Kt
busI9qfHBMUOy0ypmp1QnWM2anB7S4tl0mjR7xyCEA6Z+w6ljnLAUnZUHhQE3NjfyKp0J2tZXYS0
t+ntsJ1AQOMNzhRDexBemkxjhvdaVjn1fkMIfJPii1EdK6Ung8gMA/Ix0XN35nKsO4O8yFvT4S4r
gbIg0Oq1PyTymh3XIs+YIwDcVuD3iIQSTNk135JYw4+rgBDT3uOjrBKhh/kRFzAS5THCZPc4bGil
KOsXXi2kT9WnOHcPS01zgLZFpPDpKPKzldzKmJ+4CfLCV4hX6ySyvWqtc/62EMK6/qHo4qH42uax
QXDcNmHkhQXbHxAPHR+StP6RcKY2ii8TEqQNGOc3Nw9vD/dsvIjsr9leLn7DDyHbGB5kuvD//qDu
iWNs5BczRRAI2mv+9yqeFXHmqqThOcaR3lxfpO35GbMIoLfQH5JQob8F7zQkiKD2U8A15FNAKvUn
NjF0Q2Hz+KsK0syMITNIBjDDT+xYymK+8dinIJQAwHa8VUBcTa3ejH2TfNTv1qMI8eMUUdronQCm
QjgOQ34bYEN9a+MC47lvku2R7hkpDhUnf9euiYucJrR9iBNXX17uxAmwfjZi056y5fn3sVF+veDY
gvQL12bJIBIf68irKNjX9+0gz7T/pcej4JpUmc0fKfaIRoU1RmLqZBZpprwj5xPT7pOSH4Hsnpjv
VwpSKf7xskEK/2M9GAuAwrahBdXQtldDOxrqy3kdeTZct7tYs0acLqo6V107pWlUhjn4dSn0K8LD
ni+wuNDpSHS3gFzqwFrdEzANuejEUhr4hwthIe62oraFQ/KtIOXmnm9XYX1zaQj02T+IZA5BZTGp
xcRgn2xsByjaDhDMmn18BOeV6zM3aJzmODqfe3dlA74YQW1YXGmtF0lTeSUCtBrTCb0YpcX/QT+3
HERO1h1euusu7YGkcB6W+KbucKGWDNG850YONVSZPSel93NW8yZaTVs2ZQMsRwOutqy93llS/EtU
WYIbA9b5ZUiLEoUY1O81zsRuBrFtqviAwUKgsmgWBTUdFo99wXld2IBl40/yfZxp/fg3zaIj24lN
sOKBRrWcIiO83jrtk1vVT8zy4nfstfVPgr9JFWawyLCfLNx/GR3SjwdkGCbK3HFk4DS0oUzOyDv1
HNg9qqvyYrSXL4S79cFw96uOQvc3yLh3QQIUwXJN7GBCg+8M8AMs3f1jqLr/X3dm3e7hKVwuGryN
dAOxOzdaL/pbRxJ7j4c/gQ223T3pQRZ52E4XhEzZtqhlX3RCq29ZpEetphx/VP2sI1QnfZ9ituVE
Cer+K+MM3wtf5frLP/va0f/4wfxbgLbuTSs3m+CJmCmNjNd+ms8bOE7MYy2092k8EP/chUDlWcAg
pNgJpl3JDDE0N6Ks8DOOvJCUDkYHLo411b45ZpXozObz18jyans3Fz862LzzkV4BQR/vZDvHLXGt
QPX+g/rbcInqkn3xJv8VjQVsfck2Gx1A7ntXqc0PdzUzLPKT0VhvMkjztM+Jq4tcHmEM75TlnA7u
sta0mqs68w5l/2nV1frSel7dfk6nWzFYFn8VnpwTZO8z5Zx+srQrUvcX4Y/jbM927q2UwgCKwwfm
O3rar7lobvub+lC/cJIZK9/kGzwrukipOnsw5mLVjM/oKR3/2phPzRrX9Bof4YRUnFZEunacYyXj
1ehdin+8uqPc08Ykz2i/QSmqk5jIrLoiV1oowZ2k9leHs7tyxx8kzmIhCctNBL5WroL2JXQHjqD6
0+VyqhAWWv4mZrGl27bO6/BAUop8mAHR4tWYwi90CtgPfQxSq96C2A4I56eHuhl1c276aXL6w5Ci
auw+UHHqrIttTfegFpRaMuUXC5AbETvg5uEq9fAzxRV+SHB3d2wuydVR2DNqRA/JycFgzRoFc7Nd
P8vRNAKcs9JyKIQOIwUdq/QMTuisbY8uAD9KGPaEDT8LDA6ga0dfIoNqtjA9jnyHDMak/NrwLnZr
8sNXN9kCrZ6SYooQCcZuLrlAOq4r/iy0ESLPEtylCZ1usTQ6cL9Kyi+WhY7l3ShBcxaoih6voQyT
hqbt1d9zjpaFpm0gSlP0WrmqiWOLUFG68WrfA74FkTJ9Id+/QrIKk9oHvwD4H+PfnL6bHjwjXwoM
L6erQ5MXzNSxrTS8rsNdHqkcpjNTaZxMW9Ws0HBb8hPrOyX8mZmbgwfslb0dOXLR0rzH9UlAbIGR
2NoLlfBAxqMEuXVi7EfVOGJYEeoHsntWMBsLriHLCu8518xOyZIOuYQiXYTpquxMgHKP6X2J+pKR
OTVTtvVGrNNwHKgtv86fS68L4ZoBX2XSIHbMQH6gqxFwUwMA4IXEjPHMpBKJuzrlzAgXEm/yBN+z
9pFc5cRrys1xEV/AKDR6qpuBlx1yGYu6kHG3bx+X7Od895TyNz0d/D5pcWrt6zoIlGo+CTyX0jv8
8bbRaHHa7xc4U72YQmLAE36887HTdDW3eZVXe90bEz+Sv7iquIZexijhRx8uqDGCzVVlvLVXpI6d
StSsZOZjT5AhQhmhvXrbh76cfEzS6ye63sTboZIt8xjvS/ZUUYrhgnYO8LqcXHySwd7JPIBguvsi
narfNtC/vCxppFS/NLTd1ter6rC1qHCSBwk3qQUrfBA3fqsSLaFM0J8AA4CmU1tNhD9Q544jzgrG
18Lk2+h/UealWcpMQ6NFbRnf1In58NWROgkGIi3Vola+fs7jlbEpatB1jOZeJAVimzK51GwsZxx+
ZG8oFk7wLLgeV68IDoFn8L2NI9t7kaumFU7pliSn5X0preMUR5kHDOWCM47UHyt1n3wPO02bF8D8
t3I5ZCGyPXnzyOLxkMoCcNgmWWPjCeOe5AOxfqdZp1qEn2JNiJ8QvSCsKmdAY1XlQntxDhnkMp/t
xSXgIoR5JSzPwp1qlDzxQ8x/8Ok24NF0LUQoBeywW7D7xY9QRzp2skEBaHcG0rz3Q7U/PRRNu1CT
ic2qR1imv6GhQ97mUZZbK8Bed4OHRIa28Pm/e5f8QJaktIFfUYpSPyWsBovk9JUxanBmWwl8uam8
ivy0eWOAnB/5ppKJuAFETrIGtCfjBt+FfZzOe5Ny81jNU1ucOIE72wsC8bFY28hfq23CC1AZ2Occ
RceDtJ4jg95705at4y2ohjnnXbtBk4mf+iEUffn4QiRsqGvLRAxmXuMGz12VXloUOMH49ujsnA+E
h3rRHUS6ndT9zEZf0Lux62z5VjZeHesxMC7SvCHW7fFAfJ1RT9ERYb/zFWICyMXOhmdUfUhVOw2b
zkrvTHf6FtA3iEG6598fpvq+9LltskKHdEJEC+jlP5xB9CY1yg6wBrP181kD5ofH5N70ZV4joeYu
B4Ru6Xm5uN/a0+62X/LXs6BxnasC5OSxkX/6KAQJJ9mymn3OlPu9ELHel/cT5HiNAnlSh2wP0v3T
06by/LZlEfmeEOsG11AejLAcRtZNXAehqs829jpyPm7lG1tZMhIG8N6ifcPZhcwxSA2snauCOm6o
2SVDy52tPlZvunOpV1gPyr3BsgQeWHoihCh7ZoiCLR2uRREfW2rbmATXWFMYnWpKovETYAAgtbel
M6sw5OYs523u5a+HEwj4u78QHP5Dx7eqJlVwNxcPCYd1G73L8wnt90e92yQWzjPYgl8Pj0yGFlwZ
z/MmNZpGToON0LdyRy10cj/CNbGuUNtHUMqxBByEfxlxn3x2IPUZSvRs0+z3FKrK8Sbd6Jx30uoJ
hZq0C0PbAStJSbCnHCY4Ic2Qdu3yHRUqsuIEw5FB7OKh0oUNC1qBPstOrN9fCn0jcFqR8CU4UdFG
lp3v4oxnS3VoT8yj9LtgAxIL+g+ebAOWL9+WSKWz2xmXaELxFeAscxSV5iX2u8VbdYQSyY+PoKAE
WXo9NE13C+RuexiDc6PFEVgn+AyUn3LPtmI/iSJFpjMubE+B6s0/qP42uq4lM5olJS3nL/Sjx6yC
4Hk5rQi4f4Vn2n5l54BC/uI1z9nyKEU5NHU+Sqripwz6YV/hcjzfOw1lEXvZqkLGHV46WalVXoNP
3pl+M7jeQLStM5ll+D6CNt+WZDxHlRms4z7QkJWaMOjpJnTQpALjNUzGDJtnaYJ+4wTLf88Pv2hO
iABvpDYnqtsO9pjgDPe0xjAU5Keo2rnzOaCkv2LeyK0Mep/BVIJ6/Ke3NpnblWWIyWvK+Cp/owjM
Ax28qrgdmviF+1X9yi+vTXXm3h3s60mSTbqhEzlnD2J0CJEm4V/1gIYxbD0ocbGsXgmLeX5sja+I
BqWoCq60Ehah0Y1TaQIts/WkTMhOwd6ioG69Hg5IPXbM6cS3JbkIZ2VRrd51DwEd4i9Y3k5B+vPH
vtgg9iL535B1fVMo0dfp6L7I0c5xKZqbPpMi5L8syI2GLJndVWz5tJLncd1TgdjSDBHnDF9CcyAy
trpJRE5AMTiRulWHT/i2hFON7rcL/p5Ta3uDOQvSCOJidVYS2fgUkg0Q/0se3abfEyXAFML53TuO
vlU0JI6IWpa7yvG/lPg8I3tfIcN7OeWzNp2aez4KbjDkmMNvPE+vTADfAhkRzeYihKVT+a3hnZjP
7n+iv1KtFXMcq/2bAhMaDCGKlca6A18TBinlpcW47IBeXBuz+ccM7jrSvZCRZ30UAOUrKYwyUBcz
G8ISVsrRwvDK4DeKBuaesfGc03T3+HHjFxj6VSm7WnXq/wbLRLcreS+p58qhpdoNBBASKjwRvEjw
Oglsi7c2Gu/okr4QrOOkSlTw8knTVOXN5CGnOiub8iXz0/Ui9aSjyMKIUPalbqDL0s/aNmMgv834
wATni68om87McccbafhZhKgJAQao1iXqyEE+qZJfDD+0oqlNmH4tZiW0QHWtisZNBdGEOiXIncEy
lZ9LTYA0m9RBOp0cPQZrQhJHJO84gqXfmEOE7ABRYHjERq4PVXn4blL6LP++p1S7xlxloz2MU5gz
Pxewg6QNN+ZS8cE2L6sXAVu6/dNHmx4ivF7DL8zxqTg5a+WWjxukkJ9BcYfP3P4VEwkjTZgzkK6g
aTNSKq6Gq3wqMhPgRqq5IAy0rW0WQfP42iZCyuYLtBEwAdLA1HTj8/VRVZ6/j7EIvCVOXsg6UmOQ
sjigZDHL60kjqsMJcAloe4nGFt55mWBqdcGQc6MKTM/8Am8HsVIfRrmR4W8FWBZDmQH2t5AUYVAb
jQkiWx6uhhMDV2J0DxOVPvY3c9URAlw9E0Ad4Ov85cz0VFFJgJrB/0OiQaXp6yA9kCRiqOYofJgY
CnDZDEF2Usw7RCB3ciA0ugnl4r0V6Sd08P0lrfUKc+IQwJSW9EHLIEMFpceE2ZhO+7+ZkPBO5N3t
OW9viIcVQE9XFm3DlAeA1a2dfz21paRSvEksRxb0eNJz5fino2tHdJHlLXwc78mzzH/a4S5DkTZ3
LVZiYzdADrC+oLCKGLMLtvIMRxPEwC5jz83vUniVmOj72gw3JhGmlf98tW1Nlg+n5BYHPMfsZxju
zFI/0OpqtiMzE7O9jcZMdXL+u8p6a80/EjHyKtbnbvaoc/3pJgzCFpbz/upuyYCuopTKbe+iBfq4
lrugaTwgsD14rvoJRo6O5MeC4maXaOjIpps6j39KgW5Wz9viLb1dyuJYS3eXUgs9QtHCCxbdjPxP
t2kxQ3ttfthkzhQvQF0yYcWUL+dEzzKWQTCqHgQUMtAy8BFHO1ZrmTFBUYodrFafRJqUZFqjPAjS
HMS7esxpBo/aoGn0UMbci9wmotkdSQlYt8Ht6c6qNWddOlIa6TQiabGE3fVBsANImcTw8xR3KeaP
qLRBwwctk7KQsVjvlc70DfvDo22vCB54/oxW9CrFZ5Ly0l8/M4ekJI4JTO+DYrFeFtvTyeAoj4qC
MeFPmf2K3lMgLSDaz0SAQixnHrTBLgPlUGNpMizy4DSWbqBQOOPB42CkejpfqTWalBKxars3qBwW
de4TKCbt/PzgKDDiV4dzozbbf4rG1xqdMXh2S+afMkwqammSI6Ryvk9niDkvG6nkHaBnIV1OYj6h
iUtX7e0ggL+ir9Ma7obELvEus2qMlx8HJ/cZVmt4gCTUr/pQI5w6buUhFj313CIOjLM+jC1BFnaC
s/+1Wdj/m+eZMMh2LEAOaltRyAH05WNUj8p5yvFBFUQqwtLuuwOCLcy/SqplRaav0xX9H69Usy0Y
Zsuj+6RiIZT4wSIgVc/hGLkfkKJdCPY2kKB6d/Hn5EGbebFQ3VdASusdoJQaTe3ki9sncflcxddY
1qmOGmW/ylO9To4ou6fkXYO8MJNBMHzLZWOSlhsi3S0QKCK1P44m5wF5Am41GKXD0c0BHDTk243w
ORv8AaMHbhjk0AkVJn1dfEPFAN+YeT+Cywt0O+4RoZ5xAHseSspqbvS21EyTFmjB9I21dB2dDKMz
n6QqCPiUkVUEFQ53DBCZ92txMcadHWuib0cFiv+X4rSBaD1pS+2j6do9Hv5gWbLdIUG9dlTKG39v
MrQGH8lD+9X3eW89Z3XVI9sUSnj+Bmq7zCDebo4/1Jl6Ftg2yvhLXef9wEoS2dIyEcvCXIT5enK6
E7L3b5Htkmi8xsuJLm2w8RLYkYNjeY2u6ouBBH3wec5d5wGvPOvjg3IYXf9JmQQQyx0cYuDLG4VF
HFwwc1+xZl6s+q7T/49X2NJ2dbiVZDaSfaqwtiiPkO2MQAtkUrxOkXqChrdgZeDmjDYI9AaLdxgJ
WI7S0dHifYvVcOeRg/wXvEeMUbEN+36j4hMYUNB+SZ6JTxywAmFmSt+x8h5lDm5m0LWPxZQSVkIO
2SAq99yS3aaSsaa5vXHrwMk0PKq1ZA+1kqCRuDaSyabu6qMK5M/FNKbt80a6aZZFtXDqNUJFvIJf
TuzTFsEhgrSi7sIUud3PFEBRSrlS+0epQ2rLX7rHu0Ubo2T3V4TcO+BJjt1G7hA7yd3wSYTGlpa4
D0CvpPQ9r6JyJ5dHdXCUF+j2HWUJX/SF7pgNKdMjeohSxndzNscKNtfdWkaJD5acH7x5tW4JHH5P
suA9wnkgi5NiCd906Q2t4GNgygQbH1mUh7T0WaiqcQZsVudiGVaOjX26VhtcsmGH5by+2AkBZB8T
0LXSy/WLNN11ng2y91PS9pO5qlI3A4q2Z6cf7Z5JdYng8AG5JSj5Ket2G9tnJ9R5tCgjKZ8z5ehu
Cep5dXHkCOo/fcqFT8Uva5nx+9dCAj5ZKwsY6DChsE79zgmhGPX2+rXVMUptnr51ueIDJnTmph43
GJr8QlHxxt7K2TDu6ntn8PsFaz4wJUXG6ODJ2tb03spgKY/BXcHpdYv5ql8YWLBmE+4lKsDLpWF7
qep7dGOcpDtWzsjRsY/bbf4nMdd8AxGRfSPHdz9BSyC1tEc7vxwi4fZmjMeb0Q+ag6KgidCZdSob
fNpHJBqtvt7Qyp89KRy1zku7wipwEb3QvHGwv1BktgXMnkewmdQNP1bcBaogRm201ipQro/PlsBo
Ac5NYbqCCp5Jr+SnWaOEOAqnBKS85WmT6cIqEKcth7HOuzLZ683jucRTIPljkAVrZ3YSRmEihN1U
N3gS5aaiQGV0iAQhEPARAQe586QRGifcC+tXuFfoGVLaK2tzueBy0kDAaWERO6odAxxAU06MHlRo
TBgv4NyXnVxlR4nsy0GPOL6CBCfPZ4f28XMgztcB0td8ruH1PhfX3iNt3kVnmdccPgACdfvHZCS5
FcUXYScnTUCktcK6GHrrBaq4KfJbQwIvK4DE3G0Rf5toPrytQENMUsVx6/ef3xuU2s1EgR2sFoQJ
tJV8Cp8mswVKghdOQY/pFBLliX3dXXxIakpMvpmAuX/9ONIF/oocpLcMy5ALve5FLqwZAXiYq7je
RD4XafidXGurztzoinwojaGNs8WyJDnRVv21T/AncHBCwAtsmYjXr1kllNmJul8ipMy5s6WsRbjY
o55NBp5sX9tEhn85DcRz0Ee40vJEJE4e0gCoa02yB2f6WMsANUf+bbwerNJiiQ8rpIdTwJQUHk/t
TD91ajzbwblbDufWHshCUCh0LL3IKtVqq15TMD26+J2+uoeYfltcB3puBip42O18jp28XeGMuH8F
mObArsSG0XlwDp9NQGGvfJSE/B4fqSaF5xxWIs1I2UUcztM+VYiUn7aTpkWxSGw0RopamYjoHWw0
6yAS2+TtS1Nlk0daBVnqPFZzrGCZx/0jwF7GF20SRMjn3VImUBMXFbhfyoqufE3yLD+lXCVf34Y8
1hKnQcLAPLcN5/rQSHyrgox+IKqf/LBCrgPW7Zbo3qG8Oh9p/p/5MEKdxpJBT3Ao3RS6iZrcp9wL
TdGVsHvMBcsC7ec7p35lUMdmxSDRNv9GmP7HdQVXYr1ek4QhedblVWSXFzx6mVZKULbOFwdulg52
sF60wNahA13MVkcNWZC29xujDoAa/f8U0nCuODqTSlY2qAPl8f9ZVUcpUk8F761gbkeOBiBOIcRs
MTelk1ZlN8s1jLzaNmsXZt+Qm/LQEQJrju4XmR556FOE59eddV+XeqAgL3r8XEGoErHeu7ioyjw9
Xp/yaEgMZjeW40nODopLYNTLJt3ov8ckLdgHp7PvgYXYtmbn3umUrhnvcFB3BIc2Q1aD9p/kZ9LZ
qtcEEauCW0/anZN4fEkDCj6Fo445ugksg4AH7LRMHH7e0gnJZzP7fzmh2KQPo4qv2bri6R87SooW
pQalwE8zhZ7NThGNK7z6Dt2I1AXuE+oHfCfHWyT7jwyBPzUwKEX4jnvv+a8iYH3S6UnZJOIBR1+v
jVnx+vyscMzVbABhY8xrxDRhnXGObwQo9xihjGZBVXUMdieTrjIp876ty5MSk+KLoJ8EOEKvhB95
mn2nqXsqI4q25XGF7k0qhi6s9NoO0n3siG78OGnLbP3yYn+RurdCxILr96F8fAbGNROfVgXy4YJ4
4GoqAlXdfiG0m2MhdqqICFgJOLTtYENgIyXrmnjNhSxVVGWIFUSYi5Vt4toH+S8znFWk/V/veKWi
sLUQJLioHF+YB41YUr0odRHU44jqhvO8qcZWYoMXjBZGWzNU8BF2BbRvuzQvx1cwbJdZfQPitIFz
LL/0LkOzI7xhMhQ+6OkHeJnZTUSPQTvmpBEyU8VHV3LPCqAZklUfNt8KdhP8z1XnrlNAqAUaWnSC
+/2AZ7Bm8b8oD9PSxO6lAbYfaemhp7jQir0KXDTbwQK2ozHgq8vF4xSjQUNSjuOxXSCNQzDRa0xa
bEsazsoLZ0roxCqSh2Uktjrx0VPqAccR1bdeIHctPBtPKrYIkWM/Jwil/1oez4LETwZEcDSCeNZn
CD/LgUaIgrYa5o1CWyWX3MNQkW0cOe7DFBt1HSMLshojI3z9rAYsWby91XNKpKmxFE/N3NMJDKUC
GqPu/FCUyAENvw7mirrKybc1HYqcGt6Q5J5czR677xSr0hB6kgmn6ousHSiwmTPZ8AcD7UcL/E3U
Aisc8JbdOuDAg/4559d9fulcrD2mDRVwzEx16YAIv4l/sm7N5tOo41MRY3ftJPmeGYY1Nv41IJH2
7YIMqfCN86FZhqybjslUOqfSSuoLATbGau4/8E1Z6k7k+J628E8q1UjIMNgIXYM/DpUBeB5ImOlw
/Q3JDHuMj9Rj3rIA+DEOHzBVKdCovWrRjYn1pjBmm56vJJdAjfFRzjw7gSj/wtzDc8qczgfgF0AP
BMCrI0oo166sOOb02dnCdngjjK3QEpew4MtImcXkLC5oxew6GiuyzQ5mHowvhJWLNC2cYO68KW4n
PKt8/AhTQ4FfTt7cP+ZmByXbKLkxB0xFdnBcVzz0CQLdcnC1DbQGn6yJ2Ve533RM6v0gXSO5kuVE
8oQkYxCoCUeRyQtUL2rpTBMWI6Qw5+VwwO5vnR34VKhPAsRR7V+DBA4dOJDnxADfTwZz4YUwtbO4
ziWwqGY18BlTR1iku61kf3eXhIrNQTH/nRyanutgJ3DJAa3Tyhr8VAaMo9CbBw+mvIJGbov7MrVH
4a7z2rHc9fNjxyVyHvQ06JODUQ6sEj/clGTR6rFCbO39D6cvtRBUECUecZzcmfFS27tLGI2J4bu2
MSeWR+Od0a5AXSzRTXkY4apMFaa5nMP1dPBmxS5T+uzIDKZ1dGip1w2fYnbIGPzGMKRa9lS0lutO
PFKbLvK99n7i+BFsnfQ7r1W5QBvMGW2GBdWiHb6iMjpfGz+7WYjLWMKChdM+rQEO20WkJU6vHc4i
6E5gtxmrNvn2hEzSiWAR+r6KGGiL18CDlTwyEFFnAQpQ3Cz96l9Ot6CtRD8DtFbc7R9Oj/Agfpkv
+iK6lLBKnIPhiJPFLbVKS92ejhTGsurhQ8RvbJzEZSGfXFtgo34M6iWkxkygiVFrfgbtczMLW1SB
MhGwR7rDuF6PLJNZc55i0AjShW90/g2fXGI8u/XmMxdS+MX36T7qLK+uBmUJrx8m4x9neS3vBfNa
PnWTl6wMVe9CvVXNGWeqjUcnYRzPMk5fuVHre44Zn0iritzhRrGepMF3C7yxPEFG96iVkLvC+XPg
QqGMw7yfXhVv5Ef9FJqHbxM5k9XZPuUMNGcAfOj5IigF3w76hCZZR/FqIDG2OKwLKpakfGye/1bb
RahY6T/cwHdv19AqB733b/7ioroiG/I4DID5fYilGiLXio8hbIQJ7mqqIoFk3NKCEu8Gyowfm8i/
DVy2cOtRnydGcZR2nwepFNbkvC9GG5yV6NwN0fXuqJTUX5DyZUC1uyVrJ6T+sSSxMCpUdEQEzdf1
Sxsp7wFqT4TUpL2kqj7o+kU33M3yTOt6ncv+uEwyXVNG7dZVE7WaMbli2Scq1a5HO6m7uGJZAftb
isREDgAxHNJq9LGdnteRYNZmBVAkR3lpgOvpIzqZ+4E97ynrR5waBE1dSpDIKjErb6GaxsinSOb/
YQ3vP1wQqNUrS+BZV8nTWwBqARvyvldgxt6YK3BVEhi88B1OByqZPAEfM0PfIJVmQq3jy06Q7Zk3
Y7nRSs8kOsqyEGCYturBYWWztpSxi4JDMtx6mwv4jUcCSJz9QrSIiFXqqyxMlazgvMnr6rgpr4S1
qHE7JwmpsNhh+uJ1finuhtTcbHF5kQt1nkttdJvMAxmPKGvHbgjbXcgCDQO4AI7ImLF4w2acpMul
GpDoBMz9hZpmXhpYDp+ToG8zFlHDyfoFqGNoxH8Gi9V8xvA+KzaBsRCST3bGdXHZJJizpIMFJQVt
8G4is7GEZ6B7NpLugftbM7ixRmFhv18yo7dEmusp5Yiz6Te2qQ4KXjlwfbJ4WQPusQxqWHsz4UO/
C1anP5LJLxpdE5YwZtDsMTbGT6ZbYMZmbLNsKjY8yF1ar2lGw+0AhnOXLV9AN/XEhWfJSCAyZXz7
TTdUPkGNoVU8fhj9wUZjzR0COmpDSLCNar9XwalOMUIjJTDsq5P3Yx8ZeKnWoqfA7SGung9k+Qj1
K2PnwM+T1bEZmJF1Q1w22ORR66p9HdqwdS6XWyoe9800WTA0H9tzULhhxj7oTPE8yFl6O/0d+9PD
UC74iHCNuIkbbnclETlidRYq0l6/dpXzyzc1tPdFBPModNrFV6jP5cA1pIfCWbhG3e2l3S97qsC7
qd/ERj0gC7uBMjdD7U0WZCrWLhTy0EgGt7GDNrUsLHvup2h32G/o86oSd1G2yXEq3Kn7odQZm0SP
TbtZ3AiAEvreEH0XF5hUqWNq6QohsPxPAKCtIzlN7MINpEbuiwZeWdrHYl7VCQftCxiNEXZgikva
h2zO4lw4IrWuV8RlIL0gYdR/Vz/Z/NkLMY3CAsxG8hhCOM5FArYygGx0pNDqLC3pCXOGY889NCCR
8Y96nr6CJ7tB4IeXkmVlZp34+VRVdUDgQAmcoOo6htwpJc4Z0ADowOd3RFg02c59znXAnEgoHOkJ
CB7gaJzWwTnTaFf0vQZLHTv1DuxVK9MtAnO/X3YMJThljcU5gEZyK6XWwe1xJp2kkBSRaR3JxvW6
/cF4lCckW1b9J0Ix/wwCRNF8sMKraeI3v0lIkcOW4tJc5Y4YrsKsNxjpV+esCT58cqUsSiHAYH0U
c5auHlYIq8uUaiiZcRzQ0a4UhI4NKYIvTIJKQy1LGJucspRi2Me8nfKsAzRQiLB/a5d1aX9etsSv
8I+ct2ztUSe/3Oo/CMbqL/auT5Y3tBZFD67yqoialQsTnkJgbajYC8DRawafPnEEBbSkCEo6y7D+
QGSpiF4Ohbt8bU78qbhdSz14y8HHx/hfCkWy+/VXvnKpwko2fP2mDGgg3xBL/b6J+BD8c/3MleAV
5Aj7s239E6NdPTRmTy5UVNYTcdBtbFLLkboU2O0SBMmmp1IPrqXo47K0FM4VHb+Ax6rLqC/tOp/+
aRq2kCX5sMxa4JI/VOjfJfR4ArSCYIYehoF2CLapfH6Jd0gA1K0KuUXA3iL4Lgt4dNQEs8pG7XFK
4tj1IPPMfle5vbIkFCh87oZSKpNxrymTn5DBVhHk3Ek7HCqVeaqYobTq9fEr7c2jg3XgpEwid4gK
RMvXx0qOsIQTbD6f9he6pgRK9zVJD40dyIPZz2Iu+H+fejFRgG02icoNQcWtIV+yzkXjPhBRxQwl
C1+rnA64373whDsp3S9ntqNigFGYdD8rAgeYb6Ie6rrDmza2ZBIaPIRNGQcR3CUmPncqmKVxWbOy
erIZvqJHCR9+DUyomsbnC0SclZkLtzfOKPveudDxZJhKg+YRAafFAaKiGx5eTGiUj2pGmTbsZ8cP
iibo9zPVt6zroHYzNLthkzh0ekVMBuSQcisrKh8A1hiIG3pf0I206uokZyHScJt5lAENyRXFoGiC
N8Tq+4Nd9RuIehqwjtY/NF26140/7yv74H1U88KQpQG1RiaDPM/8WmLosJKUbK+VsnyOTK4oOmPZ
62C1IVa5g+YBHfB4uZSjl2/u5sS77dCPPjy14ENQ03Oz/QATP/RI14Cctckk0sVap702jEW+EQTi
f9hbRv9V+kHrmKyTzSH5fRE8hC+J90aVoveZ4etoRcDsRgQE0kX8ex7pmU2CFTxQVOn8jDvCLtDn
w4xtsEh3JMK90MNbBXQg/NOTRK4H3088VutBaq5O9qHwUz1J7DdAmpD/fr5/LmBGsiec8Femukte
O8jHxQMjE2AtjiKBRNDLqqvKDxnh5MEVm6YOfqI2jFf+XAzLwznZO6vRA2V0D5ySefzsS3cFSDsN
eCmzGnWVZhXcD4d4+mn/Mv+yuk9zBb4XQffzDexjo1vPhWvSHGADXCTiZIhKlr144aOBwMbvnBbg
a0TUA2vsSLG+9BWeMQ1tVXlmNmjH7u50krh4LFZdI8ItS+0PeFXZXJUBLcZWZImHmc6Kqg/SOU99
h0wrcDVqjIN8X0JFDFsUT6Mzbz29Dkf6Jshz8dI82ZmJTlJ/5mhCAHW/aicER6hYY1++ikhUhGlK
DtF177LrNkeukNVILvIOhoHziW60yvkXeFcUMtBzEFUFSbcjnBA/hq5ZPxmnSWSAm3cdrBoJF+l9
rkGk7Zz94N5xU1wJIdbttxxzhsgxt7iTyADjO8jqcZ5wYn+ZkKmMn1YtDgfEAR9TQAfoIIpf2pae
wlovqRBkpTiz85DGsDCg9zAj8ORjS72x8dtn4MlflmzN9FdJ029IEIdwmEtyuOIbQ9xQ6CvR+u5p
yx80277sb9djsTbp284OwuQ50PGAYKl12lDCeTUXCuR4hFgrA8ZBAkSHYWs8pMxbWQDn+VTS+bA1
x9Crp7QxCHZMC0X2XoqEnj/8HkzmK7NzWZUK8eVnsHHubtQ7QQ/lqyHUZgvNInf+TDATHUwW+Waz
B/eKjOrBKquRu6tNcTCPdaFtLJc51icUl8MoNFsL+b+nBRt7hmv5V5JkM2VVwYPIzr0oEvcJZwKH
UOkYgkQ1lNlTMXrqIGGEgVoATX24mlBu8+/UOnWXJep8WZ7AJ6O1kSIkwJHqz7Q6jkwEAC5FeRcu
/wpH2rXH5OZU2/VKXwnHNBrGQG/svwAmxpiOl8TlzYvZI5BWplNxpPWp1d5DTktkTvbZcr2XY137
HDMrp0LI6VARRwdeXbzhDOqZuIDUr5RIqxaTalxnQWjUQKxyVCv5Sb9bx7PPztc4XW/Jz96oDGvz
2zRfN7QjSBF/z7B5Z2Az7hEtNuCX3HTzxmi6x1dxd/J6KR6WZcXwlHwWVhjkaRJ2K5KsVwtHXcX0
+c6ChJkIoZQJKUm8IIq4U+4SgFGK827JtreKIejA9cTNWfQQutXmlX+S0Pc/TxRbENMlajXaC+6y
4/ecb6TTqVdCXPi1IycKH1I+mTaWGzyajxNPOcPJHw60PON+HTv2os/Q6YpvA6m4dUGE1flPwrTw
jlFv6NephqVRPKvz8mv5fpJggaj1R9DDwdfwuU71lIM2ID3lc3AoxVDwrYa+AiKyUAGXBvkyprmD
EVf51+IV/Cwvq/U0FpsS/hCEYEGMR86BkBvrV0yKPeAo8nEyiikml9h7M8cnNzd8NDOZMOV5KrrC
7j6OzBB59LI8AuK+4b/Ija7sYdBlNQI8J9Uh424h6UZXMDgqHBY8h2VN/rSXvgDEfs5nl/bdTWF2
1LplgIsDce8zsOPKAGm5EeXxkwZBxDlgRYgCkJ57x3QAmiI50IF7GP9rsLZd+5+ey5NGcwTfuT0A
kL50SgpjA11xyW9svpCmsVvTU7OThUjNvBFEFG5K9fUR5FJ3hx4QrwWeEbixK+wFTHAY5NedazN8
xxmI0t1L5XjF2lpAttk0xggoTxLCVUceFfpFQeesBktOMUwz3th5WyGmikLWFQH+SC8BgdcwL55Y
5JnZRiMXn+BrEqXrg0TMPiKK/zyM7jqyuqxizNijPyIwcFFHdMDfepKAMUXlyWGlUPsbF1fx4Oh7
DsFJcn0Jn+LzetXaq85ZiFF/0WmmgMQqcE82Uuoyyx7TsvYMVCe+gv4eN1ZT/ICiDvjAu2BGdx4J
9x2ENH2yDDRp3Jy6zKPMWmhzoa2eaowFdteimGor2q84ZtODk8ujGyy6BfUHwHyQK8OoM0TK0qrd
IBQsp7UOvn/iDgtCRYXL9ZpDjULy5VLSFXeSxoQVEwZN0iP6OAB+rDd0ohrNW4YeJeRhls8FFu/p
7uIoYeieBOIAQ07ftL+Cih4o2gPzKarGpz4/6S+9zeJk/fc2W3xq9jb7HhRHhRqB2dtlpdn8qE2i
8M4FxKN9KwIJwCENcOAVbzQfmoRNIxozoy3zo6uPA1QwJXxOLNDwpetiKlmyKd4bM4Dc+MjP+/RY
2nkow6X5VxpOSmVbSwXzzMDHc5ntPf8XqMmBspDSyCrUhERdWjfArgUM6iK71X7Rv/Zehc7n8b72
1lXaKorB3cSOMwWrlJOKWp1wwyUVHYvhWo9Sgjsiwv/9+Zz42reY4C+qpMoh8yjIDygt6yLIUqx8
z3Y5SqrcRzzgJAnMUkuzwzsbSeJQfZY+d3XYVA6n6L0dg8yqeseIHw2blLW4qigjmzK71Nk4euV1
U0Gj351TuvyqcTXrUAc9dxqAtKKJlcFxLLgo98eBOIZfgRygJpuqyDFUszTgmqi4k/BYhdPlDkY2
WpL6syjR/OTqjqyq4j/WWeMvpLPqnrHc2jPFATWeh6wAj4eDTGqGzBdN+QJDMEi9Sj1Pkxf7YZVf
G+6StJxXRAGwPn2Uz9MnLj6PR8Kh+4eUzBxll25Kyo5AvJnRddeEuMNRduqxwcclOsH7ScHYhTOp
Wund4rWP6yTXRbrt57RU2t+uNWOp3e3dXq+E0JUFsbtCIZzTT7LvKvRXB6mFAvo90lMdlPx7Ugos
QS5EsF6cWwvlgMUs5MHfVnUqLt4RBrjAoOgyHI0icrd/+9iIE4FoLkM/aGMiqWlYPwL9OHX4zJ4G
P46jkcJRzYMDZypkMYrNvcQ9acmjDSTqG9Sh13++mnHvVjoY7Qzor7YoU3lXXdFCDwHyVAwXBNON
WlYlQs9WWgFlogUsQv8B2kZspk93a0lp7Gv/SpC03WyALN/UvAbwTIkDHFXMUGSYY+wiNN9xqJWz
KWplPiTKYiCku4DVuwkewYQM8YCTUPqqQx2eTW86NeJoiVv4ncbLH2yd10JgH8ZEOwiowcnl0nz6
xUopnVa+rbjGM7ss1GcnGCEUfZI4gUWSXiH7Ohx+rr3gv8E5umVL3OOY06pJQGIW1v+m0IMw5ad4
xXk0W34Xr47V7ikLP3v9X9uoqWMo5rBTJ4M622MDykzM+NRd2Ua7ouu3VKFjfYG1DFDi8G+t2RlK
JoJjK4CXAfWEJ5bYlyT8Bj+7EtKRxLJNbVwPz7IjxmCJu4ggZ0Mb07V5p6rcxNayUdoXQu5U2aD/
kOculoWqDIuxkmqf/wMRnBesoYqY2YajhwEyGfzsbqZaqmvmiakjc7m4wJJS3SbsRqxOCPQ3ZIvS
qKp15dOQr7K3B2bcA4wIHaCDRQtDQJUFGwz7zD/UPh9kjJSKanF3dvr1D9mF/l3v685Z1HnAUaBu
fgtSPpmcb0MsFzfFXq1mVTyW7yxkp+71yZKeVflj9cQCt8VAbf/ihibVAS0iqcC+RPW9yUZA0vvq
Vuvo0Lgm8a8lf9AvCYxql5+b2aHZUE01dRihg/L/WY24MiXGtja0XMLo4aCVGJkNOGZjYiKm6tzd
Y+IosVtR+zMxVdJQFWL5fjhWNolcbaq6YM/KwIw9jzeJn1lmq9xUtWsqfQAKk2W0U9qlAtUXKnEh
Rq8FCxAWVNvsDyGEYOjoEp+QamuLZcwn72aeVg5eSxpdo8mATgK1plzKUiLpkbc5kaltFucEAKIQ
8fvpV990wTNtjXuvIkzHFzEz8sS/x97jPwh1UEELilriOfYoMjjLyAtbde2Lx83iGKCs0SD2vafj
OINj3jsd2JwGvX0htwsXJDPV659MIVeYNIBt0M0Kl9EPEudVz2Ta/W+D57oUbs12oookHA3QnMku
YbeIXn3pEEAaf2lsfV+BIqrTbA+mkScNiPJZ8012qEhVo7NEnVrUJtxajuKDhvpl4ynglnp7San3
HvUx5mxTJG5/SDz6LXTeV9de3BpVEtOyoPDtP33u64EJGT3Z/N5XEhSvbIlqu1VjAzfFJ2faa4/7
2dAwGKpedg2v9NEfg4Nn9Z06l5VGr5JcIbM5RhDz8jA8Mq+0Cft2x5lTtWfXwOsCVG6Jt8hGXEph
mFu9lOdpG2RudSELrKHXMw+7KPx2hIo7s8vMHH7ddodJ/n0Cw2IcoDli44BPn5bd2Q2A2rmaqtO0
fQ7XGZLi1iiKL65JdrThqa51TT3SRDfvvZsrbdhDsPPRdigRVcShvzdz+36j//lPfZe0ZKdis6Dv
eTvhgqjiSk9weYlXT1az5g3VizGnpcjw1FoX1aELJ1Ikq3rPHCvFYA7Z0z25D2rbiakJOjeMkfnM
T5PtXd/4E+QM+Mbydcx0h9xLXXbN+7jMg5f9QBUgf6s5waPC8Qnlh0HqFtcg7j74nNrmEMRsxD70
DneLl80ftmW21jh5MezAbI6oJTf9XTE/8LGxMsfI6GBDHck2M5xCfuh8YTTCQ+8QJl82CoguuVJm
N521DG2j6BP9e0YjKKC0/sVvx2wkjDJjswxPN486IimCT+WxHHfoGL4fB2jZattQ0kKV1zwRRs9L
lSNS0aYMWj2NIDBCg6bjnk514SnuHlzW918RiB15IME3MEVGSqUTtRLnl4EbyM4oMPkWjPRH/nf3
nLD2y+0XaBMhFyygJg6XO0Pt9I0JAhvugztkD9SXwldzCda0WONj1OKmcWOf7PaB2e68FXVZE66H
WSnlQ/Kcp0JjybPK3OR9e9WssOLMXG6k6V3733t3XhFOjRH7gmZFILxCU94NyAZKuHIT7quWt+Qo
N0nnn2GOs2x32bCPBA24zmysx+YYSVQlZF0S0xE12msQ6XxftCBQ227fIlOd65jEUrmatEmAveHk
2VwiWOQLMTS3qaNS3H/IQ23g9f/ft5jJG41Mp0wMHVyR7gG64XsRrfhs2dqh6bRkYQvp6jUwIPVZ
p2biBydsLngNq4rkv76aFbNc9r1+NJzVJ/rg0+FMVtpjpSW/AWcD8yKAnUMyNObCBRUl0nSJiK/S
pnZ5FKuD5TTXKNHyRBcX//24eBgP7fcRVI2ReWqFcvsZ7vrBOJ4pecPReXJqDKEinrn/HFMmssls
fuEMdK74bUap7CWkhHUoRjgqjg49LCfKXqmT8JYU4PYqlRplnwleI6rU8LAw6R9RTMTbRAjO68ds
WlKnhKGxTYNNc8SBbxN9FbAklHTaiarZlqL9P8E21DK99xnpFLocpdJcX7zeSFXSIQkx9zm/k1xQ
jeKD1RNurn1MM22tbSB3C01HwkL+5JNVeMvyiYrp8uAbUWSP23505lwa2RccTGFT5gbKuvciY9ku
9VUUGU/ABPR4oJJXXuWATTUotGg8a8hvagPHoN3v+QNfHAdtlZu81yGm7WiDubnl8rnB9plQSGAx
hylb9fhY4iNg2wBrfpI+gv9h02WPmn6NFvh947jEKToWe21NyAPC6m2BCsOVynrZKF2eR4fN4EMl
BD3SQ+EndOE8FbAFe1/bmWnRlnTjt2NQrRJMjmauasGFwhXGUmPMndn0UUgc5LTdFzQ17zb1GDC6
6w+7s3Dje1y3rXrSjlLTkueU59uScohF6RIdva++0XLMFiIxNbPBV6ZeeKBHAejGfDCKeW+odml/
wPI21IP3KNfB+LuT8KzXqI960xJcyMRqdp/qcZGHH3ArQky06e4MrXNhV8oayMTOzQZcXE8dc8La
7rVAE2/kGFYeHrmJ4jNz0SMqPdv/QFZAhAHC6df4+QhLxGXbfmMkEsTO8QbZND4d4UctHKo9vWyz
Rdj2+KnKCXrjTiWQdYNz5TbWtK9u2yRuWzXWWewdqO72Stc8Wh14qNG84vZmBHzPy9d0VkV5CYXu
F85nAqn0H59ucgQAJ3SvsLwMbE/up7fI1kHTcVz/LazpOh75DGN/Ps1Gb96J3ONuYBVIRPiy76jz
kJE6N+CyBmC6zW6nefxEyWcLeOfAXahSkh10m37bRhrPTTifzb5i1m9QK75PbpZ//Dns/FeMslcC
COz/pR36Wf3VWAsgkgUemFzl3wrUTTCZm72S37WTswn57zTA1/BES8PQ8nog4u4EuCEU0aKx5Ndn
iq5CAE0lHyapdQ3Xei9SRv75S7KVm5NeD3PAGfseoBrk3Fw3QGkPAwhiq7BASUy6uIdEXSyfbwUp
ALd9LuD+9TbGIY5Tb3b88IwcwKfc2eGewORGSys2BFYISjlXSC7cTUdejm1HZAqdUoyNC9C71c2R
SN+rC2aZP90+7i6OfDex6g3mVw/FUa4V0cBddm5Oou9rXy8b6YxGIVtzoKhVSOn3t9VAkWOEr2Gm
qBimoPVoUQ7frA2vZvRM8fGse9AIXdNMRKM5vyn/OADmEDfTQ/TT9scEjD8zUVREw+tD3losHMiW
T7Kn/g7/IhqoAL4TpzdnBFgfQxIAt4EqkYEvthZp3uYf81l8svndOAJJhbaCXqHhSIq/hvEbDok/
8uNVrmApgSFRul5aOKugYnpFotO3MXRyfOHbhGWdTQYp0UU1Bb+0rELmB/FcfK/J0MUcve+GF9Qn
3q1ueQw6xuRWNKCvj3TfyqbAHgMImK/B0GU1jelUlvcJNVkxS24EKLk4lPOb0IXJ37Ailw2cGO2j
CJbZKkRl2ZZwLbJzjK1Lr48VmT1YPozc7jmt8AetLb45N4lut058q2A3iLOJsi7dYXym1deISE0u
xav3f+wF/UPqWPlzi9HaRTCwA8snRRnJs4iC2uQNGiPARF6CXiPmuM+fI/6K7uA+sFdNvy+V/bMX
sNOgnAPObjAReJ9C2l+0lroR4UpC4sE6EHn2ee743k0UuP9OX5+xAlurUbAS16du8F552YudZWF2
1ejixJWRutpR0qtBV1flZAE+0JGWJZ6yb03dHELMOEu0k8Fb9IAS/qzHmUSQ75QDNmfaMzGKGfNq
zBENp1WOaDRLk6vxxsWtj+fl+J5VU3Zkk0TulGDBON0TAY/PpSIOmS4eara4DN5UqvHPh/wyHLuf
3bP+hzfGKIBOUh5cBouV5loqrgH19y2rFY4lfzUZNSVVsrG0iOFwFTtiFGRFPRXV4sRUd5IZ0LVA
pLncAfC/PeaZLre/z3K8ISnHX4qkrNd3z/TPCkDWUYiqy2C9QgFxdWhOpG5MTd5VSV5lq0dou19R
CTaBPI3wvMaHBgf9LVGzQeF9kkzzx/8FqC/ofvfclQ1wYal4dIPtuQmL61Azf6UjHlO/qcmMXb7K
bhJabfgSRywZgj6oMdT5Wi2o9C5TpxVsPtZyHiZKUXU/b3D2U8EapKczxLTSQT9Sfrbftf+Gi158
NQ8QVtAPPCzy/xLCQsFUTooAUN4dStXx2J9wPPFXcrnmZONR4QKesLQrH8CA5yD84hP688Zjvkfz
pJevGYmkDqFU2l1KqWppq/JNavmRXYyfm0jC0bEI8sjdtDI11ER074wrXP4jW4w2w/4N2ddCh5jr
MyMmLN0W+MCE4fiNw0jBYfzaHpe1N+Dd/ZpeXgZkHyT7Z3nYPOI56PRjH0/SDGA8ph5NcWzSjLKe
L2+IcnBEVNrJMXFV+YPlIy7UGrxHD0nRR0ZD/NbeuS/UpjOr/JJGChqmfF00J2v9ZIUWu9sFCK5W
VQQN1zkEgKNgOjkS062ceJksr2q+DwP1AgP+GtSlJbD5jXFDb9eiEW6r/PPf1Yj6ssu5pt9s8wjD
OZnXzdDBhqhhQHoCKCd3J86cBB+QR4Sr8VHrwfUGKOPNjHTm/EW6XkdjKobb+H7l6Juv0VhH6jxq
3njAYbCJ3v8oBuFvG8NHFeRZCQ+O5tahO3b7VnZsDS9u92jUci0d/6eFZcVzpkJEGLPYc/pvAvC2
aZKKqxPIcOXYzKVlU3kMIGbCHUsRxzAVeWtOk0Bu7Uurv8XNM9V6+2UjmIM4qO031eE7OZu0eWbI
dlq4TkmMzp1aDsG7FcYaXZKcjmHCa8RoYMtCBq8bvcQ0gA3JTw+oMDuLp6MA5n/DBLwGu6ph22PV
4ZnZkvFProUi9O5PATUfYZVEoPOKDKhHV6LlRmZEtvdTbwVu6U3bOhqmki/SLQrgPH2ePTky1VWa
+KXgCkeuzE5Q42d2BGOJWik11sSy6wSVkn3pJhEnfYlptDxPRt6fXWznf0jelrcotZZ85LFVpfKH
FTCuZbPHlQrRLcCWfZv/E4OEv7yJ/rQpkvrMywL5Y8tmUujlYkeU2DLffcqcSMgz6zBSMlSSJKOk
AOen+JzkxvOqwVIhWbwGCbsnwIj+c2iBktOSBNaxiWbCLvv3lcp1r0JME8Mtw9l71AEkooFguQ7D
0TN4z8nbyct7xpQCB8E1kCzHYK5bI38ptRSS3cfJNcjeI1Ni9Xa+CbHAcQohjMmMQc6xQObNDwSN
bzjnL4NlWjCxoH1flN1J7Q+0kmgv6XDdWr2WhASZT1ddOBGJT/1l68QBk5kDN6kcjw750Snm5kLY
ru9g1XC2I0gO3oJlC3kT/xxbu5OXcU5Gx6TxdWMojmyAIQliV+FdPXFkdJXENSDCJeTjTNjixS9u
UQ3O8a/koya6oA74ZTHXY6S2i29tOZYbHbwnQ+o2yLI8J66P/0Ce/J1YBX5JBZ/kSBo3X8EOD77+
JAkNqDXaYdNzZAayYF/IB7Whw1QPhn+fgyHgCxnVFHDGYzyHZZlnakPhBusR6pv9eepjwoBwzMEJ
avQTnNMTqTEq8+6SJYlIl5XT7l1JTh0W+HWyXOOd/nFm11OUmIhydLKKcOX+jxb59hqXbe8OJGBh
sZiq1BBbEu2D+oaIMk2kwSIG2ftRIxNG6WRaV9/K5mCwUUEmS7Y//7Any8W4u2QxnIeNffUgIJnA
l1NWwtnxPqiT38++deFxW9/RfAA79i4tmIi+2ANMWmk0iLY7q9fSqYSSTM56iCBPjH+3jjKlsTH5
dh59AiXgv8v06cfH9rqdW/6CRzoruXCge4nDwZ0288kUyYRuOLbr/BpEenh2tHQxvwXGY7f7RIVO
w7OaSFV4i+IvsBTDvDUVaMGC7jjqTjS79aL//SEXrzlMgbzbDXWNK9XHWGmbRoHkKAOImEIH9IIf
+a5cMcJIKrR/eJvATlu35hUaQQVcDwbsOgYWbvoT6WO24KEJBcPDKDL/7Rd2dOmJk6pex2HZpsha
mnqwpwH7Sa0KK6rgxi2Kq+4xfUZn8NR/3dXTgUEa6WmVt+4iII1wJf5I77A/+i+KXO6NFTMkCxNu
NchqxwtN3drDprWgG5gn0x2yV1ocKLKE2JITXLdEf35CokZ6xU4Z5/1Ehspp1SVoL2/XZAYujeqy
YYlTpSMoEqP0jjSKvDmh4wtSz2/iKWTPR3/lVNQNeDrCZjsBQxn/BZULAOd2UfLhhMrPhuXzHTaa
DWsaLxAULFtpFAoogNTk9i9+EM/K1AZj+r3SfCkW/NkSbIfX3HFsy46SEmFjI/cDZz9W2XZFNcUe
pxuqpH/NerAEc9+R4F8+z5p99FKYL2M720J5cQJwpkTZEQTbWayvg0Uf8UyZbPhS4Pxf2K3G3iUn
sIV/MEa5AXMhsGAW1vHSBHXgowFWmex7Vd2Fmk6qSABojYLi+b1bddNaWzh5M2STVLOoq2b51geO
aPheXvLk302D/kRNNdwUv9Y/YEca6lt0vKXQ+4aJ5hejOviaTCbToPmgzkufecgmWHf/UFjheZNu
OolLad6GGr/rqlLlMWyk1/iS97IDYTrb3pZmgL+szRPza8Log7XCyyxSUbtDcxwnUDlUbx1G8Bjq
NKRlEsydCEQ/+35LxXLBdvB6CB9yphH4+REMwlXjPCm2LCEaZsZcke+uPJ3ILlaV8NfKegKyyqcX
wLNdA60QM0OTlVU5SAAO/EiL6LcnXLMT78vbHF816vJUgn8k3LAOUs/w4PbYI4zp7Nai6n5IPJBp
vnEhP1Q2kDWnRjtuuL079bi0ymIKZeRT0i86bEETowgHtlYBeveXd5K/Rqq7mpqRdpeQAPUx6QYf
lSl7RliuAMnIWto4EKY7oW/54zc0Lwz6pBj8KbLF7JWUkubBWTS8MqC4djMgGR3p4NPB5FdWgPWg
MsJSUgSmvwySoABeXRM/zHGZRkgd6nV3x/a7Aupj0G+sAVTYQzPMTNuwm6Tn3JoACTkCoNwh5Siw
FZANY3OHJPWYauMRd29rqao+L5TZ9bKeNFEmrRtfO0fsbyDesLaPdBahZfZ2AtjsrIbwtjr6QCAj
ofufw+tD4Qqw+DDhpYt0Vox8uwIWfNSTQlm7iF67yfgn6otuDPthutFD2EVDRgx+KC5GyT0Sbo01
jOcfvQNOJJuqvV5lklf4JZjOUXvnCZ9nusjnZiOnKIrvviNX7k2KMNtZ6Y7o4oSs6bet83AJ7EVr
BKEt23klPZtfIhswkKQ60pF1653jJd6JuY+kWqvlqHoQGugcLtHM2yGF5ckkgE/jfd77N4jE4fKu
gVcU6ahzraOwdaRXrjFEqcWMExYdGys4nTKRs4MpQ4QebzumZofrWuu8On+AVfk5geOadW39tdNG
G4C9umBlp6YIa18Bktzd6m1KeXZuKCbaoyx4NlxRzQ+nTZIOuGl9CG8UHlSI76oFIee3nwRY0cFS
JSfAWIM+FS7cS0RjpHNi/e5MFnkJN7eM9/HEBcKDSlrQPKXZo2soIDeLPhLwqLb7AJZqIvbjGkau
bYsShpzBxlK+0XmTpP09HywqDPllioxcKJF0UUxQEzIL0pmchzXdoRcrPCpLB8tpKu9r7qW7Zma3
ytYcYKaNiezBHuhD77T1nL7ymmTFxFEJWD1F1mhhWWDXEFw9Wvz+MRzeXG+6pMw58gj5Q9I70KPL
vP00pU9/jw/dP8pbZJvz+lOaKS+zU180KyUt9otWlrE03vzBIHQHoh7EkeAUIPTXQu6yY3keZKsg
lRaEG0sia/p7w6gRxARGDJSWyb50pcTMU4D9N6IPS5dk+T85pEIOfMbK+HQjTGun0G2fS4k6wCJR
KRbvNT+QL3T6QSfUCQl8SwIj9E6ZSaM0+daokZLOx4TXEpR3A18n82EXl5l+6mFhxJ8CWnEKQRno
c8hG6cdXru7IGxDyXYpPykWCTd9s0RGqMKbbgQ9e8SfRFxlvAXgxWsT+v/M0XC7u4J3illwS8Mp4
EBONdlWsu6eMpmnLG5HBZqXK1CY35b0QQ2nyAXIhpWlaryqcINLBjvXE6FiFTcVvweZGKaIOLesv
coQcCzcJEzmUlTnYPvE1VInSU/s5/ClprluRmUw543yCqjifRt71o5Hlx4oPceJuAZUYrX8PuM7h
3FZMUHtpQOY2+Scm1xRmTuNLOLAX/jwKU6ME3PqjZdEJUWIe7BVt9olWc64Y3lUr6AgU+Litwepz
uPSxI9Yw0F4CYCLYgweDq+/tAcwj8i8eSt0OhiYmhHfBzqcr7qt0U6eoF7C8h+YqS23fG8HHdboX
pdQ8xNHeDTulWzF1In5uA2e6aCHxCk/+l5RtFXjM6GKNr55yDsdzDN99fNgBDqM6WRPXbBafzmEB
XYIMDPTP/tnaPTwBQzRiJhncpxqJcWSKU4T7dfqjSe8Yw60xwUYCQkVpDPDEG3LprCpUj84DSCef
nBvlzlhQ6V6q+lnXGRYPGToChUBcaADSEucBAZLcRPQ3YnGhdieks6pR3ygWrcvOduUEZqt/wx8S
Y3tE31xQw7ky8nRRUClwYugx7nyw/cqZO8raFLeX3BmhI4X2i2BBCBFw/aV9zyquRU+1B3D+IAZK
BdwnIgfFLYyMQVhQwDxU7U1x5tH1i1OnUns87oppwbMCvkANl4Zkb7nXYgZOqSiDf2EQxo8T/dDY
c1ODiwe7KF/y1Mzq33E5kqSJZ3VcSFVgbUOSMfHyxCkg+gjkfRxLmViu7xkbFPV3K6YBM8sQ1Juf
X9QVVtYEFbjk2xgMD+FYZLdH4O9obSxYp6YlbjWOvwq/v3xl/CqrA9C47AX3b0VloCN/lhjDyO0i
OaIuAzSq/NgFCPa9wVstsi/TiGbbrlyd/enD//BeMK9TlYzNSU/U25ExguW2iU6vAzgP6pvCBNfW
CDshGAF9zL8Yf8Ld+igoBAT/WTmYDpngPxuCWqXWfQ26v9mPBoyRNOovgsx9xAaW4JkFvs5kJuQ3
nevRnjFbq6y27D+tsBp/TpKeCeVbYfm6dSoOslOqbZiA0aizNLTsttpZXG8uvn8zLrdMXZ6NO/Y7
QdGz5HsCFyj0P5VNI8iuKGNfxUL74dxajsMMBSq0V5X3IbMxp3K3pTfKO6UDhX7CSt0LzzPlBwIB
NM6qRZevW1gAjMjWplLh1RFK5GUl4n4laSA+Zvy2AjBn5YiNrAi5k3Zt8CxS5MMD6LzMJRsZKMsq
DzTr/9744jR7q4AL44YUKKO5Ebgl/OcLQaG3dK2NJ6j3NXJOSACYWyCAp8F323WfG5DWIzhJvURs
0ZjOtTWlQecDZVYmRDibGb9pMF9JzYmqLv0iPgrRPcD9wCiKxFKcXPzLaP+ThJWVoPog/g1TdFwa
gzAnI0F+Sh9WSD4qI70KuOAgh4FYgEEKzyutVhou3haeZ+ETxayVXbRlass+kCL6pMvgPidRjtw5
3nmKlBKfsAAxjSuYbtp+wnLR4/6Oq1tWWlWa6ZkYdET77KaccvAiWNQ6kbb24om/3Plbvs1a8mCx
wqpGwxdPaw99okLPLRxQ9IddpkNT/IHzWavRDRhYpkJndDIBFzPp9BWmOb8BLE6mAe4deCTupSne
A+fxvgVE8Gs4wKm1lBiQPiGUySAb+mI5jj0q9iT9lShr52FChmC3+/rW8koZcCz+45tpfRG39nhQ
sm+jb7cGQz16PkKjfN/ooiC00ICLltfOEj6JmXfv0WJWgIif/Oqxbyz1khe9wBJH/q7RylwL8iOg
9vRyEIJu0uuMZ0MPTULjMB7ximUCD1uC2YAhsp5Bh2ICgma7RwuvnlQc1z9LVOUlncHwYqYH12ts
af09HBZEdkQl9+gEz3MuhL81HlvVN58kmqNUZsk/+jgjLPMNYi4o9Iz0vwtQfqfYX9ScClKh4/ly
fsY1UM1JJvJiILoBgJN8/gVO6r4eav7g/lW4Y+n1uT4K7y+CBaXFbewPgYTubrJ27+XEUyGIesqw
+YQuig76qmpE4kPeVwQ9h7VXIaEgJJp1ILSrVDOK22RO7+gfCcdnj0W2cut8U93Mja1ZP7A6K3/T
4eW7Df8vXebIGfJkqwbfq1oCkLCQzwHxHAjG5yo/s34//qhvFEQNq5BNM+OugM9C/+xJXpwYM1wI
GLWih4WMUXmMO5vwR/Ryjfeeqw2kasPFiR0mcGQYrYK1LyGO/pN/MyFtUGAE1/C/9h9LSeCN8kv1
cx51uQB+e7rptKBIZ1CPieXDQpQylgWeSJBO2pjN6CfFJ9ww5YgewIL7B3yPhilodDPtyxht18/R
2LZFVmScbRXbkLU8tIKyX9a/TemshVJr6BcLR691JJc0v3Kheps14yQuGoAw/Yyio8eMzyfA4iSW
dNypDIiwTKhjsoaHC00QqWUX94PYAt0z1X+Ymu8PDQQveU6qcfnuAwpPB80B4Nux59Y0rM2Yt/Ha
LuABS4uJM5gmcm9hxoAwexXF4anokRDZMwF7QZZEI/g6dXUP8raksWrkOXZZWoLoJtKyTOIawKmv
647EKuWwvBnFp5KcyFwHdIMc64g1C0gMib/ZS0ralJUaBg9hooGg98/8acqqyZai7EUdz5jTilQl
dNcBvI2FymuUNur2VqG1qG75golnsXXGTKcudzUJPAu9GwxtDnLmESh/DEzXwXOVdiZMLZS3+NkE
sLt0XUIf+DGODs5zuLtMR2Lf8ZEuh05jDSW0i9stnzRubEkWfjCWzZodWJeIz/UL2LBwS1r/vUoz
skuwvAahnzk/mioQNmiZv2OyllmzvydsJL1B9tX0Crja/eGX+WE1IWToG5lT/sfJELT2qtNHhEFo
mxalWBD2efJwpCw2WlO16EwJrTEjy1ITxutpLbLL6JwFUtWgpgBOa95cklJJGaKz7M3L5wsRTe+p
hsX8aW4G3+mTVljNN7bfI6KGLTzAKAaMPaiEryHqsOqOeUfBM/pQmorI5bs3xf3IMMUU0xTJTKYR
0aSvnYpySk3A8K8t74THc57PnvIlSiZmwyIy7jP0eiGSLzKRZTXJOEqecD2UzVi/Sa1Qv6uETjcX
fCVQ8+1XX9Rc9uCJrHHEa3pDFIoccCQg7SH/L0Amfvh+YZxT8t3+0MhyfdSjk9YGWWMYu5oERApU
Taka55Atlg6XIOStOyIpmddc+/5GKYfpqTEcslu06m97zIskyd35UycbY9W51Qv+WFMN/9ovq/LC
dJz8avVz4DRJ9miK6/3iqeFAbuzf9h9YrQtWOcVMztDbNJmpmecno33xCONxgOTNFSsmC3cM+IwB
hunuZx1gLcyLBkENLKCGFm2Zr/NoBrNVi1LzWUm73j3DzafqAOgDf0jRdIIvJXvezgvdLxPWxMOz
Vvhz61nCB5v3Gj8pxpNYQdLXRaaPha4TksfTxv3FLa8v1nM1XUfJ8hd8CpGXrD0MqxC/SSm364hf
kbjEnZzQYHc30bs3VLpnJ1soKyjQWDCzJ7kZaza09fTpB2/AFLpXqE1uLPeCjjV/IFuqmtKaG7Sq
dMUyhHR/a57zfL/YJlLknA/0bnOkpHw3RB8oxjBk+36kITvRK+QbcxPD/ONvfbwIyGxfXf5dFBF8
mS6uL+MvXbCIdi76ZbWAoYOj38Y+xDv37B/aEKVSsTUEU+SOkndlvypyq7LZ84HJo3OqhIycOV8H
EuL65AOrlQQ9XdFac/xUsW8okkvMpEI7K2nCI3L8sIv6NLMlOAh/Gk+gGOg/+UqGdiUEVrhHE7JV
Sd7SO5FBjoPwXioj71jOGfkfbfwx+0z2wyi/HLYOLs2tKt8JNKZZyWh2BBHyl/r9J8dT0N79dZlK
B/3mw4xWJGtBvZzspkjbl9o384N/GHMw/UKFoXfQZyJlP2U5r2qaKIhDDw10oSXWP5YU0pCwmQOr
jR6QcBYcxsa/tXQLHSt3ejy0HFfFMZeqf6aH5PWuwZoIIXqSqGo4BodsaHGS7QjnOMAlezYiA4m2
RSeMQqsbfjRZfQuBmD1paOPxHeoKF11it+GU2yFnMLISij61vq1w1ideEXbWj1w6LfobUgDhjhsn
Vw3LLw9e79rePiR612uPtdd7nZ6NW+bj3GOdt57DZev6BefBaD/yGguQY5VStTcjbUYpj02oRpW6
vcoLc/B0M6403Bm1l4uijzsl/caIG6LC5B+XXIS+7fyPGRwSD5ehwQxn7LXtbMEG2zXY2Q71yQOM
hDHKL8NheDWBbKgbnMRhwRjXL9l5F6aAEasjRutr85R198eImkvXofgDCIJz6Ksw9e35xCR9mrC3
aNxncsxdUMaY06cD5n/KRO7D2AtNbpvHhfNWIiI/lqx+7LhVILc8XE3HjlUDGkqy5M2x5BUsP7pQ
8Hs7kGE0IwkDlS9JF3Po87bpS/v6
`protect end_protected
