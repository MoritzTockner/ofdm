-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o3hjymGg6vJt2kyE6mSDGXf5D6ubqtUi/To6wr+9wTYg0PLmRCw52J/8X7xRiUuzO+y0yHtZY7e/
zOY7gX74aGsHT+bjt+UE3B4KMSajxbgqSuLi7QfPvW4MREvCFC4GXU07gZd4jqUSCoejEhnSN12q
SZMzP0Svi+0tX8DwR/HpmvVW48yNEmXvb9NPaQTQdYpmWj6GsjSdog/oyqojadJ5N7ZYqXzakBeO
J6ulGeNeb3bw3++OEiDqlcjHZc2Xb/k8D/5T7ZU6ouuNMbiz39EDsZQz6yeg4R630WDrwWQohoHk
eo1j34n4WYZRGMysjqiSQxp6hGhKqKjkv3sjPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2960)
`protect data_block
w5SsosTo5//XyEN+Xj3wPwjF7XpfpmBpKyAhQTlken/AvPEStTAwTBuzZrBRXVIM8+RU26HOeN/+
mB7toqPOtaemPOByMz1+YL1ZrW5y4NO6fzoO7kkKE93gsB6wVlv/VCDsfNNVxgW1K8TAij5uuqaT
x83FCtymg8300/X/p84alh5Z0s1bTcVDKU6DdwLS5aa9juYdeIFAPIISXx0P1m7yOIMJ2nDYew2J
AJ0W3UMHbwcsgxUM7vgoYdPgdyEIfGiyBWRABkkzWpcsiFUqbAarYK77zaN7ck8NqOyx50SN2KpB
AwMnNRPkriEcIFaQH8PuCYypJVPJNogGFZanMxx+aS2Yu6N8Y83Pt7kZb8RBwzmdkHqvAEgci43O
pxB/nsTysFFKlsAaBap5FVe2nqXxAP3JvWQinDah6dYbHC5fpuROpvKBJdu2kh9a75EDizw15k+y
fZ+dJ43M2VNsjkebqgFfwoaLceLKagdtnnPzaEF6PfGUq+uITYvHoJn7FMSx/mw3tX8bVA8EmbtZ
m5UeWD1lzpGkIfzJbs5InnUE+irTh6GIkkNwrMGPBGa+EPeYATYvHVbZZpXy7CxQjmG1JWg5TfW/
TX8faeV/WqwT67A8q+QthkHhEiX02TDJ9bjPvR5BPwv3ef4QPQWX6Jea3o7Ed7WRAbxyzCkXbhJ1
Q59Ubi5Y4oDTS+O87YQn34WWVBtyaju3iLI49Sx6Qv74K/fVTawf4Cp0FaQkAxV1KRV8YzQZFx3B
//LYC6kEsQEuRxiDt+k6LHVp3ItPGhqYLgTXb+2WeCgKnZAiuZiL66xWUX/8w7RD3cOkTw3HKqUf
YcP3De1ODriMcqiwe52JNDq1OssyjGUnMNpknfQ0ip2QQaMTsyIum1lMuYVIAQMAPm3cxqrObTxq
PLX1YaDnh0HvPk0LllTYH4Ll9mP1cySItejGxcSCcpVf592d2SW3qxnJnHHoa8+/boFGOA0StdaS
sKkuJOuUzrq2OoTm0FGdto6khtp/1ffPrr30X8Wqfy6i/osQB25m4ivIvJH5cHsth4T3QxB+c3zM
zryoAjDXB8B6YVF6SioxMqdJDhWJUP8YpaAdidR87DHrof74BC7qZlLkq2MJ9w0aqY0oPJoJJeZI
WQRydxblS2gNcxGxD1RUTunFawLCwMfUCzk1D6cTHKO5502mVw6PulCU2Zg9Pg/6UDwgAgYa/atr
FcckA2eeT+xhQREwS/lVAhGgqkPTTg3gT9+yIGebhsIeo58msgAsZtTOZlGZNEo9OFw6pgpwKs8K
9U4Wy8rFHD2Y6iM8lRjMY21DM6Q+2h+dKGysXro+jdLKcErHp+BdYmRUhbY/YMy85T7ejT+KXkTb
EN5eT/acXW0z19NzCmxANMhJmmJ/wTKKX7dOJQXLHUaEVR22QCYzCaQ0dp4ciduc886aGd3YEUqT
bjwyjYobAaYLBaltD6pXFHwGdBdCRiC1BPvj/ZEhGmdtGH304u3WKy4dVQsIbYdBXZMbVR2x9fhy
FsVY7Za5J6Lh70tSXfkuOyFxNy/sGaNXrK6SOHXt4QL/cFXN8BlA7Qtz/xr/iVfm0W2L3bKLOiOP
8sk5SNd52sWui8z5kA4ZnZy9mGGRQWHBc5j3SBLEEgk0uYoDzxrFwaIa7xz3Ilue4gX8JM7QXLDo
vd0G0EeUmVEt2m0s0G1nBzogw80we2wU35DwOh06cV5wNDSXhEsabvKdJcXtX0fhnA8a+f6MVlNx
IlvC4ONssuf3YD1FljUbSvdV6KaMV7d+is1gsLMnbjiNgg1rW2qIHG/pPlvvlg/FP+JG0vkT4Gsw
pK7loD9H/CxZ77MKGNz3sTa8ZIr0UgF9lc2SnrAL61Ts2kAqu2TO0Sh1yeKtZWE+737PMLdaN7Pk
UWkY+b8etMfbi6YOkRupQhY5+qB2/SviA3AZHSb+YdCS5DjAyZM5wHSH9AgMjDS4n0JTJyN+R6ig
dknTDWbaubWY8aquLlyVPZgxA6GOPp0xSe/rhpTMY2QcwiDV1Z0fOeKut50uD7szdm1NUI8PObHk
iXWkstMzCpYksyd9cu60z765Bm1nM6+WEpkNUMIQzUfDpkqAcOvu6m6UfCeBwHlDpc8Do0Hf2PgY
3WeNR5mhacdcoBvRIZzATFvqGuMR1oHWBlQPzNLIDTBxqpNns33c+6KEXd0r1mbSX3AD8riKdUgc
ydMmC3kRssNJkhDZq8kyI2o8z2tdwupiCbD2h3rkHFBYnNxLMo+lh67OcZtgvHfHiEkz+NX2V3n1
0S5BwZeeQNpOb7G1rR+0t3XFWh1SVPOmNtdWsD1BncR/ER+6u2X+1A22i+l6KJjhizXx2yX2rlTe
V2fEIANAnD8D1U07OPLoUeoIxbawcDbMKWeXpYdnxxkjt3OPzQdHUDzpYdU/1siOtAuEOkvlGoAf
1Lqmi/cajCWWSkfUUX/lTOvgBylCmlsM604q/rCY7NN5eHLirrr1E7TMR8DjG1v+R4RHMs5sTJF+
OB1R/bFYoYN6Cz+QT7JcFc+f5J6Uqm27YosbXoB+FDgE+uN+/4sEbBwiWjXOwhsBzDwEaLPUyGx8
TrrQ3Pws2GSYaPPHBKybi5i981ipLVF5Fjch5I8uYChKEGyBHuewjSAX6dW5+Dij7N/9ZN40+hQ0
A1sXqrGsXNmlCSkfuOV8QOKxuNmswUpYvEUIpA3pEgpjI0HS9fPCL75/4ceD0MsmZkDG2x5QzXfI
68rDdMO1rlVFvDSJQDvac52wdvZ2yprrQd1PfiUzcYf1GRBgvuUT/hlVJwn7fw7b+A4ySqaYhtRz
VVuRi6JYZMVzkttnjGIwHi3KntrU+71CmeIt0q9PewM39g2PMvHfxO6QU/+Kt1EYfPi7jJSX3IGP
acM8qKh92lmy/Nd+NRXNmy8l6IDNB52LVitP32GN1e2YjiSY9HwYY59BDKupq5BgLt52pXuUu5OG
01XObB18PWNNzyDtdcAQYOCCQlrLc82QWWk6pkQIxvMWx2FJ1AdYKbz0Zslkv0uGTvd69hFx2SyT
nr9RVX7HIBsQHOsJGb1Kr8oKxjWe4dpyKUC5Ie0++XHHFjfBtu+L8HTrifR+/c42qE2Kw7MGU0wG
ZDL1O5fd5/DIfW+x33XG5hboOu2xtPOh+/Sr6LdveFKsNhnUuztRMQJJ6B0FUt4SHOB+0k5rTzAc
y6b/M073izKO9+yLn75NGqDO4/89SkKFaXCt/+6JS2PsKf7rSNlCMKhfrJybaGIWPECmaZQk8nj6
nLJbsxqedpjkHJVBlqkJrfI28m5XkhonuNNBpsvgcCAO/I5IPt3pmX4mG223Hnpeaw0n2slnf0jJ
aWkvrGuA3TCzK0qyHedzJn5KfR2yICF6C36CplvY2l1EWzteWvohnxH/AmWsf3mkzxUYXdGkl6BO
f4J6LjoZbB5aZjpDLa879atnXJW10cgSByrev36i0fozrr2BnQQIQC+MYCkA7rV/5Ul6dWwIxwgS
LsJ852q0QG7ezyGn2Eaw2XJfD3QRikdralPYK8hbgDt/CtO7pmmBRstubUBz2RIV550jXEemVjH/
MTaLnf5HhapEaYbBcY9XofglpF8EHc/e7UxNAESzyWmCXm+js0slUUcq/+s0rIpRDO/c8ja7Mu4j
xJzW+LIBOdqsMIbq1BY1ffUisBWjyEFqvZji1fKHPtO5s5+uUnvST7giajLIJp8prGGCDkSOt2Cm
0MXrYNok2XUjkdRwtWCc13TPMA4mYK7AbTMZwbwDwUwZ2OaI/9EYitkdQ/SlyUMonDjvsIS+tHLJ
T7jyCkDzCDIyKecEd0QN9XX0qcVvPBj0CWFlw+ZLX+qZ+EJI4T7CpkNMTBJyeGlNOiGPlRCBxPGc
b43Ub/nzIMERU0nstwTM8506nqHzmtk5zDeFWI7VE0O1wPimqgVlF8s0Ap+Y6uS5zrLIdJI=
`protect end_protected
