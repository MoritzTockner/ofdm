-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1V4ryLflP2xxpkXOpAFK2q2orejKSLf+bvuslNGgMdJtwmGKLyEziotOObh4KZg0VYAyqGrmftHN
q6N84bT51VzvQ3jaCAoYmqsBTFe3qksPR5iwL1QUeJQkCB66RCTEq5oSfbenX6WIAsGE9ts1N5py
B6dJsX7sWlGM2Cmv9t3nHqCuDS5zhQl08OgtA3DqmWx/nswLNVUFip2Vql6TQmwAAAjTvNxCUbXI
S0TBlCmbiviZY7IAOgRV79I3qU6YYI/BTx8EKE+C27BmyXBu+inZM76Wr2lrT+PgFwRd0nmUHDNS
yjsQH3WiT/exHzcwdm0lxE+R0/yraIhHA/Z93w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
4MkYiWd48+CVHafLEtAeCjWmvYhUb7Y8aqVZlBz+5RR4VaU4b0wYIPoKC1OnvoZZBsgYju8HeVOO
NXAeg5wXnfp58kwtkROH2QigOGxWPj8h9Ww2Zz+G/pKPadhwHe5Up8Y5WGrmcaVZho6hSCaoAKNv
k7i78xh/ZOga1NlOLwmiZA14tpt3hK2iJaxywFLGyyVc1IgNLVzIXrFHja0qKEHqxE1j8ZNc/We8
AsUFMf3xNXk5iZKzkPra/Iwcfpwp3BIB79I5SM5Enf8DCg7x/QcOGryv7Uy92Uq8Kd6cOPPGjMyX
/ysEAvfXRKuRsPfiaU3G9/Lwrx7IgM1oMgvq7oIyqaCkzPAN546QwRVeDGiQeBStHTQJnwww8qXK
9P/WE7LWLzAMmwuJGo7YJzk+oo6ZxODCnBxm3z0QGoUEXoM79CP8A+L4SWfJWqCs+D8IEvZ81cpu
ViyW2C1/45/xs2/lgFODoZTKacUAVCc1Uicin2lHMdNvUZsC4VaB8Eezioe5xbjXhefa3R2a09qu
4wnSTa+NSLS7iDl5zbGtc8zjDPMOY9UDLgqM0dq6s/YDo4b6ymBucjJD1MvTp4Z05qDSynMfOqRx
io8PMIKuOizMzrFFJxuS6R+5o1S2p2QStrhVN/EQMEuqgo+2zcRq275HGVD4A8fG0P2IJbn7Vgv7
wqoWHjjASezRCsohcmd/X+g+t9ERUcrp1DsOL2IB70K2hrJei4uSjBkjwGHx0CtSXkmNRsxv+Tym
MCllDZfwNtm6ko/Qic4KMwoLYnO5B62v9QSEJnKHuWtW5KBOhL8jzi7YcL8tm/K0U22L/FYgXd7l
Twuv+vKeHytSGNOcJyWEAcn30b40gh2R+7Pa0mgMwwOzvD4hGA4qbTNN5+DIdneSjtwVEJj1xItZ
fnYEZsearaLoNTRZYqlN5W3wrqKiL/drwmSpFo7db6S9jDeK6VPweLFr74A+FwAL73Mcejtp8z0D
QVTuFO7oSxTUDglQz3TJV7pkmemyorR+fZdm26DrXPi0jcOp3kVIYpFIYbnQZxXMAnwokNRO1hMo
yylcyVx0IX++aagvaItXFNYL+vN98/8eJk0hro+T2CQrNUmsy6hvqO4IrVCb9+Sg7JsoCYfJLPIH
l6Dy75Gwba1oe6X8d6aKa5xqgrI7DcDap1jrCp+3E53slnZZnS16j1u2NvzdkEJoqSkaaBc1skJh
p5UjpiEUUHRYYJ0Rq0DBfv7nYpHaramf+f7wKWP3f6RrryyAKsucVpItox5RWqWKSkzeVH/c1YvE
vHzZaFZO9I8bby10O4zjINWMQByOUx5LnWdwK1ZCT3z6Z1WbBWAOiBXn8+SxD9HzsiRqo10v20ak
aUtHmrQAwBoutQd02Lu2ju0auy1gQJLZSLC45pyrWRR/1vC3OJiL+Mvzxj2l6detGBwLID1NYPDD
OGKEE4w2hp/QrPScRMN55su3X5y5DR5cEcQRrIEOh/nzedkgaMRRr52TXQD5fGiJRIPN4x2f2R9A
C42Dz+YfV8rad769LEWYP5OAAsVfPkZwkXmScfFQTXpNkepomLQyzV5VtAIByoiQOwGJmYDD+Cgp
bkgmfMpTHQ5gSqX+9NcuitoZbnyx8MiAdrJngHt74p10fFdp2dUYBXpKZAfho4WvtCdgQZLDSQxZ
61sGXyj36mnQ8+mPOi+6x0hAVwDM8ZA2CJW6dYIIJLn/jmheTUlEjoTf/RMzS3qAxim55zKA7q/r
ZMUc7VzIrXdcNDA3Othb5OHlCxLxNUARQTVnOqdAkkztKHGqem985AD2U7GUdr+AeE1ZFhcHbvpp
t7JRQtosa1f9Ojjwwpj6qktO8ZdDx3e7EanVA1tYCTYRok5YtZPCOXrueMmTarqkJWickzCCw4iQ
9Eb66N3cr/3RU7TTobZ/e/U1P1UwSG0A1JFHh+0zZFjGnaewxIiEucvni9wfYLTN+9JnA0s59oFS
BXLTKMSYdsRCi1rHK+QZkQmXhEIgnVkghV2DYSNaD0FN7LB/aDiZ9COgZVrezglHrk5GGt7o4TOR
OSTcSem3vNyuQitYPdGtDCCoJeJ9ADAQ5XoYYfKO6s5IZWgCMc0xmAl/a/j89VEueqcdFVq+Y5e+
wVa09AfwMpIiJavHND6uZ02d3ifPFtK6pKMR6vxjVl93OqvbxhE408EMfuO1KMfzi1S/w6ITNRrA
UlqXZzFyVNJi+6Dxh27DY4Q2vRcsYozjgUxW6j0HSu3klDQzRsstjrWL7nCrqhueEhfLPjCx72rX
f4kKU8tGbiP48OGb/TDn91eCuwx9NL57Z4MwW2fFL48pFQH3hJVIprbKD+T7kym5ndPASvhrT19Q
7TKOu/ccErva8Jf6jpoc7fed/oYWUo7DJxf3EEI9h71VnwGkXsPryDtNJFKyvto8y8CN9rvb3RM+
sHxUpkKD5BLS7AkPFxo8OVHHiH6J3RZqDflekPUO6Wf7W2kj6rF0IN6Yew9vfd4e1YNWbxkBEmd2
PnAst2ZMg8ZJyVv0c9suZ5x/5MixNOhuHk/gPPkIHYppaLG6DHot6dYCRENIfW61Jq+3UfAjiE5F
5VvTtnujE6gwINcokh1rN63eEGzA1qDFLTDgMKB7m1A1TzDi08Dt27F1x2OITlgg959ulD+qYnxO
YO4zfIvSEN2+adz79S5kwV14xYu3sMWyy7Makg8M2RxeubDq4wpghphLTSqHb6i+vw4NTcRqJKbK
sU0uI7Fz2TWLLxG+eoMUzWqyylek8NhsWXeX16rBDMs0eYoi+GmiCHeumF69mgGkff45Uj1FJMfd
bHxWKCKGs2GMWBNma+AvZ2SRTW2iFf1b7m2ZgauJxep/78R56uAmLR/mr0Hg2Ub1Eo42tWW4q8cP
X6+lk6tVsAcSYPHFnuIXKiCobzG3uFwL2JK9sdwgqvcPNECnlqnREL3+LEctj1fFpsrh8ztDtPYh
dLEy9o07+dKbImqm/lmgSXOTqMyeJ/c+BOrjXXN2GQkkmir5kRn+9cHi2kjwoXhobvIjKElSpblQ
NcqBUFloeL2Pg+wPE/J6aBp7jtZyw5OHdIJrUcJ0WvR7nwJq8wdqF3gVEqPFw76DKfTVPs5JwR01
Uy+cay4q3wqSuxtuynTC1th07F47j2qtDJ1GFA4j4Mciw2WDoH0tm8Dp/N4cVp+3SSYTSOSeG1AR
MdExMBnqzJdQw7oiQkayjO5FZjpnaZG/H3waQrzTRDQHNQJpFmngkZ0ugQZuHsy0cmAPDRNBNQ+d
QUnm1k10tCWanzEHUwYr0iN93CBYu8jk3p1SpjGyUevxwqZ1U2z5ht8YEiz/x2t81LyPw/rYxvUK
LaojShBJALM3gPkX92Z2vlB26S+00b5zoxZkMKWWPX0AMeK535EKfovwOvzA5yBrpuTgWJ3RuywB
x2fR+pVabK74XgGhAQwkIr66N76XJqZzsy0KBC1qBJEPtvEnsXusa1sWWSGhBvxCd2UhvmEJ+OEv
StubZ3dd+AN6JoXy5muityqb8KFxGCYz9S3CzJMV8mFcu4dMLogsKwgKcDHQ0rlr2FwgGE/sStSt
lYeUQfWx4cnvNifqGec/xdluEp9cXgwKJCPpmufd7cscgnpIA/8Bs71ELmlzk5SyXMe3CORU6zcL
4teNe7OR8i41Vzl3dWNxqFz67Wj0NoP5KnKiO76tgIC6XY07qW7UrSTrWyqnsisa6rVTx+dODsQH
gpcBmY56NBF+YnR0e/raGbqW91HT6pYZFFHEdvsvtJXGuXqV7PlmoqzvlGzva/fT6Lx9TtKyXzK2
U2vzxDIPi7SGweA+iTNaKv4FOIFSHtOdAYvRPSFTrC5JxWF79JiICpg6XOjBC5/CsDEDF99OFZYZ
8zywW0hv78/pbBLdOJFgdVdSt/pDSsmbc8bcFjHN7pJOLf9unz0inBBe806VJnIpT+xQ8zBGGuMq
jxpldnRpKblFQ6rzEc6siKYY8bzcQ/d7PBpbaMyB5O36Qm9IQ6KVLjdV6msOpacGXuLS7G0Xiq1Y
dz8Qrc61PWG8XEj4XrFjLTIcsyqbhK6AIeNSA/0mY3HO+q33x9ySfqTNA1YiLwuZZcpeB19s6Dtj
43uls0xf03/D3zieVeKOnBwOlptlHOsP0ukQ+OS/AVUBWxjZ7RbL2QZA9GhBYiQ7vsxUAyDiXPPA
0xjI0IRY40AMubDKc2YUSs+cTBBuEF9Kz9i1bL3TYdUq2grj9j7/H4t7dkqBN0VjMBgr5tD54M8L
rId2cb2WEwJz7Ri5gJ3IVcWlBdBJkDJHYpiHy+uUKbVM3AMLKxhViKLioOH+ERhdsjRWgBmqKJOP
0Mio8C9HPBxwJ4eYMZkBRBLs5tRtl7sk5iGEf87xfzPiltcGolpFaiwXayJ9/Zk6v7Z1UPeRgwvH
gDVBZGClUTy/bwZbMoZqV87fHvy43TIGqk/HqphmmNw1L5pYjkBq2SAfWNu2JZczGV4L6FcICYEQ
KliPu34Bn5QVKY+ZapIfvosIZYflCa70teoJ7RpHuWRwcCj++/Ep6axLVO0PudkUQ53q1ZlVhvTU
l2226iGFRH+u9yg8lFDwTUhZctTEi4ABpqmDOnnqsCazR/OG7PT7ZbeqayQez3WY8UlFDAbBO/hI
lnE1jxBGMtHlKBoF+/xIZPymIYXTlzpO7Qpp46N8vnKtwXw5cHWwdv+b7qv4jIkqxJawRE6b+QG6
AFqNdmnS23ksqiwTVTOZZ/ag+l1F/xc+3ZofVowWnjAYc7W2Q52SaBseC5XVzcEjp+S3GPQ6CCOK
qrBlWnUUHqFjNpumeeT05bjv+mBvG5skRHMkUE5NBvLuppbA7FQMFGzZ07GNHD6p1UtBoagDgyWb
LqOMQTPRzz3Wbg+YrhpT1caguoPpBWsYwfgE8MfMZGKwE4VI/ucCbpLync2TOanWw27PW7GeiYsO
zq15mIP0VFhBEPTJqvqxGY4eT1ghHAJG1SdUIwtzfr0fPC45MnEfyyfp6DtLhPo8GMX/exlFH48t
6CvF4UR6v4GDonsF6VEhH/91+KJdUJZz/V8cGVZbxhK8tWH/Q1GCHqVh43S7C9zSL7RFSDkyhRFs
SGDFYp0OA/xCUIlMM+KTMdFNQZLegxa85EcXUsm4pDFY/wlI+fgXQwnDjw4mGy35KklA3nVwvmvL
eSezVMxKOMx0v0IB8zgmceUaVxM2hzVgeKnbyW3rrMtZCiYnPT2vhQUcIUrd7NAzqWL52/L4W9tn
8zT9ZpXDsLfAjsSTP1K/GSbcYy7fF8y5lIonb7yvetqBDFVYQ+d7fSHNPvCEpX/SnqSe8a4b+Pn7
rxMOz8LMjCClLOUfDmDD9LFVWEL5jD3ZELlISLBd1vXWD2LoUwtDlfXo3w6Qj2dQmtRlA07gtIdy
8JfU5ZtXXErS134mPy9uzAMolHLgDttFDSXNdbZJMs3/1lP4Osmx7eE4Y1dQ27jxcfcCojrXw5sk
as6nF4d/zEQqV1M0HMe7LTrYL8hx60XkX0++AVoskFCJ8bR6XR2cTpwv7PDgafyh5289Ip1rQKGr
JVHp9dna2RjuIdM7aG5gXkvyWIl7SPcQAsBHh0YoqJCEWfMZB4T5adRD3Ow3bp8NgJgCj+/YfQ/h
TvcyF2VMUJHwzRA4HjsDH/QE+CmA4rgBkH8iD+J6hY5tZFpw1aDLxqj+Z6EaVTKq52F2ZxGz7Anu
5lxm+g9nowubPKhspf+AAvW/NeJMgAEMYdeCPpEme0ZH3MCqa5IdjzIwkE4d+Ly/NLNpMbQDRYDF
pDuDRh41pOEVQspM8PIhE/382v69N8+I53SYt9/PNnnaUfeoivOphmFVyPKNfnJTXxWmINRvCi4K
0SHLBQ1OZjNlcMJZePmnXV1u3DAfztsLomLB3ul1QsZTb4alTSxXuVUNkMlHqXC9zPsLABYc8O02
ZOphDBwUzlb968tW2f1baurWj0F94U3ix31X/tykZbgfYpJFTNnB6PepCYI6ibm6HjTCdCMF82dF
y0aX79nS7Ywf/JKH9ib4uezX7ZGhtTwY1KuRfVxHRaCwHafB5dQDvqgChMKAuNrC3j8hgdijTpd5
RcEpO4pgNHVJkRwg/7ZwxvmAn4TXiCyLCmQWwAvfHYqKRHz/A3o4PLcZ+owk9JnNYqOaGH8qtJH7
LHE+DWlGvOSIM51QhfTaJ7R70RyKSTI4M7VU2uVl2CweGS9Ip9f5ayzjvozS3zDbOOiMn72mPayl
Phwv4B1WTt3AmCa7EIRCKHRzd4Ta6FLUVtafeRXKPn7Ad+toMdWsEalaLsk/5hsc6ywMyRLUToQM
Ysn85xw7NtrhyS5lwkry0H5YsJt7sLMyeCIT3Ahsm8Vt8Zbj6nK0q9U33Wz/PHAmSQfGtFq5Jin/
FXzsjsUWK+MjFxga5hObvW1A/3CKZiakuVKqW73+h4HrSc1aEzYjnGMfntlojnOEDUgbvyGkIHeA
9nGSgNt4KTNd6Ymv46cVf4JLuydoO6fH1YSn18AZQG5+FjZ8rSwQHVzZijAbdnUHDmUq9g09QAH2
nFGm90EbKCif4hPvEOd6mGeh/ZZ0dHI24y5wI+4UUjGo9VNvULcnDUOvGixGlcjDBQ4BsSKkYDzw
gnoi6bEzYlWWT2MAXv/5B2AAh6CykuzCBaoUjoRn/rTJETyvVdgEl7V0JGGnJKZaQmKr14ze7s9Q
g5P64S4c9Plcti7q79ksgGqCz/djfvYeceVt4pqnfzYrdH4bYEeSzAze0YfgXwYRX0acYl52DZZH
YO2L1OXxsBkb9Q+1b66CIQGuVZap87jImiiFuqx4grQKLc9VbSHOb5BxynDkSztmx1HlFOMFeg7x
tD8M5gfUOk86t18Kb9jw4faAvn0PUIA52AUeYXe9Bmn6rMikXHnmlEqvSexoOsgVSf2WtCVchqSe
0F8zioQd+rbY5hyE62nDtID6PtFhn4cJMqyDNb9UWA7oK5/6a8156rVotyhbZO4e1ltI2hXlj+is
cDy5pdEyxH7uOa20QqXdBYIVfsTORG09G9gvQ0LB+XHRPJguOz4McQxk6NROyihYOEoWfEDEp1CF
P1k9/DxXc2LjX3IpEtUVTbIMgB4mRyG3EYUd7njlYGydtn/Ial/WwyZSUCZbEBtBm6KJ5MiiPuig
2WF2LTUGDmVeiHYSTzLHxFBXRYpUjSSl/pQMWrt0HHyJG9USTo5LYc7ljIdN1Ned+oxDfET/YHmH
MrAFnJXJ1vTYLrvFVCZRtXl8ePZGm0Crz2ftVrYa9rvCITjbd44ylN18mojbp0JWKbty79xli/q6
INRDBF342i16pn+HN0rqbnWGzs/Yc9rj4BGpIUWh92Bbsv9t/MMf1I9Ub1reR+KyT6ExnlNt4p5U
eFyOEw/1uu03jLCqrMJZuF0u83n3eZ00PR5ftWgslW21D7x4j9LECn7pFXljLHfbstND9dj3FMgB
f978Vy3AMmts9lDc1LdlOdcf502Xv44aaZcqPNmNbIJqrHnzJWtbj5yg0RmMzuINvqoWIERoz4UC
EF52FLb7Y1BmQ2Uwz7WPTIPM74FWCp/ChUhC3xvKIC7HvG7A8BnkYk0roReHgUXosox1tbHPllay
IKLsy6TkcJudZ17ei/X1ejxkpQw2RcVhUsiGTjiScJoHQY5+JFfgTQyeRR1/29ved+3t8pL9tUKI
M9eR9FHMC8TlAVEzALNplYABA22ZKytgoxT4KG1GbktoJ9+et0wGdOmdBcjTvy07fPRCmKwlSnfq
MF0D4YnX1btmBdypU4G0bFyokzYSyoqw1fOccNwTQD8aR03MtCTSIvLh8zMsaNsap/L2HRwR96qE
4EpzwVR66e1A95iMg9XUHBk6SMXTsDlOtG3AkhpwwTo92YOC6Nq3PMF7Gd6YOx1EQUTpYgAkcp3e
BgfduGtYZnO+jN7IY8MdOFSV1MgayjZfNoo70FpgeaO79zaFBY+icjKcuxFnwRGthHD/xTJt8+WV
/K4dKZMwqsaqngpS1zMAgEWjMWv85ZCl64ShTt9v8luLr1E+6yXAnzP4ARq97r3owzmOfia4erpN
L7IbJj26qT/LnESVSS7vdjxMQweTKbNj3lmlsWvq0DrF3Ceb2oMO2/DRiuujeRT2HIFZ3HW2nFXQ
vrDO1EfJKR6CvjaHc4MaNIM7PCjn60QFChkO5j6RtHIMJbHWuryREGzYAYEIitbP48c2Nmy5xb0n
cjWl+V95tLg1Hpe7nuohCzjRHEBXkn1GtRgG0AEdU7NUkNhn0qtPszQLJ30uqTn2lcDVZAnA9zvR
XCoHYrBEXhxDq+bK+JMbvSaJpanuBpMX9IU4dxnvLPk8DYCQ2l7+ojB8w/rIdNL/kbKJk3dUPrlI
K7jHuQqMDK8z2WuR0hp7d07CsIWEVarf3eNxxL42DYHDkdrWA2ZqfyO3+gfAn7cvleMP/d2IXaHA
43HKAdXlbRpKK/JffRdupmDWK8YwP7LMb4F0NIQyW7vR5/rVeIvVukZ5ZrDknIGVAGmwhK6nz7yE
GyL4X4zRArstCWiO73ZkHx+H+zr3zbhmx8qdySdBUo1ezpX7q1FW0ldTHT6nNRMnBtaBN1M+u7X1
ndB9VCGLYMC9e1XdgHUVgQfRLElSgpdZyAR1aTijsPAd1l/XPdQ0NOlCzjTDQ1keg6XzNNGQ7KJr
dGCnqsmYRdoJ8uglIg6gLE1tmZqb9cJIbJOhku4RN4YMzaPWxjWql4X9aZcfeWRtom/+EPyGx9LS
HPaYcQ+0IaJy4AA9Uj1dd+/DyrEjKT0AdSJfqMluxY+xLEKb2MOaS0WgjaX8qz9p1yl3WOg07V70
hPaz1JDJzsOK+o6KxpM60eIWpV1rjfQ7ChhhkOyhEc+GUTXG2l4yUPDOyKfftwtzYWUsyyBWfiwk
vhCx6b0e/3QgJ+VvQZUkPu6zWrzyYSKI5kIvMj6NhUIzIlhICVfBpHzwTyb8D48KksSu5XII3sY5
BksXBjk5m4ADG6cFuFT7DcQ2Uor7kJNhHIpYDeWAhx5q9NpDs1vTfeeKN3rPz+5uGmCP7vWZfxn6
LKYWumLtma4Cad2YmcFBc9hZMvzIFLl/QWVw3cfpVBq2SCw/ldGU/nctRDJQO5d16t2NA1gKji2Q
zCh/5B4RxcGZn2bDF9Fu6Nal9J49XNxjA35PKc32BJMsehccJZJdfbazCckZyqC52BJkE36+Leej
HQy3PwbvMqapcbIzTcIN16AooE7JsUeScmmEReMAN/MMxUYreeJx2lktnv+RWDaFztO1WxNnxH1E
scOLkIbnkgou2wOxYgR7ORILCzStsIyzAQMD7ZbBFnCIDU0EWuM50X7TL+amCA7x9nZ5EU9JflBC
XLZFoZIMYh1G4WthL5VU3YjyvqP1eDuV7m4B3dnTmi1t17QF27aM3X/nmrCdcFXXvt/16Rp13/ll
bbJjEPvi+KdK8FyB2XiNQobgneGcsQqaAsIUdVPWlirQYT9/PH8pLOc8E7OgJGyDT3dJK8JD30iP
SteXVQXfnM9uuDmOGI5wah8xddlZQF3RuDfPMi31oH/VxC9YppqVXNzmHXDkID1yBeRbKS0KWhZw
rzvAbZvKS2aIscJGLVCug7EKUdFw9A9zTqo/ZABf8afuMpEh3VoBCE6rySVkzeIurL3dqNZqd/Sf
GoXRDRnv+TCin87gScx9aN8UFgCLeqGr/qJcr7sJWumOUd5DLwPR6quQRFDTfp3Hol2WXLSCrXkX
rtDcxhV2aJBcC944aRg+PhPwl8rVbLlBEHxA/SWneiq/QNqMDrgZK60AEs74bKoO69z45fc58d+r
AwJDy2oC9PUGC+JQtE2oUkBtJ3+hJ2JPZ57urloCwRS/yImohuSJa0i9uSvWOPcusWPf2suoOul2
7CYXNZfb9OM4YhGNqTZ59RSCHVqfdv2BUjtBM7AV80c+Dr0VvUHiKb30PzOqMyhACPES6KXuiBUQ
XbHDvaeLMlVrHGTkqun1aiiVGPqmyy/W0AD77m92/nELliGiiNJLnpO3JLNAhiMwciVfNYFSwVmE
aou7YQJGb/3nHmZ6xR0H96C80MPE3RcTii0phNMevYTDQh0vRqLGTBz6x6qZt1yIQUBYnut2w+rf
0eKp2a0p5bMga1RLL+mR/mF7+BXkBHsuqM/CVKJikIvIC2twiDKu4471a2tQ+tStE2arGu251HyE
VtV7hN4Xf1YlLOvhWg1rSHIa6OQUHvPfHZcYQ3Q0CwlbjqAXzzxt9yGckhXXATuL6E2LWZ+1ukvr
5GUoOI0EKTBMO2BxQm4iZED/VdtkUGuo7HhRG37Am/sx2vyzYBFDxIrW7dYMBoIIzRHTSW6e+yYW
k1iDhX/gjmoH5Zg++14AIyuBrZNRrC3sM/BHgMGeqenZTOujqAafWXioDGvYHCT4LOi5bes5UL+Q
I07f/inOMD8ljSA36rMbFPNZ3ZCeMVx6FObNHLkr/6sBb7SQIxwZULzoMk5oGCVCn+jYDKo70YEH
C6aDCMKhO1vXJFMfh/rSI0xCX0pHQd1lL0K1GtyNHsVGoSupMFWqE6A3EH6Y0GAiDwJxTeubxToT
qt24kynmLPKqTTirJoQYNeEtJbhyKg+O4hjJFinMzCQ5TloGyilW7Tp8pc9YA8zpUsCrQgnUAM/w
WbveuOJg+yNBvjVCRLdH1iRgG5jN+/a+KVR9wA+FQPdNrKA82zlk44gbKWpUTFOXjgde5MgapW7f
MLn+YSUmQhEicm5aSS60WDERWx95BaGuGprqUmv5gup1iEysiGL35000MBo1ong5D7tLmAi0+mZO
4uQtPy58mtZD2crtBiMqJW2++u6xZinFEYGNKa1EN1CEtqrXSdFJQAvWW9W5L0oKCqg+mnEMx9OW
apWiO8mK78i0QOGVndmswi8m8rW99xiK9al25Fk5AY90q56CvtgNlRSxM2FH5CMtMBERA7XO0Qqa
Z5GUkL3gPR+0Ml2n9mJuVIbAyyx4r1t9MsQe7GPWNzSbqM8fJDMP5zPD0EBFeLYBaCeJkISgryZz
+Xa63KdXvJHKz0w/Oa8KnGOOGuu8g/KNnad6IT+KydS+KZK8xiYYWYnAQnW1571olUwBJohwqyDo
AZwPNfYaM7JhXbC0ukiAMIQKtD2vXsPrxoKdwGz7gjKoVVhcpgJwHgmkjWY10K2Kw34nw6TON+kB
IyBPtsvAtAzModAGyIb4icj8rIa4BqNG004dow/IfPBpqYxVbUhAxcnbKD8y04tqh48sOXyYKHE0
wbOb3aEDDhF1rWtKTmOoYaGiFwJGY1XN5wuMU5/ZcLxasyw/ZmThjlsfTfcTwC5fz+SzHIONOFK/
tcPPhVSHnBdQ0i67AOSyQqDr3xM0qSe3BbtksGOiO3VByZ3y62UkttIyvltPHzivgM4ZV1NSF5Gl
FB6tMVNEYHrZi2EEINECuOqPvi1B9Ce7BLfm1cLyD0XpIkayKc6vZUAjx++0GrVIBplCXFvWTWcj
EzKC58ALtB1s2c/Lz+zZOwL0IauKCsSd9WESN6AhsQGowAkGSkTQyf26HF98d11/+uR/sN8N+9DG
FvJj8xwqGqtwhoMdECMhmPik6DVK3Fnkmxvu0IQKPdsrdwN1qVEDpwJ/iuNl4/FRmGbW025uilWH
xLgQpl1qLNsssmPiXfxc56xb27zhI/WRG8WWh0N0hMT5JxOmuk6tweXIMl+Y0oy/+4SrxYkzR8J3
EnAOjURAPGbbaZBGDzczYC7tKTVmiBctj5mH0TKiTvwpjnPS6s3R2tzOA5eNoU/WnT0oQdlBU5I5
ZJt4e8S1LHEa4f+QvLbr8+GTNhp4+IxEszV697F8qlc9WEEmqxqgGlfYjQH9JxdlAkpCEZjJ3Ej/
NC0M7gq4oXOv2Jpa4A4YKabJXtqavbYUY6e/18S7hUGJlEw2PiOsofAjqvdqrTgxJEwtpTuVibG2
tzdZ07w0bKFFbS1WC63DBvouaIJIlV8YbNxtiObHkY0Um7TSJVL2ko5054zyo5k2IqHLeAIMEQRR
tsmeWUSIHN8/ExKH0tOAJ3NO9nHYOTW/xs9Fp1wAYEb9sGGxOgy4v8jtrISq6uMMruLHAhbMZZ78
6Ib5Qz7xEKJQj6CWCfK8oWpucCwu64aI86n1fOtdtNJjCSLmME+6VyyG014+yyX0z7YRouzEXuhY
t7K6o4mqtobA2PVCArnTdRSI+nsiE8cvem89+GIogWiv9Hl9RwUf6mlzO5OR57kAfAEvhj2gSGXl
h6Igf8h9c+w2zI5CLuT2AXEq+8BVXAD3pBv2zkoBH8vvrPLi8f+gX3E/D+a02GK0xy8S0d55zj4+
t0FlcTXlRXHDiv6O6gd+cYOBwhQs+kxJw1hHh6DKLth2lvhBNZP0mQcP/ESnFusF1xjVuh8ja4YV
IEL4NsC83gtT118jq7C+8iKnfeITiJz3qnBibhpN8N2OoZa9Zcocz7g5MH5ApyiH4nk8gUigk0lJ
7faLI9Vq+faqppgrGn3EkBwGwsDAB8zehHBlIU4RqmZPWPLCUIeWuTlKeCuHgKr9pvlYzYl8p3f0
X4Ke+lrkdWHyixAjtTs+Ghb0ZKNSxrDnhkZI9sDVrXltg4N6dP18S8zk99lmxGNJSkuFsPIqgd9E
5CpgToglYr6gxqi9vuLTe/7f1KwQfjT3WWG016OSXk2XkcIxJg1oB6xgqSTA356mgB+YfHbw+d+H
6Ut/YG8XtWhSDtBdscP5bjoPjSmJRug3hsIQ4WAtYId5hWcBr5Gtx6w0/tj+S6fOYoObPpSxalFa
DiPoJzq+ZyaN/piqDnq2zKC4kdoFC7jcfUkdDrN/ixWezHXDoN0+bGODdhy8n/M0UNyRzC+njuTy
edaSIFmNwpTMKoFhJzEg6wHcKKU7hgPYX2G5k3ajiiaUphYKdLqwsSi06sBBLQ4bgnnfDg0UGq2D
WImAPyxgxQ/pef9XRvyYg5T4EXCGPPOYXolnJTgXm74bTfn72W8H9WLFKmbmOfd/AIQfFpzjhrJR
Ffwu1OVbX+vyYfBRPvX5UdV47ScKmf3NVoAU4skK8k9H+0osM/iGkPZjpuDh/yCQ1TPGGCRX8h8B
yVOV9ec5v15dQHq25abbC387kXt4oPXvNE4r/y6nzku3DRhUW38xRTFKdB9y/pH4FeCHwXzScboz
nk35o4D9FWEiVvvm3utTOzBNBUoEreiOZP+xVeYYlUNbwy/vl7KadlPTVLQIaS7WwXX9uiCoMsCT
RBOmCTkMqg375lqAXrW5OMTyg869bsihwMwrFvdYqtYKsMhmjezDN5jJfcYa0SZOez65YYolgaz7
unSmk3a0ptffOODhScC/Xl4BMZ63iJXXIxL29C4QnXz21kLVOzJtmQ+gOGHnSW7iclQ/RD6tj86w
8B8Pnkeb9+PDcOhlRHdWWFqXx/IihdCxg6tyPj0UvrSiYAYkousA7LC9cbhWgHadCRV6R/TOS4h0
1McIF5zKD7V7uYHcG2VP2O4PEO9AoQ2wWusuikckjtTJSjJSUKgalZlIqYzu7o+V4b+HwX7btRe/
JyfwjvvFQ+WQSbEaV3jSFfD7CnGJy/ZRB/pR61KZDBpORoG82Im4oS6tXn/zrSM6Axe/uuFA53K0
5j4I5Z78Gb9fGj6hKS9Ds/HPKM8plPk/V5/zO9VHP05+PtuNvjO69BOeTvmPqJpeb8r0v4pn0icr
gMGxFtujgz2+3XIpyiU/BWlpCwi7uXdzbyYr0uztrLOCfuhQfZiIn7kYztLhk3cBmkU1PwKGAaKD
cGY84lwu8thRtLV33qyOqimzEqrokm31+bOqv6vDHBLPzevwm//bdI8TBm0U6yTQ3/3dwSwhtvmb
DfeGJEagUIxI0GdB7gdigeAAXANDtBvXAd6KIFhFRsCpTVGx0risz02a33V38m2TZjXFRG121JPF
ppC9kl+lqkJak1Tc2LHLIZCANNkwo1sNCcQ+y/ZHbWC4dIsEEJFXs+5t+Wi1IKFfMWLl38/Q6HZV
BuRCGmjL78LOd8lWvvtZlERRh7MypxgAcl44E6aI6QBBVhr1dfuUe+pk3tE7yBJyPZDkhk6IKSEJ
DHw2Gw2rftTsVb2oD+7f3Xael8MmA2rVem6a/Hr1RWOAr+zlJ0EXyirpFwgVytT84F6EVOp7gEBN
gCMkk6jBM+Xi8bGy+wOcn2nhh1maLTe8xPmvyVuaR/Lc45lyLCLVliHRxAaFa9tlrg3Dhui23mu8
f+cAzxmsbUnEr8qOm01gsD+FAw/h1r9HNW+ixW/CDm7LKkf8Jr5tUgr4iWKwy8g24OVivDSucWsy
4uYYNxn8NaXUPYuQexlFF9DJE8ciQFeIXfOo+q9Hie0pcI+4oxBT4JH7ceaE7Z1L2UNLydfSiMEr
VOzK4MmSavMomURTBtXSsLgAjaKtwvvU/bt4QnO0Brq1FQRyxaMn60sFPMzUAhULlDfzfL0K3EYx
zxYxxPzbyS64LIJ2JuC1n6HogjcnHNsUaC1ol3YMF1Hvfx6kT4cEFCVSicSWVWang54xHV3M3N1B
YdmjpafwKedoNm7LvUsk6K2J6rJ8s/FrG0Xp06LO+P97u8nauPN3/2/hCmMkJD3bJL/LOTGfUwnx
ADEqC6osIkSx+gMZln3Ilwz5s/4/837T8ZCCZSq7vYPZchf8aAUqYaorwAc+4NUggI1W+TyCNywq
NEl3yuPmWaJSjBY8jd83I/DCTesrgswBcYBQKISPHg9UM49fqmEfDR9HATB/89vTZMLiU6XXAPjz
62B4cLqWomqti6XHDwjRWxQefTbmLueTclNMuuol0cQerXmwwsPcywyK5Ub/zkUHLtHrJPQiIjAA
CKDw1GpngHGKE6yISBCEErhWFwfopFx2+7R7UZcgHhKhd1YQZI6u95UzQnPYtMDcg6zdA0GPcEG3
TXSSrSBJESXyJ1lR3lI6Z6Ydk+Ollcku9hsK6+d+QMZnIZ0KlprUrdbrn4G+X2+I6LtHT1exKY7G
9scOPaR1svTyiZ30ChXi3f+zTb7vqzkRHEb2Vrk+TEV4lR/2t/8BswV06a5p8dvoO028+xH+vmlu
DFKreBPV05nHU5V3VdcUJVbq9nT/mc6e2M88mZnhe1RSW581WoNqyyloKSRnqZVR1Yk5HCna9vn0
DHPknhVJq8tV5RQk1exmbPKbWVPewU1T7AEtVl+WBwu3xvCEY5GEVQxBdEPUKgBl2kuQSo8ZoHs9
Utg7INf95TMNcTOx6VEkG1kMmIAzw4s5PabypTu829TBPueMSg3U5ODCQT1DX55AfCYg24oKGblt
lSs0og3aPeMwwdGHUufXhD3XW/9svlsuOL783cvLa8dQxGb1Bg03qsqbKRstUzI8OBn/BS7vz9gQ
W7YS6KQBQiHu4e+MP/9YLLlLolp3WCjTC++kb0c+V2LHnhKhYars/+ZnuVc0d/0fyT4RCYsUoQZA
4q0kqmNIzOQq+YDFLKahBE+2uAu4eBtYoXYc19cicovzUyZIK8adUMUUfuq31m55rWd5KxN44nm8
zWtb2PuqGuPhjdNrniuxDjz8JVynfXwBh3aM3cSHpmeJCnGxukKiQE0cDzC2iLEjr9v24WPu027G
Uc/5zLBWX0JbyW7B/eFeECnJucS1rUDPei9Drqz0gY2UJBvrhm0Va/L1nY1+VA2YJVr2YlmUbdqA
3Spric55ixgrcjKUg6zx3CAfhaZ+6qzV7DaRA+9jJ7KbcDQBxYjlRh/5yB3QnGrtrpkKmRoEQU7O
DX+yNY4yuhsXY0jJsl/hSZ/XPuzOO79r19LJxN15wFwQj0ikx+t7uqNu3ItZ0uQvBVehvzBiV0GG
JzWo03gQL56rfjH3RIsWvbyQBLdpbZbQPTKdRlz6zO3SeKYaB/YG2NaMciZ7R/Qqew+lMizNJAJx
v9blSUULZFyF+N1ZbbyUVqhhsCe1Y190ekpgxAyidI7dL0WL5V5fDvfrNORI1njFkJ5lbgHV1MF1
VJbvXBYG/JHMvgt+yLHSAqU+nO0WAZobMEYAAy3nRSUnU2HBr6pwjxCqR8oKbisiMtEj62S6l/jz
L+dA8k4vsmQN9n3Asc/entLykxZl/HWkTjysHewI+KQr6jFg384AFlwg2j6lTs4C4td2LghqP2jy
wn+rKpo5g13ycFdfDqs17DB9rC4AHElegbqNLuleilVTFSPeRPvDjnJCC6ly+5ZVe8VZ2i4bDR30
WcOKqMPknXBrR6GExN0Kv2pb76y4Sx9siAeBXt6wxIkBVgc26m0Io2pZIiEMnQMEmrsyNVI7vE+M
7MdcK4T1xen8azQJ5QR/d3RjXqvbNKI/hxT/TwoEiGVw8ezwip92gXFg08iOubjeJZklDUo9bKaM
edF4Vo8eKHn+jeMFaEmQmxb8AxK/yfvwfZVcDm8g76IdSDPpUTjMJ5SxNprZVKkqB5ak6zdEU6O6
S+dN8fi8q+3rpHrV7nA2s9ETRBWVMXaFRy6fioXSvrCiRvandCeZP+Eh5QOM1EpXceJz2i4rNEUz
dx5xPcAomMMsyiS8iZp6V03tGnDSth5aVti8xoxGJOISjadggP/hvMHnUUfu+2Givr42N4CNJtQ3
EaoCKQnCNx/DkGAC8ew9B2YkE+I9BWMcdBnQ72lgTvA51VVvjJJTGmU+/Q088mmL0ulbwVhFfY1w
muiw84WG2C0Qcci0T1mVZexD/94h+gK4yIxGp11LTFl+rVMLlVEtX1WDj3euxGG4JXhWqWf4UYIC
0cLeSCGTk9Fiisvemz1hZwhEOcNMfmDpoEvzIfjPPeMCSdT94+IS9r+4fhcu1VUWeptSfSHh9Ou0
QS2nin44ShuEfLEfwS3BQmN6DdvFh1gjrisnT5dwDPzE4vSbzsZcKSDryKZbniM+Wy8coRSm/S4K
MoSIUkI04qsPXmOLwKp1b/GU5RmxMWoOWIpxhKu1EdNpXA4s6xbeuhY1GbQLfMCAr/VDIPYBjaWP
tKfq46DuSsgn2DJ/w7ScHh8EAR7B94QltjO3Fxg/pQv7tBaS/gbrfPjjwT76BFs2Xs5IAD3dShuO
za13+jhld/bRoOdUQbCBkd2+Y+0zzP1hLajkMZZPylwLATkoKYpqE8UCcdsAzc3pkC0/wLqke43d
nKSI4DOpb2zOOFJFjg1fpzQYt5OKdBFQ19dwTelFMEl+71OPtqXBZtkNuuS8A/4bSslmFPNhUxpE
XYwZ9Pr570crhsG81atdmfUI51ws8F6lo3Js0Itm+49iBk/eB3Yy/likc2XxNe74XbOkFBmE2tGG
YCjr22WzkkccwiJJRGJZ6qJU9+k95PjRrxz1qsN3L8cdtgadIJexQ8m+cjzt8qY6aMrpmgwGdx3v
0/znNYjfkEhOWoJPjsA8Lb6+3dSzAyo6SuaKevccEdLpgMJpydirP5puVtDadmMhuGvkR9Zdn7Ht
8vxi0QuvzxxW/XYqklcvoAvxF1IfJRSysntom2cUCzLzi96Vlbam1K5tP7fLaF5fRP3g0bCBwpZZ
NuJOkCy7EeGQLiDmHXrn2MtsroK3GSnvWZo7H2QMnnWXWc4QFC0AySK9fGhULhzYE5QFaZp0OfN3
iEBff+WgH9phSQDt4DYk55cq/iNWrlQ4eo2t6MVzM/ytpdPkWjhYzHkrXHjdMrSDGgvsMt41HEB/
cPwVQQD5y8ohUeKeS5T58BZ1ajuXrQ7rMJLTW3uL4PeA6lKC7Hw3ckukQkhA86BQtZJHUYVjDqmR
0zrNNCBQzhw20P96IZkKPufk/nNd8/bHcpkGd7Mg4gsmJ6wCDfw+kQeMKjVFoumZgNGe6Iz5hOl2
HTtgwXD2NuSwefce8v1EaE8SxKfSyLnA0RSdGO7EflvrKSRRziGSjlaWgGa/+cEpsohopnI2aK6v
LjVW+RhJpoUHDxcbORVv6Mfa6Hi3iAfrJrCcscCbTi8yuQZ1lYY7z7RdC5eL3qhzJ93PmH48LvaX
d51GbJgv3tBBxW5oglBJUrscI/zqiZatqU088yUkNaU9qe4nY8idl+BCjgnct3/+LJXnjzF0A+RW
B6pcR43g4f1dHW2lyESBvkiF39bsC3ZGVaHgn6B/uFbwKFdOwzlHOphZT+xbgDFJl7XIYq72Xoaz
6ofGBf21C7CfGjg2eUXvgpHAeZgrzf0/DtQfYU1iHP8f+fxiwV0h/ActtaGpz5xWKH2+qjwaB1UM
Y4FbF2RpUvLLpHxYXMzLJiocBKC3jpIcqYBDeoPGIwdUxAoowDqNtaJ9hu2JTQ0JhVGBmrzdERg7
UYjMnzWUL5x6LELUJWl3+Fp6vduk+tnhNmcMAFxS1Wj8tD+2hgxLH/qmg9SYPv1OWzQxEf5Oh5o5
M9BVoy+5bitdpoRd+6vZcIZhtjBn+Q6iQ2IoNMOKrVRxZUb03IOFPtzTmDvwF7PrpoSknRkxjS3c
yFZ6ixCdxalbpemh4he3Z6NOsQrirTGxE+Ik7C0471ILvZYBDre9s29/tLmQnwZtPsOYl+s6GPdW
r5FWvEMeHE+QR+OzFZ9QA3b6UAc0BoSHqCA72EdtnxlVh+NHhG/IXa6Vlnc53ZPU+iljlJ0KISf4
vXn1hzNg8+UtfoHKP/yBMmLBfbU09zdsfbSGpKuIS5BBCyFq7L6qsOYUnVLojU1zKHmi7sAwuBi2
0Pd2m8Zp2UUAAafQsteFcD7TKQrIW0c/o2JeFy+yGH74PHRrEc6qlKnKN2W+9zXLmr+2oba/jGOf
oLd56ImrrO5vOqlGBVEgYuJBTXCHiqCLUYhmoz0VGmgAAlWeuypomaeuHPfFc6jvODeDeW0PLGys
oJC54F42/eTdjT1hhDqxXLc06+/LAl1Ma1gRkNZCQHUnOjDXvRVB42kGdhxse7Q2//K+Gsn9e4YD
FONaD3/Q8YPP3ToYs16L5BjJL9TuEJYWS3x/QaqMeJgzLX2gLQY9Tw4RfqCXmd/kfPuO2a9oPFCz
RStMtX17RvN1BcYNjXledNary1T7D/G/8dyngxMOGx9JaQn8jcfCm3RDeppT8VU9W68boM5+PMn4
avkfwTblnhX67XHf+pk83iZPv2fSL13XKO6G3JZwG0Vcesgtk/J0ejLr3b6YxSJVZHVhxytUlQAk
tR77LVl4VKvfwvzgY+4giJTb0iiXZ539sj/zN1Ipw0pYvmQsdxgUcU1FBGJ618WckRiSvwaJ32q6
haDoZnGeH1ntjpmS/KZLSYzlaxz+24bpEbII6mL8Z4pqueDSkGfrqX5MjuTy12e/kg+ZafqKp0GP
ZwmIzxBwQsmNSyQAxtPi6KNNNRbaIbgFcL0Szmgjdi+E+I83OOGFBECKZzZMZmjtxdLhV2cn1VWe
bLG7rlGeEEcSyu2HviUYgRwdWuj66luYRzgyQ3105xB0RwZbXOymUhtf7GljX1JCIrYKw21+++sD
oSJlv2siYVFjGYAo7DJ4K00FeYhYRqZFKv7KZjnNdvyXEPe6AP6p7/cK9KsTXWQljBu/aRXnUe3o
0xbu6mhKuJ/dC9DfBm9PTUfeukGyA+O2Iqlb8AE8tJMX97uxXXfem1jW9NYQePTT1ixVvy1l3UNk
3vfoDJTFUn3ZB3hloKlVlCBbnYJT9eCd71fPpViESyx0VKzHSHZwrMTNP02fHWq+iyb5m7ivRpZW
hUKuWYzdIou0u8AERXkkZtlucrBB9mnLSglKSREWcAYf7nwwuUEbWz47apbZs/Q+JChxkd0ibcxY
9rj6VZ8AmTtuxU9h0bl8q9AQKB4HOIY+VWMxVPd6tRt6pv2+xerHjOryzCLxGr87yCDROrHLMK79
JVH6EMFOvwDCBXQVbQG31y/67HxRuwlAldhT57ooXEZj0ltdOvqd3JbbR+NLuU5gPSxhrEDikaql
rbIfuLW/dOZ7rCw2eb/0GKNPLuF+bh9OsZ6qT4wxigvBA8W2173yBiNvG/kgh9Y0Lqkq5Jg/QLJi
keSiA82xd/nP8GYDT8rOo8ywJfbFt1P8B0zYhxcZnxEv//WY0zhkGimUMmBUYDTKIRaTU2OMtYI4
CyE1ojpKKkN+6cXRS4Nt69DVrzj56NgOxUKPCshLm2r93KnuzWbjd4a+XGllRMijSPQ/FTuE3Cti
0r0h0fC/LutcH1zC6id/eHU1NCj4TLK2yT7oUR5ff5KuZlA2py/Siy0wdLrxV5OfBcIwVFDMuX1l
i6xx3QV+4XeBGGSl9rrhcSyjVKtCiNUFbWQhIdetnIPW3xBm5nzYwumcbFcV3E+MR6wmoH8ulTjQ
gLLX9IPQJpvkVoDfVQIg+oE/7eWaRtcGtIms5smrU9puiqX4U+6FTqIVZCfgXPSxPwmIt0P1djyI
dkqFbtYl2f4In4jTU3Mkvoo0oU3nAbeOJ91SiZKsx+NOOr1EhpEevreZ5ZHO7VPT9ffqvvN0ZI1S
UkK7OgWBRwo5L32gf/BAzPx2UsuNuejCj+Y0axB07SZ8MxsVLQWlFf4VpRAN6fd/0DyYbCjhPrQ0
QDaMicm6CXkgo1+I+FM16JxLjtUhrSBCfF1gsuDcAhK4DphelIq0OKUhL+0hnh+zRYwoPsJBUfke
ecVNpu4evYcxjfAC9mTnfeutXy2cpcFNIGEhxw/6eifJVzRXnMh5up0YWbOPUXmRrZ08DDOEhLFv
x/Svat7g1QBvlJxcZtqPosxhRKb01hlhKlAujev2DgckbUJgETtD5X3BlKsl1Y7CjfB9bXGYnTXZ
5vi+NCwKmwdnk+gaJTevuNdyY32xJFIsPeaJawI3toVON979M576IGqKVPgEKT5eSrFe5Paz0j9x
8kmW5wYmZqSpEjPJ5y7rM3g2p2GgGrPH/ACFebhcl+6hnI2o2+mRit7QY31uksV5xaBbUG393o40
8s4jgcK+im1lPPs28H5U93iupTndW4F1jtGFueq2kRZ97QtmWNlf4eFJwUxtFksb2GwkTI44Wh4+
6vdLhN4c9vi0eY2nJ274DK35G2nVhV82cTqZvfOg9P6yHLjYk5a/zNln86c5j58t7xgq8lIK7SCy
tKpAy1bCw2qaZOej1nzJNJCFoLcdqokOHZ6Xs6/6d5cxTZMQBXbMTTNV7u+5rzbleIx8g3nDoPT2
Xh5RCSpiNTEzteIQhhQjZ6Q3BHt8CO2aEeSP2mDIVDNwaqrZafkiS7oPPEg0imlnbcLGjH2xFzwP
71K1qt2o1ceWpGgAyxRmMsINIDkdN74bsrTz1fqGo+OJGaIML/vH5FfNrS45FrVkE02mz/ZTEpf4
hyRkDm4kjYkoJJ4vqnWWZvLMM3pleVkt+Kl0Lb6KCQUAvPoe947tUi139C9WvNZTmKihwn+VvlHh
2qQ2KIqZZrAeWjcsaRF5UEQMFwzBdaGJmNEiTDAE+qFE6k8BIyM2OhQzKHe2mKgBdneWX4N5o6Rm
pJsa0+kEV0CYlDVd7Sdfw1x7HGQd23bCC2DWd0qktmmfOU9ol2qDYMsm8CvQSmtUjV86PX5/MKIw
FT0orNEnptYPww6DiojzoJzNnn7fvyZSJB9CIVhrUpcSqiFHizQXSXrREP/utFW4xPOhUT1+/iMX
DK2tMxeLamh/G/XzY4KvzBMc0i3YlvW1ZGcpLb5RD8mnUXdPRPfaeSjwLG3OTozsAyy8fmptsmgx
sPxVSonCf00fuAp1daXfMmIQY9Xh3tjw0ddkolHWteJZqfRSX/Q8EbWbZw9TNCW7HidjkOeD1Nad
hs/jowoyllYg/F5Q65CL6WZDrRunieAtFJKwGuFAi1yL4GsKeXxDQ8m5lZVX1CWLpCQA2jvqHnyH
QN0yUcWGVEDEE4rRmu5EfN+c/iJZATUu7FUdBKOPeP9eL8jVJ/wKFyxnsAziLDl28y50+LPZDqFf
aQAK8t0noaSSG69DEb+8P7eKmSG3ejIgbOg4B22nkmEgzBykfnF1qn98MvTkVeL0q9JAIife3JTJ
Eigte89Vpe/8WJgi5/JFdkX6au04M4ynd5Op27KB+mxCZAu5yY+wZC+5ti/drXf95IEqHBjaSQN0
XXEuLcyOhP4bBkgkWljcML6Q2C8vVsGFudn4HlOReUzl5MBqRKkdIf9TvbfvgLaoshI6SY0KHf05
n4R7CsTYQNLPJu4MyO9T6iREeXAsN23GfxrUvOvf/Qm+KKpIKes6lynl0BKN1mFBoT07H6JsE3M8
7kDezqtmLBsvRJy+s2xSV87sB+DAFaqMvspqI0++OQ+1oF0Kp2AYL/ymv+aWeuuaLlmXzI8oQ9qK
+O04P3aEesne4hrAq/XumFyP/zEo8Oo0uoncA4I131Eat1FPtlyZ7avmPPkrft65Mn5w0amOhJSH
MzTd/XBrMaE+P2IorWCmYdQtl3DeYsnTI1q12EFcXF3HWC5jDG0pPdM6bdQpMzNxIxwGEWLVj24l
eZvtuUNHX5z5wPUDL1UAAIiX2dRCGPVX2MOm1eA41nJTz3VkG5TKXxR+FIFRtm57dH9v7m8js2cp
XuhyKQj9/ctJMmlFEb37SQ6oY2W63dH9nUi9UpYu9tVwn5UagMA6fh51wMuVBMHthq+YXJ0R1Y2w
kUQoP/A7V6df69pz9ja4A1VQTrp35MHUtQahIogCm7jf0J0AE0U6ck9PW85C3bud+0c3qTyWVdIz
CsolTAzS68NE6RIgL1vnJ507blTgyTgOo31orJWmTidZd67GWuGT6ALJNmwXTXrv7ox/9uZQk0tS
6CZH9hfN1B1iHZ6J+wwea6Sw0y+4ZCm3J5mTw+DL37V9SN8HRlSxWI9zfycGr+BWbd+Pz+50VGJl
GthOVlITDUrcKGyPMi7YaK6PmrJHn4q3KSz9imUMnOJ8UFxHLcvtZN+qtASuWndRbVu8R5TYo/nO
9DXr+45pwZLAEDbGigxSIBPxWWxR3pJUuV6wc3TzFreqDz166pIpsE4qko/jZj3+tevTak9Tgl0Y
Ft+KKO8e8Gw5CtHac886M7sZhS8PbRfk8aZUs1YPcu8plvCW5bhx/8GONZf3/zvkdWDljN8ald/O
+qn+ErQulwovIXtHJGOCEYVDbjOcq+TzQ/NLWiIaJ/GtU1yo0OoSM8I1MxTl/Tk+GapSLsptcyK8
vZ5/WQ6CJfZpGO+4EJeuozNCIF5bMotKVbVWgI8r+cELNA9E6lLGTPm8/Y+34QPhNVR5taURWaql
+P9J9hxacg5qi/3lEqV5BOB39COhkogNfXY/LDCt3simSc0JsfX8/oBJqytcLyI+/xSMAE6TelgG
dF/huaYXjdyCYL5F5zVI3d7hOZDNlQWYVAZu+Lv6CYOqTZ5lghS63ZgBEljnf6Pylthyaw4+LSJy
53gEh2+t4tHPWhlsfHT5D8ZuCmfRPVgxB8iMw1dRN+Kq78x4OyXcbXTUZnW3kO/9g8We2uy0CNYa
4BxNUih0y1OfWTb1JMWucLJbksmU1xVbJ7d4jVOIHVYv8m1Ky6oW/zkUECm4Lo9On0E8qTuylYDI
1cMatF88OBcDrp9iqn/K4yjEAiJKngVebp+lpk8qBmcovEe0V0cV3zXLY0V0zlVu7XTcwaqkTmg5
1HNP6FCKHl3Mm0v2eTQPZOYZGhq3mmCHUJpcBh8/Qn+NitDs4Hv+kvoT5D8YLYZwz3ms+recZiOz
lGRgCh/tavFi6Z7CXthTti8jXAvgxP9x+OqNcTqiR/SBCkjq1rHe311mf1ukXAGSjdNvAuARMSko
CBu7JAKrGW4zltAugcl5EXGr6ap1tbMpbSI5t04+QI9AJG8Vt6pERBrYWw+lD5Kr08HCe3G55M7+
S9ClmRy9nyDlxjdwePvu9X8YeW52/gvBGoId7UTG8RRO/g7aJi4vEnLbJ1+Jun1ey6CpQvAgHwji
4i3+rWrVDCdseyGs3j9cVyVIoX+exjMYso/mDIHnjiZHntI01OvjHxB9nRcLB4nUSnXwcWMGo28s
XswFtDgFoUmtjKERD4upLUxDZzAgFdnKgsiP4GJhnOIt6551UYtRPWFIQsevEKaxzlRHvRoWPoJN
pw6D7Hfcf0b0mp2Kf33vAfr0pgL1zJ7FaKgnLOxCa8Wsnt5xmbnNbH4DHcZzK/4pf6+ggJPDtKKb
vpfwrvJKhCZFmAMGb8/sYwHDUbke88B94oQmqEqnR+k8LKfcEL3mIBrHmvsLac6O8RhArn6u+RM6
CSdTV/u8Y7bEorvWplAeVXeqr04uwiwJ5of2/sIWYAvX/NnHoKDuMex8I6NEuB+4vNNAhRFONE0s
i9NtvcfCYd2d3/I86GYPawTRpz+t9oET6zadtwEutrY+BythqDNGQ0QL6yax3ihQocvAU9/rLrvl
C9sN5CmZUb2gVOk8EW0/Vk6PvbseDy3YZb74NPuJKdItP+nQrfBbljqunUFK+nIwaeu+Rf2NGmVk
cgrPjiESYb9ZgiCYYOS7zVSGNu3D1ry6fsyC4Wp1BvJnfoxyFscwI3rJLkoT3EJ9eKetrv/qDiOs
3qCIcTzPUHZ4vZYecaC+agu6oi7mJbkKPNlN0N0G0Iy/UnHvnFpKO14paqEuWZfDdEaRr2831i4H
h3YrSCBlZ9gH47pg5ZQk+SsDGswNSEoF1kqgb+RKXlnEhSLX4IoTIxfq3dMS4SF7i74LCsUa1Frs
pjKAJ21ThQ2o3QwAGL935I9HFEmNwtvGIOn6LHm3p6oI9+ZwBWSzVui8UtayJqT+I8brMuYMJoAE
F09QvJjWl8yOQbpChPS5PZ/lojDTen3kroERLdiemjK+FrwSliKXtaEKB9v3wS2RNrTGTL8q6o6O
V5Ai2evQ4+zDJeCrGj1BGlVlhfzacavFLvmJ6XFxQRoW9HxlQC25hE+ktSdPYKbHs74oXI2nL4H+
4MUwhLtc+A2yr17uyGgl1pGpEPNKYXz+dBOI96uWCWbzT8xYJndALC1wfP2sVaevAwp7/HSfhA4K
9mBhh0BQTlOrIGVe1GSPr1hdINOG4jIk350lx9OeDSuljkZn2nRkZUIck+aPH3dZXnIh1W091sOe
7BMqihzByNuHufCPQ3t2dGUnIzZPL50c77B2zopT27GJ1V91rcLRpNC5QdcTMOdGnQGnC4GJWI9X
uVG/Y+bSZ64Vbi8gWT2v3M49z3QDDhx3vEHC+DVXVCaW0/k7kcgFbhI0RRpLimAJ/bpNwdSeG5R5
gopzurpOzffxVoTRObyWO3nrtViMnybb4wMfaMCUqTClk0KKEURc1dGnIZ4bI2ftzOhJ+5p7+Dn3
k28HNmBkMeRY5Kb8Ty+MfRO/jbFUMm/46Z/imDAn1yPbxcEFMEsLTsbavD0tIZ5NxEqgx/9r3Oa3
Jumv1uiDkZnwDPIZu8cwpbGG8XImvrjp0edPTKt8YeruanOBcIClPkysPxx9aMb4byVdc4ukT3ZF
oXkIt9rrSCyilaVA4FnxaEERfJxJ2cfQK6U0ygfHo8Ts0vryy6/QefRDvn9evemFsgN3iwxwRyiT
VZdiQUC/Sau86cKft8maUBGbwDrOrxdBMkkOMfrBJNVmysbtX+Op2gH5aMht9G0BOK48dE93M9Aj
6pLGhdqvx8AlipuRu8Gsr9BB3slgvcF3enHfwmzTwSa8ZFyFTTxyHyB/6GH8lHu8/Z7cgIziYYIJ
tlTgFKO35PXj/cwdH6tB64FC4DUch563leaHtBu79ptyR+hOSjaCPomtNrrgbHio8iuO2RihEyZj
c+y+mxn8Df9sL6noBzqIbwcOstqJNW9Au4PIjBYUAmL3bVmCwQ4VFFTVA2Dll1nLrOcXH7YNjeHv
IiwB9I4+cIqeWL3Ig96XZXFAa3HCTs8xRAQ/g+bo50+ld91a9H4+8TIldM3mDNKcUvkDFTu0yEXA
URez1Vz4QpdbxrOKmQgRrwprIXReZLynixRxbJB3hgWKid49vXTUqyZKDoMJ+DAaVvoXfA8cIzR5
ICqWKvIWVnrb/f5wMxE/K3TmfEEFqS7086eAlQUKcP/0h2yLmdcNAtNXmqoiDb4Kf6e8rWBkfxQT
vh1PHJLZwHlzyu3CuBDUch0u28kS5kBj4V3YAESF2/YQnJBif539f/vpwktZJkUeQHk+TYtbcOlk
M0mKyBAafSsCroxr+aH0cPNhhSxs5PpxdpwP91KdWv603KKNKiaMit6IPiF2waXFuRq3Se148qPh
mI4dEkQWOfxI23zqmVYDOttrW71OZ2ZPzxc5OYKjtL519kCNs+rFpt8lYxBrAJzBsRcmTOBBmvIe
1FR1WHfiZRNYf0DLfslI85obTlqrWiYM6TyfkeSh4+rZGoW4eJDbIkdF8UES68t8OkcynoilccTg
ilSdpFA/3rm3iytnPr41MBdK3WYSmtchJcuyGvUxb2vt3UEbsFq8Ex//UTceH/fnjLFrVTJJpEG6
7zkMwYIEt6slmqWWtYX7Zra4I0A2BB1mOFECmRR1o9ZZSLtEcSNevtHTPgVOo/ca/LEmgKpKev1I
CW+LITPIk3E+Yerpg6MsLvig68g9HnIOUCn4FRf4IHXLHQw7tLZN2Tp4BQV+I294jDKABVD+qn88
ial9xZ0nz6P2lZ0fT5KXFdxlucAfR3+yy0/TYFo+edE3SDzWZbun2DPMquqelY2+5QCnojmIomSQ
aiWyWOS5M6tiBuvFALow+NqYyUfNJOrI99arYVWe5ACMNcyMiSRSoVduqN/5ySQi0NIjEDJCzUF4
xZhovMexEcM+CeCAbAS7gVOt2c/4X9vKz3POk1yt5sWeIZv6BxYGMESGBiGVsSnfLIUsGEeEEepN
GIsqtGMaiNwdhPDCCRj7GXLaISuSn+dahpnIS7XxkGFx+Li0g/IKQbolCDHgrUxzooDhteepFl9t
MLMPxRFE9mwxud46y345T0+fjeVPM5emaHa8qXDoUPdmoUlUSmnrFPz8qPi8V0z0dTvm100Hqq62
T77nJkyo018u0b8vP12O4jjtMOpH87CJdjLprum6VMbFKDyHsketEj7K+N7EOMRhBckeDR4uRFZl
aTuhBa49Itl5X8JhWe8tR940flFhCKfEqW3LTuqqXDiLFKJLSDYzUxF8PwhXmmcCgIiX7PqOOwWb
/9w7KehHtMi3rUCDuwBr+kBpl2tRDCxQCR6juQ73ExvX+wTYSHxUfRlSMeNNv4s0V9IRJa3X2qsD
ht4tvOHWxqZLyi9IeyEH/+oIMq1tLbg8K266Y3WXGum3sRfVEY/IcG8NlAa6alKU5kZguoYULwDc
23dqFTq61Kt4uOeRaIMu8tHDr7h93iqCcWOx5mYfG18WDqjIWNXwzMOPNp2cAY+sKXeFg4JyE6nq
yQaurCyHVoAeMe03GKhHllELPbOOnZ80mtGU6jfTndzZr80PCSz+RAilL5GeTugWzowlXAlvSonu
ht/AmL92w/FYhMAXXGHuq9Yp6Fvrt5b1w84bARRGaqWcOsUT4c0iIpZh/Y47UiWAE98B5R2tXkxv
QmTxE86a5LFgJlsgcPSn6HIzEIoW/YQaueJYXjmtR7rDRxcJgAJOrNKvWaqo8vrh1Q/rgFYMa+ub
6Mx5Vo8ICSqXA9s3GrkTPN9rGCd0B3pLgaUF5TvU3tPBjs7gDs0cuODVjTcIwVwOoBBl7Y1MGdLn
9WsXnGllKMSaR3SSZktxLScMUNNPUe48kTmFb2xKWthPYEB4c5zq2dtjrykOH5ntmm7kELWY2fLb
TYgIW+kPc9ghz6UwEcVKZ8SlRYL8fNp8kc//gNqRrg324beDRUmo6pEV3b8PD5XQJN0X0rx60+nb
t6fV+Q2xXo7DEi3Ns4olQjKpePiPHMSVPMCB/uV3ZLOEL/todyyBm0itha3BBQPOUQ4umoYDI4Ps
C9nniO201Yys68SfPYobFSN+xP12szLeWMgcvPBaztGBJiH5d7UQSd94xgYvdkhT8VxcfeQ0P8uJ
GwnyxFc2hhHSyb21JuaFVS4g0tR4tPrtHYKGjX+NrRhjn0je9onjg6+04OQ6mzuTqv1tnPus9ph+
gxhKpQ5gSE0x1IcQT5/jJeCLjR8Y0mtDkX0ONnqBx2An7AOBrvBdKzgeVJlI/Db4qktowjQa8Dpl
aVDyYRICUs89WxkTEPR2R6yo4uzdP2ALxOpuqzhGJbPuv/ylbkmlTdp/F1AmMKmaTZO6r7PhUM3L
F385Vr6f9rx4ofZ0T1nGhgH2zZ2pcXw5hAJ4x+B8xFXtZEvYSnK/I9nxffPOd0mTKkaWp7D9zP0I
FxujMlnAtgyfLJc8n+xR3HuPaWxdCU9VgtPMaVSn8nmRV5nfqSGBbyNzEYrefSpk0vBckDgJdTmQ
Q+R/5EZrTBcZsEGv+N5aWi+rXKLLuG9uYJRSASA21fDg0y15D1IquPFEYTi4lZ+CbJWjEcklRf4n
S4gq8zwD982lLgCX6ogK0fmBhMlGiW4REsJFPuG/S/wfrb8vRnfo/HPWn7VXxhuagz42PL9ydpse
xcIUci/h4QJ+b0fiz6esX/RgM9BUu0D4Eh849QqxhJk5jORKOB1vdVm8MDjuSBrF3dF9wpnk0ryv
Tc0KItEhOppT1hG8SmsWJ2tA1YGL//GE9baclW1wyAGEMFoNfmxaUxK4yLvuctne6m8MbOI6P1La
rlsR3YeN9gT7FPU9WHDDioQK6q61A2Ku/dpZN8KtFFStCfhIZEDd3OwfmUAk+egZjU9Dfqr45T0r
lwaordvKVndKnDs4IiEXMz0laDlMILY1Z4f0zARmvNyGCgyjvltAgjljXF5FMARHUcicmoVSk5kn
BJLrhdBRyiAA0kyjH3VuhC8EWfRLhfokYrptItmhtA9LLJkzbCJmYvWCuNmAlJIUqcFBSZswxmQL
rxSd4cxZavMxGvmU6CbFo/MIVp+Y7XqxmH3an0L6efWa/XkthxK9Mgg94atmMCTB2yVNZWL8rKjQ
wUeAbud2E9+iG9qbCNlk3TXNCNzVMfPwTiN67z2iFUSjjB5IfcwOQsJjBGLJZZNmh33XOy0k50Og
cU5OsVuVFWgpnLq4deR97oOkNHhGBQ1g2eOEzdCeRhT+hdJiYubpn5tkEVpM1tIkv45vUwSGfbQM
RSNw7XyMCFoPK4qPhvZLDTB3FVkgujJpwMs95AnsE0GEa+ozgd7/wRP+x357bXv0EIwR9A4F9ivD
scZGD4Vp6zms/C/kVzJyh2NsbVenZdxpi1nSiiGK0XXX3uUvGxnstbK1o2OUsPKFP/Py7dmjaNQt
tMkPo/FKEq1w9LgZgs05x+TN1ZiA+RbQjuX+G0ilrfvtaut9+SGMg3uFmEeiYR9eXhpawFAuaqBz
frBSGXTeBbOdCtRQbV4wr5kqUOz6WRAAD89Yrimn3lIFg+9nRNrxIGci0w3ex6glle+YDkvGbmMg
18QjDaEHTaBrj3zuuvMNtXIq1o5J9P1ia6yRbWrb82WNlGGk4FKugTzkQSVWgogJZKPGYj4294Ez
Z+JbFj+jeroUt0xkfsxGJeD8Bap8xWvUsU8XlCWEbtqz3X+kCKtf1jrlRcMhiIqBWLkEdP6ked7Z
wolZ2LjmLXMkszpCqrt1MQRqC3fiNvRaT7qLc2rDxRRo93o5tedylwLLZBRhcPKm4FI0Q6zLb/Y1
AmXG24/mxgCugTb2EKed6GszJbsiVPgMnZkOTEfUZ9orPKD0z2yJ1W9/FYRQ0jJqsS5ADjUorJtF
Pd0vJ/n8Sv7V6K9iHapf6NWEHfHjgbcHZYHZ3xrrScwqSJXCL1hDBlp/xlayNGXv3v0JK93Rhwq8
iHQmcYe4O16FNWg0/yVth8gdWD9XQHRLMJZ9ATktLPCj/Aur9H/2M9B+1YoeqAjqD98H3zWcrmwe
XLlNfqzGQX62f4gFVKcmK0tWbCAFBDZwO/0btEAnKhD5PbL5dwkdESz3TAeMDjsj2CEkKQDRsdZE
An07SgOFGcn89lb64qJ3EWb+wH+Y0KToFQ7d7emP0gpfLuXC37B+exPOg2pkQ+HRvrtVznQyZuet
nlwFt+h1eUPQwFcnjaCyFXMTtI/YcF2WFoDPj7c43/5/gd0xm7mJaso/xqslSQsJstcDxKNOQMhB
98Jv0EV1BdNmD1ymlXSJIrYr8ChBeATquYzXSO8qo6Bq12cuXmNZM74nqpMt4dwhb5w2fNtJybQu
A84GKJD0VgrL/NjKifU9Lfj03VqEC5dF8p/Avk3gQKTho7JTbYm6LLaeP6/DxJQRH/DCd5o/sn+2
b02kR0Ko3SV17mRwA+KiESwlnA4utKpBVvbw/bYEbNWSGLiPI1KgMEcIFQKMEZBV1v3u6EQHwSv3
x4gbop3+6JOuAp13MfTQJh4XQdqw8qlpu8FEiumQuEj7dTGRu5HHZNE8Z8IByGQxe9h9E7H9acv5
kwvMKhcl7TSu/jJ4c4vb0ZFeP4RPrQV94bclTvk117OguIZY15XxC9V4pRzIydcFxts92kx9fgRl
VYHOzCtkux+zQs10qHFbJ35+ekC9tEBpjm8gDYVv3b5CIOclt/xN5p1eAk0LGMPHLF42hSUrEfnM
W55NaIqI5r2Dz9VWxm4GQUFlveapMBMflAMhAAwctNV1OgxK90e+vzgPNNJdLHnll0JJRiyV+2Sh
LDYWXbIWwuvcXdm3rRL7T2tKVlwZf1C3LM0VaFsZ6PbLBRoYAsy3FeQf+BKfLPZthDcMGq8GOFgu
MaS/m4TxSzscOeiRUBgTXoyNv2ctAISCMSRRVvUMhYLnExGGsqBWOc7L+8pyNJJWIJdN8E2y1U1A
t3k/G8fOFas9P55FjOgMZ1B89+fMtQr0dFvDmhE8+Gw/mhvnT7RgRNPV6QP1D8MUO/miemYs+E5O
VjCFOD67LTCU2z3CiOX723mMB5BsAOK4bxX5kt0vR1PePRMwFXfKJQG/7j/KnVyyCVi9OpDdx5ja
vzAWreqcbHCLVC38EJHWE+FPW4gbsue5XvrHRAhTw5cYyJOn9cw7Pk2FpFpnxpXe9DS0IaSf3dZ3
qOMjRtQ1RjNA4ZQUWusS97bqwWYYE2Ga9wc4eh6Bcj/um3WsKIFP0FNQuCXF7l9UFDwEJk4vzFL/
ol+pvIpuxgie27yngC7oUg+aLlF0Q09RtXKiP+mrpgxV2F8tlHlEE7vU04lSVCNdKw==
`protect end_protected
