-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
h8rs06GZlRE80R2+DAeLuj21jcLx9tdNAzMAG8pIw10kgOHXkBD0TWB18XMbbzfVShfq1GELehnO
t0gOuhRUeVyqHyPNmxZPnkxtvKux+N4RC0T+z45AFRN4FD/YW1lEPW3zGfJMdH9fMNq4aTqZAAtJ
kqUptfMAOFLQvzM+D9qRGEc2y4zQ05xNwwu/2viEJajknTbpq+P7OpVkSGCB6RIaIApNEXzaRaBI
tnN3i3wj7gYPcVgJVmhL/3PaVa/Tdv2OWsjaVpC6DdpUjIiCKpWpvThDi2PIF6yUSxctG8C0Ga1C
9XG0bAXCydSh+Ijl8P9inLrKXSsxxmfLyjGPtw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
ZAI9v0npr4UGNYuEtBqS3njuEKjUqoRl3kNpbpP0KfrptZANGOZbwveTjZYM/CcQorZbYJu9ZfVs
GRvpopYQ3q5Lp3MPp22/JKCayLon5/rcbKhLx49hR0qR308H8WL5rp4/7Lc5uorNyRgSPvzHKy7x
2gNs6XzaZhFtFrnh9EIMgVIJvDpEABptpwtM0/t3RrkOJhKZuSKkp+9BKhfSyitqFSV8LPFe8Cn2
uev5sVq/kOxJr/StLDkfYNOwboGnRdjiteNHTAW798kdelOGGOMlq5Iw/wlZVk+7/B3OBN7Cz+5p
tf2Rf0gVwM5fm6WqnSABMhKjqOfUOlx6eGF9Z0qETrQAAz2mTZtzHLkreQ+n7KOvtfPGNUy3L0/U
JgdpFpsKyQBF9nrITKUPQi2Ksf8iJhGNBug1DPqFz4OjX515sUiIh/2ZVfQNnNfX5DJQXpwhZ0f2
yNhoCh/8H7hXNEsJ/1+7miIJpR7n5Vrt7C17L/iC/V0bElWhH32y4ZmXB7w/3sPsfLdULwZEbB4B
OLc+VMyt11eI/jcuX/fIn+i8R5OqcKubUOa0DyTYUvH9OCc7xeZyDip2W7Xxj8PQMCHiY3lheLn/
gg+MLtCbIL12B0BkteppccmXvPXXfVOMxmpwubBdOcYTTxTnljOFwuFnDVARlMVdZzcZa2/YSyW0
bDjEZaO5/Fw6aYZ4cjL1WhiLygHgZCO9Oxq8KMF5xGm+1nqGaXGNqAvi0eiVHRiQo621uHt01ufc
Vk2dpnD04KtP7dVgm7n+ufACRPRjrDJQRgug9P6Ppzd7G83QZYeR5CRWma2bvVchUXwmlT5R62Xt
F7/PtH/wE8NZPJ7nxU3LN3ez7h0kRSoLweGCLP+WzGn2zS0vWwP7HOABlUJQsuoZvCYIiyjqqu6e
3m1fEcc15BowQlfldjKqylHnxExtLBGWZnezqoacaLrLtAWdgY4ttOY4zM+hQ4+N0p7kHDT17bKG
931OHqjL36dvYAcrs0KGkwy+lK7xTnasP5tf0C/6108/+4Df7Cv0P6HQutHzZYmFKUSvg8GI4dsi
gDaYPEdsdstLXpEO7wyCr4Yr313IuFPRwatf543Rh30t3l8J/ynpeS11H9kEs4CNzbczt6S4k7qN
NapjKRcXmB/Yyn1avOz1sVxuBgHUnuxhBG29gotqVd9HkI21/7yfuzO+h3KqRF+7/9XRcZHvQlwv
9QvsC1OY2o/3sTfymxh4voxbR2yqw5oVDW7kzgquymBBMIVFTDsYsOy1Iz/rMqjasA6Y8k7y8xP7
7y2mC+teOHUWzktQlws+f0qiTV7hj1+lAScjL5ApWI0OyfE6f48xr5rLKTWpmjB5oWxxjw08sUEE
I/7gMmLgcD+65HNRg3ounkgXDCiNPxh2tV1mi3cjQuJ5eDotUf06nN9MUzDsuWyR5eruQWpMWv+z
NuSY2xj6V1kvXXxgC21MQa5YiOEYOdgnpQv0Qf6e22EOrRZ12C5QS74pu6I2QGvqSCQTHCDlcxva
ctJZohGZy4LxHi4Gwj/1qXq01K34ulEf6T75PQD/AzjV1ZyKWIrOCFQw5fU/JuD22W6O2s5ksSgj
Uwn39ZRhoNmMAyP4AqT9dJ6Ro+N3dLUVaqBb91l26swjdTcXgiZ82+5sDtuFDdn5OaNt7sxUW/vh
+5FqKoBZ4jRSgZfgdbtOdhSgVEmKYLRt1kZeXtn1FtDJFnBLd/Vf3EFE2O2rTXDwPFDEBkGDTBzO
N3HKFk6gsRdRPPKwXb4TlWR1+uJHvfyyPol1GO+0FORPLq3TZZCqBkpIjB4xpiS69HIPiCDdaHAn
p+oG7yELVTXF9qejWsEvH9lJHOrrcrYvVF6mw34NQ3SAycfTIiudkXIcCQgtnD+mtJSh1Ajswxqy
RX4YYou5hNoEa8Ul/uJ1HyB5et6Lz/lcikUFQPh0eNEAm8uzKBeLV7zuQGO/dUAsXLHOTN76hTaO
ADxO6Rsysm+LJ6ZagugHAfRJSg4WTJNGV7qVuJJJvna5kDOVv4hhkpKCo6MCIMwzUcJON0cSqf0t
5Ev1YFneKQckjzGL91+VPA15106p3f6vOuw+5wXcN5kE95yJh/GUGAK6H7J+4zKHzCCs4/ZP/VZV
XTAgZhU5tPHZ5IWrhKoIqQng9mYtYVfzrQ2EHbw5oX1s+nKoKizGH4qVgyin2zLwQtNx/WQz48le
c6KWu6GXtBMGBBgijH+YtMLy8IuNpqSZ0umiID06hnRHPdPheKgo5vtTFqx/1YGfIvLiUcso0oIU
KobKmC8Vu6QFTOdw0X0sTTnEmETqZt2pBWufum+GV4Dl3SX3RI/cCV/NGiFphb5+ceJE7h/ghoEq
ZLVw5FSYAdVf2ViWLr3bBhrrEv33HHZXOAiHj1zNapfLOINjm71lo3yFZGAg5yVc7/4fXfe5B20P
U5YZ/HqUUDXm88KDnE59zKamLnjS0Z4dcLKCVUh58g3ytETQkW+gv2c9q2/xr22+JDTOKWKVq8yW
MJsnXgN0TOAp0YR4OWut+BqEsAe4XWqaKXijaea6u3QzwcZ4WqcVv+LcD0rULRxnMoSq+8kxF6/z
pkm1UyfmYnFmOX3QLp9Nyp0PzqjuLTnIvhUSKtvB5taPSZ8ZjUVJbAQzmBEatE6VB3uJCZP7OjYe
KIepS8/3DYaR9tZzNsC+2yOXMCq5ZUP7O2XynJzN6Wua2Ixd+u4JFUpeVD1LU7IWZ0fudgHvdYVD
eAxepxDllgg8YZWa/65exZ4rmZ7uX+mz7G3omhk8Ti9FAL7BThcdt1fHXs/P03sh7plj7bFko1Xq
CFj1Npm3g8zDM/T5xq7lXu2XwzUZXf0u5PbgTd/2yXJ4rXtvaM9NLt7kDOvA+Y3laI+6jxDNW3Hx
tUU0KXi21IqLdOO20IHl/1haQenQhk5HxfuLo73k8uKgvw7WBj9mYugADIO2hvFX2GMn9vZCkiqg
o7m7pWcWC7kiMGLESR3Va7qlIv/NGbnUpy8rtUuOGQSSgg9V7wz1l7aBmvEsoXqPpi5N5cOOf2RS
rJTlbspv6ZVBaCE1FJpAJLkd79xn2WJFlRvfKL5kCTu7jgc51sOMg1S/JsI2Zm7BY5xc2JphZovT
eZDiLYdLYqvvCjTmdPgABmlIWBXkyadUfaWuBcihEFiDDxAimuIOVbBEgrlBnc7N4r8GxLjLtwnV
MJzZToIchljlZi5A9vSsyIwZuR/ceN1d+QSpcTaACpHl1g+5f/xxAlsJH1qP03FVRm8s9/wg3MUz
SN0DukxFsvcL6+joBMQKyWtetclYh7IZPggyIbCwkaLASijR/HXwimzRTLV/P25SXuzvogDr8K1V
ANigU0Ov9rlInqhVKknz1R9ABdVODnzQReXTntEayUTO6+5/kZmsb+atHrLzdiiRdNBMW+cQWoju
/vkRFurqhREJmrzzHq6/yFAA+GSvR9xDdz8ARDDPb9Qd2xQw9iwpurBMsIPjvoy4p3D9Z9R8L/Nv
B23q1wPAnZ2RQv2NlsaeurzK4FyPE/QWIIR+gumzCKoiEg1ZQc9juaXVrPDzy0ZAtHRZDojRu8Fl
uGZE/i+SPS/lbH4ET/KDxDdFDiIYLqvemwJiwsasRsk+ummeZfL279BpGemhUOjzJNzTD2y50nmt
yUVQ0PtN7ix9cP+YvRdWXvdNHx5bLUTAkU73G0OF6sBkMLOEiH9mCnGRmBngTboWaZPK0K3U8baV
I2guyrEu7eED9B/xjNdCrF8+q/XuaEFePN+f8i39eixIUsyXnexS9FokntLD1+V67FwUl0SRFkJH
r8zvRZtV5xQSosYeXaqEB3jPZCir5DX0ssc67T7SlfaxRNQsWzFwNlQcVR5JZGNNdeDLq3A9Fg+z
mWjq7g0LGtFtfo7mJrkZ2ZWaZXcjYk70iElcreNJ5LPjOWLLH+bIuku/UJX/sFuWi4UCLW++eXVv
AIlzVTQ4V9aWFIYKvRmxwGxMywrvTZStJhF2DYmp5Hu2PUjMB8nAgtpBNu/mkJX+RlPxmkVW78z6
g2+PRBmcLh4NgdMa5dKsKBZX0uXN9nGpgKpF7dIqxY8hsVZb2pCrbgJcvQd456Xq/5wc9MnNEuYr
IImsrnGGSClhkO1GdwZNrqVolYr8A+udB0qRZ8h5KANYCPcArRmj4HAb+ykTWT+fXrsKbgqPkkpy
HwG7JmhOENDKN42xz9Ga7WkMT6cKyy0QeUDjjZ9S9lNRVRTEDsokEsCFKyFOK3pZkrB+lwm468QA
kfQqU0ReXMdoYQn0Q0HArnDLzml5z5QXbZ5a5EpwDgT3e9RxBne9Z6dWFuJ5avTh65bftA6uTu/I
ipgUhtJ8nGLGkGFXjF7F9nLfBcsnjLIK4WoWhWorGXnLSlkspEoE802RuYG1wVA869bnBHyyfQ8P
mmFHKNCSYb7Z9ArFmIHmPgG+pmFLqIIJpB7V8+haAdMZp1THrkOSNPNL2bC2bHxKL1QKMqbs5O2d
vS76KCut7cwND3LJGkJ3ozDDyavon3t0yyFPLckHTyWJZLO9XZiwnA2qt8GtI8qUxzuCD6vVi7ap
IdioZC4lnz4H6NiBh65e5KP5wAjF5CLNUvtjJ6Z5Kf2trnS+/UkuGXXOVYUKrNlsaU7B1xBy2TZo
6Llg1AfOseEQ0mfecihMt6tH7GITF1hc3webSWTnXftr+3W7qYqPMKNPBpSfcHoI05oCqG6jR5li
H+Z0DbUXRtqcuUOGlaRhRTxwUJWXHO5ECzcEvFV2RuF9LKX3NbHRduIozg75EjtQynV86glpSNwd
USbWmJGJ4I9pZOawsb9ofo1FYHVV2cs7FLLVwGMm9yaMnXox/bpMvsshRlJzV3rcgs7VVcAMvNeX
YJx1n3h0/OKucCIOxnrzamKtqjWhoYG+4P3FGzs0BBkchq2v5Wzmxr5ZDoMWJUtgVAZQrgOkvwls
B0GwoF6Iap5skI7En4MKTIMlY92qnIjNKpZGut0Z8HA1/Pn0BaPWmAlEAw01nbRmRWnjejrWsu/E
CRBbx2cWhxfmjO4L5o7pKXxEviLejvpkAmZfhmE59qwXME5TFWGDukMBN/iAbQwg2DM6GmAReNVK
Sj9J7UjMyCNqpPixZUsNEzobVnow1N2stoI2RfWzrIqNuICusTsSn0fP83o/cjMdfCqjNJ0Vd3ie
XHwqkApS5f0LN6BQ2Z0LwNNhAm2mpAdvU+BOd2ior12AkA+SmaW2pMtc03SkoxMSnKZL5TPJLnyj
5e2GXoRTwkASPpmEsgv7UAnnCEwoOOZO4PscjLj6jKaVBvx2VqqEPS78qKa6jxutO/39iX7MgpYP
ylFNuhdHDLARhJ3O5moWBj0My8T4Dnvr5OS67WnWmE09pnOwu4At7vJGEQbGzkmXEQSpdBr2RPOy
XwCECNVyaRCCxkdFy4kb/nDwtov+LwuvdZnBkqOmtip63DY9v9Cxb1SlP7S99p3YIgGPw1ufPEtA
1mHvhhIXCljrSREF/6GkV8LowC3MFjQg1OZQJEic5Twr1Zp/Yg6r0GDHnT8qUq8aAYysKMzX2B5t
iiSCItU5Q5W+b3l/WVQYZROsqkMiKZuQHZkvfFODhA39Vx8eQntsRhIrDMckXSdFghwzQN3805Nh
J9yawYTNXoyxF9VhV8sKl40tBfgLGQOgDwLJp1kH9zs772Vot+8ncvAacRz4GGvfShrBHUupvvqp
XXpZBJjScXIx/0lj+hhdAXOl+HHeumlvV3bZOX6HeuW5y9yAMJiNJmKdkXpIGIwAcGKs6EtHPzYF
oBkdtF4/Si1IRpvVzZ5/MRRMQQuzJslNfDC7IPg5z2dQHkWBuoQZGrjGn2XbxUEg9U2EI004IhaT
Nh0VbBeoNo92huoyU/ZWiva+N1XxhUbpOQHoPUoV6uuGnOOokXDbgcqJ3289Sc83raelitX6ub1m
DeFW6HLj9qIou8osb1M1sQxCglvF0HNmi6cxRUE8hPJgpO2hyeq7mDmPWtGe3mR6jfPGoDW3Bhz3
7dvNmp/DifvfugC7RVOGUBvqkJtBHvBynyW0xWLNFsAX1fz/9uKVDTp9ulVkgGAaUhN87sjRrhig
y+McC2lu5u7l/GDGAPvZpey/cobBp/Ulz+y/nQIw3k/p8+ZA+hY6IJmVUho9ohGm6At/Cau3srTa
wmc/Wc5/ivjDmPa5V5s2LBMKBss7c2kGkLtoXfS6s/BDqO0iaELuncHX7yrhImCeC7u+PZj3gWQs
1cVhSTLPbcS6B/SjyuTV3jrEwWrU54OkpsmAtOGJ5Qcjpdtb9dLn3qYZdkKxB+dY8g4zcUxJ+aLi
gg54qJDQPFU7FanzRedtJ2FQIoHO1nplnBZ6JEKoirj28fIxSt2YrTwU+UcUXo9ZcnSv+zRxjFVj
gY2oKPNXUrIZaqpMIGs7mu29zDShykn4ZZpWh0NT3b2R4Ob9ci7dGvgkDoR9ILD6EUlWUO6hCWBQ
52kjfZrziOQKF+bS/AK8iYwF8EW5XpFMDtQrk+TLxu9V9G7LLpLai+Mrq1wTdWEM6sY3XGqBxzVi
TkfyqaHq4IopV9csC0BLu5/NRBNWeOIOIazvVyvNdU6qfc+kd7/0VtrPs8PqTwafVpVElDtgZyc2
H31nUaV+OOuXBEQbfPnE9jBzAFsX/jEDfNy4yEfGUpkMgLNT1vB9z8vZ0KIIExY/LP0Kiay+PvPb
12PF1HypgpVLakfrqIdB+ejOfiw7pB+cFRDNk+YMhrA8kLPQZEsW/J3TCKjBlt4HzkQoYxX4Z+rL
GTM0/HnNc8KW/JE2sUZ64XnVTaB8h3GnALCZGbWd+Wuf7ax6gUXcNM1XzJ6pVmwlPNwI71Mv6IOy
JVAvyiJMhtefrfy6ScN1IfEcUF4gVrl9z3YBI4xAYb2LYlNEnZSs0iraZ6OWHDFqyheQkkHf9opz
v8gLvSkXLTsWW8Vr2FN1jIPnR0BZQoQKLOawxzMh2szeoKluS29rwHRpN3aQopcJlRK4UIRkwHjU
1T8I525/qMsgZ/tsPyA5cUqx1EpKTT3M4vMXJLI5XSD3Na/dPzQktIu0tdjsz3o7sT/zL6hNxG8a
Q3oM28keBmkrfdJXQKnpdjGN2AVrDjgGzzppGLWG2Jhvuon4uZ8CUywcB9UEQzeWbawTtQJS7d4G
cLsfYl11GDbgsdeoQNLprlN9zIEou42bIJUeC5hBtljd12GienSKAuzvqHSF2DDyB/2r+Nt7Rt4B
4hdRvhOW8Qa70fEh0y5OctnwifNxmJ4/v3avbCfBlxEZe1Z7Kam3VBQnsvVQZ9kIVkt4Jw/QdrKY
ZOzXiCa5rr9k/3V+jfTX/jVj1nlENjZ/2Ns8UCToAJ9ni2D33f7mOfrvn4UcIk8Gv3yFFgWWjuho
LAhbBjBtHWEdZdNXAukhbkpSNNmcCJAf3U3GYbipet9Rn6/sDBRh60HiuVfBVc0Q2jCNBOrnprLq
gnxHiDTZZK24KpLfRCcSw5yy39bQhmxaeYtKdPVe+0dN7LuoLOdR73OI9RluuMEEtGoJFnMdjyQH
Sj4cqN0hygl8mIaCj8FM3ZFQKBp1FS8gFj0DgWcfIQUaAkfGD1Mxyuh7/siBcyDeOg+YUT4B7fCS
Nfuz0Cq4gNUHh1rkSVQrAixA6whwFOyM1R2ppGgWVQJPocV8fmMab/D0smde363X4dkupToYfuEW
rgQD0w0RW97vBWoDw3S1CD3mvJjaB/zjoRW7/m/tTpHu0iJGUbUM0D/FyBpjLGlfKEeEn8JzflWQ
gTW78d3W5t0UafU+fDDS6aYwRCsvX44FwWhiquRjcnZg+Vv/HjahsnqxH92W1TvTGbflh0cUjMEQ
RJgVpJODDhEWDUKBIE77JeZYC8MztJN9gEad+4aNRoRpRsWH4rCQ7zolTakrnP0GhEKtB9e3lL4e
anOC7IswclGKPQCpiXIDzhhDwWfOpMZPkSddpKaWstAh6sqeoODAjGfgsg3ra3mdz2KxQLZVDd7D
8DTUx4geEiXtP4L472Oew+fRYAAooZ635HX6Jo2RnbwzsR9SGhWrXHEzFVT/oFopVP2ldQw0lSd2
eem0a6z11GJbaBPxWvxFqX5QOq62e5ZpXIKlMTjdol55UxySlw9aP0qTHtf3qbTVIgh6qQRRbuc+
Ha2NJQwce2KJx3OwQaB64De+6aj8ROZMPg+oOdIgzjkg/BVhiuVHu6INWTokHMaG7tP3KHF3Oemd
yau1rrApuZguonnNWW79D/Fa01ArW/qBQ4QX8oPokO5CsputIthWec3CMTuo3AfC2dUuHGel1ZI4
dHnKF0j9e+3oB8OHF1JmQKOtrN86cmNjm+y4wu2RVvUBhRe2nis58hNA+psT/o6ScSgEdO70tki5
PjRQOTB3v7zY6iZv9FuNsDS0wXibtkD65RwMSqeLMJd8QzAaJvrpcR017BLQeeYS7KAxqYun6Pyk
rdpMxMTRs2Dsb+ow1LqFWxBxo/eIMKpThqDU8sdFHWg7fUgL2s93lo/foNvwhCdOj4dFTNQh1mpS
vcXwxSP+OTJ8TJs88Z7fdX1WmKUEiS+ivPreAY5fHq/vhJWtMHqwxDtwdBW3gNd52ohiGJ7/LmPK
zbQ3Y7uv+WNvkOLm+ioWlhyfqrYxSye8LImQWwAd2WJ7RLPGiDQi9+laJvfNksZl3H+OXTDbELZZ
GT/4wqMPGzNwGYx1IL3sPTk4Lws+TKUoQTBuqzG+PUDFdUsDXBzEW4COklB/QUDVxNladxDiGsJ3
F05Eq1OqQcwiddplHgUD3n0svw/gFRMO9URAVOrj6/KV682iwnMjCpHWqwoMcGyuP3ew/8d/eHk2
+R9yB8JMzjiupslabv7POfg5rEluTpr+NDyljlgwpY7DjCdCuHnl5KAWiryVVcyi+/tUp67Y8D1E
9FXTJ0NnIbckl3rRdZ9O6MZMBKUVD4hDxS0K9pZ+VYUUQ09pWm6h7yZ5VUoqBMjogpOQZzvnW+0Q
mibfFhZ8GTRP/rnTwTAtWbPfcUPGV5HvOWZlGCXz7W1wvwQSq0Rzo/g/7j6KL9Zb74qmCiAxg3cT
Q+LRXDcpWlO3lFZ/cofQqufmJUS6PzhlNuWHGtubPwrCAXCe5jcsgW+GO5yZsvODZZeKeK4YrOWP
cq8jmB56Bv+zTK0TQEdP9NU3S7Js8d1ki+Sp3phZlcxjT2k0TikJH4CfFC709+YhrekC8BmFzUGw
PWlDmbtOkfJXY7+Nt5GiM4wlWh+z9ZqGer5l8+4H3mMMLIHt28WFvyApSrrO5IeWtN0fBbi9i1IG
Oy04kw0P+MQC2AKb+Vuaf6XFEydSsmoLXOeuzPMP3wK7YY7MESpXGpo/g/Q297WOEVTkpTR7sJT5
MGvA5IcOcuIo8O3pkna3IGO/LuzaqGjsJerMK9lUXKwAcHDaQglcX8mGW1gQjEN3qv0KLrBPgldz
liNWvrxb3fl8tRu9ySVfPu/ZhpdSOguXSLCkyFWMjAnYWv7zLbspIDIDBRhGX00Vqsmy1wj/ISzS
RIHXM3XV9PElrJj4chaJNmF8Zvk/V74OU0qqR2q5IAjZn9Pbu5LGnMBSzVaoBJJkDZEJKNzH3VoV
0SoZxbbNPiKRUFOggZAGtSgPz7nmKypx0gUyzsopgK9kEehjHqOZMBTLqFSSLe4SODaC7ewPi+vD
8zErZ10t7x1mYM/XV/rJLs/RheTngfk2GzWLuagYDyk8z0054YDfrWMfRMH4Bog7WH4LqUE0j+7p
YZmOxduQI1ot+YsnOriVgODsX6ONeip/SdhwZb1VnQaU9X3CCm3GclRiZYT+JRFlqDJnZ4pdRu45
CmgOIjTCmrazs5JzjJX34sirKFnYbbJZutuvXy38Ss151lr/Ro+SwgjWr4mFHu4ETAWcxM68zOGh
N8AA1lcDCE/OPaITSJPiilmDJc8NYE4h65Z3H+mckUQoCSfAbuK0zcLz+ycgD4cX2Gaii0cLn0QF
fXuplR0Gj0vYEWQxO1YSuFNLTBFIwXJsi9sDg40PZ707GViUZjgKDPw9creDRfxxvMGWjm6p/2NX
AbhL0sTwB6HfSHLfuO1ELV2/Cec6wgAYGsBigyDOM+BYSVAnN3xfyacs2n2Mjr3ApkRGaE1qI05Y
AtERkycKmtM18eK/IvCsGECib8ErJ2BRxwdZ2m7kXP4bqU2lEpErDEBtsOfzPO67jeZX9sNb21Ib
WK2JvZkMjT8duro2dyvjd/0x5pU8nOxrxdA3dK1bZ+mmSGtoUHLIiyJ4P2BThTIzaDHq60IRN8MV
fwmcrqdc7AS9k9Ndpp+2l4HZqrqiXwdQeetNjNghn1Eav/dIrtApQaMo6/bnOUTDOEVu85Gvg1YL
YDfT66nf+hUfWK6LqoOURJt6eMZGs7yI/c5eDy+jwTgKl6mv1sebXNpD/qYhevQgG8K9LoNAuF7i
FC3e1eAQ6Eudv0OxitaOokw3t7YgB4R4Ci/Ow9vp5i/Op1vmpPws6yubCaQxE3pqnGsKjrmVVqgJ
06GTSwH0eo40OGgcLnJlk//24LfFeuhwMUoSudN34iyvPUSouvuns+tjVLNWwPvigbdK7RbkMBmA
ask9MK7ZOc6vD8LKoO5oDfwu4NzobIBECUsSGMFPXyFo3xrRhgVoD7V3b4fFryZbVRxm63Lzb/17
IPkUfeYoJV7KeeSaKcj/Ig1xXjHLP580DxlTl1qV+KKdE3HMD1nQk830udmTLElLF2Lwr3SP0B9D
5Pdw6Cxuf1b/9Z3OyJxm9FI+sRCpFZezHY7UY2VZinadQI3/lk+3Rm/DMoWPYpALStW5Wy3LoEqf
oPoo13vZdp+pe+x7Q+Jkbx0h/Xdwkzs364+sv2LuFs2yGUd7ezSZoJBkycrQ8JhzIhSOOumAyZGe
0lz8saVzIHv/p97FoTx4idlstR0eIoSmd12rc8nJYqH1xVuHOi1XEw9BMlvpDEl0XV+kPo4pu8rO
oluFV+T/rQFyXVaF+5S9dh0qeDUXZTM0Id48yKa/GkkqMSzP9MoDhHRiV4fU5eXpx1cHLk++5OmE
8W/QDBrZYe3B8XKpQwlkkw0e633buxJjPngCOKNXEG3b3yXlRmCrHDfk8qdy92ZIWNr64ygPwxUz
2fqVuImwVZxutP1sHS3C8VwNygMiLojeEmAnUJIoiesq1Ss9skxnQdxLw0przhEwkbR3Bne6CoUh
ZKovhSxGgSMJuphKH3O48NvH6dw4BmF0oa9xFqSCzjXW835GPwxSyjUIjBzJp9B+66//p5sJaCtG
MKKt9X40+K7RQ1OdBoZ6bHf5KCnCZ3ut665uxOg4IXmM5937xv/eAXYdP+mJf1KoG9R4sl/lTrBo
80TVE2NJfhmO6N5yw9+/addiuSuW6Ah0j6kRa0f7SZQic7HHqF8IEowZP7DquyYyJYUf8o3XcKnt
cjsJ5DDIsJTOtCgBC5Ti0l0ghkC49cUL5vU8Velptdu5PIYLflvR6YFkrIKhHeOmqVXmci9Vo/JP
f23Akj0e236DGMBzyPge3TNw5T4LCT38go/EPfqykopOQ6O8YKNKa8z0pSATXCkctSDX50rVDYHV
gSmpVY8uycFtbdSk1JV5v0qkalzYvvXrwlw+CZ8RM8BqJbXVBJhrHg9ewx5zK96fKD+oR8YFcBUH
vikuxmBT5ljsJ6WDHUdBfqpYKvLiCBQ+qZhuYUcyFuVpRlPOARI7GwyO46P4q9nXfeTc96bfGHzY
8Xwo8omxshe/Xuuw0wUA6k2sOl1f6FQOLQVxpAHGfChMMea4+WAnQ6EaHc3Kmc19SVyXi47rllIZ
ztUFQd3Wv95Od9p+izz7pQD63IhdfSLSwUzEWE8zv/tfadEciZrDCR04YzVDhapinfCzqyDQQv5A
kZ6OmpvuN6N64tHkpRjxytxgamZfRRaLCm3QK+qTjLWM491wWXHi8kcY7vh42m5Z5pBJ3SFMKhTf
j6Ka4Cf7B5MqHPzl2/RrVwIX172x7h88TiHWUrgGxOdQHjetquQnIKokBZQbpqs7oN+czX2RiHkq
wqyMW9w9hRRifPkuKtfAJtzUL3PlBDJyNEQBp1DPG6v+8e0RCj+HsbYsRcl5QCeqRPAtZH9cjg/1
IQ8nPY5I5KheU42aSgIDtiZAQe4lHCWGRhNKKCS/J/OqoI1uDW8WQW0fHLpiOB+Y5nzQjdZSJL4N
fqhn/DbCXRkaV0KUngm6+/sIZItuOmtccTR/nC5ldbuSgEE+MN9+aesgFmAXYrIXfuuhZA6S2KFt
QDi89Mu6l0sLxgDRlsWiST762NCENNA5fVO9k9YGzIGew/Wl/pRm5MqGPyFIDU8MAdZTKpLpuZBC
CGEOShG2A1DvCTpuafNAXdzhOdcD5QP1qKYEIy2ht6ShPJtHG+KHPXrMdB8PrRQsSbZBMtFBkJC5
y8qTOHsSYU1r81uwcbiNTAmXOc1/rrY8M8Da7ABtE6j43wLFSUIXUmFp6EuhGhyxs9Y4e6cVUyp0
disWDWVxasNixJIyNv2h5T8M5emCXC/ZMdLn2XVxHPekPSfbeIbGQgctE/+nqGnqtbFbOySNPgsD
8EDjk7CWdeVE0nrgjxbJMCXDssQmdrWDPcRw2rVOPprERTTLMEYpEJ4PkDSy3DY2+f0ZwWBNX9X9
YtsgJzXoxEqvCBaH0i6KSQGUIXlmNvFAipLL/mL4E3eQnT3aaXrBLLHkDGuVmaKe4w6gz73oGfii
9QbIkI52LCLrSd5oFYG9IeW3Qy1mDIShl3EsYoJ9znZEukQN6oHkAS7AoiWI+YsifVTuBSegSMKK
mNDtH3/vWepo5sG26OHzYoQ4HpK7CZzzlhywEQM03NY6yMXhUj/rhmarShzhxkrJMU5/3UJbvG7p
xmkSU6ne9Av2ivK9z1/DuwXm0Z62BQdkaUOfecXelzQvAcIWgYwUx4W1AlbKhraVOFJjQ6XJ4EdN
B3BC12lFroqGxOOtXtMrshGlh9n3tY+xN5eVtiqgr2/qX6hz4hk1fJh2vU7Uh4BeG5i5+0ZxTgNg
V1IgDysPp0NhOhRSWSwopiJeZ5BskhuMZS3WLPuSZDT0ypn070sQL1O/fDnmpuEh79St/GC8Zjcq
Kit3JQw/0Xp/+rS3S1AkdZiBx8dS9JS1v32yTWDwi/mChv5ViQFIQkj5ZDJqi/+Pq7gc85LAiS24
0JPDOMPlN6CNkUF35lZGIV1dIvzUBtpfn+b8CzMaEq6sQ65jjOQYZMTZjI9mHffhFLr4CklteNdQ
gCMf7/IyS54ZoSgy84UtpnVJdVTyEeoIkCQsRgKfxxB+zRKh+lLNuLhROYJehNBoD8VDh/wT4f94
OXXHUtj2P8Q/cwxS3KzZwxPWA76ncwjzoVMyhgL9GjPh6Zfc5V/nM9LzoGEYItaxplmzZEP+sxoL
mOEY6GDeWKI8z5cfQx9Wq4naaQYCGAF/DsZk4nO/gQ+W57AqFuk7LNjtsJCSAV83pLScRWgpg519
Zw13eXuGUItGZL3ehuNrybPYz3avKk+YzFzdCcjjOh9FQasmptDmiIZDRPlKWIN+KsYtEiTtf9/Z
7SpIez+VA+hwAmu71lkivpm2URTbOIFV2ZnvpSAGqSaHueGQKIXrtL0z7yWDnOuL7FJEAmFG+cWL
NpeK89Xqk537QOL0gT6UWzNJPZJVlamh5xWUo5sA3LkJoaLw/ixNMVesNd4C9m3G/4QAV6dDIYC2
aLGCfIKogRdlqo70206pBsEgm/Mgkh+vd9o3sc3sd/eirUfiMvFm3Ex1hWOUHrD7qk6y2i5Z+gkX
b298uuVdpe0M0NX8NaE/vARCJ/Xqy1GgQCOa6DJjsuEOtEDGuaE41WaVJB9ysejmK80USV8n7/Dh
owxsTUP2P+WD1JvT18fFXvi2+hLGVN30F59uakHxHxeZzp+P85KgwDONCO6eVLvb6yC1M/5nC1z7
c6KaeiOSrYVJ4lkY4712gJFqssjCuIRvk9W3jrepuPgJhSo1Kzl0gR/jLLho1kT6Zv4UdGTDM08s
0JGDKCAx6LRWzWgurhzae/uUxGZ9hM1qqqoH/4E3fjaGeeoUnqu/02Sf9jzFrqSQAwR0lnuvdLQF
WLHMrJMkIO+BsyARJBzlCTX9VoyvM4V9s18T78+/f6YkmwzE1JdSeO/N8WqRFyZRi+MQamJoQC6W
HE13QnFgipoqTqdWSqphCVlLFLORx7KncxXl47YqKB4TYfn0l6bJndAy6edZzPRIviNycF2d26IN
PTINYccys4b1zn9N+/2mjkMw9Orypyd7rvFzgBmYhzUTzm8OkSAuXj13iBa/iz9ToozprIlynVvJ
UEiDyWlAy8g3c0qY2qfp3zofTgkGmdSSHJQVzGwdowsV/llJxtpzhFweaOI7hjuxcRpmAsWBTXGW
xSZ54pNu7aQjGek2rWaoZa/wVgCloIOI5L3BNgKaHJCFGMuIgIjkgFSL/58LFreiyDUkpsJ6cE1m
zOJwo4SIyGTbz7EzZxSaNSEJDa7ZPAr/ot23pkV8im7XF7fiVlHSZyLUlKqaBX4yTJ8TC5ueYrNB
vqGesm3LxWOmxvIWPBg7vHhB1iTgv0o10s8Hd9wj1mysgaU/VxRaqurP0ezBKrI7JA+vV6e2Mp2L
hFPYQ0J4AA8HLOCpxbellrvOcnDeHCAgCcztajP3DLl2ZwyihjBDi9W37N6KJf8+l1LJeGnNC0FC
YShI2Jyz9ohtX6yb6oKWiLkpE+QfXaPfBKp2/Cis298pztxhwckC3gWZq95te+VlZbtg7viUgyiU
UCgWiK3QECLspJ9G0cAeij8V6iVu72cGS1JSALdW7P3+HilNYd2kBT0pw53fiFv3+bU6OqabkaX+
JrnBn5aM//G6RYgB0cSbbWX84haMYSgRf0VukBWpYMYy3OVvXWZt5qOu4XRgiyxnqhsW1eOY01qA
8U7pBwef29ZpQ+Ek7/3et9libBNquZnY+Xt4fZzqMTyMMnxKkh3TLTXZl+0g1WxotKNKm8IxIT/H
sC/GktUmJcisPLeU9e4q6H9oU6PZDyJk63EqfLetKiCYCRXs6omVNHYERpjjCnuSFw5ko8zhhPDN
cIWXtEfCUgo+5g12hvZFrBDFoesARvR3hAgdJzXv2ZZFuvjWQQqbJl2QeFtkPK3IQcf55NzJ5MjQ
PNDioXPlSyvEqeH+tPt8wlC73PeuSGLj8aDJawn8kNZvP8uPHNA07MYFRuhltQF16Hx2y3EtonlP
WPuEtxrphMYfx2F07fFD3Ebx47AfAnZ4hPrpRETRol9MFYUrddRUBTgMMtq0wsXwc4Sqza5arpwz
Rfpf+seW0KeZRU+J5tQrF09bFmUO8tnxSXayPRItJkJGSkWB1A+MW+xl/azqW53yxM6DhJZK05RW
mz6Pb0mIy4/0BM9HOE/8C9tatrHgfou+cDFHXYRzw8kiMowbUDP44UKtBcyKybHtes8NsCmRodD+
5hencpe2auC9RpBpQwPahjfugnVnfStYkbxFQaL7vx97pG/BytyVjhHMvxzeP7v7ind8DEcEeG0U
KvsiMncYr4SvlOkFI86N/t4w+PTdR/CEMKSl8D62TpXXheS29hEJt1/75zkkZuZ4A8G+PYGWb5k4
qXE+PEhBidOHXen2yHW1LijYx9x0R2bo3ESma5Om+K32bz0RKrAKrSdczQhxY0s8kLO7rhXHBAYc
a3o4GUjUUD2fhU+MPWE1fXbbhj0cTHbgYR0XyOL5b/8Yb5/RrbH8oCzFDQvGAIpi4ANfiTkWFJCx
zT6l5ODus8nzSHKpa9ABjAD8WwxxUivIzM3/NyxojfaQ/giYDa4seGWVvThCKD2rMbSo1knUNglE
2C5q+LbTpn8WltV2aSytlgFiUkDuGNlxZbWnBdb+lxw+o6MQY7gONsfO/jZpXObIrcudGwP1yoS2
iTjswjou+3oiFPNjXmxdxIU8l1RejNX+rxD9zTHca1b96Vtr5QnUlwlEwCx09SO+BlhzOcw6BOg4
0qy5G3vvACuwKz4iKVt4kMa/UShEVbGLtFda8149tCXkfNxoGYOWqbNbEfnBqFxdStGzbaN8FOl0
KS8vh4T5wyLrMEbeIZfv3wjwMvGycJcSndvy2szUAX1pPgKUKPKeOAnLkr6dM+DtilWWzCL91i4l
payQoxatO43Kf6t51DZPiLhW4vMeYZAbiJO+H53UXD99A4DNpYp56hD/eMRL0hsZuPUgxd8RosGB
+onVmZuSNdvx3nx1CtzBfZcdfEHZlpk4phbk138jvZr1OrcTPBTXlacRXxdJ/CzGtgC1uJ+wj38K
LoZuuCzfV/+6wCt4bDmKNcBdJng1dykKAV019sNXinQej6WAKq3n4XH3WzXSkQPr8yAYYvehlXTP
/45hnmxGOh5RbeDfxcS/Kv1HLc43WMBcQ2ZlgKsQkt6N2X7mDPxZ4nBhoNvS1kbEGOiJKe1Aq+mf
zbCoWjhibHGbKYn/1wN+ZLioOBRHBUHw2FJ/k9hcBK1V9Mpk5wf8zNjtdPnwp21xzXzZa9XJrdV5
PuMAe1+oet54dSAH4NPkH1uhZKTNADQTOyLe724MSsxCpBsH0dYwYYiYX14wa9OSVD3QNTBAqciM
PISjHPF9TVpZX28SH0zBQ1sIxK0DXUjCRooaMUxx7UadzlaWJRtMwyTlRXCrYq+N+QiTqquGZKwv
OuO8cqi5M+302PiGsMtfql4mBepToOOoVHlQUbXS9TTIrIRj33aro1l4f/VM5+t0FwvEfUIc+tBS
QAIbd9o1GhV/dIu7/ZQL4qDU4z+I0DYUOEY8imEyqoKd0w+RD1ebcmUZ3whIBEgG0rmEhrc/yq4l
NodbGNU771Cv9woE8N3QfDaK6m2QUji28cqdVoLLOpJHYGX1JF2OzlcqK9FQRM9uct5QN9tmKFhF
PHfpeIdGZLA8WEOR0MMFQj81GXm4OaFiiOWt4HmyPHchra0U1PFAG1JIqGzM/ShX3R4UhMfZeIAc
JTdZEkDWuLTJqc46yKcQyPGA8sU2rh5/hsfoAy3uRqVNJ/p9IsGbXNjPTClqkYxn+Nf7xY4fkC8P
ulDDQ+VrRfJFAqjMriA9olp/4P1VLprGGtPP/jC28l8PAEckRNOK3fno1b3AfAzb624Qa3sAokZQ
jEOtEAd7zgcWAjV5gdvToDT6n7z7IXGomUBmcVMA5HlY62IENtRCO9H0cQeSbpnWZrfcnQU4xWla
XGqSnFv6fHW3wh4nvCgKfNkfyDFf5L75Kz/ukvwX+wAG+YuWrLi5hmZFmp59mz0ah/TD4cRvOxxK
aZC2r+V41vTvSL5Y39FzSkp1ocT3Z7SZsg8fK2yZhIhwQ+UuoQ7CZXJttfwRPzokgWjtcJczzB1U
3edMyehpGVLG+dYsl62m9+gH4opjibRHN/FjNq5SVBZrWg8zhxwvF9QH7WQN8dv6FHjkQlx7gPMh
oFyez0SZ7elHFjHcppwKWnQ4UshcWTQau0iNMDfAEsLR5VeoYTo6XNK2cyyFgFlmATkqMF9m/sH3
w70ZSJoRq7cjjwDx/1v8ano4+VK89ht+fSjUPRejK/5yg0Sgqk7uk9jK92EcOcto+eUhVpk1VCEg
PnLbpJHEnhq9PFeEVEPT9h89O6mWTPY0DtzDU5tUb1NgKRXg5kEOxPMmavZ4gEL8I/8YOq87gGc4
B9tCXsqmgOO+KgpfiO8XdlujD5XxPa2P5J+6XyV6GWa5FJU8FcafUgML3PjCJzPnzhJzasthALEJ
MOfG9M1YzqgUdbfMtILLP6ZdMyPo3hNTehmLBYjVBLae9AXVYBB2SFfoyyvf+c2k42CKUll1TtLg
rjP4P5UQrMxUbGC1XyGc9xlmRhNDvLmRrTHUBgnTNUCnBfEpmtNLveVb2dtJjJKQ6O4wNqsSwlX0
eYPZThCev7TzP1zW1ywJ8tZRQECcF2qea1F6QZNxyUPocvJ2Ht6r943ZOMsg2uEMlZVitCYgJt2T
gLkZWPXY24vI5AHmPaAGNeM8y9lu5qgf5KIbnopxkZqgOcbpwrQp9UeuxRQ+YPz+qL7mUJvLhKuZ
FstWNgnXh+q0iaJAwZW6yyZ+mHcBHPXMYdfexYwc8IQ+VXFQ3xJ0qHgs5sE40F38TesDpEtuE6Xy
GNsODQTYi1FiLhAAXUMS40fSoJr9YVMHrFnnJ+QUb7Cfe2DPorVcUTm5ZrtedqEt3rydhHHHcvCG
R3fIryMOdcs2FnrcsFd6/u8TCR+mnZLOqikJZhaS+WNckIP8yHCZsJn3K2SETC9hgaAQUvD5W9S5
xZ9BLy2jKg4WeQ1LjB8tpQ8CsxC65giJkI/U82TMmDIXfOEP+vNUgwcGS9tNgpwj4dQkmnq1qqjw
c1tB7mkGkns+KNGLYriUrj/ZhBwcC8ku7oWWpXcp66cHC2J1ancbeRwi2VDWZD4pK29w2iLPc76c
3s0eitSJLqVNnTGsCGPEyLI1LS63Ynfbnc5USK7RTd6XTCo87EnMgNQKdm4TvKupD4BR28yM5KrD
Fqyd7FtekEsHvKqttwej2KCGZNg2k2H7RbJ5oYz9rA4IDU5ZPhg1q9rIBe/8j8FnMO2FwGPCM1no
yKBX4ecgLIocpKauzCQWpQLuLuMQAVFY9mco7EpfS14sV6UoP4yg6Uq8k/MMXtoT9hvTNVogqV/K
K2Xd0S1RzOel8NTdKNAmrN6iEf7M5BNKYCBsTlTbS0yX9hLHGub1h7L288IYZgrJQlV1Rd8zs1qO
bY+08Vn2JhHEUwQRfVfNlsKF6yC81AsmiKfYzNOjOK3FFkLuMs9w8SeUUrTQaV0oNR5TmITQAIsO
5pOS7UPOC7YLFivOuOhmgYFKmXtzEIfjaXYRlG/DgjwuLWV9AOrsaym4nGsRJ1fuTXQTr4Un3uhH
bkK52lajE8zHztR/0u3ZY/bo9SW5JbIQTVEzFxk7qXqeIhEObvFpuIp4llovZRzAaZCQQsJ5d6oI
1pgPjcP5RnGkZBWPfljwc/a03ygo68LVq3yv19Zr9BcKVGK0vmU7mvuHAM1efb4Gma/CV+FLDYL4
R3ITDLgz+XsWRw4rLHYFQBT+NnP4t7PV5A+Fvq/BX5K178057d7cJmfS9/VVZU9hl9jHSIEnXhTp
mwNcIZVAvaiOdTwS07ckcRtQT1sKDDNIYjNsKc8UIaAsaEVa09nlPaAZTB4+7RvaWsDFye4EkMqT
OuyOrlRJOSZHMpTgRmDXHw0YsWVk/T8IO44Fgth/pMgSS7QK/CEIb4P6lIBNOKB98L4rUGmKFnCG
weobF5lCmWfajEuX+IegEvSSLa1Q5WwATDjJKFha211NqB15GUJ/THWmeC7XGp1Ws03DkmmT8xvb
evp4nZv4zRoBEfsPt6ABU4ao7kg1Zk8QmsCyyg5xKebhvyOs6cLBqG1tx/xFO6JPZQWaHkxkvnG3
b1m1xkIj4kLNfOn0lMRzpkAp+/bx1xl4IyiXy9G8UOkWJDufVRpAXLOLfk4aDHbM1HlmHtJMzI7C
YtJpx/13VRO+N/jBYjjPH4jWHOudd8T3EgUzs2LrAXiIcxaceMtRcaRUEqzhpJpMOiXpeCuy07ZK
C8m8h0YvJDJQf7Sz2k6Wo+7RARMW9ARRCYpBaQq4EHK97C6uBmaOzJe8uaHxzuG7IbxZVaMDS1rh
gy51YRxz1Nfyaszhsy5AhefR+BpbVNwYr4M3XDW6/cpX3iQ1VU5JweWskGx3nty93znjzXvhJWf9
jwRvtaVdfdFP9N8pjk8+zseebMnacbLGDGk5pV+OVP9lHyWphmr1/++Zna4DqllCoaUHcNyRbyTX
OiYfzyw96ElV07ejetk77Ps3y/1JlmgCeKdCC0I/K1KTCOIbhcp6WyYDs8GhykUkk7/N0ahE6aQh
m/No+dh01lgMwSjAwtF7dfh+ies4hGSJ1irO928OMlg24y8gL6QPkI3THMNv7NGdbkHa/i5Od4pC
qlE0EbOO0xjPcS7tS0O0y1H+rqbxNcQM1EcnmkNsO0oL9xML4q7zrPS/G2Dae4k8vkpGTrH3NHbu
3u5Ya/dAhn22mqt3zXFeny6kI9yaCjZgJeax7hpiq9WDaUFXd+fNjrUE7YsFkxyzX7VxJChSr5Gc
Avr35m/JvkqmzAwsYx3olYKzy92qpC3f6mBoTbPjRv2/7h1eRDfpqKhU1SqA+oucvsZtYKgkuAaO
NI3k9cnNRO3vzRm1XRRfQ+MkeMPoq+8InKZLJ6K7BAijHToO2KZgk6vkFGSLfGOkVZy1Agd+cgzd
5+wW9Ph75+K3ZV5szlvW9u0rswZoGs0Ffc357RrBvCXuYk2SokwNqFYTFray2c0dpGYcYxELcyhM
2t3qTxGp7B7NMvMAlFlbEGtFyAi7uwBQi18tU5rMW6DQqMNJ4/1fUWFj47RTTlsQwpVk8Pl8xEAE
7e1ygawq4n7KvqWP92QBio/dygDyWwphV8brOmORo7G9dybr8XbbUnRDKLb3J7ED1l7XhH/UZFpC
pqSnGTxi7d/Un4IgbNabujrBZ+CV3X2SdOtjDLdPGHV5vUDreqWX5uqozi4T1k4tunrZ+BWGfnuI
S2G5Gsl1aCwy9L8dckCRxRzqY6XXR2+Dn0u0knaWsMsD62Vb9fKQvG9bNlVFzC0GEjrsqW1lJHON
U1CpmRWfKjskp9w82D3ZUYkSFqW3NRhspu19gZfRzQKjA4GSPaMp88V5xMEANSZ3NJurjCvQoyN4
MJQzXlLQ9iTrPm5dszdIjfnwA89UqSVn9xl45Zc2vkkDp2IQCWcwujPHsH9ZC500+7H2bYm27/Wu
JCKIIxZ0drrlm1WFKnZPhHzYKBxWayIGTO4xNtOz4/r/bxWM49weorxav+MfH9SkZty8zVnxtOpL
x65tbDEch+nJKClCip8Onz4p0kjLe/jjdzMzEA/nDSRpi8AjnvvTAch0ApTFatP5gyzh81h1HwEu
p6aUt5VnY9GbOcv84meTTA4gZiqd8rPHAX2spYd5vUf8QuIEVOKVlsx3nJO4zh8GMt5vnDGY1r7l
z+BKjwRhMNH5ovDUrcowi9txA1lBYeNmVOaB0wOeyeCRcW3OE6JYBJiJq9C8FoiyZerLkrWlhxfq
5dzCKoGc74Ay5C88OkHvwCD6CxxWlXwdKWe/Sxe2dLv8VCKZBcH5FRyU5uSsyPcnML9AdQ7smY5C
WVSk2kvH20684SDVOEB/Fl4Ch2lpB9TVaIyajnGrDRfBXm5ane9mfjbAkgtKtYty29NTPAZ0T9pb
zHeyK/jCjytEn2NOzwybH3dyq3Yd7rg/G5632V+uTFmR0fnQn0IaAydjg6smL8KuNboa/s1dmBjn
sx0bttEY3HJpFPlAyZDXBEbENgLNG+mE/vNbmFJSkIR/llYH5irCydpUfXP2PNdBLzCd2tr3hqYF
HiX2FqVNZlhOG3bBuAEl1RPvKDIBzqLIKczDWgf7NghWR4W2294jW+Gq4275ivVP3zqsL+8wzxtH
H5PR2kUriKIr1h51LYiZABfhT7rhRl1jgq8vhmNbKgF5T1pXnwIfpKgkLTpmIyVgNAgN/OpDSHvA
HFbvYWZGqK2OGVAIV7sc8rGXKYDZsnh/S3ipg5R2jEItWXT9nx/CNCcICGgX/Qsu4/sBKnB8/tOb
1GJfhEyEFPFsg0/rtiz9pBqKBi8VKEJ/AkqKK76bl8C4T9jMsZ+yTAOW2DWa7S64oUA1vU2Az3j5
y9OIBTOHr7YSB4Hk/sp3Z/th326LTD2Z9uNOI0/OOWLAckp1xgj3KaVKbuQVtNdeFxSG8l2cYf9h
rwWTWCRLpvaErmMlQJZyPwD7aPBfYWjxMkyMtVF9vBndzhNKcq6Nd1SLwvC+JHhVWqT3/XXLedbs
MU+8yCiGWvw0GbkEgs42gOLXT+PXFcWMPFtNw00SHEqDisF3MIimVZLS5WNjCZ6x9d8P/JQ68a80
SktfzrLbNvEodKLJdBd5pynBvvXkFOnYe/5Ebc4ohO9GgdNQjHSAOHisrbAo+gNP6LxXtPnR/jL5
BuN0qtzWn3wnJM+eZjJCPfdzKYoztyqFX0DH2gueWb/7dHdLEimU8Zg5zma0kmNeXQr8DG54elst
g2mXhjtWhp3JCjXwGCiyi6afqAAg6lDPT5O9nnPPBGAHctXl4ppOiHzt0VtlkL4thBF7oICi6K97
MQIWjLLpz31s4Y6GfpmfkqeMCfFR/4wVNPwW84P6I5IlUFqbfSqQQ+mXWKMzLPi+AbRIHzAyNLxr
anm5LkBGGK9Ilfmfs39av5z6Q8t+G0KVu4pBIWBRRLAWxgbuc8kxfvLdQhymegfyk1RIzMIXEySx
h39pvYjM+r9YN54MCSQaa3kS2umApqwOzj0R5aAmvVAOcZ6asZujVqx7de7ClmjRRMPfJSBrQ4KY
y44X8FjRawuhylhyndLEp2wJDOOcfJ2bpiP356UpJZaFItiUJU8uYX6t67bwQgv3Eeq0rJpMvcSo
MJIBT01Yzwdg6GGUJKkGNbGFPKxoKwx29JmKoZ7Nkld9MFxF8BRHjb6/0jrIbjub6/OsXPaaJxP7
oId4y9IlsOTo2zh+pvsfqBa+7tZarFmKeBd6a3Sd9n/zcQvnw5vw5Zh3yfWBwKkQyumE0djTEnEZ
LQFlPFIUQuogcRwb1SnojSJ1vNhL2t3t63+9TBTGy/zyn6Fw5vTSXIXTVQTEP4Kts/LTty7iEWhR
oSWgMKEk/5RjRXTVsRLZDy6wNp12czQLKcO6lRPEe6SsUNC44VDAyPUpKcwBichwWPDNGpdo3uEe
ZYFvHh3Llf30dQoLJfAMY0CdTuW90hWUDl32dDioNlq9b0CqE2UhLsuHPyJsdn2Tg87c1bG8rg77
wHNfw81fVTpsThNpKC6KDMiy0yG202nR2YMQ0mOT497qD4kUhIOUVVXsPO+IOde8fWmVS014Fnsq
E1eTlUGxPXtVlVoQopU25+KnwH4gq8zX9e1mpbunMWdtD+yiuVIdF6veKGtSEbY5WA2oXDWJSlqD
DNjw9qfbmEPdgluSSHx5juRQx+Df3W2t66ywYOmoX3JD55nfqXPR73Kkn40Hz7dvhLz1w8LS2LPJ
RxbkeQrh/T41WlhV7lp8hRdoF5hlrjd308KBENUfISfpwxmd4QDA6NRj76z4G8kBTXFKV9GYKamA
8301bDt9Zt07KXZ1ioIZpDl3oQjIXNwt7klBAAF8Vl2WEVGINqEXgzkdfpLiwzNBqLYLvknwQ7oi
3BXTLVrK8Le2a9h3i9ScD3R1hyKvber7q+dZV3WRI/7J4rrBlHreJ/bIUaqG+l0CYyog9YoURUW4
9t1CadFgOJBhajA2Ib5nu98fLHRlY1qrshUu/wAeXDrwRgkM3QpFKvmITBoYajOIB9PYjOQyuGEe
ogaXF8flqC8PyP2MEjyXR1UnSqIKqkgiMX1UHPZDW20XNwdC0Mu4fMn9SF9Hhb/eS4xTf/ZC6ZA0
IJVth4nbplbJB5fGmC2I18pY7VXxiGnJFpJtpaT4GDW0EcrCvikEqRvHwPTuMHmxvPypgRl4/I+j
tjZR7lrBGdF/lj8/mr3cujVF+i9ACAt4+YrkX12PnqHA6TQBUGHq9sMGkoXMOkL3jQgxK1iE0u3V
HD/Wiq0uLbz0CQVauZ/ATC0WJ1m2YAFE1nVwQZFs2zlfd6sV4SmbDY6YWg5bUyQzg/cz/LUKAAVL
j0ftyCfrQZfcYxEGdEz0IZiwoGpSu/bdN7eUQVazIgV3PEieG1oJ2QH1NxkWOw5fbABvqKjnuJit
isXZE/G5UckokXEYPRDNyOkcTZzOOgu5eYd36ZDn+BILtadhVjUtPkV03lyJARSwQF85ATM5lANf
KL8MhB16YwISgcPmRum0lS/YUO271rOxuYW9bjtkKh/YqB0BFx8JeEeSe2Yw0IGEVJ/nMkhgvasY
pLHDeZzLLPVCUeb/XnYZAVdYp2BBocK+czNjkR/Mgw9GUQwLq16megoS/2ubk6Zrc5KKb+l0Otuj
eLCxvhBCi6QSIdBYYpICDzuAVWvldwwxmXZ+2p0dkil939qYbpckCKLUj297xowMEqMOjCipADEj
WdtQQ1zKh9VlSE0UYCjp771M8qTC7r6hOktwhGHsiL9BipOIzgi5jEbDhy1E2tvbLtT8b1tN3aBY
5lnyv+DzcrS4LllnzQm6RmiKiDreQQo29p8LzrLn2EJD4wgoiXDuycl3d7WGianomHQGu++51Ypa
KJZep4vw1q7oawmw4UPuLvl+XQvuKQNNLenHic2zBgC/M32hDZVj3j8JnfgCc7nNy7LzqE1I+dvB
o4Mq1xyn15EEQKh5JU2B4eQ6/3yTdg6vlho66bFDDqbDI4nW9cA9bN2yqy4kRkdKNEfJdPVlWG4W
VZl8jvRBHQP7G9rxmRcieAV3bo9ThjeyOHZ95+iGkR8tVMUYqIgvUQ28VNnPy3kMmW92lDVLChGt
qPIALRe2oYAjXTlRyE06GOZSu/NgROfdbRRWW6WbuKF0oSehc7rHe7MDJBsRlB2jozYd6fT8NjAD
BAGEzZhFRx9UCAGdEgsU8hAjj5oP2J65yrGdS59ZRdSZ41DfofBEnJjwsi1cOOpKFR7uVDQS4MIR
LUesWJNAsXUV0UQq1E5k7UN862FQi9B0r5gLtlmbYL6naACgLNFfTFeLUvLNiqPzcQW1rrAETSwZ
kNi5tsSN0JdisrRvaj0MOvgwN4OlFtFmwg714oicynp2jFqX/jtYY92aFB8XhBK2hb22bLlZ+44p
Yuh3tMW4tKzGLJv8brINr2EDUqis3Esv2bHHkxIUsU2rpbvKt6Ozsmw1uu9yRvLxw/qUILvhkADE
FHv0/NQCcLGT1RkspVdJOHEuh4LyU+fdr5XgEpjcklkDE85Wf9XhMSnww6nhpjKiz1awJ/MHitek
dJzXYcT+gHj8vvqx/eTcKrl+4nKdJK6EZv+J1UHMnZNcsBpEea5ne1d/GosK6Q47R99McPz5V7lG
V8GBsdDSRPHGR0NVZ4+34Nypi6Narb2AyMzZUIOzROJKkZb4gdX9TJM+XJeGgotNyIMeB5bELCK7
rgnXoKZj7O4fRzmkoqosDOffw29AxmTQnHFKe4U+ZhYEzeF+YiUZFd09Q4yT40XEOf8mdit3oqWJ
LwAEXCQsCktGRc2SSJt8Q/OUHlLaCEhb628872+r1er1xaE9qNXX0iIjvI77tFgnKZRUBpmD96rS
4QNRDoZ+vbFHAfrJGcExbeNITGsJ/oa8lcdy/HDUdT4hi6MsNCRIFIwIO1ns9SuLwTFsjz3iqpAc
qt+lXb7/qEah5VZh0fRtCX6FjRPuBdVVxlWlmTuuJmESxeLuxCQKVQaW/4nHlI6ZeGvUvEz7zGue
yb7+1m8F5sFRHeLxPNph1dRmn8BZABC90XcD9ReTDn7cgiFnAksWrq/fmZvxrhYNADjQfWdUCXHW
yLBeBSD75n1C/mD318l6sys3UXkdLIfBLezsIPxFW4XieC47/SRFTnzlFOIfUNLjO8wzL7Jl6ygL
6q7N/aF5wKJzkio5A3li4vKHIuClWLCuWP3thzvyGItmVGZ9G+SqeK4HFc1/I2SnzUTC3jNK3OFx
yulAAVfGI8ja4WAc8utgEkq9l0rYf7lquLKo0EAA41oOFjUXNEWmf/OK7TAKC8z/nwwWycM3lfw8
rSu92eAYpxbdk0y1SIcI87D6VnYbecJJtP/3Hq+4dhYw6un00AGtlEEl78REOgHhQTvoC7GzPbFg
NUDHhWoGYHLMRLK9pR1RCpBiiZATrMnUklt1dc46l+ONNx2V8fiYnRIwObA6mWt2mV/+OVoIU/D6
RwDMvioiYvwxonW+uT7y1IL56zrPXUT42mOQVTVDy5dmVa5B8Ff+Eg/OwQyzzJlq+lXnT7hTjcy+
b0I20fuyJEQiOQepXxOwHi0q9/Aohi3pW3euGuP7TXMlwrhnZQsD3t7XaZ7myZaiIrcYaTpuO6Hb
nRP+12NiroJE1lrcdvzyPA+0Nc0LONBoORc2e7KSnkiGRW5ikJVG/mDvje4AsASEeVxFWca+rY2e
pAqzkyveZPc4Gyt/Fz31ZwppJMalAdbO1FrwB1DHQcfSnU3Hab+rvPq06/BdlJdSiT2d3qcj6b83
qs2wO5tnU1z1S28VdbBebz0knSG3qIhvKtWe7Jt0hS1FGBIp4Tg363FMdL55hVf7oqiSS9kw5c4D
IdULK3j5OLdZgkkn0mX/0LjFWyPKkJCowikkq2usN9rW8YCtR1aBk1OL1+haCKWo0gOJ2lY5RIll
f5CBk87sw5yR6AHA/KoCTVZAX5+Yn3grnD8NhUI3rAL2YQ12xyRcYShcjKzlPayRR5Lm3DYxsJDm
WiiBxp1oB4dWYm0vx5b7HpKzREK1UbVFbo8zAu4LSOiWZZDpVQLM10Il36gvbAaQtAEbIEceZY4+
7Q/GgmpWPd1NtVm8qgxmIIsy0Rjcpqke2UWrcIIVGq2VS8Xc8kQp1MCPo/nqKowxR8aX2m817MFF
wKT2qjgDz3u5DykA3Hx5tTZHfh1p5MX5UBGkEol/T+5qgLw9KGzVsR3v47ybf9Ht7V6HZc50DjMI
DzZlJ2w8JjEiX2YCm+DybGl7yQ1TqOKZHWLeeTk3uvPiH+U8HWBqV315EfGYDxok9ot0Vv3LC2/5
et0ab3K3yn75K25rntHinDG44e6AbK1pBk9WRfs+/glIPt9dbg7ZFgsxMSxi8+1HcjDqJ87Kv3at
Hc0DJrLiUs0XqhyQpWEUUHo5iX+aLLJPw+3EAmt/cVluGAaGnoyHv2CfDk/wipkGW6/GtY6+E2k6
JBepPE17lnm46q/4K1w3CuNs8W4RuvCaarHmiwilYJU9vU3NjXEXo5X7oCXlnEkddo/4TY20JvT5
FpWcpDbB3X9WkEZjH1GW/XZMP3PGynOOg1XgQM9hkUyamMMoeqdnk3RqzGSvinC0nxHveYv6WXLi
xk7Mumh1U4VJlzN6ipwM6aeNJIN/lD1/ix38db829I6Q6d3PkdNmwvDQqx+Muyc5guuhtsmjuYBI
ekZ+MtkSCwxvwVvNi/4OJoMZHPeMudweNr/2FkRSzx4O/PykUl/jelaLQHkfGqXC36SMuJSQYN1r
LM1QPAMDsDY7LsMufIyGvkBQO4I4rwrE4sm8Z9BjO+EoSFJdYr9hy4Mcs7to/xcXZY5b3encGdLm
lIjpuW/9SPBUEX7yKHcLc7U3Lk3r0bYR7z8urerhXclDkxIW7cDlITLSgDkfrHrKreexggBwYzYA
Vb6PDLZzNASZ0ys88bm1QDoEHWl0BbclQVQbS/DPhe/7ZR1G9RMCK+5yRqneusYECMSN5RyYoUnk
sG7/xWCZkKanIwiSU+LlLkSX6Wb682dw49SlnfuWds0t56g7nFyToTH2jBtcxejAJW0CuGVa5ae/
48bnkKPGpFJ82NGQa4YXRnPb8COoonmF9WWMglYTEyhuoWUB2nYwMNm+HE7qk3T/axXfPICDXsQb
s4zkUQjb7eM6lQOXECOuim77b3e7BgkEL7EzcUK0AKZ0QLI6YF+qpIODde3uSBnx4mB+RJpcIKul
pwCuEQEas2EtsJzjrQ2eZwBA+8WlLsd9GxEoKDlf7RHjvc8F21ouvvWgrlZnIWfIkg2wgT//dgrE
a5wgsBk6EjxwVxrhXRnWnL0LPVGp5VMOa2xdt7ajoYijTnBtBOmHk795olBWhzrRoN2Ol3ODn+r8
8iVMCuuYDqCjUYS6qZSHOWlreZfT+G8rk34JxzJJZVdkPdwXcGwn42wuH81fu4pVU2L8B+avkCiF
cr0Dl/aQL7i95n2xHZZFQN3I4XM6SsycqpVzEXO0HPpjK61GB4yxRpKlAOy9Z1iJC9Iq15R18yVp
tjqHVijVMdfcMA4XFLsDhwPkO407bNdTpn1W5jT+HK3niCwYygYV68i83C3nMYtqD+1JFSeAB2z1
rH2X/Z8c28tpFmTTIApfP3NoGz1gyJyETwh/oyQ9ck7y/nZk8JwUj+BBwSHYzC/cUURqUn+nTCzf
iHnDRAivZQ0cCblWuTQ56RKFnS95DJ3luSfnXJhgBBS0+qkOyKUBYIZ90ha8W/W6o7IAcp+d8NC9
7xTefjcoFB3cAj8br9KkyGR8ZpQE9sGkpBz68Vu++KW8BhLZOuR99CdT+9XbHRUUGNM7QojyXwUa
++vEv6k6nse7AVSbW2/uiAt2I5PO1j+nKWr8nlbrRHRj7brxqbmKVYcVKlmcngo0McEVCDuAan+Y
d7rXuQOi8EGwjjqRupbf+05dOtB60dTQukY+OCwo+rPNgAJze1/5qrGzjZqTVQhi3INrH+O2LqRF
MC+l3liFg+exdIIsgLjvBBrLnpyjFFrukm1oJRLNpwuCEOsNdIU3PfdzYMH/vC/NTCs0G/r16vJJ
Becgp/vrIOFPJjzgh2VZd9rztrUcLJjZ4lCs3Yro1+oLtEj8T8wbl+zEEm1g2JncXnn1P7g0z+g1
lt9q0x5YP08R/uIVOELCfAXOsmffrvWD9nKB4C7dc542bqusP8Fzd/vAM0+Ig6wQBi2OywkUfaL9
vmaslfTLv6uKy1adiB52+Rb2ePCxY9SETmj4PTSKkXKg3JpnjBE65eZ/N/vKaIWaqe2mbhWcDdAD
MFKlWJxxfpMa1UWw+vnQTP/MEtA2hSq442cmzQXmBNzUmT1LVNq0PqoqK7xtRJmPanYluz6ZTMSd
VCa3AZbrUSeEfYvrMEnFRW6QRUE74Kg/Bbp6fsnsRcpYBW3NXkpAJH8RPeQzs0g02D34FdssOcwa
TerrVru2fRS/ywSYUFThPBs2Zw4/rUS9Fh3F3LPru3T53olwpqjAtszNZG2yNMjJvO8JI/1gaqPy
/2hJ5/pLKvbOMc+8WNkgpKCAawX6MwnYoUDyNhUPXEzFpe+c4S8hKqLbIJrTfNl92hnzdnog6SK9
tmIQCSOCmZI867UEExlDB9lDAGJHVp01RK8tKhnxD5enVT8cBjaCItncRGp7+WpuBSKApvj+zjIz
XeWlRLbNR7Y2ZRQ2vHlt5qnyZmDpolt5i5ncKA61I2BuA/8LhDlpazt21pd+WzDo3Xt+A546Foh9
i9ANhEhO2b5226O9BwisBfstVvWtrXvKG+gWIcrRL9AWGu2UniRu4tClC40C2snODJ1Qs1Mw+1eH
5Jw5nzDpSGIyD+iyNTJejgxrV3BdfRFYmyMcQCC4AWEuAf1ogqDX/vO+xAzmQBAkkeIAc7BBaLo9
+9vdPKUV5MEVaXpwVDm0FqJe0EUqThzCnlgK4eStDdcgzrXdL8vLeHl1BOuS+LI8a+IEb9N6Hq6/
Bnjj/XRH1nYGIP+HG8by5dHUB+sseDj2bvngnz4eCnmL0bqIijF62jL3r9jP+wR9jyXZgCE4muCk
MFDwL1GrZbwLJzpDuzk1YD4xqScCdHdBGSaWpFaWZr/26sUi+LaCieTlhgqAfjTWuSNSz2sNBE4v
9SPf+EYi6gBVuwFG2FIWwR5BJXzphTreL81tsQ0G5tjifx3HzKwOZwktZvjfigpAUFl8hZme3agu
Gx4YvhHbnfpgHZ0NepWCcIhpGg8M3YSLbdf7oNkABr7IheW6Ha8eZl1iUl/WILuT19+F3H5/gCMu
acSpigyTXSEXkq1uqP3zGIAAdV0dE/fgUUZ25z/vpvoH5tW7mW8BBEsVKWIoZSynhPjM9YFbZhEC
2sFFHTnju4OmkSl4tMIgBGKU36FtOtlumVUDBRRJyAwx2zygOc9LJsYIDZXp5FtrG/DFkU1P/B9N
82dSd+ubWD9FxSql5Hzf6fIB1ET/uyZb6ON0m5P9IZ6dxJAYk/h1X7dkyHjDoVMHTIggG33vWm+i
fKbOi0bHxgRnJeOHr7MgyyWMQpsqzciPNRajGotXTpTqmqjgESRzYnKU5jjaCjroqH6hbS7JTAg1
0VX7+RAPT8vEfr8TqilXWa4/6FhjZ7TOdEfoKv4c/AXwS2xi+cdZj+bsH99L6vdBnc411bgBy+Fz
M7ACLOv3DAtvhSrdZWaoxIym4vDV+TDtDP2LpA2YSO5a68bAyGuZqyrCWl9SmrFEQ+jRNlUIvIfq
O8MpqcxybuwlMfitIJa6ELZ4KV0MvdnICZ0mK/TQ+JQ9LIOA9xyWptxBb+m8vc7y46/AlK6/9dW2
t71hz1cnUTiv1AD0fOGhxeR7HIrpxr8kc7NtTx0v0s0kL36Qg6st2eNKE97csP7GO3MOrmMRR4Fy
anPyz3n8xf6ACsRnlEUvKvRVQrrVfSMaUvTRFXkURF+kcVwMaJoBX4HcHjkdu8M1eRoqIRYL9On2
dDWVl4QUG3kgG866KjExFCMoveossCEfDG3Iq2ATZTg+a7pgY6AF9NGotyXT6ZVR4XOUnQlV/kvh
/+h1HGGCRoMWLx1BebXun/otl3aiVK9nXaCxUd2u7cTF3Ei1XdB832bbY75zHyLDCmCUFzNaBib4
7O3ozlu6sbQ2lisbbUjWuDkjcYbvyGUHAFgEfApIdWd0gCQRd7bPkP+fkTi8GOBHzMS5aapkg7qp
Nz7lHmnQrK0JN5kt0dhm1kbbcLdNLufhF95BVg+mKUmFCw563p0E/+WfjwxEl6EzTndlVwveDeuw
UN7JG4CF5NBemcZ8lW2jGNWGsi4nH8GxEGl/oVrtNKjiIqWN43a6LzkDRK9dwjXSi0/aaBeryziC
4UOaY3e8EqUvAk/Br8qc/pnbqxsxjQvhsjTEvIgrJcCgo+UD2AUOdzDNZPGmhC11WN/pPYRITKiX
Av11udAoMHV+vUZTl5BJWBt7r4JRVjI9+ZwKJflAxZB1JKelT+7cvTjqfFQ5rSxJyWOgVL2eijZo
iE1UiEGKjOe9MpAZNAaW4f77NLB6uddRYd9wzZaWheQEjFyDbuKH0aR/U0sGuumAvbqhRINE0UWA
iBZseVNBBrDCVkaWHltWbg+zlB1JwWS1tev4v8gL6rBWomjEv7b8ntniiZUtos5houxDbgpkH5oY
7R+oYQjHvRKgjoyksPVZUDDsxe0P54d9lzYMBmaX8r5RY7Z+oRcCmB9KVT9vVXA7FP5+3UzHBuMN
dGLW7CnrNzv4NUj+I/qoQbBL+lFupKL81f0Gt2Et8/yX+t4WKwnbc6MvjwtOdW+m5COO2KfxA6CY
MVzACeVJlT4kS+VsM+BurW9h2HQrw44Uumd6CMABM6PfPmuu+6LG5hrfhlq/oppAqBYsClkIsUyM
DPSy19Dt5LH3F4M62eO9H6EPYMVRrPZi4N7AdX8M+UaEO9eQrhiAEuaoAFjri3V9/diLErr3XW/A
3KzrXwx5P1uYUN1YTaHHPpLUm1G+5nDhIWH4/J6kEQU/1ReO9VG2Q32ug4hnFbzHldRVAc/G0F/F
Hm+Xx+Uw3+P6XzciVckVXw4D0PUnSk48MVXzmQDUVdvpIJTJu109j/77F1tuZP4DioPAe2eRrTxZ
sYjVtL9n2o2qnfoPYDY7BSTB/eXhZcXPqkA95R0SQQGwQqIppdItN8305Tg4aczoOIAdxPY5XJMj
G3SK2wYx2BCmNYKuX2qCgktWAL/GG6uWbdyvnYs69GndP4JP+yYCOZB1OyyhIIq5Yud80FY13DVw
+qH061uZlYInMcNCkZcELpTm9Qa4S9RlRm1f8lyrEr6IZ/fmHLBt7Urqh2eSH383JrHCf5YaaOdT
H8tcRDJ6ivjYFZt7pbol0CIBmug2DY0PjZ/LmrKb45iqfAsh23OfZVEDoC3SrVv+cfw/NJYfWW9k
t2BabCUVJVgLUlgUWv3OQgD6yJ9nOYd3fn5eAOEvRQlioPnfJES5rnWuYRyWBQ1ZC0L+TTbUtCJ3
Mouve6/BwJK5fvSO2Z+x2NijStrfHtFSmb/0BX3fnu3e9PnPO8W2gFd0/CabptXufIC521r8HWfn
iI2Se28b3JKYCB0tzCUzakDvPDiV8gXdMTG9ihCLlaUsEsx7TgMYDiIzwOElNGF3hyMVKKnulO+1
WC+3+i5svxQFidxP7Mx1WP0SX96biOPqHCyp9o//s3NF7abOWIw04e6O9aXLjcw1kQqwtMAvz7/i
imSlDXzQSapHvDrpabL7sUFRO/99KpyFJEOs1JwpW0PYEcb5Uk98KdTZqUacwyheMoVSN0xAzKyQ
2AUw9fHDe3B8nnn5hktTEkZJbSw3BGi9oNEDB4FE2rVnkM5Id3jBDr0QNV/Vyqn8nHZlwoV3MiqU
8jh5lD7XRvqvtilEVmtWOqUrkcVDsFetxsc7APLJ6hI8/exnJbIJWnFKGvBhvOeNB9p8qewEj04H
3ydagY3c9bVuvRHwn+sT8/2VfQXYU2Xy+wXZc7QuzUm8u2AYEsgp2Z8q73GiMUe1m/kTOfUjusB/
n7NGTwcJEEbDzrOpb501smfdT2LjA/3wDMSNqIA58oImrhgVOSqHwUY1rOedJ5tqQvsOF9Xy2Iq8
aZLBNtzSyvUQT8N6xbsniDxuzMoJlyc3GZ8r+WzX+VXmHOE44tYeXY/ys1qvYS+g9iteH4bN98Bx
hklpb87Kl3laiFTR+GbUtu1pnHKeLbGhzHcZbFpnZ6LGcmPxp1yKsjinlbFIjV/J6melR55L9/6+
am3P/3YuSGwYqe1nxGYs4Aav5sfUqMQXZ2IEkgbXuf+GPVbHdYMGDh0z/cZhRkDMOhd8fwZL0n8L
B9JyVM0tsrhg5tO6MTFW+QX3mI495BTt3/IgFlfxVYka1cv2LP7SdaxhRc4LlXBRVGqbmex/mAHn
OYCrSf+AoIhkF+nChUcqKx2/uibX5WDCOri/pFf/Xzo9HlVChGQ0xDFgq58c85yrWznbk3qNyGkO
u/kd7IuFu1uZ+BWAOM7svkx7hCv7K8obVRVX6GFfFmkZo2hBoHjWOAYFbdHLV5/FbxtVKgQHD90G
s/abOvb/pIJVMyTe+hXTQn1BxxRBYZFrThCgfZFMtSQFn2ok3Wb0e2M3+CECyF1tGFMrJg0zw/C2
nKCP6L45tZGS4ER6Xz5/6734bzlHfUQ=
`protect end_protected
