-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZSeJ7/HSdkGTFg0tVmnjOvn3rqAWA2/7YxIMa682s6ZDpBBimT/RuBdiqEopewwEMwyhGrivSxUr
LrPJPcG1gGsxmtNspsOnaDXaEvbLyZhJ/XBJBZkXT/oomnDl0PQGIe5jWJVx4tJX99Q8w1AVeyBw
BI9b65IC4qr2jWdZZ5HS2Gtkb79M6Cj0SPo5uA9ovo9VHS0Mi4dZycdnR+w3AUVawpDYz73XJZRd
Im1cP97o4X7hQ/dQ3HLJHSGzkajmyVhO3A9jc9HFvntXQcbbE92E4KOo/58ZlwHr5Td/Dk5aiorP
8IBWkQpYJ19x+d8vEV2+QP5G/DXjRyvzA4Fomw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
kKcGdPmrFw8+sEcVxfDXiMKzk74mJc8c0FORfDwRkp1nXXvogQzuUxLgzQamWiu6mdy4GKhi01WM
XvW8zg3BzOnIRxVoXu3qKRNuxhHjKutHXXZDwKk6Hu3m24OI4J97SfEhw8CO+5qTsOINae4RQSgE
6+ZhVZSAiT/g6rYjLfRDET/haTnb4pjmzsSSgk3ouJFPWyjEVlDPmEe+3eA3wYsfN5Z+I+/06Cfi
4WAxCwoaNNTnLYMzTA7wOFjqxUWbHBxxSnMitkZRVgfEyB4Pmx3BhTSiOFCiOj2uQmWqRqmwQRO6
45ft+L5pLOTgfxSXMJz291XeqDtMd3hsBIKEvfe2Hhymbk1VEteEm9yEIud8YFcaoo7Dlz9c+/2b
VZgq++P8dNnqGAl0V2K5ychrGK4YJmT5nmcE9MKMQZuggGS9PXlzLa4BrDD7+LmHIVQQ98n2J9nC
C3tp1IJyvj/Tx68l4d9kaP7WAkaTjXkBkrMzg98Mnpnx6V6kzLCyCiEVK4w5Aerr3bG6jvQkVa+c
GZky2Efgip/RhWrzwvOM7iLOsJglH3km/UjsFVBhVDNuwlTUGfn5fju4pR0ODx9qjIbk+hl8tjPc
bgR0ffsuw7HGr9qat5+lzVzAiw7WfnM7X9oJgk3PzgTS+FPgsVdziHvgGdbCwxogl5UBKE583gUv
PoXubBPCvt7F1KZjv/jMdp8nQQzvoGf7K0H/1ZHhpn7jNVfaqJQGKBlI+99vtcgzFyD+IWv2RPvW
bsP7qu8s1eTMWFCmuZ6c4PN7L4t+lNvQHiglzEK+HTSiw+Zon667k0lIA3o0ywTTTcFbzCkKI5HK
/gliCA5VzXuC9k5nRq5bLjT9+zBG8whZf0S+23ZP1Y8jbUAui2lGPthwXzXzRQm3z5hRmdmmCbBQ
6VfTf8ifN2AIJuplbMQ3IDi2vt/5D7iYYJmoQrBHhZJ+0dgZP1Qh4l8PL7Js1SY9QClodZlW0iJz
GK5+DpNhs04qrH8mO7Osj9Rdb5cgWgC+eNKE0oe1xKpcSI4YW3xPQ6Bgr1b5WiB67xVPkQP7NSOB
LqxfcyGDpnIYtW33oHdb0UbpguKn92oD1jP1QqNbIg4v7YzvbB1uY5VsnF0Qxc4x0J0Ax2L5NJvA
55paKJvHpUKxvMTDHpUr2aMO7jVWzVlpg+MLM+dwhjCQaWsGOW44LqhyDfBY0fsTKe/qS/3uw/UJ
d61h9tJwKsDkUNc3AlYFWSQNCAvtbjNBONsmd553Eh3MX6NtKK2cyTgqnI5Rb2esiXPrUntGwlGj
uLyoAxFJ48ig3vhyCXTMTkjhR/k1z+y6rbTUXzINPsVN/tUONC+vpvEHPP+zG0LfNdlbCNS7ENVh
378utNnfEvQjNLvhJ0oD9pLw3jBeq3Fj3QdrZs3m+k2tIu/f1y9HzkfbZOHyPH4jUURSUaOhKFTL
mVMsSCLjFiQ0EkXK1RLMyIaUnGvyDttjPBPUt4oHXFqvwEGmymjJiV6yPiEGEyTKwtBxK8WbP8cp
62zTdrOdtqvvLNI36y/LlrIwmENIqZ19NzQu02RYZ1crt4k/X0DNkgxAg9jzZVeKOeL0DKQ+o1xP
0MdObGHCZ1chQ5DN/OHV3X9wzMHGrc38gtGu5ML2P5yPIUgiwdxMBe4Rucc/9HIN2I6Kl/gqkGe4
QIdEE15Iq9P7g9Ag3LQue96tEswPeyGH76IG1lt2jtzM13zAcB5UehjG0+63JN97OyJxB+jpQTMf
qHFWHshSkFyecCECt51xxFJrxh0nwFtlwwU4gYYktv7axyfGInjCLxNcw+THkYf0Y1iMNn1ZF77N
0JiEAH2AOt58oml0ZDW9YhpSlB12kECRhGLk7nJq4FgWPkFhnqyFx+sdLCtuuPNqIZXx4gTAW+OK
XyTv4vDQKu1XdskDFR1DT1dKP6mKeP8mLfHDi/QyURfXfy8UyKRRSTz6yWB/Vdu52Qr4NHVqBghW
ktBcbzv7OnrWk61ouOdwSs0cXnYxORoKnmlke0m+o1vFsMUa77wAXk4DzlZCDIIQnoad1gWmv1uo
ifLptJTNTsxC8W6rYDa6tOerZC99fcXsrwUO8EgE1AHLad60DMj4Z9G5YIB4Jn61cXwoVRQHI5rt
FLSLYgLauD02/92/rjvzH9F8VkdKaofYTaORnoNZRTTcnVEbxcQykckvTl21aHXwmsQU/zdfIe1Z
BtlD94UpDqwcdLj3lhDHh+3os414X3ahmnYS+4FMprcLn2vaA154BDJxtph5D94LMoOlIdb/8TZW
h9+HQLJhDI2OWWdaNedLQd1rQTRyYg+JM6wSRAM3Y+myKEu0ebrMWkIFc1PYKIvja6fktLB6+Nfj
3WqGTu5ExlDEbJGRI+0uBKKeuvOx4nNaLdD8sZKIJl5ZLgEsmH8AwKdWamnrtH/Yt6BdsUweu7ur
AknTOWT4NmnkljDXplLEIpTL338xlg2q3pYS43T5ElAgyks4LHmxCwiNQ92uOOmJ27oToUiJJCVF
YWGZ3RDhATfnzAMfkt4T1PRNQ/NgVdboXQTOV/0EB2DEUKT3JtbfQ8HAUTRtHt0DSV6wjSsY7jib
kteyRsxbvWyyaOkeiGtg1sh00O7ZFsfFrOcKua8VOrm+vhnx7emw/oy/hFJ/Bd8zTYaQq16g1vzt
v2et64vXO4cjWw4+EpzFZ3KgCTu4kDCp5W5nyN9R01Aae8epH5UxLZTKwl4nY3M4otqWIlCoYsRS
tgVYse429D3ccHXWCVvlvYVj+GjqsS39hXJKLLXiPd1kdTKtcw+eA8uvkRAaHgNdPPq3IGZvuGeH
KlWMAK9GcHPNmUeufYN7tMx5fp9F4pVM1eYvMxe1tLqEOBGBZ+BxmHj8qXs/14tM/y2sFaUiolpf
IOCEYcAs94uPj16twkh8aUt/NMFHJFZ+CqENFMePDzcVbTcIZBs5Uzi3moeuaEKcVRPP5dVLnY04
jGd2+Y74UcDqSNDkE08CvAalw40PmV8i1azDosuwUkyXHZ2Q3qHKB89Blm2FnoRX108TRQys8qnw
CdlIhRe4xw0yKeDcO3NIlyltjvuLpdhCp05vJxoWkZRiPkCNGLvoA4RxMp+eYCfVm+/ukBzCrZ/S
UBJDDYT2fd0PiygcJ4Vyy5lc9Cnfex8kAMP2TPUVr2SKz26+9hg8y8LdNkg5WZL1ypjNn9Asn32/
qrUsJg6LFLAQTaIvHMuCygsBJu4Gjreq6fOdGQCwDiplX0IaUJZcDZ5Tb4nKlzUGCewljduOYhx7
9kO9V+AXElM7XGLXItxRpGt/m+GaOvDwAJ4QwaZietw6wc/cFpuLuKA+knJhFd1/ql0LAxiLdyQ1
LZ6OV4H2TqeoiVb8BssTiSOJKqJUU+VObq9eB+yVWgPi7Hh29Ubnm6iub6HH81f5Hwi8aP4IJdO0
lLHQmIT73nHWvyaPR8HLkD66nMUvDA+SAkxAQG1DXzDIZZbMjRnHkUrDU9mLsMDwabIvpIRVdaau
/H8vNO9AhmFxYeMZXxDvxkZmEpTIzGyBYaVci32gCsbjRuVgA4wRMZER6Csx5r8QNHT70d5PTXgb
DRIclmEqtJmNs59GiakRfXCBVgneGqKzl56qufrIxydbEoP9bDqx09v3rQaBCzERmzHntB8I4F6l
RT4iGAXng3ZIvDoOriJhX1FzteRHb107Tw7LD6WRnf9sdgjqpUHqmxPTYm/Mi1Az1bqtQeH/6Lj5
3tMtDG70FE6oFnknw+StCHn4QywJnbwhfmK/VNYRLClq8+GUVMT/bk3dUOSf2VP98KlLIcajIA3z
TBA+QsWmSHJMKl6BZdkjN4UZuhok8W5SVaFCZ5ui2VRR0jAC/isCUJQSNEj9xGPEAvWoxPw5KXsL
6VhT4SVYHEgNVROcc85ZgocqxAyD2Ri2TMor2Hstf1oE8mKAXQu28rGYDhQ4c4wg9A41DDEJbuXa
UCg6eFj94Oh6OKZP+NVYd9Ri6g72V9qcma4B+V4x97FPiCPOi/V0Ks6kyty/R9oTAJDJGow1MYRv
P1GLZcsA0k9KX2SZQm/3MG4oZlNfiYCtaqHcwncC7nc2VUMLPb1ViVq6wmPUIAD/8ISG9ZRTu6U5
Oy3EvG4Q0WswyD0fsBrmRZxYWvVQnUMOQaHQORA0LtXNLTyws3qxlwA2RmJRGtZXU4oU6xPe5Yrk
qZQfHuLfG7r8hjL/QOi0SSMbfTumVyigkk7iBX/BoriHY/hohLBmHwtNdfse9Fyx47Pk4SIoeS/x
pYRmeKR2yWqcH4MpOuuMGf3VlU8aLUqiZjxYVkNlVQqKv8EWB4LthOJwyB7Zktt5mWZI7Jq7rw/j
ZcR2ida0arTYvCLVugx+7C4Ku0Ilg+59wvekLHGFnhvvZE4ZwPCvc9zn3h0YBfV3SEcJc2Eld53t
Ea2k+ZaHzRTu99BCafwmWIUQ6DRWei9D8QtgbYTT/l+MlkQL2d0p3Az/7DJ3bqWGksI5sVy1OaBm
ShmLS1fELHxx/Q7YJbdpw9eVTEAsbSwdgfxuvJwcRG2wKkntBsJYs2ElcDQwvW/apa2U9BQsqZI4
CLbKFrN0Ws+XnNbLzYMwNMWEiza2jl+FeI03sjte8kXZ/WyWClL19Acq5xaUy/LhA/IHkB9sNeVd
fCS1pd3dU0R7ffCxPiujs+Q13g5Ds0HbxMjfjb3UmGag/xb47dzfxuwoS1fy8OwP2Ip5Y9IApIYa
LrS5wjMzjyem7PdDVS2CALn6T/BENhupnyV/tB3XpDqfIRb85Hps/sLiBErzXR7vXN0KbivyypJz
cMQ3HBigEgVTuzziZGL9HIM/hN17HA/QuEPKRLCMWbppUJE5vUHXL+M/583Y/KMpyYHZve6FuFNS
EWQOdR1AcHonrNDc0nt2eQBVJ1Men/W4fm1N+wWx7EnTceusLmjYaSl1lf7zzSqWHlLHzDCBoJR9
59s28EpLaUMq21j18bgt2uBF0/kUfavFKCpmUmtSYecu/fmiGPI5VY4rLldcgSmJfiwfNcxGiVpE
phWrmieRBTKKMlHMzveNsqpr+h7tKDadSnLdrbF5ILFc92eDBys5qrcNGaPwKnoQjbg2eKeDdfWL
MMAd1agW4Kp1sguiwSpFJl7yTkQXMYI7uUJf6Dq7w07eo0gbhVWDJhqbpkL3ctcWLCzIzXl1ByRc
ZmNW7EhAFlgwvRwVeiQp5aSUo8ajPzt02xzuDGl0cWU9LeC++JKEvzhOGq7NY+eDOmpF7H1m7Sty
OUcI7aNB6QR668M1P/vFKx0l6iB/6xjmWgKC1DPW58DnDE9MbAb2v2lC7E31H4Llrc4fGi3N8M41
KET4v4scdFz22i3w9eXNxF/wagVufe74uXX4nhEgto1SkmERkVcWTL0eosGo254FjK9FNtIz+ARa
oxMKAMacyW5D8g8RqEr1u7Ep35eCygiZFQktJHQrbNdznPgbug8IEavx+0L6diMTqDafYkbvehYX
+2oksxq0zggUIu5pWItuQKm9jcw6+0/37rHtzBqie78uxjP/APOXfFP/7NDmk2oSF2JOW98DwUHK
sq2wLgygI2iLYCFfAYuJf6x4KXOQkly6FHssr/V1l5IXs6fGIpSWxOlN4Pz0HtTGvJ/ZWKUP+847
L9Ix146/cfRIaBbPfHbXIZwL+fsJL5e5j2WOGyFdkpvEYLYQ/4kzJ3PY/dnnj+/qAoqxjumoYA+/
sl+/r5grUDzvxWX9t7eO/3fqtL3DyYcjgHusxFRS8hvJQCIHO+KbenSOAVg+ADpI9RSqoEif+XuA
W39IUjKfg7lrZpmk7bDMymw0AC+xh4R2Xxob8zDDMrzM4I/s2+v9Sa722iCE3L4wt9wmNXqyl3mc
zMh4pybmWVGojZSMj/PFVKcN2lTvDbBw5RmL4T0ADYsQ7S6ksNT9cNJGHc17tdljUvhZL5HjiN+F
2Y/GghoLtFlf2T0llgt7JyG49OuQ3O3/Xhy1iUW1ytHtJMx8onpiqUASBhJ2tuOhKu/K6l6jXSnd
73Bw8Trsly2f9ormFPifLslvcCXZr4otyVAE/i8uBEB/IBuEG7VQEIM89MrYS548XWBNyjxrAwN7
iG2U7knZvSjjTY+45K6xBXpV+pkMwy4oyF8zq5MPcgwP58CWY8eeL3PeL8llaD76BUe5ZhpZiDL/
xwfuBgTNXx7CZMIBP+4j3f6PtF4lu/JiWMvy5qy/f7eH1hlMlR8iFS9uspCII/2qeAlPqSUqaNpG
98KD5Ga6K/POs13diAOZQn+X9AcEAYZE3017uBcu5ueAUr+9hGJlaDord9vqztg0b3dD2r/qRM/u
AolZJFI+4aTvWbnjnhRL+jczdLqo0SBiPuqafB82dnh2hydxKs2qXqQDBYk9wNsa0fFkXMNY7Rpn
ftM8+EIPccBffZ9op89Gt97KqmoKxummZPAKKEHt8m8TuaOy0EM3HZ7mROfyNCipUqHsOPTSTWxp
0Td3Ccr5G1b8bmJeXJeleq0C3mWnqB8ecpHvAHw/snrYUXIcDmeL2pHddP0Hakc+cKFwjaifLnP4
NNQSxiFtKX9j5S3CfntC/sHKLPqJ0PtFhl3cl3SjELF9qY2Usj1XRBIfqD+bWGjOhGai1ThyhyPu
Jg60EEuJlj7FfTj/6p9pXWQtVcJjFD2m8suiq5M3g7iiKq6E8VAOVHiDI8schJ4wXl9BfUAUch6n
rHQanYF9gUe4KoCd+g2zb20zGOwwqWuZ9TE7mUNcFnFki42Z9Lv7ZOuEZov2GVLWwPCKmUMNwEHo
PL05WCOf/iAOmQZWah0W9LVEeoSfvtoKwFDlHCEf3ZNI2H5McW47R5oxo7i+yJaqXAPtM6Gw0q9z
sGMXM18ZB87Fg+YPbftwGLKVpfRwQkgEfDHCeU/L8llaB+9J4K6ppRmgF0GHhw6TXHXHwgDLDhqo
ny7iNU29gIDbiPXwOIdU5ZmcBiR08Wte5OV0ptptx12m9ZQVqcuqTHgsuNoTi5GjSD0BvTAV3kAe
fa452C8fcyWs6122w99j3XlDVdbNiJquTkWzdyuYnJKlMmFY3ws/lSqhNXyvY5zjjKcPJuRaThFW
P9mRkAVRNZRdr82tR+hH97NWGsIVMkIXAVyUZk2Dk6/inczxrp5/Nc6Ld4CsE/vW4QXmhK1rxmYU
2UQ22XSfprb0JpqlW9CO+oMSPYeO2fH/Xi2ZVhvUjPpirnEj6JRDJVoCWeMzGpRZKJdyg2lPuZ7p
5fw9sWaTXU+Plo36lIJyd12O2Kvyx11lChvlOE4c1wSkWI9qPW7lAEYwX5FD9X81jvgwvf8xKUfn
Fz+nLrgYRC4m6FJqyOjLfzzTAOdKKBgznvRXcst1O06sA1UshMId0yArudwg3J2wfVBqakE0DlY4
Dpd/rvqDZh6kguvNE716kt08g0Ovlh9Zb8agj3Aej8XvEGWH2jOXkWNgCxJWngIITvS87FOsU3X5
CFRTD39XDdx7BYXK6nlA8mbG76o9t6G8f3MBQhTv6owkjVKEIEu6S7fsPE5y6PVw5xSeleip8TSw
HoVHura11pO4qNbUnCJJ/WHMKfjLyUBCuriV/2qSx64n0cfh0HqT9fUEUGZSUF7SPjo0huNAXtDW
NHdwK8O/yItaFHMCwUSZl5iNPF+h+wVhXXUnOyb+TR1BXLLp1aLZE2YOz/d3FiB90mrLUOTba8hv
mCCc9WF0+iPOBbug1QPnlQFzKbPO0n8qWUot4enjyaOMqKwaqxaIcEe5KXcXjdb8z5ot3AybZSIg
kK2+lEFMMUBmEXSaCcfmutCJt7/A7zuLQWXK8Vw31I4RPCgFU7qlDOeJQicU4W6L7cSjZ40ZUSfs
BMV6qcMaSz4TrRarOeUg+OBYZzJF0Jt6ELdGDsowsaFmkus3HzeprkN6QRtOOtgrwMtU4vCNNcpX
pzFdGmZHBn0IqGZR3fuINyPZU3shBqUfyY8qhF4c0YsTYHm37fkha+auwrcmtVjEt2qrbz1ZUl27
jnNDNGCf7x61ob2KiFAcwp7mECAi9B+2uTm44FmGJ0RjAnFiYew7v9XjrB6rqSQF+vIcTiL2c+OU
VusxhjvohBmtCySNsxasSN6mgnkFxDKAGX0gtx+8Kz0+G5cWiGo0l/0IuQkNr4WsrvNSLks5KfLC
+NyRQUbkZXoPww4H4WPZvR1JVoGeVqmtELJLwmPm6cymjiX8N9e9xXv8H/ejJY5gIS4+ack6RZEj
084i8nuC1JAY0he56IAShz/5eEm19BUO/aBBZLYM1IEXWva5RZmAEgDIjMF7kKG9aPC02nsr30Ve
BO0L8ZL6NKfr3l+tXa1iRfj2RtTttIzS1vp8aGgvoVdodBY1J9N9lVmR4pljGqPF3jrhli4tLtPT
ep2A1ey8CxDcGqmiOV8N88fUenxXjRFGre46WM1dd65sLBDtknPBcXZLMWuokDmaFyTTR0LYcSrO
36PXfltSUjRsD0mOh3zoaU8B/BcQoxL2P0rUwXiqoLmq3vKT01EGA4FDI3V8t5n2rX5p4BlJtmy0
CWNcR9f40UFAG2WzHX+Xy1JW0fza0ebwgeKvSXgm3vpq/bj+STLL5qJihVXLowArfaTcFfYtOoZR
inNQl3MugoeiUaGY9rgv/DwGDr6Bz5yWIFwlogwzBtcEVUv0Mgz46/SHTvRw2qy1QBjtgHkLafhi
My3U2ec41HDrqItE0C6rP0VfRN+QwMWIwI3eF1yxPOCDNWB/ao4Z5dHqGbnTy/ixhjWCcYAzDJOX
IUoG1NOA4s6U09qgx43rFNSE5GvZGJowxvor1Gs5Fhf7jQs60asa6hZKSf6o2L15+WUSrAzg1s5S
4qR9fiXv3Mi0sS7VAN/SN0nzAy4hWLNaAZiACh/DjnlJmNhjHCWmKvKLHxPNXOmxHGHwxgHQknT1
CQ1fn8XzwYYnTopkUf4SuYVLffQlNVkv7XLZtFMR5qXgmM6QhwSFodX1h81COcKXo3gzMt+XRidh
gBZ2wqhib+9qD48G63gQPN+asiBIli3ktOVjy1QglU/wgI98pLP3lACevQIF3h6WmyEC2jbYqGhY
MA==
`protect end_protected
