-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SelB/tKQUSAWK6J3zNcsq23kLKxsdJFEKyKPX/5xlwZWZMRG5m4AXSZb1L6jy9c+tziBT6t15K6C
0bPmQ09Xg/Y5PG/GSF8C6+dlVwm7uHdCw3VlMFkOOSHqdzrhV5OrbZ+73l9saqc0QZ+tSZ71zVOY
g1lOcdqh6/jknNanLSEoRvz3YrQsV2OnySwVULE0hGRH2mBhfK2/cyA5aC4sLdem2LZ459iOmyzx
bcOdpdk0wLhJSHVaQ7bgQFHKlosSQO1yEiDPZp8LoIV35J8sL8D33k9NIkW8Vf7yAy2WtqqwhtnM
aIZ1zVsgivxW6bPYGXc61ZQ5q//BpVv71MXnHg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
hmouwSmacDyEo1ECSDvGsHGWtrGy0LXVSkFTgpn0Cwb7UeN151gsAWsgaTuIDA8SF/2crzbJfsQ8
NbN+jcSDwjt/rjQv8qDguQG6v6jpnUmrybGvSgZmPWgRckTMsHD335w01fUFigfNRVawehr3vDac
VqcJGNQtUQb+a10acbuiNTW84CKZyMe9Nnu70Ucs6XZJYRElxyKs6iH9ujvMd028uHE25JU3M8j5
+QnokD6GC2Ej6kxNlV6H6Ubz8SJX5QtiObE3Tym+1+5U0UCG6H30D4tTKP8AC+dJ9JMWQI2jYWgr
Y5IOLxsEnLKD5yRvOfD1T/6K+oSHIW8OJ91HGRCr/eF1hNvfL8wqEjWL87v03aHVc1RFGdoMHeGo
royzawbLEX4wQeF3JyDHEtkSkaeQZN/UL/tGF4Y7cDtWE/6au7Rehue9qFnyt7lAw2mfvCnJzLVt
vZwK5Stms3mitJD4RRKdogoDeUYPW3bt5i7SCyWfkalKbfXTQMIqQZwxBnuIV3OLb2IOwl93udwf
VV8mmQyG6UwsyUbZNZ340GPXMLtsdZM/0pkcbJDBr4Hi1UeM64U2SOfBVlysKzjfsbm7EWxwlCnM
/hV265yRuiz93DtdK9yVvZrfU9UWPF8ukwoKFYKx5li/OaDQP2UEuv0oC9oY4rlRCg53KiC0lejj
LiU9xQkMYcBSSD1JTGLiYjCKxvZro5WviaD4gRRPo7rbVaM26+yVt6K+mwepNgiQae+xSa1yrba1
eYPkDVUphxVn4WsmhI8DhRHYu5FWjEXApMyp8dn4RBOyBtmYkHmry+oZLb31IfFQ6dg1Lz9qhZNL
4RfSnbM36F5POy8LnCTX6C3GRu+OJJ5TQ8z7pB6b+KcIkP9PGJBEErgIZ/oz/NeiAla9PqX6QPgW
dVRplKvaybJX26lYo6fuVoLAhIwNMjqvj6dZtvVaBpWiXjCklyl2923znR5WvDUQjzR/q9ucQ1ht
P2b1wSJ6F7N8VHGsnQfCJ1yqSCnU6EIIC6uVCafo8Z/KM7Nd+/MFtrl02lXSJ+FnZiLlbg3dndUX
ohQIWWXv+a/gf8f6Om2krEpDkuovrbb9zPx9ep+19NtzGR+MHiP1PcIScYVVQj80VtorV4894qB9
jnGVSboaDHu3ZWHDPyuOQy64/+r6jyw5L744LXrYehOqZsnKQsRB3EBfuwGgTra+xFdRaTku0cVn
qW61xxfwn0GW45R7wFO7oEcT3GOi13M0IhH+26XtQQCoipbzhVBXS/M/vQoqknsUi5D3g4V7IkxM
FoBIFh43xeJzuw0S7Jm16llek1UmejZqoacQ4rQl4J7KSdVcaDeZkAoO+nWLcL7uVbHhmOnWr+QP
QtonfUZyb7n1Bcep9OMrjSUfRp579mMC34jyBJzqHRj53HpUuTxjpic4StBaPXenw5TUin1GRh3k
QKLaQhEnReZRX5V8efvw3+p+LIYcJR3s3jFg5Ya6DFU85mxiBiKDwU7JPqLzc6ThMSH3zBZLamfh
SgFqt9Ph5ZWIvui8H+SBjXqyg7oOSB0oNRKSeWJG2Ui4ykgbL0wsqJAngUAP6iCM4OtFJdappolv
Hcf6CtjD7y2c1up2T3CC3YbW6N8KyVamVM99vHG40g0WLkk7C45bX6Ue2gfONzaNPX0JTo1hhL/B
VUubH6CQK9QoRECVhfhX6AM6DVztIJjeyIZQ4tRgi8Bmueq9z/8aBBLupOqlflmXHtmHvEoRP7Cm
MZifP7dr1GLDuicbcEkgsQM49xvpVrGwFwc/NaEuzZR0ZmLs2BrCtoPrl/nqiJrDvF1VGkeXouse
khP1pWhWf8l6ntKBykm3nwY0QIReX3buV/VSTyOX50SuypK5BnNaOJrCd0ImKPB4fGQviM3YyF74
ulxKcytpNlwh/FD/z0Egzkg8zmz+Nc0PYPUNNdu0EHtzSJ5T1fO41bw7RaawqZko4C7e/qdpj5CL
U79kDhgDlS/2rqF+Os3guDVDitckqgbV1Fed1yfQs2yBpMeIdCCFlm5c9fPYTN6p8eH4sYIZEN4D
ETJMrVFREQ+Gw3NePfEpiuGF1dypbaipfZFC6LQixk+OtVZNDUE8w2aQeihLe2W78Fr68rK5WhUR
Q87WyKLd95NQ9KPKElxufK3/32l6eFBYn4Lg/7s5EsNR7CduxUV2V0TthOI9GFYiA2GmrL4z2WwL
YMH9ZcryExs5RJMkzZbnJucNtP8OPgPhpoVYcWNAHUz6U0PQIzCV+b7NL58xaM1N2PUc6hVKC66h
brpUo1qLoZMU/7oi8gdVXv9nT1pPpFZ1HZmK7rNvfyE1GWraD9GRixRvXz2ISPeYQlCCnEkRe7MF
xmo+JeL4J56DtMb5PrhNS8PyO2K3fHX5CFGoaEhCjiM1MqqvjHm8i+q0qqMzaKGM75yGXsSI03Xr
7FP3hwLXYBIN3vTxTZRBn6MZxUI8u65lNkuKdWmMmXOUNouPHoz9O8RlCt/a0L0Djk8rxqz9vpEZ
j2HpHExt4frnhq3tPrjWgxhbvGDdeyoJKhU6uJuP4xSbZBE3F9KCEeJYqaBQ5C0Y9cIy/Wuo3gAC
JLfwdx+zRQxyJKCEiX/Pn31jJh35TzC9A7ztOwjNyeOj/BXvFW9MMPZf3vhVkLcxNCyPzhAbHtfx
ueEnPFMI7DSzh51P14Ss8B6hShLW56ZaKFkuZOr5GerNiFcXFpcxvalb82Hex/yYCTdpD64viuuv
VT0Ps6ZkiX5dmwEL8PsIAmD5qVqTVv/kWlDUJIbZz/wpyTHhBUgw9017h8U/Zp4slU9pak4higtf
gK+sNR0KMzSMJCRBmQ7ydN6D9InmqQ2MBb76cC7z5BjXKwRM6IzuFnSI/GtX1lPh4jmeA7PLLVd+
j8LeADbu986lgKvY6nGXh/BLD6BA3pVJRWYb9FgWGCJYq+07IAHb15UFCZDBmOXsQwbzUX94eMzZ
qfIZc92/Mh8p9p02FdvIbpi0kpktSCqI60Q/bkQy8YSc1UdrAJwsUl2AQuZ/4ojvmSTy67KJxcl0
PAx1NE5MiDwii7SlcrM7u5vq5zMtWkCL91Q8BOOj+x+lnWCFLLopuGUyEIPTHq+P1o631yMm2D5P
OUPzLAW8hwSZKaKZzBYNqz8gnt+peJyGflZSH1DB6efSmCezCQereGkFCxScElr9z7J4JbEbaljp
OckUonfVlAcf55yGl6zxlgFh9CUrj1baj/0B11P6MaqgtBb/Ysssm75acnnO+t/ZfMXc0KFYCWow
un6/yidUIvSehbG7Yp4F64poADdrpFHvF+b15FA7476LtwwLhySbH/QTa2hNDlaA9+oOaqD2GLmW
EKuA3NpR1721RHftzEz5yu36d8Uf5w6PVVoMcO1iXVixrGf+WO2+6WDeVOJ9tfC90fNQj4goZ1WR
Fla40L1gmEi4Pp8u71JuNGLlkuI/8nHuJrA6BLecwyIpuGHtqnn6IgAL1mq3kMNHz9BnXI1Cucni
kqzsdld+7ESaOUUuLkP8E5C8Qr8mfcCncfJ0Jhq8jAy7F53QcCnCgli+X1vUNd2G9WfxlxCotjV9
PMzJot5JZo4e5C/8v4n5K9I0aZC/9BofeD19BZkgm6M2PzkDwobH4ZII2yRkQrHubZ3MntG0r3Xr
hUzzlDyO+Cjs9bSCznBsWhjfWNktrdsur/0ejhPIsFL9TGNc5jg2YSS2ekBzK2w2NqSVHJsNWbWN
4GQ/0bFApf2Ku3dG+cmRF43bkwKx+MPHl76hqImTUawZYCNNU7h5NwYGJvpxoyhklY+u8VqrlKg7
rdD2SVhh5iQ6b4UkmZ8A2qsSXZ5MX4HzC9hnT7FcfDQagoTSAJXcSAVe/PGlKNR9EFTDS7LIIXf3
iFlUImOgjgAIXcCYaYNiYFZ4x6i+Jw+XwsqoBiHc52NkZmfcUWDAhmBDzwoakNmtMwyf+wXPX81E
WXDi7KiB/EwMPdQVXFv6XjkxdymSVIaKBtM8J/JfgmYrgwME5/fklUkl7te0JGhwCEdAsqdcISuU
hqM0RPCp7FvtFFPTD+J4BR7hpKg+8YZ9aqFRqH5q91geeOAEqiAyjsZX058/yJ40ePY/einKb45G
jbBaRrWWVHUz+EXI6/oW7XQAZYmHhYxNQLIG8/4imOldAYdD2BvTw5qM2OnTsAPcqa3fYx7v0xOe
J79s2h0YP2WM/INlZakzja81whszFyHr0t9M98cKdgOyLs5nezaiA1oDBZ3wNWgH7f38dZcaEVd6
zuUPbDMocFXEjgl+5VIWdFWTZB98399JlwoMeIzPBHaJnzVZMDHnmEHeN3CY+VAwNGDRYoLV2XOU
drSrG9mc4VUbBHBNpUWnTWLK3/YXPP9pBoJhORPumXfcLtktXYcq7P/kAvp1wmi3ZP/6gyGC4g+f
Ork5mEsH8/+EIDvRi0kN4HrHDpAksxcGBDIeqR2aOEnejSL3vuedZCqil7/t6BCm1SPy6ZOA/VhY
ehFSp142G9WohBUe6Ht4c6FTpZRBp69IKuU/aUslQx6ScYuoCxmBMQ5OlDw7hDyA5uhtTZpUsfre
Vif9/cSFXcthrOM2o/FI2/jnpjUMZUFDQMCH6EfELM+ClC1rl3ahfaR72ZUCQ3MY+DpYulHTMsiL
5XWB8GajY8kKhdrXiM1+hESeSeqFmZx261dbntyP0bd9fgx5lR0PMEfOAycpfKR3mGJHsbvYuXxl
AXk4ulz8C2xfh9He/qgBYcnXDAc33UTqa5BDwp6OboM+aF5V9Pdo6p1blORryGUQlllzxQpIxIDW
7YyzKaKs3MkM4U77FReFyD/qf0RaZj4UqPGtDCvjY9DK+y8z7ZANIlar4RiLM3xeXwiXWYh1coYQ
QC0zgm07to6v97Suh3IR2lNPbTCsliX/o0T8WtTbiNdLEJHI8J/W7fpkDSRm7DbwOJQbueJQSyp6
hUAy3vuHXqa6ZedL2PUNT9RGdcEIdhqhSh04rrJe3fIM7adriQNBxgUV+QMfN4ptFxuEwVA+jqvS
z/WKCJVQWC9DGDmpl8lwmIpKaojlXJaXzvX+8xKmB8uUnPnHh31Lwwe/Xu707u+R1ZV3kK90YM0h
blzmPTPx29oWzAA7a/VjkMrNJiQqQQ8Wso197eRJVuRLOwobb/q2ULCm6vOzT3DTIjUYAPG2ik5s
Jgrm1wvucaBR1/19PClA4Pd2imApoMoFabQ0d9r3/SyB5ujuVDxyijFS6TBLIIG1cO73lEDA1+cs
jKDfwgVrEfbM/zD1g4mLhR9GwBWtz+htSriPuMlg4OIyNsfJM9QX1zC+Pq/JKbV1QMi5RRsPWRob
8rvMMlHc1eyIGYGZo0TmogpwNi6/vXV0ghQ+2uIx/1wikAppS55xYhL3tI3nJbbSCnIPVEYh1Pm+
WWDn2xzOw+80BKToQArbaDWGxq4GlMgD8o4fM8YmJWGJ52LYxLGAI1jeogqhSybqgPOibucmEC4M
Iokjgh62XSdoaSbNqxXgFL6g11GKN5A8GjomnNKgT37bC8MIlX1Ft2FXET5AzNILMi2f5xy6rUVe
b+NmgEdVcIesB7ORPdc5oFCBPrNcns6SnmvHYP9+e7swhTqmbsEIkh9t94VJ2k/M/vHLFFE/DRDT
kQphLavB3JcEb/xqVI4keIl/72IdJZ2diWnclPVN5QnpWMEscbi8gdCfBfMx9QpbfFePzXpDFHL2
bX+Sk4HUl2B0cpKamcD7pApnMAeRMtsKs9Byfxi2OEE94QnMPBt87NaoPos68lqHmdKd2yakUx5q
rW7Ss988tryfu6dTi8sp85t1E+wRvkxnuIjdXjIuW30bgzJGvcRWVp8FuejCYqEhKpkFOBTZHu3/
91KSlbbgziIyS78RirKTCTLLpE1KgJHNBsvHmVBDuoyXpOtSmwlofhI40NfVGVjqZiazG2/N1mGS
jUXh2EKcOKke09w+S8xEVjJ5+peP/MHPgxwjyqqKJHCFAhuIwpabl4w+zCIMwmzIorvwgVf/Hxty
jv6wKxH3bHKEqjXc3bUNImy7oCe5FOzedLbGsn3eoaYSEawtc1Pclk6o5K7z+LisOuSkaclexFPE
xHoiIc16aUxTfh5NUZ60y/sg85MHTmvn1kb00nfmq7OFnFiegn0qGwBUBIJNxPC9PQzCUQc4l1Q1
7omZbol4xvn3ivcDSts3YW3t90KlcekvV9nJ/PW2oR7xOSJGURtqp4KxKuFfgnTe4do0tFyPZ/Qj
ook8uvCn1v9tKZ0mjG3mFyNv0xZswMTeVvGY+Hks9x2ornNLHgYHmjsMNyzHihFEW7y5Zpez2ns/
b5dbqxCFldZRMfIhBOb2/j/qC8+NndIULuT6VLp5+MZ2RtWURumiBZAzMVW6UcyJvmTD9FMkAJDH
tbfdKyz4MtnGGA5YD267KffgwhQnHol8svUqzoinpj0zFEQBSr3y0s8NRfmWL6GTzPhrvDyhBh1/
jocXEde5Xwht+XDQPMKlq1qxP8GQSpGDoXzxN/cEzER4jAnNKw2ISGYDimDOckEQFmlmejm6G3VX
1dmcvocSxc3J6YRxNNqrQ0cLfXDmGj2JEPogQ84+Q4uesQeer5a+4BWZiJwhLqvQkZL39/oa9mJ3
+yQDunUhhn2oLauotyEspAm1ztFmIDuKnkIFsar+D3327h3GktcQR4J014G6e+dzLvVVssghrGMf
PTc0o3jgCklhG6WvdPedGelD/xvw1Ka190idevzDBXxy70Xst7kof1rJw2aJJQJhJirBo9CRgH3s
OgURfKtFmcScQybHA5mSNP3oUvl6VX/ezdXOTb8W4/blNXTp3qYaQA6la+26L1hZAU5Qk1M9a5pG
LLySiM2An1slmRQsxzM4Pb9yiU5Z91/sFN3/EKvJRxdf03tvgPlv45oWk/fGMdDPOskTUte9Reti
eFT12F2NOXkuHBZ9j5jbQaBAPZh7gTv7oh0KywHvRndh2KRsoT0GZng/RFsTz7zr6dI+45rQZN4g
OXtO/JIa/JdMDt1izPUOoRtfG0XO3Ovny+BzibtiQtEPxPw3auWmdYXPLInocFNyQ67NdplqokPJ
9kQrnRa4eZECjb0Ek1JxcS1TgaivJmStrg+MnHVHjwNOw2XXQkjDXL4PvoOEaVJb9R2DnoB7HOEJ
okcNMnzhrtGwNa8W4qf1xZESL90WUjosT5nwLCr9xbdN8DC5ov7QMWiquI4+jOIaCONT/7aDfRCM
t1famk5p5d/mjSvrbYUr3gsyNGkcIBVd4MbkR6kWZAsPbJM9UvTPbVwizJ62ZnGhxwrF3IvvayUc
LizF4bCJfutAaqFq0dIqiC2PIVScKIPbQS/9vQtZAtBLVmhz4oCKgrzhHMpLYQE/4RrNxXyPskeM
T3Fzx45/LZbwIKVldPW86LuxI1AAO0xfA1WEvpVrr/5OIxPhwwxj3kshvkKTvZbcy0TEOAFPixZ9
h6i5PM7L/vsm29zxZ68zL6tox3CW4p0cIliq3AE961BL7RBTsh08rzRNteaXkDUdTw3JPiDZ3y4y
fW47JUjZF1N+yU2CjfqVoCiTItnl0fTcnRFoe4L4uo4fZdHDkiK1mXdyaId8Eyr9JvzgDOGWvFie
qc5BwcYTR/0gcj0xEVgw9B2pLWSHYF5dBHlDkiUwzI5zsdZbHNpD4tNwR4ndFjqpmj0xX2A6pubL
97RrGDtTCvsGy29/QhLiPqGGkd+0d6uty4xXsnyKMsEEM1GdqyKAHjrr0WVHvRd1bqww+K6rVOzN
p67An0MCZrM4LmKVzZM+YNXDDATwoWpt5cSiF3Q+tOhVmTZANPu5Twq1oZYi7HaXoq0Ft8R3F38H
DIxOV48JbyneY7Eu2pau9+mupxSPsa2AvlmTI8EOtZJ7ciDjOjm0gXznlQWmyPuARNl8olrHt9U7
iv/L/EBI7QFjPtCMAPJDZBQJkLSO4WN8Le2CErl9gtHHy7x8N/cGCcMMGuysd5sp30R68ZK9JzwW
8pqfOZ2zlZYuhTmO5PlRdJ24Z6K9cMm3Iemyv316/ivZcSyamiEpSfQ8hdU9kU+8uzCq2OBzNYzx
9egDvJKmKR1Udr3YLIj6N5lc8e1CpOWbUjh24ujqEreib/HaUqVgjdMkexsqiu+Tzoinup3KokK1
MqMGvqaaBbRoU7KoscJ8aflmoH6uhtI/S2yru2JyXnUh+JiSe8oLSalM0Odb8UDvSYp/ap2OoBwn
rnm6eez1q2Z8wKf/e7czCf24fSDpnk+EZ+iKWI9nuOL4f719ZPZxCF2YN+PaTKrXh9BPmjqA6o3c
UgDjB4mfO8Av9Q+HhqC7PW1B343fK/amK5AT2u+B2zdw/bM+wfTluhWXL5/kwh2xo9EyacgaUWZb
+EKnt5809sWVAtjq2LPEgq5AbeOeYEwBXQMl0srICM1ykxxaQemj2atwvkDVAWnAjFNiUuIj8YSg
koSVdMSEusqhATDdzLjj9SR7OExqEJ0Or6BJz/ehJ+b17yhgale2WFko0pvptWhhIc4ppCjtFLQn
c4hPBFtgEUZx7be4B3i7EhoUr2ffU4C/e1nT/eW0xVmC9JQiyaa6BOlLN0pCyKgX+mn5+eUt99f+
hqklEYU+vj+hN1YT8iTFpz1Ek4zhbHaNLpbiy8fCPZDJdzVR9fi/0hf3qcAkbBKLK0Zm5/9jxtcA
s1Mi167+WI4LE+mZWnep6bsexZijN6ZdfKdsQ5+B72JqWiDpiQAzkRfrQMDoZLx57NdeLGZY3czd
+X/2Sl+PTHvWn8Y+W8fcPtvhs8vGDbm9YPGGHkX4MJDmhkm2ff3D0Mo0sX2e/xtrN/hchQzw/zy6
DzlIxO6FTFnbiKGrYA64lvd+RJ7JOzk2x9kwAejYiLRMpYU/3jvm7F0Szcnrz4XXcRSER9GlZxe1
8fUJvT3esJFRTbX1KLRSvQfgWstLhm8G2vQT52ptw7985UA2diJ4nKH3JS+gzZKLV3KQgcPAcpS6
xsXR9RGxAfBY4vAzBX1YVFyMHCg6xndpPW8Baz6waTdJ6+GsSXenM/uORx14GbUvnnS7eksej+Ep
c7QiyRlH2+RrT7hUx05ktwsegGm+J131WpRBlSCnuifLhW7iw3UadlN6WiyPj81an7a7XWH/g7z8
+lTByOvlDvUTA7Js5FDXHHs2w8YZjb1BC30thBNguqlJyrXS5bRMmZijlwPZZB6FkFqvPpdKnRkT
Y/vTHSMn/sJhVBqMDpVYuM9s3DcoAwcB9l6aRo9EQs2abSwOxRsWMriAlMxJljLLiQLhR6bwJaRX
EF9mFaH2jTrgTiZRM8R9k7qe5XtOC60v19XhD3clwFpon1hRbuQ0ifUF1S5XaIZoZnp0S+ctxeys
D2hMrN7gjHgMDRcIP5yvS62yEestjsRdtuIYCD3LK40E06Y50Fvm4tqXV2BodTM9/u8/4AhFp0Tv
AWe4JVopWDSXwyhAwHXrPLOFwG1rHIqtDPqMbHlFEyzOX+w0igQ7tVLNArBqVwZ83Nq0p+nVtOqw
SIgQFklY6hWBsVKHhLBn5HLros1138o5w0X0DFL3QVADxMf7VgrTaWvkJXGldN4T+CMeZ21qwjQa
Pu+S2s5aJ8bxnL1Bxn52lUtXesdaHV/TMuxfT1ka95sF2NrQ6KaXuGCNtifmyjAXvtQWCCl8BJzH
JZJK+MO4Tt27LuodKzRgIL3CBD1KlqxYvlFjk6yrWWYXkCxn6Em85Wsn/y0QkLZ77kHdBBnRzYKu
qqFB0LkMo+45e09atDx1wD9WYlO6easNF37JFE+2Abazpy3AKmS7D1Zo/Cd8bbC/WsqzoVFxazOv
bBIjYH+7hwGkLE33GMCMyiSyi5u9d/FFhSxTlL+6vvrWLEpoFg9hdXDkH2zK18ri7Rjhiko8jxcE
uqPlSL8HjN5j2R7L3YBT8Ix8gRB5O8H6efAMcMsmoE37yQzeeZyyfSq78g4RR9S4AQyJ8zzdzwGv
1ZMXdESQVaZc28roJKozzbQJeZa6tV7/LwlgMNrcInEi0dtV3wm6t7Zb7IRjP6KrjSoyj49Xwk8E
a562FFntp1QxBpFqGJnwQeQITWLaPiVTtkf2nDc78m1owTuKBvsRpZVRKijgk4EZF8dxZv/2IOmO
VyNFLaB6RFMpE5fZtF1LhmvlIIN+8lGOaUoilSL0RxhbDuOzLh5ioS6C1nFedpjSS4fKSEveWbnB
SlptXAcPy3exOJBbTqVLltjZiap6qs7ibJuStUlRHuGyYPeDuTim3UErjjWEaEFXTTK3kEfNPxNB
fk1guaCU6IEHT6oEzmX0e382nhPcJ8yj52HliUWMjDlYv9g7srN1gWF12uscLNR3i82KyAPrX5bO
I7fG6EFxGvXI5hWsxBNeGexOD6BRvii4A6ELeTqBAf/QXJQNI6b4ftDfJ21iefvhlg1E25AjFw5X
whLxod4TpIpnpBHpaZc5WL6jxZ4Kq0iCxtRAJal0cgXUl1TrnpNN/KrO0+4/Q/8cH/JKQger+iXc
FsGiDiyDFk4x4UMcIiJ+TUawvRgxF8C/FhovIbY719YAC00IK2blfpV9oQRqZGCQo+Sk45Qq6VrV
cShKvNfcnunO9NC13G7qHq2l56X6LDkV5x9IAM5qAy2cgfCc5U5umpUDDuCGEbRwFguR84uVThMN
tsidN9rv2TAiriEESFoqpVXbv4+UNSGGUx49+UYOLghuClvtU1RONxPeTfwTHoUU4lF4fdcvNrJm
sKPy0d8Jams2xdFORJVIC+nGBiGTIvBoXw5pWyPHVqZ5tKf3LxNJp4tMoF0L2K1R37lqtJVrsi8t
3dzbpkqKBk0RpnWhGuizU8wlDDZjfUPnVHCigKzjj0puY3+hLGz4zlH+UC1RpXrlZI8HUY40sfKu
BDEhTkkist5xCeseyeBiIy0sJo+n+0j8wLA64a48O0Bqe476xkdFtMMCwRf/UMZwOTLBX2H4UyIU
sUl7Fu8HbTEcD35JmqyyKfhO/AuMJIWqd8nGhVrlDgzglP9OOTbL1PakeDBGETh4KqydG7bMAJnI
WaLKbVVH1L+weuwV9PrdtuqUcej69B/LACMcF/3FLPYLlaUjE2y+Ue0j3cQry+8QnAXd/8Pmv2t9
AF52z4qtl1QOs8VPMmhqefH4gcHapW15ufm9SHxKN9b5cobjjF4SsJHHgcSw/p4xw4HSGen4gu+i
Dwh6PGt3JMvnMlsc4Azixi3u6nrMJ0YWkMGdM2+KAC54Gxo2VMv/JgAxvUlUGfgMdLL9tICBnZap
9F8IY/pEMPfitESv4NADhv+vBy6jrA8gefF2bIYOnIGJQmwwmbOtCo0IcABGESXQjNYh2KlyNkze
rk7GewgFUx9FQERIlPN/5URqxiSBcsg/rVcWHe79e65yboGYTldxt1G8+kN5D92pi8+DyktxWH3/
cpLFjPVua3q1LxphL2rgCKW7draS8traz7Iv/J5sM/ImbfpLMLPld/zYKqoUGAnywLpnNNxZIJEf
yKDDQVwvb/7JYz3anwWTJxRPFQShwY7eFU1cXI33/DHRfQVukPxfhpyN1+FKCzuq15+geciQTeXM
9yCXc3GZaUdpdUA6v1UPk4hfn+v+NDq1NdpegZV4Pa50OuLV+3oRBv1JfhveDNXCtByseg+qWVeU
DgWZ22wVw7DiL/tqbb77iKBoSXKHVSpeMmZLyj96aw963tdoMEGZi8+SmgdP5vXHOjo2VrhMlgdb
0B0VenXlB9X8JP5lxAuxP7UQSUzSZo9KHnwwsPIWy3x2pg0NHTwrFB18CaHPMEoNGyQHnuM7P8bm
dDuTOA6lY+8znLCB+Z7s2/wD54cEj555TGVcim4zHGaoNVufSqy/Zt4Ak2iFFtLrRGpcYbdxSVSk
eYE/+vbwMakXupMgAcw2Di0pxOYs1qEQJIz7GifMxVdayOco69m1RqbiIaUQNAWjaXW0g0Wg8H7Z
z2Dvu/EvGGTqaF7QOxJELqSTGuU7ySUSIhwxtTzkRF8tbJPK8X3e/6U8tGVI325Axe/MsZ0NThdy
kj+pzbaxBIKXCMUl+ZVtLdb90ftGHXNkBUuWyafSZZsie1vvTnbOsyhPNmu3ktzYLM2U3lkfVHH5
y6T8Vdjpzq8zr5PRH3KCI1TZQ+TzQadtVqGzVxoSEpF/ohjwyGHjRzguOxkos+jWDme2YoU+JRbe
253AEhscsa+UNFl/ThgtLtfzWX/CyJSuK0Qp8x7fK/6G5MjUyTQgw7yc+BZbI/ZXuIHQp3cjDbq3
G5AHrapwRpr7ryTYcRd7PCAIgPLu9G6IN5OLq5m5lmc2kWP3HInU4gR5pYKPCQjEZFpEMVA2vs9O
yFqtBzXKWnTEbOjkKYaYJo5dlXJeYUW/NdqblMxHnqjqI0PJoEG6X1gkOuBtnGKLETCMVjZydg0g
NbH+njsfMOGjPfbNgGR3zXzB2+DlijdSix3Lby9gQbeJoNh0Dw0sGtbhY5HAxs4O3Ej1MRAVwHwv
fMz6GU9W3VifiaNRaFF5w6P9sUMiK07cFiro5q2L5baLdXYZsDFW1O+PUdaB8VfCcFqOrv8C7fjB
P+AmpGqb00D+zkUA/eF5VQyF3Dx6Xj4sCZiVeuZJBrL4R16W2odu5G9qnUXW/GOrHVGaZ3wbHFkA
FzWg1H5mnpZW9zKbchryeMkDm9buVgLzVc1giGjoVc1mYZGGlU9Bz8eqkVHfrfVzxU+rZxiRbG2Z
m2GM7CrnYmCuYnu1f8/ltCVzHr1dGZVBHVyTLkJySGT6635Eq5deL4lUnoj5EOwxlmY52FWmYH8a
DjJ4IKBdOfMEbPyGuIuZwOeugYGGErzut+cJ1rFB/wozjVi1k2PTxTJoymB/xLvGrXIOe5Yoh1GG
CNTqmoDfwLeWWVYYOpFg2yFfn5TCvPfnhztGod1y/nR/Mq33V6+G4IOT0HaBFOLPnYXAI6uuaS+z
Wsbkt6AWSdMZrbiUePN4XVO8H08AhlciI9e0jCmsIsFNjguPruWrw9PblYAt+T8P1L75gMgPV3G3
gJDs1TGTq4at2CO5/nrhZiyV7qfpY8tqmeRjMjCHQm63mlNkZt+NhH8/0uIf0VWmq9Tpdkuq9gU8
4WBYpRkmsMwOZl3MB4Yq8U9TjJJLa6bIg2EhKMKETnd7Z5xXEby5HXOtCFp7mXtLbI0tRX/q3nOV
VS6/QUu+wzMPt3n9P6ghG9H++/p0Vu6/C0Z/aP+UKkvSN+UmQzac5056smUq7+dsIA2vIdLH+1yA
9IllQFlTD4qVUQ0AmYnNnxsQYcLKji7z5kdkNudiundM/lwBH7dJ7GunwyZzndMYvm405qw0t8iT
J3ShAFJSCDgbV4An8SI3XQhhcW5tILADwg/TWObZn154rS/OvXLdHHwc8SSwnPdQpRJzsy4c9ohG
T7rJNUHBP4qzZfXTRTptX0RQ4aLyryYRHd+VCApWKWlS0EXPzK7lOtu69bK9CSaYkwDNqwdNkXnC
0OqMJmpAN2DafcDYcEtc187XAaY+htX5DQfRIsPJcLE1Joc8pGNDPQkNHZ7ZMI1AvncZ+7J2Fjgl
Y+UcPPn49HOHKGYkdpm8eHXMFXBjvDa0/btKsNy3AGxgcJ4GFXLoZdcVquElpnwaA9x/Bbu0u2l/
Yw0w/BBHhwur6LJ0BfavGr5pLgFs6Zr/z9OECJUEbJFT1Z3F2zwXKk1MfN0UPXJYJroBAZLfdpIk
sKLMa2HXkO751+Jmn0A0ysY0s2o4vb/5cYXsLfM970zvJ/ZOuvhtNwlokmK24n3ZTQypYtTZCUgc
8Jr4YUs1oYbnT+EmBZRWvYLNZZLW/3gZqcahMV/1HR0Yjafk74DFxmzWboQzFO9sBMMU3ubT/BP8
H4skye9fhEdq6961ixP3YwrD0+FDjE15MspOYNoqp9SN/KlUZQXXakGZVsaF6CYIIPANcbVdrFWy
EDHUaQLMab8RxkGVv3N24bYLpCYujuAhGRrnClDD4qDwseVIZAJ1sbAmVQS0x8UuDr8SqTG0I2OO
rWGDdUXJLl/FfbDd4r8o0HhjsaLbT7T6okmIuPQOO4fPSdsEEgPlcz9MCIMkg0xQ3pwZimHfLqLs
HgF33nV9cCXQu8B4hpExKy3vDhjlwuN4Sw1Mt4CjYzvJN6ERoehcdyfw3qnliVuPLIUAtGTEWTo6
B9Y0vP6VGlRnWTZaWM1Ou11+ik7W3x5xEX7HrgPOeLnuxSO9UGjNdAwxNSzrUSLL7UIV3gB4+4pO
TF0O5UmxnuSJUmsanHI2MuUL0qrQtKDq/mBjA+Oh58TMX+gYf/ZMbqdR37gD6/6pSTeGv2xfCwv6
gAoNdWJzdWGQGZpMl0TaVvwVzEKcLqb6KSr1258O2+BI2Gv5XwwBCJ0Lup3l2qfMRUpnHSs0j2or
JENfzJN/zvWu1Q0A5k+VSazza6uY40uXoF7NlHOQqI7mApsEr6vXy3D9IiTWZB9Jo5HyJAjuO4Dx
EsYMkNMFxSk1g3UKQsY7lQEsTaN0dJfg3dl2fIldH+q5u6GAjMGHg8jwQonHBZoWNyrDF1TOIwu/
g4VdOhX4PlUxvIDMLFSL/tJGvD01Sq44F0zCfMxQnZwbC7u8pMTENTfqyZcpK+hxi2etT9TVcxVb
mcEUQeFxb2YvZ33c0oIqGVfQeRFxJBK6BtGCzC6et8nLtC2xHsf0lNzqdW1i9WXZbObSAtnSQZ1s
YRy/HR3E8nXjUxxQH3+3xm2n1oEawv3yFQGn4m83fFOx/fj1a3i05sjw8y2P6OtzNDtq4WfBKQ3I
zI0rmZsEImx/KPfMU09tzJSJW1yqCpIZF+8Uad1aHPMBtYj/rx0ieeu3xJOy6/vsaXuVPTRWe37B
kMLe1/Ae7ETCZfShu+WiaoQ0DYTZfE8Z5PgBE+MEVS/p07v3haKoI4TvVHp6cUcFTqbtJdd18GQu
Wn5JdtA7yxAzDzAFrtGOAphrV7ogdgOmPJfj0m/GcQJhb7eHcJ1VcA+2gaOmi3jgWwj/eX3/8iJW
Oc3x0jPL6qw668oQp5qsnYLOP2L6QP+06qbMVAwYr/5wVZuKWvEsuz69F03E5jyJzM+g7zHztfbC
ge6OKq52XpQ2dtUkXW5RYSBDISXVgxhoXlRxoDaaBeG46ZcdNqVJheHkL3H6LO5O4n5xksbJZo8l
owvaXad4y49zruS75yyfo6gm9Y3bRmAcRVDphdjVEiHsVuB0OeHKDg4++9sDucySpPdcvmqd0XQ1
VgdHRCPwBNdVLawovqiLVVnuD7EF8/danCMVyK1psHq6gJsjuDQG38Hnagy1+EInZjB5gxUtp+uw
aMOTyz8Te8iyRHODSjlHlf8VwkNBHVHechQJ49Lzqa6pOgPb9Qg1P/YrMCbUPCpvw7cjduSMBmLm
5jD59oW2JvJE5aLNagV7ji6Lqx0VbQfTahNT+l/F3oh87IY5GtD4gpIaHBXwXG6zxp7DBYLORQLO
o+noLJwFl5+klu0ZsamvmSG75lX2wF5gC4lcwEcLHtnMesKoepgW0fnd6Vrjy4wE5otl/t+RVoD5
kc0eevpuYcCG92Nu2gFyC1xvU/GQoHycmnlx1+JL8pDGLNon8o/S483dwKt+dXSSch7ys+FQ2bDV
IrWznpvCbKpVH5m9bNi03h/swjZiUU2ogmIDlikfkrCL6Ez7bruoHZOUlWTniB3W6kCVbkSN672j
OiJMbg7UgeOtnQMCreO6TdzcCmVnVgU9fmDnfLR1FFUAgTdW0wwDT2HGwUmscHbIRhRBK6oa/gv5
oDCOecLUdFMOtFXbO2h+CRiivvU7mMwzEJjEaLfYlGZUVhPsROFTNwrAliJ8gAkz/r+fN97z0CEt
ct2RzW2QqTp63CImQgVG2pvclYzr97Km0BOqYNcygkpLUAGKLFKQtzyry6SXb4kEvM525xRSGEfx
+6KISViSW1mM6wz6vJIsC839VxxJR6oF+F3rkWz+nW5Y/LtRbqph1OR4RNipavB7sTqSOufZTJmj
dVMeew57L3FF1NuGyTPPs05bEDOjxsCuCy3np1q/5GEYvrtazzuElf8CY7n+YHrsrSTE6nlqISOv
Z8aFuilblAHJSmQvHA7x1m+c4KpK5+8n9p/VTL6GQu/7f5ALt74zlTx0TyRomcyiVTnA+76Yq4JL
MTtHYDu+uiz0r7RDr5l40FsDJswjmcwNjZZNvjw6nAyfZkFCF1QJ4qq+/usrkwuXJYhGEvlBzu6q
ADztEJqlqlMGYFymEWmpgqC7j20C9TpKmYKVkN72OUA4imyu35PopO8dynG70OKhVwojX+V7d/li
p45jGfqpnUmsQ/sFPLjP/iGX3ZJbCVAcnwj/N12wz3IbVA/Tky0ABsRonwOw57uRvEIQkZc4Qt24
Wht2uj9Fgi6vaCbmjp2s/ilWaihzX55x1h/6+476Jpj/+S9nxwPJfa8y2Ps+ZJIsbflpYdUb0T6J
cIGVoCVDffcuKyGP55z18ef6Lb5Cf677fSuDCbiy69Rz8kD6vBukoT2Bu05uJaf1C3O6BUl03/j3
bqowbQicu6pRH++wd+UBhd7WSrHffkRXHiIbkCBB39qgWuu6L8/NTrYFlyqZBTdugG3x7sTOwBX9
VvbtGgY0RCsAPGiytHmTpcWXquXJUOmzW3tfdgbIgfZHI4qSBfgiOVyJb1ZOQdZSJwGnfZu4nR+Y
gIpy3n0ZUi6MtXSYdcxoq+orxsBZpBu/32E/472aGAcLCu0cy230HHFuo7zkPzoI2wdTSDOIf+dr
NWJ3dpXXjEl6Z3Z3DkXI6qwA9Gmn57P7CgKLW3tkVDTDKJHQseV3wh6lJ//SGOu4DPXTpnhJP0jA
rR4YeaNM9pLEwYHPPQ3eLiKQAuAA/LoeApDC3Xqan54LeyxBiS8CuT1wBzrU79St2EnvCCfcrWOc
ovQgT5dRfZYmdZGsqFtquLBTI8LaSGPhulQDRwoX3HfA95wSXFznSzuSfORgia77YspdsD1C2yIQ
dKQt8jIhAkYjHnOxjlvnRlVARZYNDDuz9zi1jxbB8C+/FPNg53yhuHbsDgCfEO6J3mzKRQpneZ9+
XJf4sbUhbgTvYzLUlL0uiZUEGo7k2DdMlfhl5SDEg3FX0mfQRuJVKw/hngb9+X4DpLZHzTiNJQ0F
zuaBB8BxB2AKu8IeSUvECkv2tilPO/EFB7eFjBKPRM0CgRERgRkp3lYBrvRNFpUTn1ZXkPCNEwB5
7uT1spYGj8Z5UTB7bMbPL+YVUqL9jXuzXBrD/GlHexeqDKAs+/1GwRnmHEninMoUyWzZ/0j3MXXd
MPchDJqU3qp563/31SyAO1MMLaicEobJqtJZv9slLNkC/1SwEzNOxUDWeUgQDng9ze4vBzdXUEDc
DkqMWEB8VrA5hNFOwpleub8TgkSi8T8PJA+a7ra8LRqfMbgpVYFBJd9+CL/qeWIo1j5EJrQmjqUQ
hXt9wOqkNpcGGY+gLrbrc2T20Bzv1vymMuYEeU6+RLpE7ro3dCtE1zSKPvynjL9bRCAngOn3vYwq
xlwhBEJ7VzRbM6AVGx1fW3VPcQgliV6RGumE5pF5hTgpM6bftx+SS+TV48QrLweP1kDb8QGzsH5M
/yc8TzJMS9vgpavKVnhYIVPniY+E7aTZaKhC9HsMzknju9dwqDEjpb/jyLzhM+iotwfE9fXb99qp
P5c9Qyc5g5MFswoHJKLSsQ0s7BQtoW5/HSqFHqe9yZwy8rJbaj/sSGaofWux9HFTnksCtg974YQg
xbcKjS2x1+pTrjHX0tv3DIM9hSMDYAgrsiSz1sNb9mXs3VwnkVVpUbQY79KdeZhuu+koY8dNWnfu
5yjpg9VqJ6vbpf3R85+JljZc+4kCO+b3PlfKkalZV2GhOOhNP0Qn7yRj83HM7uIqviTqvV1ILb21
1kfdVhrFqGck5zmY4ufkXyau0v5B7r49SgczTYNx4ENHZbnP7MrOUNIe3hNQr83211OQbk8Yy8JI
s03Q2Q==
`protect end_protected
