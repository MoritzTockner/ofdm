-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0u25Do1Mmb9h8904K8Gi0XVPGmqx/bfCp9mQHfXp3b9NNXs7ItuyHlT0wAPFukBusfO/vL6T1tg1
Si8naPjjtjP3XgsYtySlPcxJfuqs18CuRQGv8q+fn4TJyufOpHzm5lFBh4bu6k8T1TR7Dk1RqkQz
nJoL63ZWpJ7B/zxX8bth6xDAcrDrBQcgk2/nx1q8iLasA/H3j4kWysCyggDTNaZa+YEJP1W9iLvU
Pvw73A1ONiflyVtmKAa0ryDd0sNMFulp02YHgO5CWlXMYXiNJjQlwy0s1A7hod3xW1zF7FHYYIn1
T7wXllftsezJJg3WR86kmj5RtRdZSu/az1xZeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
gj54EBt7l1AuaaTNHmUrMRuJf22u1kIyhhuJOCccCFRozI5sHPOIA2baYwjme/JfBXgSL4RKuR+z
2JjqMj/ncvvWM0XJUfcXwr3pNgFciKAb4PHgFd89Ig/lUHpnQbg7ler6IVKxN9O0DQ4QTRHh9N5W
zLKkZujrJTr36DRq2xzIeJJRNJ7d8frANFTqNl6pSRxFgj3s1SvvJ0uZ1+GtSGuopJc7sN8yBhNY
HOdvQhor0tPK6sb/X5g4PhLxfJeelxdDGhWhtn2dNFccqhnPTPTWHdyA+P7YFn+r0B+9c73zhtEJ
T+xQXgeo0x32gu5RIrnv8LVBj1xOkJPlaWBCWf4R/+a1m0ZVgEN/iNUDJ717hz1ATTsxtDSEZPVC
h8XEX7uwd7VDF9JjZarVqLa5+ABRurtt5Fy6C/ZHQmNpi8MdP4SDbR72QHbjj7pp5mXdPCelW02t
MgWPVURhnphbrZcVWu5nuICd4zwqbFXw8yKPZdV+IKswEGh+YkDAHWrFhcJDonm2V6co61GIhw7R
JUCXEpjP3GmmxiL+qq6mkkfbNUpKDuESnRM8rRRr4vXhex7C2d7BJnbUaJV6Sy4fUU9G9L9KZc4K
BvX1dEKzgXVR2C3f76Sm0iHCGJAWCxZUgaw4EE+G1A1Xa0qLdDHwF60OjmuC796RLkYxQwltoL3G
tgO21ezGOlbEm4MglOi7yel2vuSnp24t6QmKwwd7uer5TR6G7w33uY5zqgdsal/ceYKljDWevS5p
iV69IcLhmm9sW9hNJF1nBH3UTKYklGTmzd+CQ8KyOLg1Tv1fDc4ceGZh2imqwRhRgstzYx7MxPzT
dsL6D8ptUZEd4VZynGZDIBod57ZMNdCMZs0DB7O8GSn7NDn2YElDHE5ByIYAAlRPXkW7Ur9RR/O2
CzBwPvecxMvrxIg6lNytenhww52ROC/p4OrlEAt3u5ETs4ucS/IFmR2DYs7BBdhIRz7E1iUaK171
GIxTVphUdb2rJq+OgYtTFpgOkleAi3Od4k/rIaMf1ET8a9e7dYueqM69qK9I6bN6Y3XpBaDqqFzy
c+ZqJANB69wYRpKTNvLTMl+XC7f2XOyPGxC3sqzaH3tkurxVA9oqny6Nj0nZhR20dZOcyJbzrxqX
fSi8O0SO4PGn3Opaz9CVs0PdfvFn9LmjcRXtGQ7o2BJ0FPnqU7HtTA3BG58RlEKwYHDaBbdrIQVy
Tv3XZdcfWLgX0hjPyNaHrdzANabL9CUFhbe72Q87wuvPrTgLTOVZ7ApIMOUvA6GjbwuqcLgtkWME
nILK1sWL3FSQ8vjpu7VJSsE2QrjF8GsAqmgrAxojpC2L2TYdoW8EMSB6N0pzGV2ee0HZEh1tYb+z
7Hdln9p/7aPpddjnO8nHIs4sBLBngV55T553ZaDWRL9rQDdJXJg9ofrmommn1pERLmYctezpqZkG
wAiRtoIz0DA2PYnlmVR5m76ZeMVWQmVyvwjtAQSskonY1+h8CspNcNcXeXsYczTIG6ddtQpQPVyR
RlqTJWWSJj72RFsBk4FuNnd1FvijcjQZB1Q5IzNBpbsBiXM8QifkEqqKrXzOSdnvJXLXMn91xGHB
iMX6e9r7frxGbHJhAT9BwmCL7GrPhSyE+Ca/aFEvSdGqLSGAlyzHi1WVS95gycdidmqlEfDvNktb
JdNq7RqRB3BUiyXQAUT7vHAWHDmkWtPSyn5Gt5dS3+2im0ewmIyVa1pFsKch9hJwI3Ks4pYn/uZR
dNSjd43B0B7DoWZIXxV0a0H9a42ruHnOPYlxYmv6i1M10inlvt2/Bnzg6ELpymoO3GvyfRRpLg3q
jmRnKWJ+PktZw48e+MEcszvMe+mgtmJDofXQK4soNhbZnPvKNj5jpatw0jRzjVchRpJ6Yzcd4IgX
HNQ6xooPVBtFzklUZFHOX/xjy5zNvqD/pZuPWILQQnn+ClBLMpBS9GBKZapJScS2yKAmTCS9ltGU
SqfsvZJHZifs1qisg1SmmDX8Nrl0J8fcHY7l13lGU0ron7NqAVj/HHpWXwVEOubszLTITv2tLIan
r1UyngFBosZJUN7urA0S/fZ0/VXMC4NY+3SQf8TQOEo3FPv+UBka6WUSM3TCVdVtrbDShqD5NbLo
6ht4ObShn4DCft31BkLu4AxK+y2szz0jZ7qqX8VNnkfTDA87yPC4kIfNEIJlk8Chr/KolOgehgL/
kfGwgngXJ1TWG6is01Pnvtp2gNAQ8zzirrI+rpif4uAZjjOyOBtyNpp8VaF/+sxFtLf8wdR1eG/5
d1lKnis6Rl27cZlaedaN/Eja3xV0vELk2WSRKZvoher5q2dyYq+J5ud+XWjlDBELO1fOqBtRAhak
jF+AMcJXAaxSXDCtaiG1cGN9zeuymv8OnYlk3Halx4/8OOE7mP8/c7ezmhiBMoswO2tP563VImKc
F2olEpbORMlacQ5R8Nl7Crx/DzUcmjd0AsRyolwXW3SBWaCa40yK2EF2CpO+cs8rvAXC391/WQeh
H3IK3nTYqWvyHiOO5/lROTPwmwGglPqXUdezUfk8eBRccrend1ck49yO6Ld34cl/zdYAdG/XK5CL
qC0FBHNRljj4sfY7jhAe0X8gwcqKu2MhepXzCrzuG+o36J4S/oLvqC7C2VFMjC/qIr6tEU82HuNS
8AiEVWriHl0d/mr9f6D8KgzZpzvCsl8msQ8mLks9GlrA7MNHlNc0wDPpcaRElyEMgC1ociJi/E3A
ZCiP0Xc8PHAkQuidd2iKS+RmdXuSl60Io8lloqZRMehPJpAYxFEOzpy1VEw8Mo8p7WKNSmai7EDV
Ta3t6Uv6wKVTTWYtN3UMxgOidmFsIEfHvS05z28T0udGTPAVXMOjf+Ot6/cFbDBmD1t2g2cKoQcy
jOtiqG+VDxG5x5s2AKagLzwMy7Ko8k4Zsrzz8Pg84RbvrrYm6WL/TRrk3SDL8uXeIMo57+BFBL+x
usyqEt5LI6oUShdDPSrhiJiO+35mApMVUjU2UwKZMDeFc+gXkzqCcZQ37dKlmtado+kkQybXCBL3
5mDXg9vCtohg9PnYTtEG1Qatt9WZhXXr7lTbpe5P85uySpIbQJaWKi3dvAH1Nb/mtZf1+GWs19m0
4vWlZYsRRqyahWIEcIRqAs/jHj1cypTvT7zUFLuzUMrrvNRIlVIG5EComoumcFfKi3Y56tjmSNw5
gJY3jBtWcok6se+gRetXexo4fhlNLIn6cEnhu/QE0F43YN5UZJ3ew7G5122uqylw6RtuQKDySD6I
+D1DXqlsqLV5iLtvGya2tcnEX7IWL+QqNxtLi5bl8IDJJQyH8vX+OM9FV2XjqiTXW122NjuJIqIH
I/zxqDUKrUJnBRssOTTFcOwfxEvVyNt6zRUBB987pTxop4rgA/FqeCKzQ7DhpWTz702jZjz5yNKX
W91N4gjiqYqOJAaToohzJ50f2DOLLE2Oz/4DlNBbLL7yBDJOeYJ7p4s47HCFquai6Zr0ozdajyc6
+Qznmpbp/MZKtzmmf5GT9+q8g/hfVtJc+RplO5c9heikWzYqNl+fHj6r95Qlm5qCUYP5HDG0YiOQ
We1NyQW8xRgZjWZlBbI53W0fUHzwtx08l6fTWG9mFaS0Ut/tJVhqkuQlMLiBkwJj6+7TizZh4uoT
PcapzMKWZLz2EVl5DSrWCTRwsK2k9lYoghVirHEmaefnfoWNsxdP+a2mk9+9vkR/e/IqNElNhzmh
C42MbFWUMq2EVBAwFUWSEz1EAfVUAu1sMbUvRnUbb88oaTp4G4cQ9hKIZ0ONokPrbM+VWtCICvlu
n7amWKdNuR3irmul3iY/vcJxUXw3DUYAuUfK/6FZel3drEKeo0/fV0iLRaRvkH6W0/IBTa9Jr5QV
JVDMibPY51hUfZ39pUd7AWutiRn8p8uKLI56fU73FuvgDFVznzpkCEgF75Tv868Ygxpq2j2KBLIy
lP0ha+NrtzeRgOu0oVmD8QnXSsTNRsFmL+ySA9GhLiO2lDWxIZEPIOFIuhN1BOV0/FSfnhzxwFR8
RcCKAnKLRQRe6NwaW6OsivC8OgJc8nw1emaRv2hMRNeX+i4s0x4/IBind8v3P8Qk48nzJuFjLvPq
ECv13GpplgUIKtTyd2PyyFBtbDzkyJhoYSXadVrgyQrCVcGO8UUH/rNIyS+7F5Ej39V8kTJM6rfA
DV1va7KMtjWDPqpQjEC+9qzl9uoDRyZ/W3idUbRlu1Utke7ifeDo40IDXrYUvPD+6HFzai8KRHaK
fPlJ1gM+RQr1wqkOpY2cx2R7dZfausZ/ltUFJWIl0XQtYICNADQdNCtRldP0dxNKR1MllqRam51d
vHSxXBs1jYiyCa77KBhHNwlnSgVY9wSV3I2d67eWBcqZ/jv4eR1VepNU/+zeoEyRCDBO5KYskO9E
J7PwyKAsjUYhFQTpbSsEN7A4Yn5vjlag0SrqSwbe0LEPEUdHfNXJN1Rf5GC/ZS4KJyJtWodD5GeZ
CyfzQvwWsVzrET0oDGqYttWu9Bedzgo4TX39jnZqkc0DR1tzZvxuvZ8VQ1fYH3j6Q6G+j1BeMnd0
ppG3kg5BwCsPZa7NGL6YsuIjeQqlcu4EGoaIE0NhDhkPpMggDPW/Qzdgmm6dLY34I9JD3Uiv7mjL
dMUTHvq5nW8S79mciZ1JlrECSGt4zX3rUspd3CDghjkJ0GoNQhzr+Azf9TYoCIKsckioo6Q+QrGL
IO6NrmPvC3MPZTnJ5w+zwWbmzmlmsIYmKjGqd+zUN7r7ly0wzLZV8npG+H7gU20R5KQQGvgR3SIG
culTA39ri42HejqIz6iaH5INcY9Tbf7U4Mu9lladkln0F0BiNEq6DGIQ/4TklNpIL00mj88iKAlb
4O22InkH0MuewwsrCeI7jTIrP6Utk1PYCCrFFQklR6C5w466SFWGPiswJjMRipU7iguTzBsxAdXk
tXXJksPZ09QNIdUcJSTWcgbIQB0FFnMYdXvkLVdaoveRmAR8vgKwsEqDy3JHiTZsJZ33t6XmpbUK
IYVAzF7npfLwDhWSUUkTOeVVcIywAM5m8IK6Xwdy/AtaP7xoGBv0/IIU5EJDwXm4TIdwvZwO8cE5
fTS7PZSlvS5VR+QTDddCNYnGWgeYzolfUVMpSFKTYkxaEfrv7tAsLpINr35FrTmYukqC3JmRqqiv
Vv5ht31q3i6NXbn+RpRswpDEaEZV5cVxmWUW+JsJl9B1iOKrmMkm3xegq4orfb9bqP2HmBGzVf/7
pe6mlIdFDrVP534bhaZLh4lJ1TaamVme/iWUrjASDf4PzcO+RrwR6DVpVOPohTSq9o4Ol9DCybSm
MRPkdbY3kVAxCrc5q9bkNCaVjJ9S+4QKx/vnsYmQ5GzVn27KlZvbY1HVZUBaN0taeUopaPuPF66s
h71CxufUq/bog/IBf2p/aF135FLq7y31REXZOnYsXcCxDW4bLRkayTQe1crez48IFcjY4DGUqCX5
ouSrawXLfYZSz5KlHz9EsnZ4g8DRxKPCp2JfOahG0LQyaTih1IPFEtZXtsBwJmgOdQuc1WGtudQA
8ihKhvI2qsHW+ntEzsXTCk7eYCe9OOyU2U8W0F8ZSNlqiKZXLQb9My0gTJQOMWKbdUHlEJ4dH6L+
8hlfIOqa6yP33DmPATN6ev448H3aCI8lwKhdr4qcOwk2e5vtHW+lKXu7u4STeRYz8MG74kAbdUp9
ZsiJMtKfTVp/CHhjljveggb/8F/W7Q9hNMtdolZYVlovln/Gt3oaoq/5eBgidgK9zpFlNgv6M/Io
BsTSkV//sbnyBX7o04Xf8g4Zu/m28R66Yr98gyykPCqZxa0LHcu6bcfp4UO/x2jb52P8SNRRAjT8
f17bmrT5Jt5dbCO8EtAPA/e8Ki8mFWEoHwKP+JpCXf9OwQJ6WNDi+LP283a2sgGiBC9gk2QanuQQ
UR5ItrE8X7fzlBTtbRsFrMnslYzdhq9ID+DgVYUjoApHc/PF7KaGvtWWWeQI5nt3sbExO+Ck3+Su
jImMHyeThxiuQTAfOUpdxk5C4bIcTm4PgA4dGZM1xUbkAaRkVkhKOlRfYxeM4WbZi9a24K4ZSJhC
hlxaVe0zN9ZmGzGoVIYIAnawZe1ym3NctE6X0rWUl+ZG55rqUrL8hnb40R5zEMGjVOxR2wzAxfrD
TSwJn+KW8ZbQU79SlGCAAs9MmVYYS69zfT2id3V0KgrBOMu3u9YyaH/SdxegRrK5d2Sl1ylSzSYy
MfpEBa4OVae0g/xiA9t0R49psL1UUYjDRWlom3SVphPJZXTrMkK+/At/J4PK7kK37VDWfMZapKFx
xEQTVho0wgkLfTgvLzBUoLzgIt/+lHxiSNFCeh90KDPhAmFIaiLVchCssSe2Tv2ZiGcbt8Qoi5IO
jircAllT33LZe5lsl/nesFt7N3ja71vIoaxWeqww/KvfolRS5mlJ48atfYQkhZswZ11cP/zXJ72p
Dc0iuSgjg/G7aR94iaV979QLvXtRZ94qEaGC0eSsX5xeWmYUGV4/Io1Lv3TU2r+LrH6V+HdNs4AH
TmGFpjAEy5BGrXesTBr8O175iiOXvQWkSbZxC7/r0pvxzotMDN7JRAMSFNu6lKQRHLxSr+NX40fW
qE2ZN/L61AOB5NQiiRQfzNYpStkWKK1rw4cCwsyu1Y9pJlFD+HB6JGoxf8UXLks3LwDfviwECOZS
rRmObV59WfeY0pHYaULJPM/VgsxDt3fsR4katpVpDG1rhOrzWkRAAFJICiEHh2YZErIQQBGsOgVt
qi9KFmeEnpwf38+KVdhMkFEMyRF/hoTSLAsiaDBci7+T5/t/CkrAZpqiZKytQKmoYAx7MelESAgt
c7JDvvA02aLCKFTi+MbLwD1Qb7UiciYFuI8POcgVnWesAFGD1QB6xqeMDeDcrKjZ2IhHnoSZeZaZ
UgbboNAg+wbmtuGpbR/sSAyoa/iTXukzyQ9YjPndTT3oxRpPeacist0DSxmc73i2wSJhXNc88RWV
1YABBVZXNg3Qx/dcKOzVoUGg6ehiXKrulQnf7pRE7m2Hw0rI6ajxPq9cU+jOn0ICHmGKpxezjLuc
URW1YcmIobUdJ4VApzy59lgKe5bp7UMqVoD4RRPTNPfUhYNtfA/oxFH9X8/kYMWFgK2CWuikhl2r
4si4E7blRI+7PpJwPl8wu0YRrXfiIpFtohLzpuM/mAlFfUdnbyKA2E8gatUISmBhE79j1ls80Vgy
X6Jo3pFMdg605+s1tH/fYgCQ9zn1NJdpsfj99U3i7AiZEWkbpxL652WLp7pKRyJb5p1VIFZ5Y0yO
FYXQaXzot9by3GdR843n0wIEfS6uC+mlgksXmJJ5P5WEZmc2acBObiU7IBQ2FB3h31kl6t0yLEjq
Q0uYk6OYuAhi9ehIx732JTGz0+qaywkapt3sGoERXQ9QRLCckeFXbhQ8b9Wiy20E+EQkICAsJDlC
mHjs9csDVrnG7LuOnbYgPZVuES4pIhcs9xfH19GYJrnXQyPHKK+BY09BPhYe5+PEuJhOpOEPXSjW
UNUlHAPH2dtyypwqBvRigJ/7TY8LHNk6wPm4qNA0uum+bpWoIbjh4vLAtwrpLCV3Mks0gYy2GxTG
XQicnRI4yFtmvX3Y1tkSGI7bMfwkD4OZ2Au5jKkYWIKZZOhwQDF3OWdhyzFP2ZibodLtou82DqX3
M0zcGlqnuTg5W9VCxLKKDW9NwR9dqEvBZR19RqTcOZpmp5SlcX6k0bT2GTmngRruL2Xksh94Pbl6
dRxw0FzH1tpPJhA6VRwyq9Q9DdF0Z5bfphzZhP5sXoSTD9bSKH3eJy8oTxlOkyJPGHy3vi9KbOi4
fkKT+JtwWxnfztwFpmwzIO/tZp6Jf7IQLg9pQ0Ne81whoNpyB+SHFFcjsgPJHrFhlnx9e0LEoPfL
IU6t7UYnRiYcy50RQ9lt6De15AxshFbEaSugIgwFcwJhMiBfApphczHuKrKH0H5k0KyeZW2aW0Zz
/vrS8j6teA4n1yT+h52R9ML6Bo9PfuOYc/ujAnGYW2Czhnj4xPRzYPChbN6+cQhODjaeRdMF+VaH
vt0UurjejKx5pL5KSdC2POIsXGy8x9ngy6S/geZHu8Ut1wKZ7Fmog1qDcoTp+/YqO56UNX2V0XDM
ARxnxs0QJyWd4TD48ic7dc1AHe0hi21GAQlQ/qsGOOus0fvcY9ebC1ttPsUodTw2dfXR0+Wz7LRN
FXV4GxHSu2SHrALPJZ5IvJJIW8/rZna+uItb707B2FiUzxKa9jjhLJeM4mq2dVah1p77eFnNe7AX
nDnN6veCyqFjT9jw6RZst5CDuZ64J9vNHT0RaG1qnQt81rbu+WW2WmHoTdBw9R9CciuW38JWN3vS
uNcmWd3CDtvvQucfiaIRcLDkonoOLUnZlDikS2fuA/aB3jXjqsRRmS6EItE+HuDwvLdQbx5SJwKw
I9n51vMwYEUPPRYNt3eTxVXa8OWtrR+2D//bot3A0QC2kIsFAJcT421bPtfM0TLfHMVqRZWQdie7
BZoYPxcdNuE9u/TS28dENl3hnmQvZdzJHZyomMwFI0xAEkyaxwkG+ZjB62Cgr2OHA27RleokbaeZ
sxvHI2LPXrLW5i5qMPiTmY6hDwlPPSfn0r0Zg13Uo2hYkNYGeNFTuq1mrJyk80lqfKSOVwmpGlsC
WM6qvks8FncAZt+teukQANt7HKq9g0w1kDC5DNSzO12vIoH1bQ/b8JRdKtqI+aVdZlLmQyFrhfdg
/qJuVsM/FHi+6uBdiCCfF95ZJ7ihSzE+Jwuv3uQHmvr3O9LLFpBkkHAnaL9qu2V8cb10F5C065Ze
Ma0TWAj+W3+NYzj0NeafKzrVJLfVzWxcpIgkUv9oDwm5ovjWNmvxonhNG99DPFIz3rN9mrkklzIE
phg90NNtXmr/gT1bnGw1qS3E1PW16YSlVDcyL75zPzIKreSvUBA9vZ8rRZRD0lthwafVPz4KYjqo
Q57nyzmG7Z/q5akDxKuQ2CtXR+I8E1Oy8YfhkX6ul5oAUo8hc0TEvNf8YZ4nJsgNLmUNK+dro7St
XAVerwBtoidtuziFRJXzWmnojZz/4KOTzlzt17arRJS0njm9oJyMaZcNEHwPtguV4VuFxZmmewV/
WGErcUOyX+EwNBrBWow0A3UXInvMn9gD1qEAL/T5VtsMn3ZXeivdHl8Qbh/adSb7M1VajZxcV12n
Lt+9QvUrJWWWBWaZZZY+R7KtxqtajdqBYC/FY/sT/J7obPouEzVLPWk0FFjMMESwqqT2xlzAaFPW
QQvxmOm39qkid2ewJ+4vYWPdLuuKTmT6Z+1b4Tl8SsaFMnn2YakSZSNoHCyE17u+PEa3Z6+OQPnH
rNGuP5QylDt67zrq4frAbsTQCCRA7EPd7RZHVgji+5nXEQMnEXCNr8jhCU9FFb9oOFTY1bnSCKli
DM8UI2DS/VQbs6GpBDTwm/JDjufEGw5jOXxo4x27a9xBxLlz0Z8+yyhe/aNLl4Pl6G3UjqTQCeTf
daD8ChvHuqp8Ve0wppeDaCKSQONpzsf2KqEbUUw47keOsM8WRJeDZcA1oycueKqAl2vqcBqSL3HW
OVHF//xhUK6TwvcCZD8uXAV1ESQCS5ZzwHwMhD90w/f3da+Kv36Du9wpWHOWOIA2DDqtnged6NUM
zNFqCFr6vD9k88WH1iuLpdMd/RynTUduk2y/JNykLg99LdPraU1RITE8mzaG9WU54Wh/K6oGZJ3O
okfhYEcG9bVRF/YI/KydgCHfzEgjIOvhIkX0CldYv55YIHP/wTlTLRFTE3pun32tTMWCFPL0oRFk
/d4YeJ638MOS7oCtlZPdGy+FyscprgaaIsGvMBC2Fy9+qNhwDlJrGlSoS09m+estuPydOCWWC8GQ
xETXbYLBvx+1h3aJWXybLuralpwzB1bW0IL5j20qNd0f0G75AOFwrN66mMGAgsIFQvzA6Jec3zKd
BY4KwV3nEuXy6v1gJJNKdhfam5ELN8FT3GZ3+prl1Z+DyudIIcyGNSIb9NsZszaR9MDN7btkxJu3
49T9I9Y5HyGQ9KxUyB1hsTX7Wsl8oBulq51+dgl8B9FAtgrTlk4C2zp32MiOQD18PJl44lgNP5Ms
0ErwtCFcBGnDHOgvhleG8uQOMmiu6E5LykCuIE9EktEVDHT5BBZesi17MjH44BUWsJyfQ5603kJI
7WSmucVnAHUDcVtnfq08WOsvKUSeTY0rHtzizpxVmutnMj2VbuqpOtelwPQuBFcf8INfZuVmLrmg
i1nfbg7x7McaACrFPSei9Ildg4N5tV0Bh4Fh04D2J58+2RYWdnCWLtX/odmwcVN6OdtJMmfkCdIC
mR+gJx/vsQhaCWrT6hH+Uy+jdpcR5x/DkCpKVuu8ITWsF2tdp9H75qloiem4DfdsUKIdye8S2Rs0
5ZLQq5y5Z5Mbth7Ov3u+QI9t/lLfpbdeL9X91Pfq8p6w8CA2Mht5lW0EtFHvMMJcVAHtViscw+c5
bfRhrY1LhuZ6F06ghVz313bFfRSsvMKsf2kylichNAcf1axLMnmu1nBtalxbBUeg30Yvdn1rGicO
QOJ0AsSrWMccQmwbpjs25EFrJzsV5KWVCizdqQVaY9niS73b2LcXojsoDMtP1Zuh7gBZek2MJG/q
T7eXqhknnX7jlv5roDQuvmFPxAoRSKdrYnDCQiVq18vUWiG0Pd89R8yGiUyvoyCgIlD2+KzXpAim
HlUSCGi15i+QMk8z6oeIaJkV+EZTG/GQ0CS0QYU8LrPwFV1ptxyJf0BfRJD8kezvGj561JJmuKDj
cDB1pnTWDO1zcy1f3STx7bq7So28pd5X4T9xCxWPhU06nldcmYxQXemmzhsA4jrP57/MhrvYECTY
VznOAtwV2eLuIKkt741uhrlL30zcRFgqGuhDBA2El7fwEMJlo7GUikixImwf+MDcLkpaW66OiIU9
XWJ1ImeI1NgnthN4qOtKiowiHJ64+yrl22SFiojC7Pp1SsOMR1Iz7aXhQ3RD2X9iG7EfSkNs8Azn
sJR//flcpXQ/9s3S7f4UqJV1b70OsXPDjD0yoQHQWMYPuo+FCoZ9Bai9TpqzhkPMXxGmFJoy3a8F
vJBsnPUPLD2j2ms4HsKYTYEjPqnCNYzscctzrI93y+ODTpilZ6cpDb+P/4MZjd8HSzl4VcysZsZ5
hwU8NJMmt/w0b5AM/hGy9QdQFtxpVemg0+/sawOzh98JvfjZWpItJ6UHlF9OtwnbJTrjCfEVxaMw
VLX5xEwXAwqC1+D7QFdl6nIWtehu+NqHZxAQVh7hitr1eJrjLIcBoMc8b2WFQwRtq7CNntqMBxQy
OxlYDEV6x6tlMF1bw88LLFt2JzerxcHMlfIW09J5uAyu7GxfNMNG5EuEw//gWp+/PoET7nzZLzu/
YOJANOA+9X+PHRL3A7hQfQ2u+FbD41dblALL+/LionEaxmkxbmdort7xsDSifEQHQN+EmyD00yD7
R7xj2U5celGU6go5NNIgjN7abG5YOsNJ0F0Yl7IDJEmwJxwsrwRpQmBXFMMRHfUssIs+V2lT3mNF
LiuDrSZ9dLPWfEMQ4rRZ6RTthFCDVRQZZ/WVBLKgSlPiLCjdHGk9nde4Gnjpkf4hW9xcExn5ZedH
ZfgZbyAsOyGEKACLdjS/cwdoLJROJ1kBTZ2yDUiWD4+c4h2u+sjBp+Zwwp6SoKeegCuflgE9k6wJ
nbcM+9jm/Pb11WVqBebCPhLXVBOu4RrXhpqFOw2rlLKE5IlUXjLPx2bn8R2uBMBW+l8Y8LFxPQAa
83tQgrp0dw9muLLwkgdLHj8t7sJ9F18jI/f4ICFRZHVugTCv1hsfgq6G73h61DeXVy/+WlKsi2IT
OCc+KfREL1VrkE5lKrRe0ybXG0eQepi52gJFQ4wysokoUNuPzvVUP7bV7dX6l5TkF665PT9TVRqG
FssZev6ChJ9dPA7lufOlaMcS3bfxzlJ2v18obu/LcnNXO+3Bq6XacA2AvkDeb8KYsLKh26ownv65
MVUrzFdj1IHPDxMZcaKXgKhmLTxR/QtJWFfk00TOB72X2+idqwICCkvBHfqWEEznpa48FV4rn2DY
uSht+SPRtIM/5VRTADwOsW4h2EkyMj0HJSpg7RPA8hA6DRumRBvxabRzyj8yG4jyL4MmKMk4HB17
1AMorgFuQ3wDAAjmkwlHASKHT9wHxtDuSUs5awrKvOR6ziDtOaDDlYJnHZqzfDeB52ngChbH1Dcg
Jrq5eQqtRetbELq/9Q+PpNeBXj+i2bKZGG1bl0clGl/nPLU9mjgVt4F47WcV8+JECeAZ+kdyvCdK
/FQNqwr1PiXGkCIzQABtisIuNDUnEbx10FYelebqzJc4azQmtYhTBTWhbgD636gsfRME5JH1uOxl
MrMkXUwBGToBnBOqd9ZjHLUkO6KoCz3zAZi6McTR5iTgwZIF+qEBkGrv+28fXpGUvcBSVyBD/rGV
UhMGv48GguH/rAS4PtkKberJGt7T4OT7QyptJCyUDxDwHvPc0hrjDgIz98pFHuJRyCjy/b+EGqWm
hbPBY7biiUjgpa6mYcVRKXXpQA==
`protect end_protected
