-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
011qqZyeYOf6pHtn5wGwBSJnBFZc0KO6wxQtKltwFn2swS5eqdJoRUHfcFR/HMTvWPkNq2q5TXAi
fVDUZhSch18Z+PSRh/Tkhyx9WPtzG2X7pmwfHBQmPOJesghJR9KenEEg6nlsmZJm9b3pOT2erOGR
ASVXO5EU2BOL6T8ZyJlL975gZLgev9w4v2pD/yFxRZbiAw4bALdbAyLFZavUMBaaP0XQvCvqeAH3
L9IDe+JwXh1ISWmUg2cHXRzsvtxXEfnPgW/yjSH1lrmfCy/1qkjagv3OSNeqYway2m2q+Jvza4ny
ME18ZQgKCKY5BBhXr9jrcomstnz0YpObkPsj6w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35728)
`protect data_block
bj5FMhsIAK8sxZV1EWkcqLJsICgrIzN3cw1ZarNXIuGrkWqZ/qRFdS4ooNiywWfqr/J6zbIVnCNr
ZJe+Tnr2z15FhQxeWH3EdFVfYlP04dfq3M22ZrbgfWsv7dLU/CzehX0fr9ogKaqKEiOqdwA/ClmA
A0LXz10XcZGa7hnaPkNbhBOzehfjMlfGUfSDGuRIyf7p3snXW9ONtG6MNzcI46JhrcMTYO/TTWYO
iuHpE+m6+ejuIT4ALCNrhj6mDTES3jJMyBZo/2blDdPNlqiRHHWcscYsJ9gm6k/o3ZQ2ZKTy4mR4
50836WU0nqlE3FupB1BuQ2Sn+Idzm/IROE55zp1gntf87hfQyJQq3jUEoQPswyiM5zwpfmkwHRkd
Ic4YOuXdAd9a7+KVlR0RltMtyB8AaRaOpg5C8QrYxYt+YeEYJlwTwLbK8Z25I9Y7GxNeZOgkYIDp
17duaQb6D0M4w/pIyx95qlVoprz9OAm4g1Rt0hhSbgX6gcseolNc2Uv6WSsGLytwgpVKh8EB8nxr
+5aiCOqC5rvsFNIvrlqfnE4X8ILsTTAArHagbTR6Jxe9ye7jVfnxy6VmdJSnntLP+QkErxhwvkHR
Iav1g0xGNWZRfsb5Lcd5XX7etS+EwO6eOcUMpiCN8aBhJeePjqLrsxswxoDsx+SoCbm/fG0uTP3h
T0NEqSrEAOOQhc0zZxd3lzLbb3p/iJH5zDS8AiT3B0rTaqe0yJQWSUvzUng97fBFK3HJ+N5s2sLu
ybsieQNgiMI6qlnVaOxZima8CLOKhgdhWMtiYSEOAm4ozB+xkSIBjewUjxFD/BIeDogC1mqRk+gq
aZwAN953kwX7EmItW8NX4ZEonzQcm2dQhWl02EoyOvjllPYgI0uf3RUvDB/nklCBa8IgASAzRtHu
x7JWuz8PZe2d9za0jJAwFkG96CCVWjxDbFHQSf9Auhq0eZszVJNnWmJoEp9UguOlzg7k6JDL+SXy
7KX5zUH2akzkUG4jIul6GsbWwJd/1tIfynyZD9pxrlnZ95WcrI6ic1IB7n04PlL+P+yq8Ft8Rtqt
GeU2hqODNsTlUowYLthnjeialTOYRvreRatmx6/X8+iShihzeC/hiQRhseIJzWZWsc8rgWRyCnBq
90GbGKFxpx+VAoBfeaEyIThS3EWDZtEllLU9JTLUphUUoNCS4lJbonseThrnOxNj/cNOaD6CgbNw
hw+L2q3TzWEvIsW8bPyf/02uMJZjmB2VDHGX2ZFxjnnHLEW3l7tMSknINTUSKbts1re+IB/1Aevj
TzNkbdgIPOzryF1JkTtwF1CSao7IAzCKDTcxtj2anPnDS4imQ0O8r1ljiWMgldnhqEqeVU7Px07O
vWr6bHEbmrmsLu1WYZ+73CnhmIY9K3VL1SP9QLYo3S5YXUB0jPbNHcjYAhL8JfGg0J7Cv+jBA1AS
PAl8cVQg88EWNkSsWzdl/veOtMFkQj+KieEUHd1NDh/yMDd2l9Iq5OWPz/cmjMglNUBN4qM6pt6/
Xeg7OnTi3RzgjAOXa8P1UZkCkTFm+H/nJkEwZ1CrXikmJs3jh1i084QLTK8HWpSzFFfBtKfD4XVh
isVT6ceUb6ZKA56o+oFB7oHbG9EjfpzsEEe9yKxOqM5Y3tBJODSC0HYam/XFc8iFddjA0hSxIwE9
RbXF92b5lLbK236kIpgriaUZH8NySOBOzTv2cBgw5xkKOQkRpbKg6lww2VYRgYwryexWwqD8dGmi
Paqc2Es9NTBm3pjwkuv0gb0H+pNnh9EqL+tkcSKmD+7Y2PIGRKRtFWPSNrGMq1QzgwsyYjzqhFur
r6jLxrAjlcv5BxMwYcjxfoD6j32tGZvUEiYx1K5s9w95gq+3NZkgpPVTIGqRbTUFXo8SexfuEhkw
tXD0VgCYzqBcSz6Ym3atL7Ix4o3CheqERfzIfCy294+aeD7BpdjkSIkeLdSq8HG7RZvakYqJ5A3j
iWElpiL/7ojsqM9jebrKoQ2iA1Cre5wZNTC2JIliWjgg3f1wRqGRklLwlz7jghFsaSrxz5PrrBYJ
Rao2mCUUqazY2ESdCffF4TZw3fzbG2EwuHuNYzSPxgeJ6mwRIjz0Ts4i/u24fcJ6HNLJW6uvsT5J
6HjtjagCYRHkOqVFfga24BESSNa7UkWmJDybV8D5gqMAemTsxC0uqgJxJx7A7FJrjpraYMK2sOL8
BZnFrDVlu60ytTVYx7DFmc0JuzAnoYX5Vd23aBzpo4pbUvjfLGGAu1mfLfWfguik1YiqAGqmJDSr
IPmOfGjFX4dbJ5jTaHyMqK4zRgCAaLVFKAreBpBHq1GFFpl5CHt1F+LGBoU17Dugx0Zb7xq1FyMV
tWwUmjjNEbZd66AdRTvSsUr9QEpv4ekLp0wqx1HqlwLgpi+Imo2qWtafk9AKEAZzrx0V7SWcHn4R
1bd2JDZpspAzDQyW5mnCDvm+QJstMOcsIXv92vOFz3dVhyZHSyrdnXx5mLa5SVqwk2AMcNYmNxms
avvMAQr9zmSgfSFcCt9oDWOudYK+tXtgoEdtcuMw6Zw7H3TasIVBjSwNY+wZ3Nc4nXHmPsJ5DDMd
oFvQA4CAeTiVl9qFi0i06F3Ym9d6J63L9yUDXvczCpX6vqUwVwwCpJg4xS6sLfVy6kndPuUeuepT
iyfuiohXaHcAaSxx19ZL65gvyBGeIe66Z5NjcM/UqQd1DGcWgJxc70A9C1TwukUCA/cgMj3WGaRg
BeyAdrGtq3vfeBM0kgsSj2jBRlJ2V9XgmiPEspbkvRqELjjpAMiRddTiYiculZYa9QpL+8paW4d4
/A5sR7K/JoLb+Wbk0vs1BhTK9HkNw2BFT76cRj2mxfv55HBYCTdhW47yaWOujpxqEt80yXMm+vEv
wz1xAVGgQcxVL/eIJLAFDd9XaBUs4jggM84b95c5I9XDHimaUWOn5ZW5fAMH7MbQQLLmma8RHEGR
aGRl29pS9IZrNAbSAsl4R6zSHSrsUJ5EfnECK7YrlDUzhn7sFjqrIWMxSgv1Z4bUjFU1NGFQg0kX
RVdJuFSpCgM2nf6bKQlaS1UkBAb9UZH8JSmtkqr6wfeq8VJ+1dewd9M6Ue6HY8SMgIzpTTUVBauF
WYERyO7WTSTGh/fDCRjG0QEAk5JwENqDVw7OuoUZNAlEi/m8SWY2sWXrMTCwQqZWvUOW7BvU5pxG
mZDsTAQvbRvcbvDeYl+pAEFiG/CNBGqrYisFpCaJhOausG6nelYJvm2nbDqWJOqI43bAnEZGDyHD
6HS1dnbNrCgWpCAI6B8td6Fv2fLDH6eGOkr4flpV0lt0rI/z8JV4TPjYPJ6IUyhRE7iieUcQB9A6
P8sgrVEzDmOWSs+exGvQnf8LPpPzkpWX5a6grcJO8eet7ZLHL6gL1rEs5iNgy9R5U3GmCSW2LHWl
P078V2mRx+R1gwHVYLdfg0nLo9LZmdz/Kgew4xNB41ccIVwsfB5H2B/d6P7g7287l+ZNdXjtRQQQ
Je0bjCT0vso39yiSP9Rbg0rH89pwoxnrCVZhu4lhkS/oBcU+NYs9d2WJ8p9fFwHYrccs4FV2NvDX
RKB3jTu9sqeF+bYkATGlXfc5SgkVwmdZGRkbfcQk5vGZlMQrswmMiPxXiSOj1x0CW91lX1OW/M9y
9PcK5/jOW/JszAmeRY7sEeNIMsi3HXfCT48UNf5Deb7fH/kMs/PKDbaOlw1rqfsJ2LNjNU4ORC+Q
TFxvrKzNkpK3VSVXYpC7bjmkqjovDV+4DwXPnIBkUBwX+6x9guDg61zV8w70JYOv0DE8ZcR38Tkm
6J3rBxdTNm7X/RyMwpFPdVI/ehVuTSZ2OlyxUKgpzTYG6pOxe++KsWbjS15uu3qActvwyqFCRs0x
wHDhBESEI7jok2coPOCMhpoS9aKi1tBLJBuNNjVftQAKCKnmBWf9RfNHberY1946QUS9QiVokoAb
WF3OThBkocUwHVlO4RdSoDbxW3HKoMGV9+hIbW3HH/pg0NtWKnXt2ys7AzJSBB/1Oiz4WEZr/7tk
aEKUhez8GlzeI0JRFTPiUZHOK/juF489nST3LMwxu40r5pnlBm3k3Nynh/3uwZkycCh/AtIdnH8x
/1K7z/yrFHu+glCU3L58swAAohk5DlbxaxTYPepbvFUfbw41srVelol7mQA+Nxp4KCUvNYo4gxDv
c5i5QXxhLQjQ5T4UYInd8bghQUbRsi+Y9G2fcPOSw/6Eft2IUfUTDd6+98BioBcIPRWCWvhIWOTW
K5X6PDNtdKYEPoRWxjQoGoIhCxihfKqWRLDgG/emXEJsYQT+AOc31fsv+YRzWKdubNP81rmROXJu
BQFkoWGeeSqemi6yKRxCq0L+dKX+qPUXBF8WE2rquclJDV06IuG68Nac3PgafILnPc6HUqCjwlOt
zuDGVdm3iw0gEkm3qnCDb8Z9RP6gws+wAu9BLqqZNcc1+srWuo8AB7rzFsXBjQqBeFa89nUDIqXL
GVdsafJafHeDd0v1ORfFNxNFtOIkr2jg0dm7TCNrAVWRvESNctu8QbY2dJ7gEcIpdotFFkZkmmcm
7f+p/zQOPaevlmeIw9E2XbFGULgghajV5p5FITd4ALPNNfJiV7vFBAOlPBIvKsnRPQBhaDK3AQ04
N6SJw+qUyHq/TD4pjIkM73gKWfcyvOZHatTz8qUvrbvv0kjw7cHcvHIOMnEQT+YavWE1kib4af2A
RStbJVlqHYW5gwVNb1PYgW+CpwaqHPT2VB+t0QGQkpu3Hp/94uRcDKjuQGszgJ0rNV02ndzogoQF
c61zBf9CtmHD7EIsun5WU/se9ziN08vTqG55yqK8dvcdL0qpKZ1Pb3rSzkcQNmYpgu0cSAUbUNeR
QT8j0Y91In4t33byYglwBLDJNvprAxBmqKhnKN00gOqzjhtphTGM1mvL4DmeLPEO+IyYybSQkqLX
Lhptx1iPG/lSdHdbyTaTQLQjE6PihcZb2FgKqn2J1eGp3Qo0Atkxm9iKekeK/mAXc2uVMM4yZkj+
hsr7SdLLbHTQRnlzvvnANj+VQ7VatveUGo5zoOQgk7mGSvcDcEpysGc2J34B3FrLb/l+fWCZlUS+
cdL5DPyv9n9qMrwdIdwiJv7lU08JzBMiYBoc2/hRDfRGK9MprsJ4Zveq54GdZhQgH+qRpx0dkyXW
2AOPz6Tvw0kAdUMM9+6wXKgs5wJwdKNdM/WTeDrXySZbXe8Oj2hXjEZ45HubgwCIxIXEcXXJCIdp
In0wCW0Pnqfd4h1h0VkO0i66tYaDQONiTIX/uC5QzJiyS/O5pP3XDR8b24luofNAWGujZbBPAzol
ks1bSmeuTDTLVvmCqujTN0irOJaRWDozU443DD5lIVk67aPTb26WMQsV+4xqowAdQSPa9Pc2OXUP
c7V4KOH//Rlu60OaOy9OoiOit5SgZxAQiURA9DfoPejgAdSTttysORA6S7/eM4uhiXgIOQn/7UmN
VWVjkFKNlbNr0ES9auwIR1bwPgZmMnQTgYfDtoSO8eLcnbJAFkzIRV9KjjrA/2lXmTmTh2rzlT3y
4ing7/zKaTRo80yN/1jNp94ECMsWqBIaL27WgXOH8DjVeF1x1kPDmgmFrz2/kKeE6cdnv3M2sRUA
m5V/ToFwQAd0bdMM6JMyalwUbSQWzIKDGVGyxlPlKRa2JyhXpoGBPSv4IZwoZz7HcekCqtoiJHSd
ItRy1v+XWBJS2pV4LnOyW0DZ38m9C95tJJ5iEIjvxRwEXm6y34ar22igbILwp0mG3w7gUYbuDM+4
6AQfzC6ILuwRwBR6pN3azfBAG891XFS0DWBuOyjkSOMg0ibavGTNZencGrjRqeeRrb0UeAdKDqV+
mEgEbdBGP4V6tHh1U8McQq+IU08EzEQH4B8UdBMHSZkE0hauSh5AiGbEy9/g1cO78O79XXgovj3h
VxNA/qYFx0sOVN0CLHRUbJi4t3MvDJPqzSZFnNSDKR8OXdhuejOKv0Mq1595VjUlHdsnx/QtiQLN
NyD/H9bOAkhWdb9oLs0SxYk8ftYmhIlvRmcF/E+/xotHZio6RzPpINYfvLtMvEKEbptr2SvGp1Pt
jLCeQWsLntX3IUEyAygQwEUu4a1H8WIODJeln3WUb3UMCsMq6Hkx3b1sv/asVkrEF5QqjE2QR8+s
rItDpMuqzeccpsBUNKDwhTpIHvDku4s8zg+Nqf+VQJQq5EerLwkA2ZeFPjQf6PfwZCy6qeYhr0y4
dFGeEd1Xsj565S3dlhkpxU9dQ6Pq6Myma+wUL/bK9MPH4/xPljxhSbUEOT+006yz0d2ksAGcdiLn
wdicBKSXK4HqmnrogG+Zf4VQj9l3saTHLYhYb+xy8dDZuP5LHtHecwlhBwRXEKudzsuqzehDSrVO
nha6fpiOHf1frgKmBvbKKIKd667EGByEKFP8gEp/ccdPMgAditTWH8nJ83WWexW6RW3Car5Qd+yK
Vag1wo5biVInWAE/0tUJRX3hrTpIRWk4QyWKwfptVkSDbv5jsUFNoEbGrwt1qPd+sZpoEGou5Uho
foBfprRA7VcbB6OPfV9KkpdHZDjmOnT0pbLSeNR4xbN5ODavegNyzha3GOOpufr/K6hGsOx6kL6q
Owm2B8B0FeqJA9eZK3s9oAPWypbOsPXFsPftghjtbx0YUVMhzpCqpNiEuxPZPAVwNnEbA9GluHXc
W5Wh/eFLO6kYiLEamsaMZ9AyAt64nSxHOc09vosaEuhX9grPKUOTS7tBaHIl4o814D7WE9JwZO7d
3ziYt0rFz+w4MnHKiPcJqfLso7XMgen3XywC37/r3B/nb1kBB5za3QjtGee29OdHU8YOZ8mJrR9u
2i2A7zcIG0JEVNqag7s0qvG9IDcq00T7i0KjgskXMZrGKt11Jz2cRsqry7f7pP+iztdgsgCJ6+ck
MNjbzJdohDLryKVQLMd+kIm6thvc/T/S8Ys8RBhWGiMa0lqJTakDL+anVZzT/OTTMy0oRIfW33Va
8liYe6I1D+EAIM4F2Xr6fxUH1kry6bAkiwf8B2TiGAcVjCUHKzdaQunXNMybtmSV9yyjxL9qmZA6
aJzsaPq8aA57mQNSZwO872/xtH/Vtj6/xobgc0sTL+pUMZwV5pMGp4OMkrLxBAQg9fPguAQ9esjo
Lud6ZViXROg11zKwHTHbKZC+06qgTrVT1RQd6Du2vE4VtPRYpaQA/R/9necjgV11aFOnuCk3Jsan
dns5Mtns9BT7R+H3e06higgPNQ8TP3A6DBYz/VDG1vDI90Ywrk+kxhxMN6SBAdp2A7hz+uZJfGiO
29W+Pea3887/k/X36NiR//UofDqV9po53PvLX0HO21MET9DL3XPQk81XtBXVFuxajxJS7KrNpAWR
DKgdmveIvir5lfYGmbN7XWYwlCjo6Hzm4HKLHk4+zdUNvGDYldSso+nDDzUeaOxRs/s9Zv+lKgYw
H4oQ9sVFlEpLO9xS8TdBNVNwtkll4xqOID9L4H+elwn+3LE1Jye1butyl0Oh0bxKNalstkMezFjs
rxj8yPELy0UbsMzkHkjWdTcPvKVnD9ZmK6d2whanlVUwho8spprEICujrmIU1cYpyAcKGudE2AAr
1VSm/xsSVklX78zahnFQDsOOsqYGf9GpwOg3JMFJN5DiVXZ09hvjgl7s7mRGutT+DLJ1Onhug9hK
k4mdV2wvoYkch3/1xM7JgMK+FV0T2bk2U/F8KY0H9MgA9BblV5JKdbF74K9YwKXpPG3YSEzPPo6v
4oBo9xAZo0JgJNhqm4LQAW9t5VQsIcIMtVr4TWEPpVEdmATHe19McusSWVpGx/ez6vgvhMKPW/r1
e0qY4cPxEBodhGg1TvunDKZgmLf6AWnQ2UA51eTJWlYc3Rkvlegw/RWgLEltKRiB+UbsemViddkS
8ybB3POeVWqJs2g2MCWUABgUk+8Fq7fNA4FMOmQADuzZSPMgoDXhJg54jsOu4a90aIxA3EILq03c
uuVbLOn28reptA1j09jnztCfdQc5C+n1eq0Z1PP+3WaIsNnc7X+yOtXUcR3TGEqM3uQyP3eAwDp8
EFSggEos9zandpYWLsHyJCwkGucfDsoeMsrAQmcrG4yS+WUAF5nZhoGx4qFUyPQjq98v/fA8YNg/
B0zpMazCf61y4B5UyTBMuwjOe1YDj9HztbCKtekwzU4p+jirYyMk1bDvQf6ke0vvbTRTQnUwaZjM
XuoYw3K5Z1tvEnpokDnxu6DaUCGT5Z8w2bcwrX4Nodx2KT5GE3TD7aLEsZFaroyEPKsHv9mJCImP
17/CMNPePGQCwV0+W/iaatadLr9clCxaCLih2GJVQhncxwKAJcc6KohhP0tXo3dYnwKC1lbaxgWB
zHCvik1+uF9rYwz6wsm9VI/ih+6GKDfhPWM7mJ/rtxBSDDLEExoHszDV9MhMWOdYdrA7yY1S5Bu/
vfO+xz8VV/LgcfHSBN+Kq08PpFiO3k8jEfxIRG6u6Dike5X8jBbvG+tSh/VYmQCahqpbDABfgvAJ
vuc752G1KBUzn4PgtvZluwNl8GoE1s0SEDOCSvY27IK37NiMQokTbD5yt9a46mgQDZjp6EjcD9qv
NgXCACsopVal8G0oRXyv0gXLs9eRQSMIFCryLdgqK5vKmKQa9mGB6bd03Vr4UFuBuEBWKYTRpn4t
tN63UBOmHd/fvljC8arXdZ77hmW0md9cjbD0Og0K09ohPtTu12In0Bkbmeq93QJPoNLaE6tCv3Yh
25koPdfIBPjHZz1XLgI4grUWtyEWewi5oaaNh/gQnMENTNFUX98iirIt39uN3MU6zf9hyLWU4uD2
YG3nPBgRc5DrbByKDtgWa8Oj11FIdlxWl4naoNlxYxMobKbtEceGL6ItxO5EkNmXW5oUZ0lsmMsK
OU4nntIeAu7ZjOBHJZtjvLsCKEWsU2E3iIb/Xgq42GWP0PcDKzghwQPgxE6NQbb4a+AmDevlUGBF
C9lM+nG6CN5mx37y7q7SqFQ3RlbTML/8WqC/o8OJFJddheGEHpzcs8Yu5qudxyQld6AXiKjm7vJS
fbAgw3dtpLre4x+kVz9EFstML+cffpWo0JeUkhThllp1gCZve0x5hwWu0erKy/SdIkakpT6O66Q7
9k04IRNIcK9QHHg1uTZm/465bRQf4YQ7XTaakXeIdbQh4s3d57c6kADTb1SwRPr6yHeoz/A+VjyC
oJ0nREUz5PAQcGoIGVYlPC16t1GTTG8yq44QpNmGDXc8b8NxGH2ZmnD5vew+6Q8jT9YgGl49lWiw
8Bg3m2nXgTms35+12Q00ZN6xJWZaCw+/Y6RDuIU3WD5HWCiv+VjfXhs/ZwN5SPYn7zgfegpx+SOY
POsldoXCpY0fz94GzrM1uIvuHeYnNh1rfeQgEf9fCLBHLIg2vap9fC26pNcGXUi/m9v9D4KqTTTK
k1AlnWfiIJkAvzRlRzlwkhbnKHZBPFnM5WZgA9f3LqHzcLTKgzA/+HaXgonHI6FNp3BeJcBIRz9j
dzDJADuie7Lv34zdfpV3Ex42zq4HwUHglm8AppyUqUOWPj2sUwfMOzaI8eckv2cBmN27A8/psgJi
lmsi+cKBeih4HS2EmB8jDkmBf9IJl7BQN5Rsnr5l/zQM1qU/RGkqKDnJ+1eM0C+8fMZGhgFbMF3o
OW/FNlcdJng85WVasPBwEavac0lswjo3JRKsKdm1V9I3JT7piPYqmhrjzs84rSeqwEAuWLVD4sxV
C/8LbwD5uBn1Ie0PYoeYqS9PoyRdppSqUukJsQpYMOhe7mYqkN5wC1j17cJ1K4aUKfZurCfZZIzR
UQXN72liLvHFoOUP6dl+ZW6AWARqH36K6TzfXyHQLyC2nwA5HEl0+ZL09DsZuKkLmliXKFK4KJCC
90pH1TlhKM6KccW8mSN9k9VPJvJUH3HlcLQjFCGKrxJs0YJpLJvUfLGG5ifu0IMu6j/Yd5X12i/7
TUhkjhy8CShg94G5PVzlhOWgwmcaU44/Y/Os2MIpv7O7HxqaVDkjhWVkOo9gxRPHuHxis0I4MNe9
U6Zpd4+3RHmK/ehln82PgLx+Ak9baSDXI7nieZYXe+U7fhrMBXV8Bpk7JP9FVQM+uBTVLlvlTFyA
JE3rdKkSeNpZr+Jz78NWr4pkCFbVubLSs2btMEc5JaSbxTzqUqX41MH98e4zlkvWB7FtEvgIcWMc
PhJ8hDFG44fVEJBzX0cxkzgWghDTSyjoVRg7RT80F1Ben+R3sX0egzsJPijm1kXjEV6DzGENPjT9
58Iowg2oBmviXiKg4fsSTRHV3aKt0hGSqR79LoUYsYay0LsQY087yKHYwFuquOwe03JJTR/1iou4
oZB3xiUKBt2u7iTTj8Ein/95cY3YXwOvefj7DOdO9q4d/vRWnnVWuucpjsz9o2GhP/oGSs6aE89M
EkjHGeEMpOxErmWVla+u/1LzbwX+5pTkVQN6TQJFZg/gGgrtvZ7fZvyl+Rqk6PqOke2FsHJe6HCg
84LBlYytmEnLMb/+lxUQsV4kCUIRhvlTU9CC+KwhueNY/h57BGBx9OmMGMsQgMIDPBBYsquJVLTh
THkrw6UBGQ7svz/67/B1mPEPkd85ZOJ0qmp8ewcf3PEV9+Gb9YteABduBHAVRnC32+F7H2VqAhtT
15pFQJ1BLFmnZrznRokq2VrKQUxpnR5SvPHmGxVmG0N2rj+x8weOKhlDgEz7tbOsv1j1reR7jEdJ
Svx19OvB/F6wYgWAnPHZ7kii/4G8q84ySAvDomo1PeyxyyQXbMVfnLj4wnwq760sYl20DfqX3r4/
Qbn/iko+lmhrWRvT4e6HVaqgmnYa2phxXul4qT1nBZ43JTmt/laNlHW2+eXqauKtm+kKswMX5kFS
Y3lRRj8y9p9ZEnPd3g750Qlz6pd2otSa1PnUIhAZwFB3rTAgxCPSLiHnGv78esM+o+8I8O1+OTMT
wQYZs9zJfR+U3EIw8s9tyM1oHXjyxygCNJdMbP/94Tut/EMbbkdov6TrtkmmTHz4HlKl4Bu1bUvN
RCFW6bQN4ReGZ/nhoSUJl2IbmY+ZKAZJEJkLN10L2EZq43tsfQlqp5mOJgHE3PLZdpbgp1w31cGL
mJFbd4X1wxbImm6z15Xcuck1n5EmUt7NJqF14Eji8sV6bNDJKURlU4TSXf6qhlaU6WWvVYjpQjNZ
0LcObx1flwNr1CidntGU2XuKBG4TJ3NkxNj0u9nAcmm7LnH+NSQP+Wwqm3P9S3O7JrcEVlYjRMBS
In5ruX5ZRTPn5oCGkt+794JbbPgJAxH2fhmVJw5wBIb/AizlQoIIcdCPRZFpMienhx+D1eScK2Z2
iWnnAGZB8Jvos4GHNDBXEpQjn8UERnPjLwLzrR1pXHQQgg9AMH0/3TX3Ao27nvh+cJBJeBHOzoPG
aPLc4THkT0j4aGqhg6x7PNPbSaHHjwMUlEXyMirrr9EXgGlDy3rr6u4O5Qs1FWZG0HNUoPE/mpqr
aH7yHLH6vHAXGmzjArQ9bYlavodn3nuoArwXZXrXntdJYeW0baZHhazvZ881Y1+4T4dWeYp4LiNh
1NyJ7fDgfu00MfugI69U0nkpDZGVmlXLoTMMbC7fF2LfkHciHcKW9lHRlFwlLBOhvYcXOe9DCyOh
wb85P76bsVH5xZt66P0YzJ52gCcas7LNHFgFRfYVxFM/+AzQVnmPOoV2p9ADuebYlxn7xPF77s+4
nDHyT9WYP36s0KskRrkKHR0JnbKknYKtXcdvughYtmZDkVEQr6WyRQQfPR4EeTLmQ68axOvzFau8
MOrGyzmybvQHsqdzTqwv+UOIVoXITZWCg0pPfvP3paqGZVgGhAvjn+NmFWBpPW5Oep9dtxVXjUpy
zkfU9uAK1FdU8N3j1pyMAGO/SFHSPr/V/0W0ZfWIj9Xt7h9h/1xROzfMbcqUbqAwezvL4AzbQqaz
Yk6wtHoWVHEME8lH3w+h1U7yBo/Yz3pPmpHudtHz5qXxRyMy9niEi2mg2Yi6xUJy9eLAapcWIvT5
wiuKO6p/CeCznFLBpT+RlPZsUdDvV4POTtEyhu+BWhPEzF76jhwfI2yZWd11Gb2AQ1ngfSWnJs7w
TslisfaVIDwCgcGNoJ40YnInsidehuksxkC+6g2vAvIJp7dgvPUBrdAK6os+vEm1V4Mtb7tlUvkd
gBDa6OnvAg98l9LosMUPRqolbB4nGofCApoSQ6x8/poiUpk5iwq9nqxmEJKcQBiTOEA8TwjT3Qlu
qgWg6+0BnVtuknm60EGYBJuF1gzOQAgY23FlthRoMuIepkifLO2/rOWcOgRHstM7gMGZg+EetClh
jy7/E/gZFPoUi0hbrFiTZcxgbayif5V4U5fwwygazVoBmfWZouLk09/YEUZINVEWBjajhrXhOMCg
VoBIQCWuW4Jvzft6mS6ztu3sf7Pa/LrX9uFYkVp2CoGij1oElBj2SyqZdiSmzLVrBDIU84h88+vV
LnYl9Wym6osbCPOSZLOoDQITXSYZwoa2ShQvKyBXc/dWN1QCoN2lM6TuOMI/9kA8OA7zHi1I+G0L
+zGw25KL032J5tvSkqAo0wXiYrZ3rhp7yjf+Ipc5e2/Ls/Fu9iVQDdJ+v+zjOEX4H01eZnDFMiW9
5YkmcUWTgjm+ahpHGcdLgkCBuNwCweTipJ/yEpTJCO84fR3ZdvJN8pgDogn7PSNrX5H3ZneFB2ux
XcLNktxzTO6d+BYy+JhKIFVJ2Ksjyh1AQchaWbBqZo+qDaAjdG+Qew/k62J1DZXjV4sxIsq6jiDz
YZs6P5k9JTlfL3ux/iMZbgR7nkeRxNwpbDlMRoPyPXPyr2y2ybSntMTzzbFy2ogCaHO1skL0aJHP
c4DcDVJPXwnIeYWksxMV6msm/Ngp2xxc9tHQr4LwGR2Wp+KTZc1pHVPsEY5ajY525G6rh+yQ0+qU
mIiqDs0OXCAMnjFrgIoIcjTm4du2fBVnM94JyGZC1ad5+FbPv/UZc34Kya4QcaAHkCahuzaH3pFP
UH0p/4LrKK9vu5BzBYl5aYzR/MWJkthEpTeA4H0b7zV57tDE/6RLIhz+1yD0XhKF/E/Hlkpk88qx
RH+mOgzDqLwSDxwGCM0beAa/xh4KAiE5Y8ukY8sHT+9+YnEwK9VreEEsN2XKKEHU9vhS4zzuQPob
yPUmU4AKi/HdY4wmy//P/nAdF/Xo7GevehW58NkugnMJul1Wa6AaKb6qduqUCBXaX4tfG2pYXduo
SWDhLHvI/SD56gzMVkvBNaN+SOdVsffXxCgyOkY4jtQ+sFceYdKAomHXmqFo8IYMCHjrFbgVydB+
ht1opfDjzqQWXHmsjKSLm28Ek49FzYQGXAmGlNTd5pl+3z7k8EQlK0nTQXoOEEEoZhBeIhhMMNPy
N8iznHxr0allN1jHhPGmwRmk27uP7N5jesmCGrQhOgaHk5PCu8n1g7TELn9bjNEEyS6CAf/lWOAC
pZCeacVFs/bgun1MBCwaIY4KOtndeDbEKAguaKBfgfAEryVORUjbkPSUNA0KcZQHcq5BXJdHrd35
mXXCXKFpyq5B6i19TVnwe7Gs/8pldJ+kLHufO8FA6jvNXX9BES1jFeT2jSSrtaeuh2RP4Dh0dlcQ
8V848GBuuSFlP7gfBtzoAUbGbcXOwGsAmvRIN6psb5XVwHgIgO5zUAPnLvcG3RBESJziHbFoBVHs
690/E2KIH4kkrCQpykMoS89w+4cNGEwDMPiB1AyGHu3Oz5DaQ9VomlTl+k057XhuAa0Ay5sN6kYN
Ui8EDEFsDPRH3RJY08pkeQKE5P7ea/lzMFR/crNoTSqBzw8P4kJX1xNtlvoHJPYymsMW3ex/7thB
NrIR0N61OeiZ6VaHtmEOgmFw5+lwS6KDLIcy5EQe+DpDRX5eJy768WQMn1zx/qCQQLt5siw6PzLT
Q429JK86OmbTewZPG9SBf3RdVqsjuCHIqSfKrZfc6g2Mf87UkaYlK8xLnQvLSAfMqx4GoV1JqxtD
GEH2xpZTcgDGvaI39AtqNPEmaaScdYRSK+Fo9u2QdcElwNjEv5nPLrCB2IYsp1xQ3K8wO2oLHAei
eAhljrJWAoQZZSeh9gWiBIFdF5FpVB4DY+yFAHXhxc1dA9r5Zr6aS+zJM5BnalqgvVyBoO8kAtPx
sdzTJPux/KpGKJiIpboC53R2+a7Z+0TKJ1DSPpy68a/YUOh/N3b+scNT4wrzHpfKR/prvhQd5HJ3
V/qwBKZraSzW6+bNQ5f8ZCOIOjjNZJ4AbD4GF9N5B7UGHroUUdqGdbliJf/pzO6iKv6pUq/Uv3y7
a6vkckKGMtWgp0T6AqNTyPo6jDpv5crI3ivKztJp7JdBihAMlV3QDan+6cD5Xm8mA8J45E4wqSZO
ypryjeZJ7qqXj4XFoYiDH/qVNa/7fgsd3ZOvi6FVGn9q3R0WIWk29k/fxJWFdVuBZE05rw5SHUR7
hUy0XtjoCe9+Wjk4ZqfV43BXHznh4QZOu5NHza8UkfapA1Qg1s3hGgpBxuAN6qObIKT7tc7ULNkI
uy/S/ZIonH475LPuIUC5lQPpCxuqE8CLV1vljiWA61XVnQCtn4R/lQMiV0mEjx3e+S1z10+Hl8T6
7cbQvJFlIoYTkgAbaYCT4Ls0jtUntw46H7xHoOgz8+7TNCpKU+FSHRMK1Zo0HRY6lcVqak3i8rQU
mVn0C5mYWJRyViQXdotzUnWarV1Bqz0F7uw6ZJr5iTE63T0vXkkXVlZcQTiDgwBDFVWr/nDh8Rjl
r8Ck8hxZfheOwF/TjiuP69/+Smfsp00SPplN+hexqx4+S6X6z3kig/EQ0bs5T37kcv4SSMEEYyUM
AS8vW9VcUjQ+V/O+tiblrTBdh41YrxsGJ37gVn8GOyqNMWOUm4Tur+CqK1tpx0VKFf+HZerOmFl2
1j041OiwO5BseIvEPIObgg/Tntd9sQy4G9GuEshUTxkqpbfSjZcZY0ho7ATE/ycJx40z1pu44Lou
hPpN9XVUI5un+NMC9oW0OI/4uDiCpMm3BSD02bwGL925W+wsSGKP/5sXv4p9cWgARo2JH5meix1A
O+N3ZgULgh2msVi3hWQAdo8heq8bjbkyySgKrinUJiTiAhHlFm5gzV7Ghh4vJTowohMGmf8MKgGv
w3hcxdCBukGho3XoN1KnuhzMX5mqBgfopN4QuX0huMDUlmQlXrVDzzaFDKt8d8+oytwJp1iAJI74
k+9tbdZi1zjZUql1VP3iVgbwnSg6u/AR7F0CS/LpAhpGa4c40AtKRsxKeMgavxvXZ67ye1GOTbIE
Z/40t2guce8hBdaQJJv2Mr+HTU7KbPgEKVjIWrFexrRlLLOtXSinqmGfj7ykbvGywB8ddHW6OPQ8
UddmJxjlX6B+/Wv3Y7ptWxEgWo2Ckss4Z2T8ZQ8iH9NC1XKh/1bybKTJ0ikv78TOvjkxOFIcjw5X
20Xw2NZxow6NSYOBt5PU3/mZa5JIZaxJPyCHhVcizTdeyDTlhvVFwmRR3CGHpZag5VRY2La22fyd
Qj8UzDMOEAb/rpaUVXGN14r5bd0VzO7hCzc4+aWSE1Z2ipt6KbDnAi6znQD17IjmiIAfY20DXGA3
sIrNxdv3XysIcSqtlqjlp1I/dh3SY5H9XBC/T9uEKLJ58Augz5h14sz/FbGeFHb6TqO6fWY28HOh
MDY0Puf8DUttn29A0aScqFx6D3m2aOHshlH8CeyRrms0YFFMOg+Gz29Ps7zy3Z/QYZjror1BONnj
PbYEa6N7MjPbZtts+MsnGna12bSSCV2S+r0gLAicy8JrnpqJanV+3jsnh7Jw74alPLt+624v9/Zh
JO3UzD/uHFQyghGr1FFbhaaQz1qUj/bTaG3wdnqmuQrjSN3tlIUQ2fN8DhO/1TcHB1CI8+iwjA8U
6CXArD+bxlOjM8VMDO0gx6BANqjpL1OjfxZuJ4RmTw1NN7+6C9AOm3dBuU/N7KBn1pu3X9n9W3Eg
ou39e52ujduo4mK0X1vBBrt3MUi6trKa2zxak0vN0e2WPTa1/oP51KsypV8bc5G8m5jJsa+yGbMD
SQcQjtqRrqvOCs2iJQ2y/JvBenQNhRNpCO75RpX4M6SZnYhnLNiQhuMz9LiJnlzOaZZr8YN791Bx
H73Y8zohe423jH9PgzIwEPRZAD6Xq9ISnU2W+b+jXrYpqc6azN6eiw4L1JsLeymXXm0Xvghw6z9o
OiZBHu+gBuivIk+c71ettoHt3Bgy6nk7Fp6ccam8M7n7S64UgGHKxox244ZLfl234eNGgFs4jL9O
YMZWYrKBHoj8Rwfu14ip8rF4nAyksl6/I4Eb/56RSvQwhdfjGnO/8QaCL1Dc5gQbB0GcaBmGiZ0+
ixAbGMw1+Ssc3FoWUpF+8BeiiJR3vEctpKpTIkBq6ODnmGXvYBhjIb3Y3EPcSOdWFiLCkWn3pJCv
QNqa8ZMM34tMoGmGgazLXweoOhrnO7ddtsYIGjZaLuDsZXtPfEqQGC22GUezgUIkYbgTW1r/0Jws
s/eJeW/+Sa90IdnYhpPQ3FyY4/TZEP75rfQJh5c2y4YKWR96PnXB2C419z6FH4SQYunAmXn98LlR
b4oGqgAdVStT0jK0MCwLZw9BqrSuzYlejOyhMBUzfxxl630HtF+cB/z9CLWBmFHpviHBc2zO+wDF
0cpSd3zT7DVRne94qY0nxdv1soDgl9b3txJe2ovIpT5EEj7IZ/kZO1gkZSKTebkm5qePIAsTnuIg
Zj+Ny7Rt7AtldIuPvntReu/MNTVIpguezM/EVzKc0TMqt4c05LDXV/TJoFrMCWBnO+taFFglsIOZ
boB27Qd4papKmJtLKVt0cpD9edylIXDB2pTgTOtJEmsxVj380aCQti30Eds+oUB8HvXvP6i22r/Y
k9Huw+ScUPJ3W7ogu4Uh1uGMsSHXmzoPl+OjcWBzzGKEp4FnF/++lhkhCIHzMvZw+AV+zhJzUC2T
7cviu8zGLFfVHFWcCbg16EYcE56IR+Lh9dD3YU/erFCBfpt/jffDP/dyYn9ONZUS+kqqMEQmx3oa
IcetTAeXXmCEha6Y4ouCDaN+KKi0BhmdOsxDZLKBihXWhVm/Ei85MDEHatVozHEVg5oFxBWzqnKA
CpZnuCyjkfiVd8rqA5fE4t8gsSm1yEdq40YKSMpr6K6hoGbV/l4POgyG1JSJy1ypkvAWfZaSq3zu
dhQgXP7HQ7KHLq5QZPjSFULMrCYqd5XnYtvCKBiY7xrsNOSJZd0U6I7CsYbMlygs3Zw3nRaw++Lf
1ag0iSYc/Ft7XXl9Jcc/PGWHmRuD2uBKjyOziz3DU5giyefipQR9bQg9LKs+2iRURvhhe+rarVO/
7G3wvayfr2YCycmYWYk2CTo6GIgfEe5Ls4ecbjWjQnxMMkqm/q/13j5j7/tpIIPdaA/ycovi0Kwi
7q/dC/OWlSfgQuHhRpDSpkH1b9nfJLFXSHUHibIGaxDyOQFs3s4jnv7i7lov1c0rq61advzOcGZP
nSD5CrYU9UMVB2aPPVlaBtiWZmi1CKVo/NmnpZsH6NXbVaEyczXZBH+mN7uudzO3Tw/8MAoQkWxk
53ZGiwqoi+xCqVZyUjnINvLz9cYe9eCioGoXA0qQ5mDkFrj+vwwAhHGzuaqXJ8/JkSDfQameg4fu
XplEbEG6vviY9nh4HXNsIb/tYJfJd0pU9n968I095wxys2H4x9lrb6JpIZQJz1robO/iBOIXOtoQ
QlucLnFpKV3KtTmoDnesBoPBG3LU5VTM4AsN0Ixm5jLfGjBzQFl2cUE5TRXplhPm/zpIEB0IB8yN
0QlcENF+pMUpHbezEuQOfIoiBwbW1MOn9RMu7WOQFI9Fg8I88xKHuZCO3dQh+u82sap+GUwO4QMP
9kD04PB1DQWq14pors1awjEG2DY2ZnOXlA5Hp8mvCzh7PI4x1rEEHykXnvcdoZExZ18GGEt7XMHQ
fQiqNiFP05NMAbqBGpnE1F0eJtvOIlchn8Q8jC7/gvjH98uCuHXUAEG85S96xIqZE1v6DYCUl+oz
/St1BqgixlEYPDzElbtQD0hIH/qjMAIWHXjzv86jwUuaoDgrUPXg8/tNaYICLG1NxuxutJI+crmv
dtvjEVVGye8HDJQHRS01BPz7MMi8e2RTt+RLHwkcCvfGLjwoAU5xN50fMEa8Y0GwjkMURT66vof8
/jAT5z8rI+uapKZUByPVl0r62Ic6gEZ2OJt1MAzy+zstmCFpMphBl4fTSQKUVwMQ3XNkvZSRnjHJ
eKQlmzLIwVofgxJ39gE7q4bFOcoLQ3m6inO2pCphYjfgYhkoZ0LAW8v64/UBL4dfVI9EJvB+tgJg
cDnOj79vUYQjf5aQXZFfxOL8XbSHC8TKLVcDLrbmYESYf9whx5SyAKuR7fPCC7taUgj8q8WbYt3t
1XdnwoNbfayPbWhTFwDoyRqEYIgx3rrtObz3EZ1CEvIWD96Tu+U8+Ku+pVaXonmv7DLFf9ALA/0F
8lhsmuGprKixUwCIWTF4LosKvzn0JtaefMrC99pgpmorsCEdoiCNm6AL/anvmBf8Ms5M6Gn7AM4I
6U0xgBL+aS+WRv2t/0CabDXR71zelvbMF5v2pDfaAXSTtgOONAm7anVACNt+gYyZJfPf8u1mXuEF
rqwKxObUllypoi7rEOTIPHDYFkLW311Bh8Ww797j6dKhbkXRMxnkhp4ob0WgVKWUyb+vO/9ErGgp
XDKI2Xo8i3n0hAUd2HRR0NZ4naXJQraeElix3PtzsLqDi2Rn96fvBbLjX1vFVf+S9eL/vUwhznWV
bJvAY9ynHK4180LI2f3/jiiTHh0uCz3DvHvzEo5zr72S2pL6Y39PCaqjtQrtQqTmGhj7/xM+RkQD
cHAWAWFgBYf/wIsVtbAQmCXolIgzL+Nl62Fho0kYx/y12DA+UuikJ1UKrIvOlN+BCwBZ1yD2JYfQ
RcRgkB24rBLRZA8nPzBVgoyD1I1rns0SQmrfx6Qo1HTIIgZ51qkVLnTvbtuHWCHnT9pr6Qt3aNoc
28tZGgMleDNqJfPoODBjJQGAAPs5ZR6XAXUnB1vJ1ztCT9F9UXyEFp/roN0iHBIt/DRU5NTJsrSs
5KOiQMtJH6b8W1vRzSU/y6Uxrj7+NhPeYsRjCfZQW27e8tXhwsS5G1tXbnKXJX221eMmJyXn/pAE
w3S7URduZKFiexARmhvR9t0lDJEOyaKZ0dXPVU2B7yK5GCJAnTj9545NxKcz+YcxV7wRHGZfdDF8
waEsnLK+iTPV5pp3B+Fj7edeFp+pLT2Ye9VYKmaSvOkb4BSTNtDUh6zd1rlfZTlWR/SlmF9kjNyT
crQbxcObGk2jUPHAKebmXdpvdYOqbHCiX9k/TdmXYaIQDXwKuwYXhGcPRe/5cv0mR2e6Kq49V0kQ
Mu/Of6X/xmzAI7eTdeBYK4jacYETFvUBRRxr+BXL/cWkXV8uvYBBV0PDk4F+5z5jDydcVfF8uf1p
8kXC1Oz7ULd7E6VmJzGNM9QuNKqIkC3iHNBaehsgOtUacjVaIvqFgk3Bef62fKMOjXcjC2KDp8I6
q9xS0EJeiKBK3kVOil3PgpCeuFYbRAgr9J45IGO1vw1HL17x08ZUxs+TI9eJkvaaFBAc5fKoxyci
HpZqnB7tJkc5rIMEHY0f1zr3O8fSibngvGMAiyJaJvvGJeH07WJhzyuKY0lkS1kZGIkC0mxNgSy7
2NNgMhhNkpBttLv29KH0Hd8yvg+zviB7zZyaA84rP5DB3q2Y/URve0eR+s+PkXgrdCn1X7FYcJDs
t41JO8VOaW3zboAw1nDIzHAbf0NWCM4jWwwuJMU3ns2ZQuIIOmgSkiJS37MHYx/D6n7tEU+MZxyU
zFGuTJfcQS054W+VTSTMuE3ACIEvez+iXzYG/4bqkw/zdbp8kpXNVZgke1M9NAjwyQi+tGLRLdy1
inff6wQSSm1RcWlY/PKVxWlbZDWrXXChpGjYIjOEKgdbbmOe9jdGS6MPP47NLfESV4mBY2p/FzGG
WnVICCrowQNghm3AGd61bMIBgjSclISC5NIHO+yPI0h4fc+Qaa/wqYXfTT8or0v99o8WTgwrZ9/r
c6kGhl/PTwd6r08wR5chImHhi1fPZRiGKJ/q94uT3flV37tIupco8dNnIM51RzYyHW5XIDp80Epr
m8birk0j6Zlg+M5jzhRi/HtbE6nTFYr74Z+zNV6z8TtYwDmlKDGOwevMqoqB0YUp+4RIjLN5yjrc
NVt3CIDb7toFW78mGFXZ8xlQhvFE27Ku3Pe5bdnSKr5lM8PDIdZ6KdwklDjClGdE7K+Uuh77bNEG
tZaxg5QLpWedFziL1qY+/hg+onSU9UJJ1jgHydi245uUeEkR49653k9SCUlyR+yEApuSgZc1hzF5
bjJQePgQA9R9zFBnYhVWkpNpFc/w9c4GHPuwG2Ek8SUDAip0CBcnBuJ4w6FzzIeO9mimTzpWtakW
wNQtvhNOKkqi5au4aQfv19zm+usjVrQZzzuz5cgREV3xlMzshrTAyMts36CAQ/DIweB4XpTSpqOG
6m654OtRl0iclxR/gj/OY6NscWhulNKM39lslxiJ5wgKPCo9jMasRUsFn2LjdheFR5IFrid0+wn9
Wrw91AZwQYUe7JTm+gFgLy9U3exJcMqOKymgrEYoJYxocJ6TcGPOZd6pOPAFDFuK7jYjagIJIt2G
E/Ol6lvNUVmXx1eYEa6mRTUmv7uFkcXvNmxiZZpWRlv6ZTxLoyQ67pOdj63lwwQtzDLXOs8Z3sUd
ygtz/1ie79X93nBYUQgfMMe9FH314/3xZg+XSyB6hnX12vvJo2v5I3NSrMkWJOYnaV2j2wQK4GQc
okc2gELRSJvPOq60XcKK1k9QiHhrm5siRYHklgRaLhIS7v+udqvwAHc5jYuAFiGhNU+BodGgOLJn
nTASDl3EavmRNkg9E+Wm9DH9iQr7UNaH466Y2O1aLc8ZUqwTl9dhY8Y5dJ0iNSeAhXr/VwKgrF4/
W75LsUuf8KV1TkNtnxqWIbQQtojrO7n2kbfZemio1j84n1hnErSReTRt9QiuTMuP//CCJLQ9oGQM
4+QpruLRak1wWWPY7pLMemIqlpXsksPFhAiJawCx5bvBZUcUfnn9ibDOyhzlwaWmI5u0cicWhwHd
/IgM+4um0/XtWlnAUHDc8z8wbA4Ms1b3SgKigV4Q4/5P0y0VdeT9YqI7JibAeQ6SatCDBRzqRWO+
U8fbXFySdNzdDChBNVaeBjB+YwrLaJauPBjZ8OTP0mTki9dbZlP8bFuy5PdPBMADP9iXshi3EiX8
TgdDnesWawJzxweoHAqkzrsezaRtMMsOXbT++kv75ZhsRRR712lUj93qWfVEzPLxrC+hgIbJbp0i
Hix+9RfpFz45CMFXUWRX7D9o70MByWCkkRbCIw/uYOePSEvdFz/IsmM/838MmEVUk7Ln3g0/2DXJ
161YU2B2rUTSysxBgb1angLq3UjzBVBWl2aMDvHuWoxllsIAmnxgQpsES5Wix9EsIv7fc/kC6aUk
XHwnSKSK0okQf9b+/fWRATkgsL6sxYnphcTSrZ3rIbcWmrSCIfDQm2BO38yyWte9j2SZRpLWPzi4
JLLuxTPc+pve669WQBiAU8d1crJLyv7VAHUFmOLX0y/gr1kQNQlWeR85g2N5wqMwseTHrcE7sqjM
FGDwQYqVX976vtkrh8rBaycSozg1FxC9efBcqJLNnOGmwXrCGpeYFTLGQQJJ2wULVwhlFFkjM38s
9tZfZtkiG3Ddaf2c/KRoYW0Ih260cxYHgxlhNXwdCtC+pbR31LCjW4XVGITNtcD47eTEkb3wkeMg
1UYsBHZT81etg8aFH/pAj3RB73UucHtc7igQ++NfvKqxyHwNJl1udeeLnClE77VGaJgjrqHqB0CY
Aaee/04D6hVEciCLvJPFyMMTdfeNZA1iJoBthFaE4qNQf7hpnp4DxPrgLUbvHFMvHGcVxgdj2KAP
QOcrCogoNiQQU4kn3s2VFdozQ9bN/HzaQvKiTZhdMStk0A4ScyuYhvzgQO5MS0URMHjLiYyMSzMO
ytJpFDVrYiyclOWvRyT4J95ElQ11S1qPsfDNYbtFWdueOV1KHyCqn0/zHUZbd0SPjAYGtC9eGOKw
vY1EQV21EaSbTvNr9lI7+IPf7TmE1SOhBWl3X3ujoFVlbHNzS3vmtbR/MlMEYw8jsQqsbqv6+DBw
3n4UcG6d11iyBqORodtOdjKAknlo1LcIdED2093lg8YAajYflXQDJNF+YMXsUPFTHPxFlXTLI5/q
vAqeBXeOI5ROEBe5YOIV4Fh+0FZJjyPjqZQ64DIA5UxS/1rAH81iSMzqZ9cXXs78MDgKMRH5D0YJ
kqAK0zojufdft7Yu5m/90BTwx8xr8KWmWN+h+5DMjDdj8SJHVkC2ysV6qBBk5zhpzL2Yy2TqMApQ
biEA0N/qdWANCQHibl/T4LU/M6LfaBfNHCuiXzKw2WGL8c7NnXd4GO5CPC8dueMtBqRtB6Ir4tUp
/HsRORlpRvU4spuH5WD5/hhYcIKKHXs2evf18bSiw7DWv3KR2iLydgyghPHemzz53LARcDzIohJV
G0/LvUjALd48iK3LzAlML2Rv/asaTzdSbLOPqRwMV6hFfCE8eLMLSC2h2TyBV2PUAQl/hWufgCIo
t62ghCHyBYk5KufPDIaOc8rWQvK7EdO/UYlRD79A2oRwLjusLxydUS6XclY6zr+bXWw0V4Jv7iVg
J2ScwktILyuJsm/bDeTwl9mGjdLxvY2w/aVg9TZFssrJM8jAq6YKJiA9D3XW9NSyyv4ULv/7WYUS
P1U2pDslxRiuYLTmhCdjSAvtAkO50nwxu4AhO7lmXNXJf6j3eiOgdhuT41ATzJVPwhnRZxghqZWZ
L0LHNuXdA/H3lZyuIS+iF2maL4Ez9x6AZ2FiECMwE81QKLz0LIt9CcfWsyLLRDJwwBjSTYnlX0DR
CPKLl+NuvHQlZiiJ/RB3R2/AIdGlRO2+8rry65w/H0hoL7WTrWdPgHQ/S+JKkcaaZaftPRNGS7VL
/NFrWss+MJ65AOaI51mbM43/DIlj/OefmVl/uf7TaE1P+8tGnS/VULGo4QLO3M6if2WoA/G1len/
ex/Bfwb15MY7yeXacgZV2LTos9/cZZdKRNXE92IKAd00JNN9ttzZbi2OT1MWwoqkq5asv4kuODk0
CP/VFEAlfiE5a7DN3k8+ivnC8r5GX1RQ3h5VvNGLZFf74MbbV+aUGZEHQfEfPiiLn1BSPzTQfm19
KSYDgko2IwSsfJLK2acZ6do2rx9khQ74vApa0k0lb7LpcAZsbu2LF7yYbxHCBzignv/aqbABbfN7
Nce8Eyk63nMOv8tA6mM2znzN3izQFZtDfi1EFpeiji2Zrw7x/vZgykcQzqxCdBTZFdf0cVojnYIn
4NIl2QerdpB9ETTaorkBjmvA838jfcdtdvY8zBRL1vOlFJ/jR6NGaC7oLsNeWAysqCAOJTicf1zv
MWxbKLv14uO2k5WRCLgutPSri6DKbMcLJw9vbeNuhyNHJJfQbvJMJ+jx07zAVSmpZUEd5SQo/5Pp
OWtKB/crvJtJkYS70sWgXDoBpFVWWCTWZPBOfvHqR5EGVHDXssQ4piAOzEtRKMxkofeCMkSfC92R
QnXGSBYslGxahNaxAB5z9iX69EjOFXgK/CHJViHAG8z8Wjyjr8GB/zgU+9yN6kHDhGh41WuOj26a
rDHxGASJFm7h8CWyJpubakLxYyqYWgNSP4KuAtBMkVJtV5VYofYdQdZ9wJlk8t5Jvxd3uAga8vYH
9r0uNnpQfkMeqgUGlu1C8o5UZIx2tvAjAbuAvxRjWlLfE43Y/zUME5vMwoJJwC75OdHLDwgLXCFa
82kuboR+94nqTTiPIxpIZQUF3MmUgbtjw3/XUKMiLCj51T3/Gr8Ky6C9nMVkA7xliJvsXh2q9URp
NCuDWwTN3cH8Ye0tQGmFnSaSbuPF2GEOZ1XcsGwz1OU+pAwce0akeldPprXKW7/tbyGrPg6cMsVm
XXrsKyX+YUVXZdjotOwUNrt/T/UL3jFCdaacDOdE8hQFOikpFejjjXkVvovrBCNlS1W7D+QTGLZ+
35fAeixdLyuUnbcgGE6pYWLMM6oXMh2AW5MrenfCnh0ydpHXybAFgv9EMuLyvMnBPFW9i2JftHkn
zm4K0xJgU+B9scD26Uz+M55TddOX+ueqJgEswESgDcMmfys/mpLQoyD+IyZbJ9mLpgt73R8vsZMZ
2jjIQQNOMOFk6qSbWQaCHrjt5ihQOkc/k05X3Kq3mmWeq9/5gPb1ic/k+Jc8K0ZgMq1MuVUxETjO
caxnj1WQIsTtRD0fI/iVm7w4ch7qGD+hlQn09CjSQkcdgOuQ/HgB4q1djg7CLnbBKbbMGgWWfTPs
FeN/fZbcpOgHXhTmsY/qmN+tNfHoC7PPine0wwDHMMTrUWfxugU15g6QP9Cbvec9Qei78d76OQPa
UtyW65SnQOdVCP3EmJq7ol/pk2wODeC/vLYp9+1EVeajSu/n6Y4swuWZYHcF2NdH1UcK1iKzF1xU
kwtwx8WhgNmO5815n2jffdye+DY7n1eUthESb4SQ17Kiif7jS4YwUS/eRBfyQaAa+J9xYtnqEr4t
ZipuNlAnlu2dE9ESBcI0g6GybSP6FqDRRPd6T08C687C20S3Qih/BARarHd+j3WI41+7hENPvi6E
+BZ1GXk6kc26W9oF3mc29p0xbABuxMcqwi2212nshqxJ829/hdY66OOpK4GC9R8LhPzri+fIPkTF
PaeBF4W1jtBelM1kQrNSBJbhNzEmIt15Phj11ZbPoK9ohNaevuJKnfEeLZGtRGC11zcx9/cc9Iqv
AHEKnZFVVTlKQFFRUYXQrfKMa7CBWpYKXL9+3P42Fk1y75CydLdY73Akhek/rcz8Yki9+ao6ps/H
uE3ETD5py9wZew1jTGMrI+A47MSS/hJiw4hBIXsF8gylqbLn2lHZiZe/0n9QAGlELxL8W6Q0DB5a
Wugq6TPx7lb775mgWbEaa2jPg7MUtkVWBNUBQr31pvv9qXgEXIQ4nenQS6p0dXMBc6QOnxYKZ6tQ
M+HNPGLzusVfRIXYp8DP1R/WtN4x+d0BU2PSD3yj9c7UmnQIO01y+DVTEuVrJvHs8KGrMBl0J/W3
9/IfRrt3gGTnorjAIjeqyBWPhDoEDL20vd7YEDCwkqt+zeunvz8RIdvF/1aevslsydswZ+zIKQFQ
nRraAp8AEmQKk4K0A1uSaoUdDHU2dXVXsakG5T1OkKcSvU5dLErxHUSyR/zsJN+OXphx/gII4lwh
7KMGtM3wVJF8X+bUn+UIERBZfD3A/yjHdW1Uw82zDnO09gVuWGX07F4pWxIqM3Pi6o+1p+3QzXSR
Kqy+wIDcOiSoUryMtd5ix/IxbXrR9BZd3UNbbENTWAEn5nbhInMesLkYxN9MPJz4W3kwFKdksHxD
8a0gMwk8YKQ3bLn4sOh1jvFWj5ZG7kzU9M+pIHif2sDXC/kXIzgn/m/EH1pUYMw+iGzCFUFJheB1
52nax9exqdP2fDxm6hkVvfaV/IE80HqQoInTbiFsjNV9VgW/IEtRtbGBYRMUuSpJN3St/1g6xpAb
IHrMjPhAwmYQrFHhUxPiFPtuiRQeWswj6PyazaeFBjR4bDwrxx4lzH1C5dO/VqH00GnFILq60nfK
W9YIoaIqH8CPoaDvNyHnRgv5dCsoMGLmV7EddWfkBc7CgSTlmPPjiu0Jy64NKZDJMYqgnbibtx/9
A44nSI+IEGHRulgVL1tZTxRuqBQIoG0atPfQIEEDZGyxH2h0bSDfWSRa+WxoFYkk7In7xm9wMD0J
G4yzEDDVY/9rtGgHx4zyDILqphn1Y6qDsIntTPNewpDnNyfbqN9YyHfsO2NUfnja3JiCdAxBLoOt
WYlhzSNtVjbeU6LWgd9nAehV9x+Xp8Np8wlNa+WIhkrM+xp6+slVycM0WYMkF4QAKqRfVsux2NbG
tN6WCasJbC4R4HBRZJH3YbwG1+WGyKFMCHp0sJObXRUdpIck4CtmHp7Mc7uPykvSawdy+g4CmMw4
9vWYlceZNw6QuhrYgc7Yb/CBhseWlgLeTeBhJNq9YbKc4CcEGyJSbB0UBRg6/iXf6DC4I8Awdzd7
qA3j9g3rdUyQ8+qMByIuRU2DThRkqfsLW21j/nwQ0D7B/ciyrtaVO5wz/DqJngkm3LkRTsAw/Cc8
Dm3Vaw/Iwk/kHi2Cdjsr1ELb4gjpsq471QUaoj5yq+/3qc/tH3caocw428kXT7zKv5kpktFuCMQQ
yk4r+WqShZyVI/j1OGPEdSzg6GLLfPCC0W5N14w7nxYsQD8ogoIwF60JFvGyjvY0QzVGPMiq8dDv
hsNlTmnm78LNKxqhBN2GL5xiBIrITZ3sst2M/42AS+kEEzWJqkv2s+l2eMCNJ12HaMeQb9q1fhmD
qbXRLt8GjasW+mrDaO1mvouWd9v2M1loRBDw0Pk/3RYb3iY3b+GxlSG0Yz9B58FKEXFogEJEsZjA
POlhoySHZFS1ZAXOcEBZcG65oRw0DAO/HljoSfDRZQqiRbtggYC71IdeIClf37ZXG5pa/HjNYTyz
bdbC3HR227+Z1OtNL/MmbHpHx13WlGVfmdfLD18w24hUjllkGZuEN7LxVVtv8p9eK5GmMOjO+r39
VEMKyBvrG8kAZRIsJiM100lHm/qnxcb//I27HLLzzRdTItWx13FTqJtwnzBz8etEgtFw+71bKlXd
tCsCanIER/SNlQdbVdiV0oH6u7bDGd8m05UHWiZ6p1TswZeOk1xmxFzWbe6uyXYrq8wCcJdIeaw7
2yqG5lvNYdLGm2TJumV2rpwjt/2k0gmJw8clTsT16JVPLxhI7M1OOHcxUL4THkirb5zQ1ceX07sy
OFpp6xbMPj1KbC0nqA2Abe0qPAna6mDtiMTkdoaChrZnu/L/NGO9wpTyRYBzpBE/yt173wvMXkjv
bVsMh8+CY5aJ1xsqgelf+0ecFbMKYlXcoQg5BGYsGyMqtFjSDXAFLmXO0zLEOWQD/DBgPI+LU7j+
MkBe/Bu/RFMYq/9hJ1K1m1nd61uEg/+5lldNnhE/T8bYKRt0qFuI+gQp3tulSgX8zc/vZa+gAkGf
OIq5uzR8u+2Ie5qozV3TqtTycGp+jtbgc4qk6GNEYANRLxuRkmNpAAXVNPUKw8Nv22FV/9wUKzUP
Xkr4TYKIItbksmwa6nlkDs2NEh+6oNmajBRePEpIsFfFqbkTKu7oJcnaEXtjClMxxrzfza91BIJQ
yc0jCxnpfgusyeAYfeZc6glgpXtW+wJqcbM47I3Ahme0ihQX1YArmwykJsDueBGB1O7NAVxX85Wg
/LfLpxMDkMlnXpltB46kYRUtRTdV3+7lENxG06SCFctqbbB/Zveg+dZLiHyv6GXxW2lguzBv+Noa
AmTL2Im/PxPeS4lSNYksd1kVmXAVXShT5mBb919yb/XWjbPb4jLnp+TwLjx7YTT222tFB4iPDQxb
wJDMwX6SX6R1YBO6WJ08tNPwNe4ODh77TkYtST/H3oQGHXvXuScbKEX+UEHje8ZYWf5E2NcQqyM8
www6IB9MImc3a4CKej4przdk2Evf5y3vL/KhA+BqbkGUA0dDFUEvCUqagE3WLJVhb91h0fdK4rVs
zGsb4pod9mO3LEa1a1pp1rC849tn2bzjJjiPK482/zkKudVGTjSN9aje+GxmVIqe3GGCb1c45Vm0
flTI5Ox+G2IyHaEvCYQh83cAopuCUNdfqfx+0W9hOGn/XfymESV+my+7ALkMotpyrWD9DPG6hPu/
rf41eZpApGGvHy5mfwt+nrsh04Wzx+CLU+Mx27mfc/0OyLLcttJFo53XyfDMrKsK/HzEMAnysj1K
/uab13xStXBBTQFYQ0Imzh4ruprU0Tuv5PSweVb2Y86/tux6QsB9kpe3hvOvRikGy0bOYVUywvtT
r1542dtCK/I3hRsyzM5QF7T9f+z2alte0ghiX0B34ua0Tot5BFHs6Wh2WJXan6EeKrhSx/AJLhdW
NqzB3S9zFdHoXFljWqiVc+TYCvRCj0pFXMA/IE93tyfiYcnN6MQhOjkDsgg69cmv3CDejvgXXg8L
TEHlDKY2iDjlxX3CTTr6jJ92/AtfPWiE3QU90X7L7BMLISUdxd7sVBV250ZKo3qwOSbY4yRbEJ0F
o6Vv2G83vOk4uLFxydOChZYi5NaiYEve7ooCRh+KHBDjKE4bf5P3fmpxJSiWORZNF659sB07suPA
KjThnhhjiXImx5AkXzN67deHvNUplnMhT1JiGFoBW0rGUuDN3LsYfwxodNk74rn9Mqjg0QOOHygd
MOP7oZD5j0Yl+DppYCfY+ig/qvppYX97QAEjA2aRGWmM9JJdOqze09BUE/CnjZDlnaFYXJmHp7In
WmYxu1hgJqqtwnRXOHtqjL++UACbJ5MwreY+doL0eKwlFZkWDDZhYwkyi84Nj5AIaxrFgURtVFMF
dhWjP7Te3cxvfL3SToMOzITyqT4Xs8rzMNM9a0/6y8AsWV9+dp60gEGFcATyzPhxsFYwNgXilVYV
LtjfIFJgiFocwRKbTu49RfEUVD/UEJ7hkjFyrhZVig6AqaYZITCvzgidgK7IBhWZfCD1M4P9+uMy
OhJ7Wnq5NrVPQTI/JndYoubPFYUe8C7aRlpiMcWh1nafrRicZYFaHkzhwkktkYdh6r+vkQ7l3qqE
Lb8JJZiMol8nkmHvMCUH+8OpqJS/x4JjBokDdRE1wxvs/lhI3RTP/kMz4jMrXAazkV+ux4kYI5wb
oV7xGfXuHRJvsviTLLt55m4MfO/ChFmMfva1ucNASyQn+RcKcGUIrYCd3fwj3B5IOL6he2Rbtf0J
zMI0mqo1ahTA7I7Clh853IXtv6HMU2p3Zx8XNBXdOhDVwioPLvHh1MhJuD/aq970QqigqnSEeXBX
5ilS2E/Y/+B7Oaeh4WWd5hqNunE8fCQWb3Tg2lRYuYY1FJ+sKulciGKoldxHxEHVa13DdIB2bSYw
kbQIyUS6irigMG8M0GTQoDBtu3d9izuNDnS6a3za3C3DSdrKg/dA1fESTJLtn238+0aELkDuAmDA
jNWDiFbOum5yyL6mZKBMyluVHlX5/wzCHU9WnRz3D7Yl66/rTS/Zj+vESKHG+LyJwGZ330pfTJ2g
H6dVhB+ycudPoNpl4Jyq3cB8cb8pFL/L15aetulg0m73qE8MwQwcZVS7Xg6K31lqoa8aqenZlG4x
FDoJiuC+EeUeE7bi53npy9/riKBvPWT8kVpoatVeJjrqEPefm5k/MZ8V+ZWnqR50sBd2iDNsf8ok
bdqoZG4xXAj7Ub2ieUNwS65gRwI83aDnNzlnixQeHj49AUjmUhPWPNZT4DyZah/QU9WFKGCSbtvY
XabzzcKjJHcajnOm3m7fs/nJmRl55Uys7N9RO6Vl366nfbyTCJD005aECu0S/t6Zdu2sWvZIN9l0
YJi2hxECaBXBvOINJ2RlSav9EHYRMSa0xk7KGcRSra9z0wi+efDZInxE3GLuY61TeuvQBNMdVt3z
K/w4IPk9LuOqCeagg6XqtZA0KyuI4qPz4Lz1CbsLen7rsV2X9Wj6T5UmEXbjHzKcF+QOVUcJmleg
hb+Jb74XyZB69KgcezPE5n5o8Y7i6bn/b7TfVt6E7i3Fba2QY+VeOj9CIQCSDFBOHNIEdH0MezyG
0Fz8b70ntTJC6Wjj9UdCF9DxxzHFXAQeYvJCGr3ddzreS4xRK76BKA/E3CiAIx1gzZIlABiD7VP1
zcyyn6IiN5JdGxYG2TpOhuk1U4aty4JPtRBg/Zm8soHxJ9yyV1pmTKqPNtRhENwvDy19nXvkfeWh
0wWkuX0Kk2D8XyGiOmXRe2F3pst4998m6FVAVDWlJI/VlEX3PFbkrPuABBB8NMR4xJjyNSe8KU3o
ZBhoOvZrZnbScJUrQ5Ey/4pzqvqThhN3RQCCJHOM44cHVUbueCEb/YW+LEcL41VHSXOyvlabPfCR
orf6l5bQjFRaDuSpKNBqCiOsRl4j5pLUDdoAaGwm36M6UHMXB313eUd6UhQkvwawfzmbJGGk6mUJ
YZODJA469MIkj0u0I5UHFx/4Bsq26pBAYxDQzibYTzeD2xRlmA5SY8VP99Q0jIhRU5feZEou5EtO
vkXb5LC7/kPzJIcXgfAK/0Ahomp/8fnC1lK4TaiXff/lpFgSEeQdZBgrJHMCJwJeGVKFLquU6TR7
m92ijVJhU8zD/YA67yXHMLI7F61y75kHEzEcswHJHzWgHE+b/KArUma8ccoi9AMLhSMNGqvcgats
bertfOwGRB5SuEmmIbZt8boyG2BvYRGLC0mqVAxXXGgDfszYqH9y7RqFPVIm/fUTfxjetd49CX4a
9r9rW/2T/z62FRB4/jLHb+q5LrXlJ2MriEqM3c7q/6u5R5awuBVH7lPfTVVOlsE+Xv5KkpAUUCjf
psep6SKIJ4bJfC5542jBtER0siqWfGVA8KFPpOlQdAuIUMPlwNZX34sU/eHtxeW3fll3fGihzRJt
NK5jgsF40w4+Q+Ove7KhekuX4GnUqb3Kn21PdyBCI5BGGWk0k4Pd3i0bP9X2mBxz2jpRBHCGLSXR
Zn7T0/XHfY2uOr88XCLTV83lYplMJaUcZIVtxeGDusJzGd05x6oyGFSMaOqGRWLXBPlhfdwC04zv
gr7KNrB4pXb5ygYpUDyZos38yZaYTxaE1lPAkMvUJyDwsUeanYMjA6RPa9NEYn0vIVlU/0pEyMCV
7Tet6iQsLoS/odHSd3f2HSY42itg+bQfjihI952GBC5fCCC952iWaKG1Pdu9zxdUjaeK5bid0ycO
s3CVI4SJP45xLKA9XScr8haxsUviDkuB5SrsfOdkt5SIgP8NJUdq1qOg+DibC07ZcxVAXC16Lu49
jodXuPnG+pSqvK0mytKCttC7nkJHV8ucCQvy9WAeaR0YZHJFQK8SXlxPwrEorNE8ApgVyefshYZF
PbW8hZSxtaQRJSYMOxR/t+ZhU9r72+1jzItOWMsC/0EtlKcuOt0qPVQ/nXjOvQnAtRn0DFpSa3XT
duh/0itUgZ/wupltUEobjLh8C65h6D8+pjuAUz6Uoi8QEXMiweDdIqFDHAdewe4TGxUaaHvwglYn
7C79aGfE/O8G0kX/PKnso3CeMuAXq75BuB5hQKpyjbLxfojZd1FCFMQReh1r5YFS5MgL9ph4EeW5
KyJ97QQzwUCVnpD+kUufhgWORwBaI2QT7JZTL6UDAR7bnPYC3iRIdU7pdKb3dbXLW+ODAuj0E3ld
07ggJNPfJaAtDPhV8G1eEvLxi67SVilP350LrLMlC67hiz/YMNMjdvG/2mWt9SuxI/eC/9K2hSqi
GQgTOXnrDtBx3b9Qgkgpenq4fAt6stTtvZJhT3zG2fu1NJCDTfBCfZQW9lRW/L8fwplGJDWWiy+F
LnwyqIbbubmTQhu3ZPVeSwYOxJdjWnoQdtpZTHkEyoJW7lA72a55loEtAfnSZrJTI2P4Sx0ts9gv
0QZ6PvevCAaboxRHqjKoujBtnmns+vhXKk1SX3aRMKDZ1iJ7+KhpWZK5pcNiHOa+AZlD6kiitcIm
jAoGTH7pJQaswilFtmU0eIprnQfwrVWTs06jNQMLrj6hGjWDR4q6CHucSqZziMosEznuo445GErJ
X8V66neeej1azd1Yy7TVIpFQHqsZIeCVPY8sKS5YL8yaw3AKYKB0kphPTvz/1U9pTjar5JXhYQQc
Ndei8qk9ZqP2G1DM+Cx+q7vtAallZGHYpY0GXWQRxfbW0O89Hu63u31sHMXlXEmkWmmOunZ8EWv/
eQfJJqm4/rsIkrE1lID9tLhOCZn2FMDUpG29TgWKZNNa5uuuxvclN25v80Y486JpHBz9SS87aKWb
Pu7+sAJ8TbA5fSLAZpb8Dltw3kK0pXWO/0SsMXGQkM5M0e37ZHfNcs55hx/m2V35QAo0D2TYWtYV
XlmTcKWjjJtUcfpOFlWrwgL+vDu8bK9g2DJcxlga83gVG9AbXVAC3T9FZmsTfiv+SNHPqQyq4hIe
vaIeNapDaLgVR9ZaUdKkiBSdfRBExuyqL0aJhkewysEJxL65GJtuqkH3KhUpBuvhulK/equiNA9J
WfR/uUZ/FbDGySSPWIlysr+l1BlRQi91Ui3gm4ynMIsUh1LGtv9O7wuOse0aG+LxvDdBZ6nAClaF
o+eGY9YffvrOlST6j3mBiM4wYs/wc2yIu90lFFBz6W520xVjgnhipiNKspawdQDK8ym/QzMc5Xnx
BNbH5n+QZANhmIqonUTCqe7mN36fFgHrep1PiyzWm8qb1iwx7ci/SjPrIgYI9G/BRbgMtThgGcWp
TPIsCy3GI5UWRIYUI1ZUkJjhZx7dGkOdtxkgTI1IJ3bH6c+1I59eRVMb4u5UVnuQn54kTLq1wihk
VCJB4XdR1SH/PBPTqXUNgURTKqsUxsCFEAfTSH560kjB4T2BvvIHZdk79JBfE09lXi+sO5189mv/
2YM/rH+ECJz+ocSdhsOsqJfjMRl4g5Yll411oFkidUdt2Ni1kTJdHyNq1h+BL6B2oWU2qhRWQfpF
APGoqa1fc54/AQ2eI7mGoHvBNMF5q28mddxFlH4NbDleZXv175EPwEPUfgZh0fsnYixeYQpxKEcd
NfDddqqkOEsQXCpYw5g8Eb7TPxxRMX6H+oyqjiWI+sINLW5RzsM8il9btytPLh6Oh5I7MRJG+uPr
PgwIlXyIJNAw8neSQJQaV4M/9AQbkujrqW6u78YK3DLgyxPk0SWXez6QCT3U+OkmSlmSdkPAb268
a1gOa6528QeQzJ+O7sWl4EhyboxImGoE5qCYx2kwaJI9HynWtMg5vLfyQU+cfkpeDLBxsa3J2Ua2
MjCOvK9SglUVOK1P2n9tgU40iOixupZELNRYZ9jvYgW9o4vImJGWN/8+68f4fS7ANrrGmSY6D818
EMEehIBblUL5VphQBzu87qK1bhIIGGAEM2JMPkqGDg0rdvVq4bTadmqouEb9NErgQlvRUXvWeUSH
jyBgYk52Us8Npk+Akzm2JjKhW0uANHf0sZxfgFf4N0Fc1R9/dZtcsy1QwZOLhIFyHTm9neT9mRDD
LwHe4gq6wNYQMiubuQ2QormJrxFoUW7sWGHe5pwqopHHYr7HCs/VlpHTvSsXstnEJvHnLJJdO7W1
F/SeUjup1eAktHeZoHoL1H8lEbik/fby1/zJZuS/oQkTjS2TrVHFxXK0v96jGI8L2Z1C7ipshUhH
W5gDlwvhQUkuqQBJUuFTporOV6gRja87fCo8EBoEXDBq1iIxG08uEds2kaGUzx9XLrCoqFpTyDB0
hZMWBsDd0wXGHs+B1l6On8a39CU5eCbaTFeCt+zH2f+v7Q4n8Z891hAwiZTNhXEvJlpI/AIuMAg3
7eJ8KfyFRMZSIcwcT7BpYmnt/aTqlYpJ8MScdBEX2mG0SfZT46Up7yP+LpyzaUt172Id6l8pc+WA
1RRqOX9BeKLd1KUtXrZqCAfgVUove7WNUVkW2Xsk8JHPoevD8cBqGEvVuglHY18drq8ihG0+g4+y
2+cIDmc7TGAJTGVo/umMNQBbvpnVJPPKQePR3/AysBSn9Ggkj6S36ItkSjrJyApMiJIwaiplx84l
QYVAFGoJIOFzua0QNAQMKeVDHNsjdE7/dmYtNmdBF0/9ce5dnUZNg3Iba9vEjQY+U87VdRIEu+0j
y1zFM0XPXYPCRCPMERU8+RZ9MNS+sjF14AP1L0Gabn8rGupfi55I4M2DecUdLUZ1Rt0QQDEM9G1a
bSDHKDDkxJ8ybeaCCeoFNJOen6dg7L1lRMR4yQW1QN6oDOf8J4ad6USZ9LDnsJmEli0bqq+g9qvf
Age00HpwDMP+JQKsr1DKZnKPm/2/qGmtEC56KEH6Piuy/+IwoTQ5r6SIXKGRN5uo+t8DnsddsBO1
8Brgd4ziSKRnbJAVkaF2nH0zMRki+uMsshd4Zlc+iGXbCLs3aWH00eHuENIWQ21AsoJ54Q54/ZPj
96nbd7pdPXjBVJpxwxPZFAmjQhUA6+rkVs4AcqCVgZbFrIiR9UUt3IRTZojodBidc6fphlt35Ke5
3FL5PNQ77OhAWmP0FlkaF9QoiSoj2yzu0ZvJcJnw7LeoYexkvFPyxh0z2Gi75560s50xXrDslCBp
C3Xb6ryw6JRctE4efLQdp3FXHuD188j6eIM2b9ZNfXNnPhbU5bFMlq+fAlPchGMl/RtzmfHXz6WH
sZxyNfF0kyst1Jn9lkCX73MZd501OQ1EH/BRu1kBvzQmRqcXrg07C2qbwmPgxsLG4ORk3IGYwzDR
JAeDI4w1snrlLtFWs7ftKIDXFlxg6StWoU70scTQAkpTyVtPM5cerQHO+h/f3ATGCzWnLPKptX1C
x1CGFWGjJssJzR4bjfgVYXVPGHUNr9pDop1qkrDU5q4XCbj2FeH1TPo26nvDkYp9U0ovIkWdZVj6
pcsWuNRevKIIbkfShiCsfFOGEj8v4PqW5HlJJ/VRUGhJbpqTUZWEkH9T2z7gfTRUG/5sIPb7ehQz
uitmZ5i4DrSOLyy51LyLBj3FdTHJaGZnHGPO58oS0NNtIcioaK5YTymwTodlaD4xpekHR3j8MD/X
/wMLZykWXHLGhDmJDZfeSCWd8XmqLQQTlQ7NfriRtOsIZ31PgS5D8BnVjDGKHXhstTDFGtnDcfRU
pEOLA0BzgeUqJHVvXqOm62W7JhC1QGxHv5RgGDUEmm943Il8qvpPg3NKXNxS8TFv1lAY0LUl4miV
pTqM8yhFIyF9yIaibP8bIb6AhTJM6Pnkpn5+e/v8mmH0HRPJ22Yghb9IuzOKOCyMEfuBNwMe416W
ac7iegfMW7uHZq2YPILj5ccCV9vvudqWok7RIs+5zBljFDm5l6aX5VhJmsTMnl2kDP/0nwy4DpSM
uHWzWwwEUEv81c1mC5uYou/3RGbGRXm0UYvA2a9PYOUIIB7Jef1fr1/81HM6YWvPOjgryiSN8HZw
esBFeDoTs1taCsP9Ug7bfxNN8S059b0XCKYqH2W1+wB44HXxQq3H7jKMfT2N1RFOkpl7QYJjbBoT
mYFeloFIF6zPIUpoEpMflLptLimYGIFESN5CQ97vol4kziQeyTIq+bGlx9/bRlPKaiKhdqr2ZT4l
TNv2WGmkkwDXwxSCzMTz2xmk9oCzLHfPPyCtWovUWeQi+CGFvE10kPCwC+426i516vMbhDEcRcD/
oDFyg0lVsGw9BVP5UkcvQDF4MMfqadlUvK2TkhMLv7ZJFviDJ4RC/I2Jp1yI0okLmhy6STkQIgmz
KgJ7tnxzUO7Hh4ilJsz3c78L7GonHGnWsBzseBE4WzspuSIIzGuYJj9Y9rDnRC/8yY7q1j1OOY8p
498RSf1vSnoaTDbIwDSc3CwcLKJV3rsV46dtRHTJjA8nzWUTL86FNDEOarhY2YYOe9y8YTxqRqHV
6s8ATRNExZZ7ZuSVzrdyPup9kZR++d/O+L3tQQgZTrVWC5o+Rnhk6ST8CAVNsOjos9pZ2QIgbYwR
MSFEexXMFsg1IyRPiNo2RYafAOPmOpQRNm1yKigAinQ0lHKYoYK5lcckW+BaT7hozAuM04rrGszX
C/oQBuEezfsq7P702vAkrDAKJsJQRo0YyrApuiJWRLQYZNZT2QNDcZTeQsDGvtc2bclngnsh7WHK
+VY/HeRfkpaL6swzxeiqUJeLgWQ3hOjYO9tAlJlqlnBTzIoODyAbmWxsXoPVNyz8oLW01SDPGgqc
JxJbNA09hJPCG7tyGyg9XtllNesx7lJmAmtcJfx2TI090ei08AoZfKmNV+dAUA2KuP4maZ3pfR52
FKkPaQDWLeFKaqesiUG43348oc3DZWAzj7XoqoBuBZNYgdATX/g7XqMbV2TtM8pN0xjucvKwIiFI
U4VUgaI6MPttIv6j0U6xgyl1KRluRp/N0SXCVGOm0N2KwcRR1NC4Rm354CbDmzpiPEEwoLVWz1H6
Wx52K6nZTO497oVL3e0p90w7ZjKSNqZaKwgLp9ur3TzS13KjwcGOt3OqUHkrZRz1AnoUFI9GRbDj
FsFU+Ldi6FkPi4w0tLErUZyXQS+Z/3JZS2O3U8UtwcLEDTHet7t0MRYjBNu+wNpzgaWPa06CDVxH
GVmNN1n2xDtMzu+G90mgSoHZJxC51FyL8VXAk+bOzsMlzY2ufAXQu1BMVHRavhru3IiEVOYWDpGr
qWikYt4PqdKpQevpR3KdMPo+qmED/n6MosRYAPpxTwNjFsqj7/wdd87Hr49jnBbIJP2u4vH4eA71
7doEdf8uJ9BLKoTiH2W3IqHNz9vNGulPh7OCSkKMzbFCoWsSc1c63W2aVd+CNJBi+cmq9QcOEH2y
6t+HGz3UeSblc6klmNG20sA4p0FTszXg3NtsJFRDZX3iOWrN81qiltgOYStygaCgtz2mDGV0mnCd
ScqMHM5MeBCmoIP1tZN5Ll+g/gtysrbtSCR1hJtYigRbXvQvXicNwrzFlFdqJ8G+gX7zxP9z2QK7
PdsHt7xrdrzIURn/wJq5bChXm+RD9NOzfvsvaORv2IECirhDEYvzOk6XagHQNDfhwaAsWUyHzIgZ
p056AFrrD+tA9EJooZGqjAldfT9+2LNgfXYIqqGzBjMJiouif7/WQ6RTbI19nIm9CVNh7xByi1XU
YrvaxBS9Lv4tFJXZq0qvE8b5fOAwkjreAvslA4RCIOXox1Sc5HTIZPYqAiA4b2b6HdX/265ba/mp
fdhOb8l7zMpP6ZzShuuvDnmAknJcUM7xlYffXnPqOaC33eIOdcWQi3m/73qR9G7hIVLtHACijF47
VvQU+kOU6tIm2l9dbACEVYgWDinFijjpxKE2sSpvteMXfq16yC/Zf3mrBgaqAGLGjx5NdPJoPnuk
dhAW9BKwuOQX//n2qbFG5096ogMDE4N9TkQGYJx0u0ZQeBIbLCwzC5iYf4vpw8+E5IcZJ7qY+Dos
pfIGZuIHVfnF2Om34FHSCOe6SSetPR/TBuq75wM47qOb3klB9XlmU/LorP4uOst2Uh/BaV6+mgmH
D5DjzRtSVcZOijpH/CqUyszPFbxFLnhEoxJ9+9bAw4gMVZS0FAycfOrFO3rAyUFBWy3JDlUX0MFo
BnxzI2iAHRnKZm6+oB/tcJJ6RfbKLYh7ggUz7SzHsEbp2VhYz9B6xDMRnSkFdMEtsc79nGzCJGrx
r33zeUTbr4hLBnG7pUe3pCOJ87eYCmPNclmHFEcT7VlO1nk4lTfNVZHOSOGseg8BfnSQw+hUDx1h
TRCN0S4E1Zrp5xJZclX4bbQnCddsx7HwzYNMM3LlBdHgh2zykPidPIHJqKHlCjQReProBm1v/yxY
i7W6RcVwwcPM/DbmJwE0xICdopXX67VyZ3NPlhNpgWlV5XuyldyIL0qSGPnx4CMqjSjF3Qg1ZF+n
4uVd1kG6jFblF9i+SZO4dz8pdVWJxTGpNrSnxgRFCCi6z9PcB1KVOs5O+0y7Nvx2ITkfKIw3Zox9
Ek+Fy2Is5EC8sCENNnIVYy9wi4/RLrUebpJCV2GFwgPzctEHqWh5gp91byiVRnGlTWzMJzqFEW3C
SyCGFjJ5sViqELb9vA1xZAvYHfTKr9Cd6zZEta5g0u0R8FE861Tcy1UW7z+yDtHECpsIHuWg/UsB
HJc1UFNK/SHxRBDJAsBFY9FE7b/v+YyFP1zpHRZYuJT2lT5M3BLj5UJJYjrquvInlF32UH5W6khY
y+l+mpnlhgmorz4QKhrwXowhb0ploEP3fAIGQPGEKLfW/O+PeEDJcx7VfOBZXGddXojDnUc1UE69
aicMU5xXrPPJQj+1Fd7twroh3t8SZzivTfaKs4zkzgUmO/1QXd6KZpb0Hq/hBe+dU64X1aIGjaG8
wMqBBjYOnoKBl7KPHHf9G1YF5eH0ER4kpYMeLfvoiHE4MGSE8SITbK1vxNRK95jTi260CFeR/TtK
T9hOSYlpQZ4Lxtp1Vy7JydvGuP6uGV28UfXcQbMUvzH8fzi355061gxqwZoVtvlyGSeb83Lwju7v
I6648E0y//0HaZ4dJHevxGmQbVb92ZSz9hIqIoMmP/3FrIUd93VRjN9ebgJWBuMpIWpPRNOdw2yc
PORk0kv4wV4Ktis/EXRycS8CdeAdmBE8QS0qajerZEm5ZMr+FdBEt63rbqh27ke9NsWbFyodxxoq
yk+Q+Q2dSZ4W7YBs3ISzzgsGr78Ojyt+hRA0Qi5VV8Hq5hnhSANo2Uj9gJOcRcbNRAjA60ILM6p0
xiTllpPJ9SnLnGGCfLH/PFUYdJEn5yxgSToNNuG0SUfyzNjFTW3owblroGrKA2vcRm+uzyC2E0tw
tFGg2TYaOFsKgvfVCStY58Y2ezV5ykR2njj3vRIaF1nvkSXmUYyGv1puoEmVPYoSwYsu76EniByu
36PB39IPPAtahLGETN5yed0qKnVz+ZPMrvwR/oSIVm1Q1k5SZVC5BZMIvjyoY9vsz47wtuOulCPj
N2/IkCFNKjncn/mEeO36/7R8t0qgXQSVa307coTXdoSfLLBSR3J1YoOmlRwbL82lAwrvJ0pz1kIh
a1czvrms757JfgLNeAkQGF/6VC2otG8uR3+BLdmmaBt7jf3VZdipg16ooOgHXsKhxYJ5BnCIdYXn
pIvuwS0byEmTVGcS3qrPWTOGCd4ndoQc1flTFuM561ROvp4biExDNst2iFKBQ8L5wRVlWPqm0TRO
NtHpVJD6itQb7bTtERe/zcRWCOTSpjYb5mRQKREQULYRvCJOP81vQ4fTkrqK9BaKfvB65cefyMR4
wLgP6KDqgn7JDdQD+pFxrhrnq6tUQxG2J44hVPx0hiKXeQpJHa7zHPajfDxGH8InqWdQrIuQXs+8
fdDPMtBy6u2SaFcyN2gIl82rUXMg9Ikc0+WjfUu1JcwzGN08/HGUibDodfdpxorGiRk2kM58gi7G
EIrYMDVbbXEGKOYiWFD7oRDnv+zlnQCCHrzWCcZkTbsK8Rn1SG60Ry9OyzJQL230KV2+8Lqnd3bF
ym4eL5Ym9W8hrR0tcUG4h1/czLlXT9Z0pHhYD4CP6LPW6PguhxWxIHg+IDERL6VMgbsdiTR/ZOc4
CsRWz+LHcHAj1C8N+VAQ0Cd+XoH4n53+ulu9BurLsUOsaBK/+tr55NLcHzFgzPqNP/ltD3Cu2B5F
EOi1f5/1vqlNXhIG4alcARedyrkT+9Mo75FDVFWPsUL6lOS8+8i+MvVWzBn+nl+MRk9219numChb
W66RiCQC0nvbBe3NFu91X8rcoSj1psRITDo66v9GGNuRFEYfyAT8Ql3eIT5o4yahmGK77QWm5kzE
Ox4/kMhiUORevQMvIz5XCMHtq2jxniw1GnPkjL/NtYRXvYcducmvAxqbAvRcH859dsYKem6ifNug
Qs74FoamlDfgIHeIvIw5NrlRXecHNGlVnEmwg/XNoW95zvZVZKKhzRD656o9LRRoGcU8qgH68Cq9
ksokmBcPgfnKt+q3e0oOOxdmdidsXZMMT3SYYxkGvK8l7uu/ePLIOfKpS4y+y2NluWPuIj1Mo+bJ
0t1d0Yy6GVM3fiRGcsFSCVx4RI/MFP3CMQk+VdMPBevJyBqgPtwNXdR+xicPXlR7ljlm5afeHU5Z
zey0YWUszgNjSUh0suS/gsbGvCawuUqYyF5Fle1Bl8Hhe6iwe7ekoAX/rrGvMbh/8cHlCcvWhp+Q
yddrWZx/8MKndber6QOxz4dj1uAK7Bi7NfXezXx2xF0TvtDcYVQ3idp+L3yH0YAgtJ9ZnqJt5Q3X
BZ14srk2YDfEKQarTx4Zwu3zRoeerEr2mbZTUXzjYfYQgFx3Z1nvXhnzyVWin9VDCYxHsi6ReccD
5RXGqJt1djDfBQC9uIs06qe3oeVaH1g/0J2nUtEapdXXX+1vU+tQ0LbXAAHoVcGpGS//BTgVRMTx
8fbpRxG00x4gVb/trvpl0r64qzNpfiFRpeQS1k+vmsN8rXABXliU7WWYs0tv6Y9TPS0lqqdGUzTA
qEDv3VJnR7uLJE9mmHj6foL542VQg2mW17VQ4Qrb5ojtH1kq2ayYEFxtrzvJ1Jy6lGW3r9AvzbWv
ysPu4KDvCSpEzJNYX91II6iAD8rw5zri3YZHQpg0GOzmoMwzLXuRQ98VaP8oRtlfKyVpPK/9yr3K
9wCJxWYTJcrEoUJHEU14DCko2g43l9CeY1WcsZLCAmDYUUp8PVpUb0coiSQeviAvRZQoStpaqwLL
TaF0OP3JPNFDJSA5Vffv8V394WPj9cwOwUcvaKhaTSXZbiYO65YvRJLBkel8CFHK0f9jT0potY6a
joekNPmGyDIguXtpX/AAq4wpss288nNhCRuP+9SKpY+KRPXh5/cI75AqYOSUsCV4Lt3GN9P7jPeS
Cm0/sRpTAX334pFOzzwxCnn8FgGdGgrTZvHGFx+992GlP8f/Gg8lkvFgOu3LzTxVRiHkgw0RK1ny
psNI7kvK+Y3EP6oKIdYdt01T42yTlU8DG5vjeH9Ds5swKFUIWuFh944XVge01rsl0NLjst3J0YiT
fJp4Im4lUhCTBc0DBIGwf3uCGXIC7YjjVuGeF3xI0+r8Kt5ZZCPaAs8JdtDlzrad9Tn9vUWqBZeR
rxb4W79yCjh3GZUBKBiUjN7IMV2OZII+N/QKdkJhhnNBwOreUouLv3tvQRe+YA3TKqtJwrXX8sV/
v4j/P/NyqZvuMkuozP6Ji2Fxz6gEQi+MU6fsQGmhCgBspJ+DZWe5R9aIo0EBC2KObQOo/B10kCea
UWxpbiF2I6WY9gy9m41eQQB0gORLBkTiugC5YKHoGo1LJsssx5A/u1Wvfpw0yOv1KFWqV6AVWjul
Fe9YbD3/cy5/ZElzQcanCJRNqfzDBOUgPqMK2rlkehohNsN5fr5t+HsApdEpIapWiMBFTrTSeZJ6
eJ9lPbtyoAsnhSOHzgW4sfpbVN0kTOYZEpr1VK9PaOtKCgRbkErcB5Sthg2279Jjb+KozfE6jZ19
blkw5TEpAf5pezsNFR2D9b9dC38UutVBOUdeJPfOQjTnmPJM7WbBbl+sgUIw+8hCTkHYl0Ydj424
Lmv/45BolkDDuBwKyG2ncGPfRrWf7iFXtPeDen1+SZH0Xk9WWQRHYlZZ9mbudnsP63rAsReQKLiC
MoRijHnynTUon28bBuiMcrSDsvY6tEBmc9uJWsmZ3SldL0lhtrZdC1pPSPBLdlsFRGUIMpheZ2Wv
5Kjm2Gsud5zeRhI8A9IniDtHUT7mZjtrSItfo2+igNr+ihKVgwokpLdxA7lrZn+tVB2xZWqC3Wob
8IkmKvqGElPS2yYV/WBWIqcqoyAF4fJ0VRIXJvV1/JMQ6TXUBI+FK3Ws6hmKF/H6JhXNoGEh90DK
pzTBobZEe17cf5C5qM8Bkk3zWu30MMIOkCRQ6Iv05qOz7xnwTLRK8W2TIuBrGFYi0tN3dFQy+AXs
cgATSHnSje+oT15kgUWPsORaZe2Lgf+McPIZhWUil7/2GTn7MWoTwtlCZpTZJkEoTK49jVwUnYh5
eUpW9YnNYefuivyJjJhFLb4nepUmoQiLw98NeijIb+/cCic/JVDzDyE8qZKRuGSiwf893wluG41t
VXai7ivb6F1CIyBIcyPltoLZjibrxZ4aV+u+jl2SwhevmdlM+VHvhWiTPQfncDery5+snK7ObLzp
bArE/ssyW+tfZ9JEPaT34Fl5jaPyfz8DHHxSSetgIz75cO87xw8N4RTra1GX5sPFfTRM4HCoV0x6
Qmk7dsF+qsfhEmlfB4DdV3oc7JAFb4+tqBfIISqiYLUA4aceGvZZekFCrG3yGX7xhPFS4ZcaWwGX
Hp1WNJmfXSWCSs+tYP2kGiBhOBNQrfDtPe/f8YbBHIf69t7Ju+slZaV/7z4jmD3Vho5Zx55zLy82
xqSjDHQ9LslHgbVd5RjEs+wvBM0XGciVglbj26gnxry10T30VCWaPsiqTsjSh4ixo/y7pmW8XQ9a
2L3GofxsZd6DVXwvRwc5kXwdH/BsCxnXunlz/IS78WPE5IQBGIVcP1PpO+rahSK5ryFYJ3/ZMow5
llt6WOEcblGDyp9F0I0xd2L2U1FAgbzcR3A3/Z3ccsOgcxLUh/8z9a81jtx7jUKgrEsIcjs4zvcB
nNLGphYW42hA3A86xKcWO0DK7wuruFwZbGlIlLG0J0N0Ki7XmtRzQLYRagqBeuHmp9LdKf7OnJpn
WXcIogeToOCRbLy/MNs+bV9qjEuLOOZ5Ue2Tz3M+yiu/QSJyOCyRFJtGYmJeGdAACKi4CnRGRxkL
CEH/WPCtX00r6KlsXhcHF+ji4RI/jgaPnxuBEv2z9QFLW1Mfhbvk5zqfuLl8wjVcQbzyOEY6BGGr
OVuh8Wmgx5W/zxYB5S+bIkfms/LsvPov7RKIEiQFbDfJDT5y3ySU/8NWiHnYwfl/D/zeMOhZkpGI
+yLyW0ev02MZ0NsjKTFueqjyw2MUSIluI3DOvc93YVyU7GRSojWGdIMjqXIpllvgCcu4ucwJyW6l
2fONIftiOcEP7F58sIkKT5LSr8dMg9GwAaRYOnO8jGeFLyUloQ1itZ1aaQpJXCPCCmJNFBxIL+pn
fFJuNT0XVPXaVfJwvt1z3m69zEIS9yMW75xjh8icGPWCNnLmQdiUksuHuCAqxmpbd33m637DBwAS
svqz55DR5IFTnqJSDJ02v/4zZ84cWhXzacwRvcYzPNLjXnHSNbyudYqhriRIqFh3G+66GLKrLY8u
QGt9cbpNr6WkdNYxI24S0HCIwNYK9QCvpPZAEVrOxRYRRM4gALGFFD6aPKdDCJBzfhYZi9DLMYrS
WesawJ8f/2mvlOxXTcn7doq5nuGYvHs2fY3o8T0BcGo9lzI5DiBAVBnRWq/l5A6YbyHoTSav1OEl
i9Eo4WJroumfs0fuJqwjuuuooSu9aBsoPaqFtMjH5OyAoX8CCYY+HHMtIFDXRxUdHasJ17PwRTvM
MOve1gYN807tbCsJL2jLnRBkmtTuFdzKWnDTgFY/kDQU5T/zd9NUIO/BZAkkX9ga/OkeG4sNsdSp
sQa2Gy/rmxjAEmlDYggOHTxqtAZ40E2MScJ2VXesyS6gcK2zKwCynrRp+7Cvv7eAJ6RvUudVk7/1
5Tf6i0Aw4eh+sV7Q48RE7/v/DMLaU/uvPCLagi2774/E8K22lMUzPXimPQ19bVdqpzRY+WnSkWE3
aFcuHdtB1gsOJO3QIDQURpBNw/hAQGB1ZHE5OE2j1Ry1o3By3JUbxqr4HDEfJNy9Qnfgbv7eenZ4
bAN2V303T0ApmbRA27NHCSS5566OU+A/QpcBRYJLJ+wAKQbR+BZstsPMmJH+4WHrLM9PXLiX+lA8
xrtDmkm+169Fp+Ik7WE26VXRWHTQYoNcR9Oz98/34JNHrgCEUZDGh7/ROXdd7Lz9my90+ikDRuQL
TbGbFYEbnwL1IhHebxpi8G87PNLpzvvQM88hETtegJVzf20jKM0CozvRW7xyRyKP2y6B00d8m2XZ
tkQLmkm+ar1W2JqLQxb/tMLFoi0n0Tbo7PbVIP616nTFZmhyt1KK2nuqLYvIi0iScrbWGMQbmg/8
MBkp3HerWHruxsttL5+Up2FJQuyhrGTRrttaKeHhhKiMMZOfVnrrbCXYwmJXOc5DeQi6FiKdnJbe
LqTnJh6lw2UCSUXy0EvM9bdqvFRiTRmYIJPKRgPbydu3bvrNU0OUdetyRXKbPK4ZfiZEy6n51W6i
s+M65BuXxopRytx/sldQO55q3By7r7jTPD3T4L6CnK2FWjvYJ36a/FGfb7gM3E4hht1N/Tye20rz
CDYhR34y9EIcx4m7C01AAhQjs7xSEXunQLMeaKytqk3hzvsIaSWAn1eHZmbx78taCMsv133g6DcX
h6phq5jiEwwi6hTUvyhj+zGnTcM6iRABhpO32GMyM9+1p85Kj99YxZ0CyrKXvzhfnYPTITaFcAnQ
eknEKulvZDbIuXAUk99gGFJKyZaacu1rRRsvM1YKOkJwnVX/dF7bJFFZ+V+Jjd6LYgEZom6n69DY
t0EAJOKiJlvIlMQQx1zgU1HXspfvPZVTouaAM1/OwG2llg+ng05MYdJ8D1gRT5CNLpOgF+Ye3f2v
VmTSY4WoI6EtDjvSGO4aqNtz7vQDPeB+9TLBT21kC2rV+EcZS0i1DI9trqWve518QJOgfGfnpo/R
RKB/J2HsPTgnfKyBHaKkwqpHvF0LMgufn85P3oL5Fym9D48kc38JHU3jcssU3Utc72I0CZ7uAee9
iwH6Qds0UoP+K9GTqxBys/LNUAv3OS2zskKYEHgpv15vn72glR0BIa7W7IZtemD2BpL4rtPiYuoo
Dtq352GvPcbiK/MfGrYad/7Abf04kiiveJl6j4ZVLXxxAS2oeZaUfTq5pxsFHHc2vJImRp21Xufl
wQmgztiJjwG5OJ7cPbMLp+Wh7Xd5X4BWvvJ3rX/fndwTMXAvRbMKMrGiGFbfwlTSJ33kbMOH1tMd
t/MxPFH+OEi+MC7x+bEg2xY0XOt0V6Dk32mYC9HxBo1IfemX3+DGLH6+9vRzApe1qQU83lYiHrg+
nsoEqV7yKRyxoKOdYNPHfR4sEw6wSLdlKTpK6igQuNDVJP3AUD62s4WhQsHiJY4hgIoCU5f+QVId
jifMTLltUfQy2h/01psJrEvlGRxRo86CF9TO1qSGzq/s2pMBP4WzXtBHDf7YGHNT7nZBsdjLsjdu
RPCxZabQ8YiTTScajStGaMIsp385cGHUBm+5VOpquReHY/s6mroVnvw0xP9SPwukQlsdrcnqiF8k
8EyR+xFkxbUP6mGyH2A9TzGSpvAt/xTMdO6xPjbuzGOxQ4LGEvz6UJqUi3FDKkbvkZenh6RXCzRX
eglXiTRabRf3A2s4uvm5yWMXg9QBuzon9Hr/YnhxB/ikULzagYV+pdTyB+Bt7e9f/9vysDHvIP3W
CxVoZM3v34Pn/1SWohXuyTdoKQKeXDyl5a+dPoLTaqLTt8/cI7tmdzpE/od03p/hcQo09fmtar9p
QMfVMl3KGP7Q9L+zDAMlPcSepGfw0NRQJrWgOl+jXQeY2B7TyTlriG/5BjQGNrXrtfL0oy0czhUz
MrjYhQ+dTPraYalrVHhCmnxRtr9x6RuHSYAvWsdQ9bykrf+/xFlUuplwP7C1u+c1FS937/G4EUR/
QtXvl/LBvNiWDw2RJ2od4Z5t3RiAkMZ5ZFv8Su2uuW1vSucCox/snwgLYhZmLmxJSdZMNf7IH9VU
VjUn3RyRQOshey6S8m4aZBA1C9zspdHbOlfY9dQEYWCIe/VDMZrxgbpfC4FSrdV5/3tDo0Io1YUp
OjInxrUlzmzHbo97TFjOO6VQN1mpqrRJDGgbjdRMKX7so72BErRUiPV/Kj+sfFY+iwzhi387pm7I
hbz0/8YP+RJrfsMiXM/Bt2iVfLv9Y4eZwX9VEN5VkrBq0PHj2goZUmaFEMHsNSSPt0VUEmul6i9C
OOYKr/57Z27kXVeFk1Y5qPRdJBVcO0kNGdZzXkSXpui2qcyhi6m1Mtj/YA5Gqx/4JvF9AZn8XR2T
x1hg5XwtSlyBendkbyKpmywZdWHk1a38dS1WlLH5DMbl6OsclfHrW/j4MHgNibTVJ4wiYCGqz9gI
QzhaLZBf24SFH2VV6+80am96F8l0p1hRcgFy8lzMxZ3zFZphfXFwM6exUl60WVl9ApJPaeaB81rg
JwMkL1oWuEnVBeMly9dGdfDXFaOxKj79LnOpiehr/7f+ZeIixFF6rYzS9Mu0V510a6xGO1CnmdQc
XDnadmCMcPHCAkR74RPYzE8twl9zZBihS/hhOcvPwGpOccrG0AzKaq0EqEwjAvV79Whgm/ghHTpv
iuG5n0lq0yNETfu+kahMc21FWbQNLYcbnH6MYPX5SxMapWhyo2KVQWSP9ViOGgESvehgqiizgLX4
ONoiMpNv3AxzkFxfg7eVhx8TcH43Kn2mxhyR8QoJdRymUrbqd+LZHnxIcEAaMb50JIf9/rMlFZeG
gomMkxFEURC7GwdAMomn8x1OWYf4aoyYQvzkp6vkedG9tA9AjvCEV6qbfBfU8fGKc84XkOQWaT6m
kwnLz5ljX/xfkHu8VzHCxXVGgQVMqLrc4OlCrAQ5SkPFpiJo4Niabw5w9S5cPZMkhijkvC1V+AlW
TuEKL90uKxqNcOppd341kTjjsliWg+3aACsHOZ1++FXVu9trBmAmXlBWiGbcS0crueM6apWfbWRE
y9dyHlt4rPyn395d+62tUWFlb6wDYE0YJyFcnx4+ZDDzDM+uav67W769THGefjNGyj0jYyD1AtYU
p7oj8MfoRa+/0cEe9Se0N/EMNwmJ8xmYHCiC0D56RpWAv7WKXGacBhuSd6FXLovok3y9R6CPM9+7
GBPIQo4bKwizbBqitEzPd3231SPB2GUw6VIzGp2f9rsCRz5Jo7AoPUfeMDMH0mOBOWBLKq8GNfMZ
t5SGpLtdy19ISwIf8usZJQ7yVBX/wpEhAuu1FgyzxtLpEIf3EAoZNdqXe/IoBgEPXtTrD98uCwJ4
UddYSfkKpAFwKUKDKvDtO/cZ2hcuaiQh0OEtFDSlUxk6m6svb0Iuj7czEUoja9eGWwzZtvyP77tN
PQ5ez6PWW9EXRg+gSGcAFl96sktd9W4gev7K/FMF8aM4jDrzNmAXzfSKFgw1FN2mjXZ8uTJoYxBh
/cOraTH2DeK1QaZeYmb8bsmnno0Kbp8POkUMB/+D3bEvpLaFak24kuwbvaoPz+ERn0G4M51GykPG
ZaTgqm4AQY0u9yVP5OsHM8DC2rDzNleXp3CmCIsw+tyKEzIPzBAoENgY7fEDssZAQ5eoqaelRxke
BffUIFbdDvHgjKjTHU22600UhL8yESaUIMNGVrvP0A+n/O/uwSXb1H47OwAdbdNFCr9Bl715GAfU
rCP0KXY7JFMV1L8bsy37PHhMlwY8+7k+06zTUEmOaA9o9e5o/CHTconvxiBw3YKzbGjbHMIdoHfM
mnGijRYdlgRpxVe4jzeF9ZsOZdkdOzS4XtS2ZAJ93W9SPoHh++JmuFzzu1SHo3z18bQVGkzPy99Z
UJEYKKfSU8VtopSPTHXFvP8CCDHibF2ZtSCgVPRgGC6q25GHCuYGA5BMzDbCNJYnr/rmWcMgQ9kC
IgSl+0pN68ADeuhos+iU8HEP0Hbk8Rux4FwM6uA6yY5Jss7YrNXLKqZo/+IsYOEE+EAiW28ZPlU1
LAVDBM8VCh5HuiqR5PSjcwYHkOu4kBJnLfizuiv/1TrJ3Kn3lHMbN6AVzJgG+yXf5hejXN7yaURB
2mkbUOp6NFm238ZgWx5maYdth9awhuLbl6zpRiOtP+GmWEaXtKVIM9BHRH9f62K8Gb70RKHMhvR0
MXxmK54VVaOk8L5gfr+wuwMjq30oB7TbggNjHx8Q+o8eoWoJJf5XupzRymCvKSUTRFu90498hlOS
Kq1BW+GwbzMP4NcKsQf79RabdPKovNtWl4f8zPimfjiQ06p0ALn1I1pVpiW013vTrEzykNPef1im
22Wyx7SgDdSWmXoVZkYwT8khcafg7EhJj3N9KzBYzGtV446T6cK42ZpdYQ97Yw==
`protect end_protected
