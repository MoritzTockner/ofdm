-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
aQvyPXjGAzzRHRC85OFnS7FhQMXscxw5yDYHjbnenL8rxgxVlTluSRC2Ah2QGbGZEPIoxMbi+xSu
hZ0S/cmPS2f32hRf5YAsL8RGz7ta3XTz0ACTL9Wok3bfsJo6L6dceJ5L2BjmyQr3xH6cxEdYxq0D
MeIfO47MIp/i1vM2kjv0Vift5xat2cuHxUGVa9+vm89Iixg1p2KpZ5N03LELc/5hVhY+pAIlyQVU
BO+MdenSiNegRapt+z9OSZVjEsq2T7zy95Z8fGOL0kUF5hyql/WFhHtBrYgkdoTZGLFdDzMjtl7E
aEVgMA2jZj05rDKfMiusnP7B35W8RxzzaBhpNA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
EHooXjc3eENJw3eZlI3rQIMWq+NUk7gdilgvlnQhRrNnHKCg+5p7+6eYzvr0Jty9ayvVIF9Sj8bp
OPf+LrixwQw8YqYhaGQ6tz2ZKZvnNmzXPRm3OhL/FMq+fc5lncYcbRHm7rO7fonD352woCHlaLvm
szBgJNzJFcQN1sGH1zMXr6JIdmrOz21CrkIP9JD1VraQtwsdFsgv/7HzwER3jApbR/SGbirEiDW0
lRH/J6pEslk5chAaUpURyC4w5QEYW7d+C/FnHrcKTVrJlGqyIos+5Zx1sz+qgMFDvx3mXNNWdS6k
2ruAkVZJgyArevMpWKDthR5k09zTFTem887swLVckojFzJ2pp55fGVs8jptiY67sAU7yTOXM4hhm
1Vhkt+RcSwTT2aV2vycHNj3/lu6/2fdjYr/2mD13jMSG3MwsYAeZxS4CYaM4YYMa5eQaKmhF2pP9
gtdw8cCywlvZlkpqS0bcgA1ykr2FDmUkGuy2AEEvGJo3AoARKARzn/oRy3IFCQZrRQOStWKmCSev
ufV4ypxBAZgD8yrgXPAaa4IgwL6JcWPX5rOVC3RptNw2+hv5sVvHtdzYp+fRGa1NQXhQ8VnggYlA
/BKj/PZyeLoGO2hu55seN9rXbiEd6Wk3s2gTnOK4qsPbR5TqPZ/aKGztR5WAM9iTJyUwU8dGLNN2
VimzfGWjTVfkLkayZbHkwl8MSfBAoQk1fbgh58NWStjZ10cdbyH9sGAfJAF+XQ9miOcKac41dy1w
pomTCebNhNfDsGuhoWICrhu1fnQ4Aj4cUVw9yZn/1wq55mlqRm6J3zEo8PWSxMfP4xKYQVUhvyDZ
HdlcyDlMf47tIykPq87D+MK7ciXvvheYpQlMZhzgbVrmmqyiiXUMxPkwUpSdosisD/oSYEzaoA+S
lCPr160ND1UIp2RSWpccDbocTCOGQIjzt20XJWZ0eHguw+MAkBJyFUp/MzfYn/btOi8kMl3RE2Fv
MuK4Y76gBOBXXhdS4PK+yk35agNH5octZcjVoeh4RUVzI08ncS708ndo2HSCpl48tpxblRvhOuK/
jXyJKWvILMITR7zUmhEa+agTZkEH2YnpeM5LIY3UAEE5reV1wT7GOgeCP/I4x0KM0Ss2ZL+TqrDU
3kHX7+zLg7QubcU6wNHny/47KrvP1GKQypZatc+pS15zZABlDvdJDx7vg6wcznYlzebunnLSBNxH
ubOCTFZQSTtljGvHhswsRLE4YMWa7HaRTB9MLWfS+OmIx9YKXqLuT1g9b4Xgcftq4I4hKkGr+Qhg
AsIa2hlM5gXmwUlWk69fyJH6SIXmHOkOPaECSitd1SXmQEu07Su1TCatgud/80LwMv9GluMCcrTo
HyPyIjFmOycqUqlQO8FyVOvNvaIdowljNYEU9b59DYX7yLB6uIl8SNOxW1LycKIErR5syichVfbU
qt7faMaJa2a7AKcT3QHriQKjpyu6UX7GaKUPjfe58kjmUP0tfTLZ4Pr5smXLYvnxJqYvNftzexIC
SKEquE0g9BoZ7fqdQaSWNrxO8r6Ly7EgzroglXr3XjgVG1F/iC58/mffDc+uuQaaqBrLKSLgMYdf
+/eCAF3GTeQwmZtVZMBN5CTFf2dWJPX0tLOnWz3u+0orK5YE/B/kM2pYIniPuR7DDx3WPHrw6QXs
SwpMqbV43gsn5RLU2a2FDTk/OJ+HhoKAUxk5p1lnMMmpT7H9yguCSU4Ej4cgZkJ4XsHN9eduOlJo
dLb23ttXKvQJhgjNhyqsOsbLSOmvD8oBa9YT8OBInegygePp3e0g2EC/sdQz7yyU2x2ypJJ1gtbt
WrsC9PVdFq73TEYlDm2IsT9BBp4XjAQ0dKH1x13ING3AdWqF9qVuw35zRJacO73rsg1JCU18Qxyr
y1HRG/fIUbJAhuOEuZ7VNMDwn8BZe1mKdUVqVW1Du+0kj62eCf2VSt4vSvh0M0inot/IgchlcCUB
890bXNC9/4DosDYRyYDNlnyHeatlFn7VKvvO023GC0eoPyQXmLbBPsZF59uDfs/U2lmbVkpQTYXk
ERMtuRENWbkjpY51LER8nOihrCVwsKbBYdCIV+bCqWD8pCLNAe5Q9kt0ZLWav/tcFU/RIFQR8UL0
KtxJlx3MT3+1oIyLBjC3LVnRT8h4bZjeY85kpF3ImCAbFUhzxGkBAGH2zqb9pRTF1tvcQa5bFlI/
9zuhUJH+2NgGgGNXoq6aQgFHpqpoQ5ioD2gu7GMgVSQZAHC+31sbOOJ887IHXtToWtUbII5+ArDo
FaVkU6zHvIuKA9UZhsgJoBKZQSLsbRyng/VWFWF+zJ/Xd16RavOSKgd4rpmYVy6JHSFlvjDzJ0yT
8JLj95evrddhQe7+ee3fXql8VAM6o+5rrccKtpeHuKGaOqV94MKnz0f/Fs4cEzAnTITVUiVwLPG1
lHWr0H6fF3VtsZS5Lp2SSD02QVuMH39mICXetlYaWpMc9LlxY2kesk5J3YfQcRXscgc80SPyaivY
PHiwZWJS288roupGei8t7UGsSBlmjf6F5Gm+OGKO1uKA9IaFzUxZXA0ea/iCJvwfBsCHo9jkRT6b
JH6vsymzX33opUGdO5M1QBgqb4cegj20485G/bgvGQ5WSe6dFkG7/xv3qM1BtB80Ou5vZqC+QnoF
Fz9C2n2/gLVmGKXMGGKJlavtBwCnQO61x+pFNsO7/K+MQODuPiDnzbSnZP9oZfuDaB6B97Jh5Zxw
otEreipJI0RDDCTNcBSGNhrmcrzzKyH/U1Yak5T4LERq4UEos75y0F6YM4MKD7PICKM4Oe/dYNjP
PySWi6kkD0PGcKhrkNKalspRgMN1vo/NMcKLHfUNHeKRnVCPP0cwukqhlD1RaubLoyDlE47phh83
D+rR0fwR9RoRwhvha4SnMCoTzNmfTzsXNheiL+XhSO8MtR1mLaOjgSN3X8XeeHUjqXw5n9PBCpPf
fZQDCO71nGX5mmzJ7sqVmO0PKmkk2kXTu47BirnFrUljE4MFdF8PeZrr026his6LhegUzNWTfpO/
1QHCyS25ujLNMJJPaqH1aSF2TsKPDClkBM/FpXJEt6tUeN8ZMt6/XQkcZ62ixNXpAPJX8GPTkbU8
t8keWH+zwyEEL4irDMmcoPFyPhCC9ZtqlkOeHCHonSMurJG5VlKR+dgOLqx/o9uDSarTF3ME/IBK
rxmzGGPxzO2uUra4DcpDKEVbgCnOgj+Vq1kuq24Lm9xUuK85y2Ecz3Aq3MnOCcD5IOdH6PAMUbDK
SRv8hMs97nzCEE1r9vCF2WrVVEHEYtdoqbbdaF0JmFVfEiKTsKAROf1s+BR9O8XVgjhhgw9lTV1h
cUF09y+nMyM6Jq943aJDjta9Zb4qrzdU58ihBYbguvadqAswVHxiv+p6sOg1un0xu0Xuu7NrvPxK
KlN4TdBLmLIaJ5doWauD/AQRJHwbAedEXIQ6EOSXHr8OzXaroULQ+KvjUT0cMnPQxBRBUcWHydmz
5IROUmXL/KegKZeXUsrgZ78tuOYdymLjbJ0Aynol6QV0Fiw4HZUmbD61IHdWlsvoyLntmajLMxjc
XAFQOgrgFz+u8P7xXltbJwEGHrPM6HMvpTId4w6Z59NwMYLHTrBCV7dXHCnvOoKPzTAElbw/Psex
IX66TDt0ziRTGTwfrEZlUYe9tEujEShLHCAnBfSgZy+uhusASBeDwI4UIwuPQH7qUKVnU0sSg36o
TN3JT5AlTa77bT44pF1N5Gz9sjSiSqF2neEx0Gkmf53uNg1xlTYq87JkKtcwLWLVrXk05DHOdCMg
P4WWeAQsImis2T1pH1F8T5H5la4sRhJYR6XWLz0SMbDoJz2vsJeFEHUKTdnaMmNB7it9HQk/Qo7e
gbokpzNw8kVg6nNQWzFtHe/YpOKyWYdjVPEJDwo8O8uIaynnckkLNShiCay5UZ8dNuClkfrUI5t/
MJCpECgRbSUJbSctx5t85KTW5csNg91RatL4g0rCIQP79fZjHz58yYx0C7KlXuQQvLzwPkBG+V/C
+42DzRZFbCckpdzj2JTteRiQPU9juM3xGGQNlrLQ3lOTgppsL3lof3MQbdJMOo5fgKCLqa6OI0xk
H5or6YlOIjgwKS8fl3U+bgZIMrqpGEw7lEDlan2OBmOcX9V9jEvF+UvjGsJL0WsGFOAjgLdPIvTk
IQUJm2CXgbL0TqT5u05AFyT7D+/OcjdLOLagz/tJek/nJYezDaS1+i/87zpuEt/0oFSX6LM2+6A0
Oze3KSHlMgY9ak2cKL5TFzDqDsHAFK9R5ymkwJKc38IydPl1U5s5VIT1l5EqyRqSMQShNuaybR35
o8B1sg6vrQeSmMadzBlwIW0a5hN/7Vc4o9UM9igtfjE43qfAzZkjZWA2QfaGSugDqrFlaehHtfhV
/w4USDnDaCxFbmImNo5RCPuhe7eh+N52U6Ll6a7xQpOrJ09fvXL/CNwR/PIPgQezOwfiDTnaszJp
fxOtwLs9I8uypajRcQN6hu0nhG3YTGBn0NB5f22SchgEPd/33qrVR12pWgQ74ufZSUU883MbVJNB
L6WW34hOHtX6I8n8nk9yqAbwHDDEdLW6u7hBjcbQjvk+sjM+DkFSuecZ3tlsz14rktCfgpwDfq5d
CObl0meeMnHKlKazd93xkAglKm7iIkShAEvNKayms46ZM5hm8g+DpHIk3qEubtivZihwTEjrqFRy
6gIjieW6l1U/GSdfsX95ZBC1rmta5tTlCW6E8+SE+6VAKNa7lz3AmEr4RTlVNUgcCeqUrfsnB0f6
EVWsO2HgXltstszZvZzj0sncP6NuaJQQZazeIYLBB+c5XWnxW1n1UbJCWMxEzwC5t82+ecEmZrRM
g27BQ2mW5IfQXM7+8ygDqoYGL4ed7Y4dSmg9qF7oTvx8ULreHg80AVS/yUYbAglRV+Z7Pvs9VeVE
Y5AQiZD4qdq4+ffaL+sqB1kMcDgPt/eC8c4Yg1pbyDsN7enmmPNi1sNkMPgivUS46AngtQHBDcqg
dadZIpN4kNgWNx3kSNZ1mSlg6Q0pprn3DhpXUcdtA4MAlWBfZzMflEU93dMh5tb9ARWEBPRuuTOa
1QgPeEcl3ng5k5QXBR9JHut6J/T0Qim4zTgJ1cTf7Ym2uTM+ShjWy+PRZYSIOlxWsw0mtgEjVCEO
5Ti9fX2ru8RjcyVn4ILLPSn6T39gFTEbEUbuo9ElowKt+bUbmXchxwNFYK0J5alryPmaOX4DCx5F
x89CM+DcGD2Nna8uLvcSYnDLVK1jT5OO0VpQuEgw/m6edYvgUMQLUq+HF+mD6/yOZwntl2vHcqNQ
LzVBzrxSeP/W5DyGaK+xsR+oS2wizn6TRdPF6EPLY+4cVTjfpLyyAvmVRMuN3PMep9PUIg///DXp
xD5oXLVHSmdZiqMsK0zW6Yc3Z/9U5bnhYBOvFwF7mSeeP8Pb9JbPU1shIY8udTZPtMFNWqKIpyAG
gjDgPUhC1LxMVth1W2uLJRfTnxTqCb9hiaw2KWKBzOkgtf47wBOB3s1yQMYazf32OBbqWRTfRWgk
Fy8VjSonm43gsSeXMX4a+qUfYNGSADihsPpNLSOy0h8O2kBP4TpzVTL+wfnNS05rGAwYc05aM/wu
n1Y/D+Rbc2he2GpAdQPAtOISyn15DSTtMxfiP1NYQjwGNWYpJgO9ngnTCaTYFpxFls+0EGezGurA
8aEOvY4PHsD0Sr/hOA==
`protect end_protected
