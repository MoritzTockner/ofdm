-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K105E2WQZ9CMZsUHHOHFOgeHC6mukSX9rvPjB46DHH1isNQ3O90xMna6me4MjAWPDHJ1qh+1fvYK
E2rfFIU34u17DJmasFVMESYcj5pe0PREfHFGQRfdUUwIjbFqwBWfmTXbqX8oDxcAbRUFcL4M9pgf
GfAy5UXKA30gsFhGZGjAqars8+c9Bfd6m0fsvLEJrnJE2mtwfjrJiigulZnj2lQvgWloFihqu/7t
eokOik5QZPOuRhwJ0NHWbQEolQN2+j0VxA348/W/ZlOsDnbFxYQYVLQJmjOVzHnKh+hE8Epwg7Oq
3lwCX2zrCNCLaC4FKRDQfGFKYS9h7QL8CHbS4w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35616)
`protect data_block
eSlJmXFbSC5SDXtIKhVfAQ1NkQiuPxLDLg/qG+LOM3P8unUCkQH9C0tkLmVaU+FgfjhqRQawDJz7
Pon89TPcJ3jdeI3+Mj+nnaYOKMuYP+9ugrmlnV7dGvd4zQY/6Xtt8DOic3FIfqhjZgqqnBs6epKc
b9qw5Eer7URqGoKhriVdvFmtEz9j85BCKYjc7ZS/tBjI6AT5uioFl5CDpzgkiDY3SlFD3yxhiPOw
U8z0xmJulgL6SE8JJLGai4Gj1XjHbbcKVRz+tVU4OFILguvFdkixEFymKTleWAWIzSGAmQNgDYKR
FKSMoFyNPWDraVQk9zzDzKt0q07En/3V+526sCsFDWmKAETFxG1WiWK69/PG0+l1Y7c7V8wm9zQq
ibarmwMWAu81URLWyfRqryrGckvdgCKmZ3MUT/hK1ZYgRwT6jMpp25mtxrjBpq0rOXqdfJbvGwXu
xGcoaAVUaAypOORzYGqyjbUyHobcwpqU8bik6M1tmFyJvf1PVtF96lYg6126tbEpnAJiz7WXeQsh
h6DRurGT3rkUq4T/rNJ6NrzTwu3Dbdns29vI34XRZOjyBo/I9VN8fyMMptksf/tbnN9JOhRmp4dS
pOE2lJ8UsCtJ8RhB5Ar2zw4EkJpV/EeQYGaVM6Gzbk0bQWT5621wt6GayTrGJbqo3W+VSLnrbn4c
tIA/RZdkzvVaJkL9JUnbGXwZ5jJf2jGZ3LeLuJV3YVb/rje7EDzZ1C/5iaInr4CwUjpsSt/ZRrxs
KS6DQcF27N19HJNepC35j7fNVlhk3ZTWAY/rgfVZXLZ7ghI2T4TsfdbQzZOWhsLRaIWbWBIR7WeC
rgn6qeGsj9QNJeNIc3/sDhlgW1W6Ng4U288B0XUTX266kPtcFx+L3UiNb+2tMhb4M9YBLAX2vEvW
EGNGkGnfGYb+iQ0G723pfIbfifVW3rt2UQ0n22BlDC1oxIx6PmTEt3jitt0TmnDNVMLzP8MNle9T
OYYZWobOSy3ee4C9UjC9mlZexiWaU1GLgKZR2kncotMrc+2xuW6S0cTkEEirYkzk6R6cQGxPVeFI
U2KhKXM9AUC2MD2RXwEjGH7HBSj49xT/xy0bMOpti/lnG6GUc3reh4g/z+wa5IivS1j1aZPl07JG
+gVpKkVRBybBtZKtozFCEfpLPndccsoE3mSO1maFFeh++3Vq0dDSAocRTtcRICU3u+SW5ExrVwXX
6VK0k+RSeCjprypB3sWIWYxPVX2Ek/b4EjCHVv1wr7BwP2jDDKnpLjIPjLCKtzAGmNXe0t8SpOPp
e/Wai8m/r0NAsVtGydx40SWfKsqoHu2xxPPFyYvZ016qmUUXgkVp/VSKtzgYGZng1Tp8sRX7f2u6
3oJoGc/kYNIazi3XIF2Mt31ov0Tr5zj49pSeuOtE0rHmrDHyLOjhnQ9kqU+WN+oM0zYWC1V7+O1a
fk5G5u2mCVV2rsCEYA5g7siu/bqbXR6LhhjvZ9koZNx9ifgjMsuq5auNLsvDEh8xiotwCHdcb4I4
UjFKhZac03tNLTD3EWmL9utuvuPWEaBm0LcJtTCzvPUyQ72uD/2nlNGffRGxLI9f9WrJgaGxPNyl
G1y3UZ6aF2J3LroxkSrRvIwde5A0vXpJ8/JkQA9vbKWAviFmwp5Vd1w0B/H3a0qblnDTRJ3u6RLg
qaFYJ0NBOH+N/XWk82lbWwqK9IhvFL8UAxt/4XG3B+RlpyaIwv9Jko6bwGvcwCurzUr0tYYmOqhj
ffH+/Ipj3HVncNlh8vTQMAAbBSo2h67AM/nYOsMrJq+GefPAftQWXVLY6C/FpmStdHqCdE6U/tVw
zQNK0mBBuZpGaPnMTeTaZDXAuFNK25YqaWjjC3VFN0ziAx/Es7Ee5WJJz0bg2UOZLBccKI+KLzBF
d6UWB4yxyNK126s7W0YP0mlrJKJYMz+cEgfPj8oQCX/DT12MV2Dx+OoM347iXhPMfY/NZshWI0Fj
pSnkg5mIbj1rh2uDFY2ob+eQbgUXRebxJqj6wXku7r3/2yM7digtGUummyFrA113T0ogwWC7WJi2
gnTjkM191c2uGYudRSJkBll8UkvEdlT6tzdO2MwvRTO4uO7ohMvBGbNTrtGzjw9kSd/ujBtBWK0+
L9W4QpxhA/3gPlF01MTjL4YMbTxodgD9E8jAzAhTsOD1x3jTnNDaDP/4gPVQmqC+uldO3P8fQSLD
pFA/WN7F3exmvLwQm866zynn62Y+unWCqiettt6SPr+1VSw72bM+iH6k1itV56xyyKRti2IGSi9N
+d81x2WJVxmhiIZdan7tQN3R0SY98K99mWvZIgX6gB4oVbDlJI15+q5Z20ozUNiUdvo7lcL1T/0E
FFNaVTnSmk1EE0y8ybqkhUTxA1RcAvmPAf9aGpq/dYRC/pjYEJqi3OlNkCHCQOp5rHcCCC9zBV8Z
n6YXLk37zI+IymP5MDI8OkJIpgKiPs5Im8LeuYQYQ2ObcUQenglQiIUFwTPGtXuyJxA/PQ2uXd+p
aQx/VI4o7Eg7hyQTN4nkwcnmAbvgOR4LEKkuKlvoAb9qBQqCaezHgO7hSDlmOLCwbj1JGBVqHdgW
lmYSZXV/k6x1x4zjdZ22tiLcgMO/w6v7dScJk1Rc/jhF82r675EPC+TnXSIc0IhLKI7sZOzpNxa7
Q/4puO+1ryaWCMOjJ0iCP9DmcgbxPJXrHSfCGi1xmh6JKjYbheHaeyDT+sEs8soV833fR/H6k86s
OsIkcztqpejd1GXzmhg9j9uMppnpnEqTnxCT6F1qDnFIbJk6kMnElKdpI43AlkvYM4bkDgwpgtUb
x5mtCXbR6b9XgU6YhQ9LBK8/A1dEGS2lbLOLZs+3zWufzTxOF/PE2DyxHKRsy5tw05P0uvKb2YWc
SWvsnFTxgQwVYIm9LNXy77Zw8C3FeAVJyrOt2f+Br88OrtaxSQkpKHXWaA+Gn6vcurGeixcQX+A0
3roZKJbAAUy9vcOOgAllI9It3Ne4blW8TbSK756UPfjLwLamjfWlCbq+Rou6yzo3MRcraOSwJVRg
hbeh5Z1m2jLKnyCBLJYgwfxgiR3A5A9Vrcx/DctymroSkW3fV/yJM4sESmOrdChPPe65XCQUAFPx
vcf4CkffqoT99cVXrR1rE9P3oZr5KbXV2hJYPWpGTe3qGdo5fRvFpBi/ciJyRPMG4yK8WMIJRkiq
Z/KSOFJ78LmXmsHo+69sXdjZQB6PN0tY5QGOdxibV8TefnnivzDgLT1O5BsVn9KzrgMwWA8KW6eY
jPs4ln43S0uRM/BmNcrFvOr2jNERNU8g3BGJ7zlmLxkWzDlLiaapmYFQ0ErdDJuhh0tdoUjPZomL
jocQuS46hiy2DUeEUAB5bd+2LBGHYaXDdrChemM0FXy2Tx2kfeBVAucrchck+mwQvyfez6jxqGnD
M7I+vg6/91DzuLunQmPwkh5CWv8dstWvhtMDiraTF9G1DwuniJHK2AeUpJOGo1buoLydbtEVGg8I
ZdlCxzY2m2ZFa/itKhhSPnHJ7ldHNPHdZm2tEaMWF1p2+i05UKf958BPc6oqbkfeauWKseJk6oRp
eDc5/1qr2SCioh1Xti5lawyaVqOzxqRIh1h1GeAXXzpEWtbCfjWYMQsVSDn5YwMNHx319Zy/05fZ
tI+gaGDvGCf9WZQ6YG0COwLicioX/REFLQcZg2Co6P4iVjkJFQrb8N8SSCz7fKAtFKS7+x1R63AN
SNIWbSfauCm1cOUgeHeBF+3TTCiHXLT8ETSkh8ZYW3UEfWAk5CpRu2V/PFhBMaleDfbILSfmPKX0
Hz7WfqgkFyBXH7doJjEfjVsv09zlplmWoX+yT4/yNtSqkU637k/Dw+Hv1bd0yLmIaq8cPPMwosRO
QRvriznongWPcGauS58YRn3OTFeTp49A31pA5as4sFpyNiIogXXkqMyS5xqbLCbJpwAo/ed/Bv2N
9Lvu6ObBzn5Yhwixl06gzdiU4skwiHSLBR1I2xIenv1obvhgZdn1d1cY76//4gPRGNZ/oWbZuzs5
fvDWcJwnLFOcuqhM4eMCWh8CP7mS0Kxy799dXSbPXFNnPJT18Qjz5pwPMUhKA+zJ7e2w6hyk61Aa
1Wtd3+dgIfH/FOG3zv3JiH4MSqnqaQHudUs3wSNR1ofOStuH5fz7LbIM8gxRqPsraJ1yVe2Qudga
IMwwEXuTQw9y6RftZv31apmu3+k+FOvl/eK0Wq1whBTqat50zLIY8taKEmP2XQYeY0Ow8d5wjvuX
pc5uudvDIV6gJl+K1m6MKHJPNevnxhs4+DVPlstJAjaetwDvwf1MCxrXOW1OeQc3Ojcye5b0RdV8
DCijxq6f5Ua2tAWUiiyH93nozDy7IFyc0Egs4UTRlfO3EX+Z19Zv6jIfU/C+3l6md2LZe0wkizVM
hhbBqcEre1jmPdB+fJhsvUp4qYYElhgyynPyFopNTOH7+LqgSxRb1MCjWCvteRsyhwSRpum2+EcH
2Fs8MQdi7tdSopfGbeBW2y6b6Zp6ChBnX1MZPf6WbxW9Sq3uXLP7axdqJCHwJkv6NIQaqbLfX1tp
qjNZtT8zRp3KdaYZoKntfPHXLsuFYAavUkX12uzGoagdIOpTC33YiwIbY9Y2xX/IadmhsDsai0VK
I1ISmxvg7SHmwRNg7uqY/n7zHJTEt8PA0avYeipi4njT7mgTMIxO+Cxw2WLQ0+TDPJG7CcVrhMRf
DvDAb6OvEk6RZ9QlbC5CP40RfPBe51i/hykJRdgiTlheTakwqIknIVD2wvbuOhqcqNVSKYbiXDIa
ATFEnCjOrS3MiS9uK+J8tjnTK3tnaAK2ptUpwazdY3U2wYzEvhM0o5p6vE2wz/1ZZyPRtmKzaVFi
vvqFGPdPaPccvKJvTeuNUIzTgTWgqeOgpXK8nLwBW3oiB2y83GqhHhSImCbFF8Rj27OGYUp58f3O
9+eEPbFLfm/WjLDqDOQrolO1vX3WYRPeOhy7pMMOIpvATZQ0gVnCMWK4omvep8/ILnH1/jIl9Huq
XRH1Ij7cxagTtkxQdp+Oe6irIkKXPgKRh/Ht9p20YwuUU7LZfUdjQach6wrpnF3ALEtSVLAdT3Q9
rpijlhkEEJ5g5sBfTVp06tObno7jBXfwpQpWwIEyShS6Zp+0chTVjtxz5z9oMVvaR48QLSZ3orx4
PNRn3TKluZtA75x6axup1LRwrwKfQsYxihd7yt1kdXWgoHPquJrKrkyZ+aFNo7HSHgf6QzEnysCZ
Eq9TP+0DlHbQzlpSJ6cFEXAwjSHMvz5agRQpNGnQIPK6Dgfm4M4CKuLCsV/NVi68QzkuxgqkyYTb
x6WtPdIDEOPzEHAjcwfigQPrP5ynzUnLBZqABfyLudmQ6z8U3hG15nSn2RUrGbuTosMdu+2T2z5n
7AhUCIT1K46/gNuhHLILU7QN7VBFD7XuEfvQG53zF/LE+LHVJpSd6qj1dygeCe/IHoo13xASF4O5
0zKFDNVh9Ll3i/6idTeeG/b1RlcmzzbX1jst7F9R83mUE7eIcnp+2Hkpe/chREExuLRJfimyKeTt
gm8RxZiRIq0W5QqA2MW2B238PBvWRhsMN9cMH8kcVreKINKwvkqcGLXDw2h7Lp6lH/f7swwrIuAA
5nb3gysvVubaDV50Yxc9eY0IaWkjMDdDH7pke/aDH/0ZG6q0O4DHggn2wpOLfY4DBCQbO+bA1IyS
RYf5BE+sYYU7CmsltIXEwWXP+uvbQ5BMJsV3aSMSq0vwBizYj6zUMjzaZ4b9DWFK2+JNhyHXWT+P
sZwVVSQZOsqgTkI7eF3UJ4+vDRJX8+Fvlfr6aqgfow2djw6F0zNx534aV3syHJtZQul5ud56xBfr
gFJAlFq30Ir9ACK6GXbU4IztSf8nd4pyeLXeCv4n4v7uyEB2tge92240N4KiY2PGERpRRZ+6Ozht
5d5Gt98C7Rnrbr7WnzvQ8HP4qVfqtji5OOLmt31EmWql1ptgrB+kpdrLGTuRKIe+oqSxWcQX0EAC
RqIBen57ZxmYikFP5Rh5iA0F5hgohkwkCv9PWF6spiq8F3MUmpmyNFBCu7k9RV5liljUQKwjAEK0
jMINFJg00/klr1Qk6fdluGxOZBY+mKx8/w6OD0giw+XMcwOwSBtFmLwluZFvzmPJ4SeZuencGLEg
Gvpqs/oduUN7DCVBTXpox/mDhDOw6THCqbrwtl0XtHRSu7MHNX0YjPDdzyQoaCt+1gggWWUOqDSr
CgZYfOQgugX6NcfRbtl8MaP+Gilu1NtQCwpU1VZCPB9Elsdyi2AZ17b6J+dav4n+vATTVEnPPDXq
fnD/4+QJz2Hf5K+M9rPraeGNApRHrQcP5bl/X5CXbBds4i5Iv4f+WVECLhNAFtXc9oahkN/AnRP/
N3DrNu2ZO9Uy8BiFaJ5R1J9xAHAtZGI0PHy4fGIe2Ouae/RGZ7A0TUKj3jZoae+hMika04RxHXQ3
tnInp9sHWtbP93CORxB6K2NgzhrvV4wTL7pclMGEEtUADe9uL35oUb6YNq3PpJQ7ATx+ZyyWB6N4
X0i76XoX8upDgrXj57uP5MBZwqbgsB/3hsbswuB2ym72WJmAQO025oCFHc/4qbBSon8wJBWaqSMe
4swXFbJV6ru/f0CArrIn4wahEQoryUJKL4nJhgXTwuOQ1H85W7mi+IgDo5Zd1vv0+sdkbx2AFtbF
ORez1CYHcNKm5MTVCxAq2j0p/KZDPtkaebYsQgZBi+j1zjioK+WdDQDir5f4yzKO4PF8/FuLPGAL
g8P1MGmvRJWmKD/MZ0U8NV2O1K68Jy2/zVjxwttLUh6ftfw1wB161F3xZLpLoT96qaflT5Q21jqH
KWfKXVLtj7CZuxcWDCZNu5V+nSKIqoOj/XQJ17EYKTxgYQqkQn6Jyf0ychIIbCFujgCW6pgC5RH+
0P9R28R0BAySmQj0oNN8md81UPgITmaq0pBsxr/FQskLgTN8lpHcbLi9OayJZH2E2DwL0zE+8lkt
h3fI5m7qwSyNRdymjVxx8AidZ0YACEaNozm4mI1A2jOj5XvBBR8XfihRmabzS3/Fsmsm9wjwUg/Y
8lVTJLAVyJRruXX/9OCqM8cKDMY6WVaUCXSs4c1ynlc2oolneBVig/DsSzRtmD2cvuV8IPuK7G6c
nAiRfgv3hsXGI5N5CmVYan5ty4VozhKP05gWlaRMMqC48i8Hq7yyeYLZPaAJPC263QqE5raFJOJ+
ChdURJQtYCQkGOiLQNw8zI/c5dHxzEI0a0JVaInlxSOL9xERrvg2Oj/lAQH/JGnhigtI2LZyO513
FMJBgUNYjbIcv7kV4Awg3aRWyj0UFCIGL8Me6qhOk91qMtRpX7s2Lzi/pHImg/yhWARHxc7pQ3Dz
odJYrmeXRyoxh8cxtTVHdQT0yjns6lmCTq+fEmrOMrCB04ZOM+QTUoKKMSjug/cm8waODwUVjRBm
Ofz5/tQ0KTWLVE3ADNtSS3+HQLjZ2nGU0ETGen1s3+PUC7q6O4v6Oz0RhzGLaV3pNzOW5dFzT9He
752Ve992/Tn6SQ4u36uSu+rsz46dkR52JCUt+Fl3DAmVKlYTZ6YcyLT0Cp3013gRRScLuX0nTBgF
C25eZNbglm9nO2ogCrwf/O4isRxKFZmUzIGFgNi3xz4ld+Dm2SE1TAYiBZwMK03hdsk6TIwTAp0P
U0h86wgJNXUCBxR9xcJUaeXxxda7Nbl4+Pb+wdfafneEQxEnYyYrHE5V1LBodbtQKG5TU3C43H3Q
yBurEyqFm7usUWmSW649RRbtIpNMC3hQdsyhsz1kvo0yQTtxPuRJNpUXOmViraFZYEuzZwGrT5CZ
WRMLGjXBTi3lWq4itZFB9ASOXBgdoECQ1l1FbK4IdX/dlYNlev/8C1hJTrHV9mNaXQOBTLofKBx7
Hha7xgkY+27BAnLR+9tnsvjZW+ks/HA316SMRqn1SyxAWD6e8Hyo6PKv46N3LsZNm3UFMtUwwlwS
nPvRqpGwdAluN6QQwfUrUvB0Ae7s09/FTB9Qf7MrBacWT12hfWUspjhxHOsuv+zt4ONw4CKdwji6
7lbdpWIY/JjTrjdHHHz0b+yjBvU3FZjxC/s9x/a+feZfvU5jrelKzkMaau6uSvL46iFeC5sfzMKf
aZiIB+C4cOl+q2uGBtlty4pKpx9oEhfcUw2n8WRdn6bAkGyeffumhsotBpPSdv/wD7WnnVv0Ux91
bFKGHgNQ3pv2VH+xUDxNIPvhielXv68X/8QlUk1lHnCg2tESShKSybUQHWC3jmw3+4JoSXjQYTir
7QP3QBbutZgjsIYVs83ZFiRJCh0w13q/dsf/SJyFzV95sHyWGAHHRMIqoOJno2nUqMAfl1A46W9f
EM5xtPSfKcfiw5kUyBNhK2eVbEJt7xCxeLO8Amdzf5QeHoxWKf6mrq6CsJ4XsEAWjsl0hDGe1JJ/
rHS4a2CfAJVZaVeji/179eX2mf4dqGZuknxmlZAoyeuk+DVS2t2MdT5wUxTmIDGXhQw57ff6rZ24
zQSOj8+EBoZ7BuUtTKFEbLRwAfEcyuUQjLfIaprUGb5dXTnyPBT4Z/l0eQJMtoWtvJJUjlLY9+c0
O4mF3W5ZcmdnFDHAbdz4oZSnDC/OAmbpFkwTS6/H3GXKNIc4wJExOt12v8l/3WaHe0WnG/3uZYyW
IenANOwv/R5/B9Vo0Rdmz99Eqw7tlhIMNeIu1ypBz8jkiq1KaU5x9ygctaw2qTjXuN3gENaTL17i
CjdAG3AHUn4RSEoWyPUyG4wp+Hcazv1Jo/6dyP/OIRomx+05DXwrGLgRwggrU8punnoFvnx0wNml
N7xWITKMsT8yi9PiPsj1awsVFWlamsdsaSgAtee6MGkCBg9pYcsedxXzsIvsLHhm2bFICy+3cLMy
9GABlptQ08cWbpX7Co1+f4yCYHv3/o/I9+i+Lk9rRPQFpLzHrlqVz4WtMwPYkVT7AR9XWdTxUd0I
cNS5MGy2wY9ihlYeBnDxMbIsv8D55/QoeNZNqcl/yctdvmlqrHrkmEi/+bDkPUY0np9dD4NWvhc2
92AYPshyBDYGUShPwuD2LdbCWIe+sFqxXF1i1HVcqSC8vP8AjLel/qel9DiWZtmPn1nrPSMK+z36
Bd03NqP0XibDrJ1H6ztfUfmkLAijn7WB8QSI3Ut8iLyRFpebfZJiLbR1oiUvGTgMzBhRgxanoSQs
IDz/TP//dQhtMKZCZR9ZB+CkNbykhcBjgnpNsa33B9MTXsschX3F6PlVvNbdHmWj9cOesl7qDZ+O
yPVBddWDyuUeWuIyotkul9mqWHr6dba1TVJU8Dfa3sAVc6p9psoOS+mse9oeeZHqoaE89DcqIb5D
nCN1cD3nO0N6uB+RNwVXo46yp2x6kUhedtUoj+gJH8ztaJqk68Dl9llM/teWW1bNupBVZ4CEQpGX
V3d01QNhjXETrrodGqw2i4npObRpNwHTJXxJv1kHEA4MMqrmo6LVFLcH0ebWEPT/3b5q1F8NHuWS
EC51GzCiTTHuX6jZc+Mg3tjv6+0cEHEwClnUAjC9Yl8RamjJ3zYi/RnlIDpKUOp1iTUviHwz3Ldw
lbcJkVRc9YkymBVbDNBmgrSFQzvJIJJwZnT64A1x/LwU6HkM1kM8iY3rRFBp7l+VelzPBIklQIBf
MuyNI4n1Fnh9+UZbhVUSItyyeE4rUW8co4316BmU1YPQkjIvX9nR46gqUSPqBtxs2SgCyzYpv9YQ
SXB6SkNk8+TrOwAXeVs/Bp7tdFaVxbPe9scXQttZnK5+eFbEI7FJZiHv33awy6YeGTEK1f6uK+E7
34TIkE/7K1GEsbW6DQDE8zkCk7VLi2bwzuDgg33krYfCNSS2qqgLbOZma1gKWR5LMhKfVcZo5dSy
JcvjbmEo6V8Vg9Z2BgcMqAILyC3OReeRJdBnjINDDyLVEl1syMZLj9RLfhnGzYkkKHa/ve+dX9pB
0F8ex4S1jNm/nEy1wfMiGgGHeoKvmuZARfXVGYDI9ujCAgHfwCIHkwzCQ7p4Ysdgyw3v7O0pRqxw
52CNdyenwpop2jxQerMHMEbNPByGwIDyyqHtMr3AVIOSYnjktWvJhgtC0KuwtRASiO1NSOeTJoDx
3JrXxMem8zrnuxqjAbPe35iMwcpKt58QcdPr+otNeISZ+AKUOEG2ei245q29jm2RxaeMwkEdcWk9
NMqJd+Vhecs+d71NrQQG9f9eVzfg1wxbuoy7tBCIkxEspWFuTO2ahUw3LBFL0NUoOD2bYCx4Fwg3
oechTTEGM8L4Ie/37maBxDDoGM1uEUJM4/jZVWCeRIjzIq2c45CuPAhF0hjlSGZlTpo4sg5isU90
wmnkSGatu/ao+1zeWTkekn/5JdW7McOLPWXRSuM9vDF6b4M/IU+PhaSsGQC5R1a3Ui4R+VK2I3t1
hb1IDpATNp8mwSXRm9dQLAOSbfN9XEqYXkNR1zVl+7qG4auruETNETFlPDpW2dS+fY43uDSfR/0d
vO5aXqlI1A5WzQjFz19rZbDA7HdB6p8V8+LpYOHeUogUaoNnlA1lg+7i+R50gdUfnqjAHyeD24y5
6uWHcJ6+HiYp0TplXlUolKLYIurrpN7Vmuh+FYrVglHhPnKfrKsMf28LUKwUEcSciiEAyGMIFSmG
71Xh8hA1C6JTMT6c0GmjR4936SCZOZt27NYgBW51QnoWBuKnUIohnnnlXrMwuYzkFIrUzjZtHoRA
KaTTnMWC5lelxeFDuphNpyIOSedpKUNPAz1c0tu3mG4qg6j6cyffrm6/ik/lCcoyE9xTCcrMKipk
NMITG2HYwEea9kC1voEcTY/W4RaSBPfSybzVG7nlf3DrzZ+jYloaUhrnxNDO9/glebvJhf4tWYoK
ef4S3/FUH271pwt6TT9FWKN4hgVFotjgmbkA809h+yivUfN0WjaftIPsLsyTrSBDFqpSoqeBNWIp
Xu3+JrEpIhZctIE302FqS597K0w9QZoZtjmaqQYDigwQ+00aVBJqDZ72Ng03QFWwiF7GT53IUrT+
oADfmXvJ+NG2B3fiKkFkKxOrq1il2zRMHYzt8A/KiPnkQ8XBazan4fFvAdIo0dlPtSLEZ/1xlV/4
QnWZ1rE7YGAVo2EIvxBpaLLCLrL4A5xa8rcghbtWnJT9WerMBtHwO4y2xFp6xNEzqkcXXu5zdVPU
z5XkX50bjVE8Fi3A/3jAG2GFSTuT7zOXJrnBlExEVyoz8lKIUfqwDQsgObB8/t3rC0dC3NflCtjW
UKkT/vB8pB9SFsDvj5e/Ql2Fmx5Wy1urmTL5HimjN4Rwhj02uQM/l/zALLeroHQGo6QQiEEhDqyS
4umRRZj5x1AMS82YIidZSEpHiuD3kS+AtvLAGX9csm8l4HnkqugOpYtcTGP3MinLuY1i97WP2TD8
ta0G2pSY1PXdFvhH2GHi3Veql1mj2ERDmls6euKqCHvijJ6u8SGw0kNgBFFo31/Fj6ghze5QsdHB
KApTD7DqLr5mk4bpW5qw2N/LqFdB5DKjqZlvH4/6yMMC1mfAgS+RwEvX/k1ZDjIA5A6OQOKekdiJ
haL6my3MpsTbrCpADjap43ONaaMBEpBuIN3PukrXOtMP0qdXxckilOkT4Pcch2YVw0gSb41QaX8y
WirSDf8L1u7TeW4AHD5n8XLtzFy/s+uhJRUM7Nsl9CPgdmaxeygf9sLkexVw5wCp4fSH7WsZrC2D
huZiaGt7djIaADmBQmJkKOYc60Lvg4cs8OjMnkXRJcspOE6ZPCeMq2MqmJKhx8ykDDu1Q8jZugbf
aJDattlAFMk30OG+7M+FO9pML3Bbhgy0sKjBzKsjsf0sDxn8r6t75wKg+pH/GLFEg51YHIVuPVVf
9afk3wmaCa4lBExKX6RAO5MnN+iO7W4ER7qeVNLl6qkmde1nMqRyM4oihNG9PACENwKPHVgo/rM4
vzKdq2GWJzlRlkYdQjVAR1KCn2HAGtpy7rz+nkCqF/GSmNhlJmW4jbNQvplNMPvL3lxqwnUCkBCi
4/FO0yoCDwZ18hxTB7ACnlP36VqhI5JR5ElckEW1oB4IE4morcKRPuTxEYS5feZs2ICA2jJh8iFt
xa9ROfKXbm6qsHINfwnDXIiLB4DG34oXEUbl/QFpNrJF2SAxkPTGiSYKt2TwRItwiDgAs/l9s2MN
CZpKEL8mgGigbTeqn1rUzBUqp9Sm6PN7BYAWARgzkHlFKOotLp22B9e1d+VFuzW1UvzSltyYLvZ0
TJGqGgyZfwZMKHOqF87xOOUytCrVfAtoYSTn7kJ/+B6mYTDo04naT5XaPyggbfciWBk/NsIhwtdE
oaOtfB1OckaG/VB+67iKR+Dtz3fANPk0HQoVoXYphvxYvGAByQP2M5y2+wl5l9ZPbjEH2dNGtKUt
qLTtDoXt3CQ9vdNTl6NLCaPzQjCumeoV0iYG/msoorK/pHrV7DKRYfeOYR/5QNvaYD8C1vH2ZdFl
han8mx20YThb2Lr9UB1ZfNYVNrXcjjgSRTh3osHjuYOZ+XA93AcB7T5oMw/NG35aLBqSDOpaLZjZ
KuqU3apadjVRUQXhsNK3r/9b4i6swopuG9pZq8+DErdlHitUXF8l5u2DvZ9xZu5Ypd8w6lTkvBRf
tNwGke/baq6wq72Exgh6JaBd0EUvUfuCLLqaaQcYiXhkMHhNKQcPqggaxIcX1aCCnWQOe9TUtRUV
f4TG6pyvYj6A1GRzuTBfVMRHA1YnM7CNDaxuceJlt9x5d0W17lzbQtih1C75iPAQgvF77qF0XecL
isY6DzMDb45zYTEsaSSGVDHUustY7TWV7ANtsDl0wrxnfzajlKZqWP31ywf8ZAgnbcsmcl0ObdwJ
DJs/mJnzMcH7jJvGUxXlc0CYmuV6w48socYJE3iOWDnlp7dulNkfoURq07p+qDNLpadmmI8Cfd7y
gBRP+zl4eBditlQVLzowTRpuNybhIYCfjoAF+7Cu+CEcO47bJq8gRNiseE+2p1Sg50XFzUGY/d94
kqVAKrJeX9RPVdXQ97S3aUOJjAk19HpYiQlOklrTdBS855JrOJmcPUM52XlDP2mtxXCKSje0sGQk
1Lowk+/7QKe9HUK2XnE/S8CJKaJGqQJ93bzb++u3RW7CJdByfkK2Tv+R2jz+PfKZXrHrJ3ZJjOJ0
fmD2y7I91bURz/Axqa2a1BURmkjv+xeWBIFrGmWHxpnqbPCjz2Hntu56R7OHTrnG0m5weSCw4TFB
PQXclPZhtT+rpDclpA6+15PLK6rq0atU3QSgrvRj0qgcGdrLwxBtf8WNpbVd1gAfqa7sCGJxyssC
dnqcjxqEfaga9GgrSh98bEG16AVlxCBy4B3Bs0UyU4RTNDy7wO0rVJTj8x6W4pqz4UdNKJmzhjAg
wcymoRz881j77MAhtkNCN+GKwnu1hWewiUT4L88pL1BeO6O5WRO1g60j666/Sg/SwMVS7VxpgjVu
n1sLCA6g73kjOUCL8WhnRSN+WVIQU2lY6wcjDXbIC+iw+KljU4ei2HLN4+ZlFzBjwHEHMua/DrqD
aRIsoUnUkFOT4EQFXG5z+NoyhroR2Z/nwiPasEYyK88IkOKtcy7NbjKKjsYXKNuFqpevQU2A6mjv
m75/Q2HIdempOrLr/QPThenKiztl7q+hFyn46ODEXarrMxrbH4HSx2oTUHU2zuzyLgz9UIaxqiaM
RXX/B+/jgWiKsKzjsKNob5Jzpkp7Ji8jThLB7TQCP/CsDKxKrDuSlRqBPvxYOSEHBH6bRQYInCzU
qY5lqM61k4eHrYv1iIJU0J27U9X5p2CzAetn8lyTRZ1l1Y3Z4s9v7Bq69ki5LCihqxoCFS0rfPVl
Froxe08WA/7QviWF44a3wgQspsXMsBQK4icUI5g2BWuAWv4pkQHm8HNhfBlydPj38j0npt54B4S5
ULTMu+/2FBmsrYXHJX977Z0QC1uFkfcgLOQ2o+TGd0rOvm6nEsxPTJI/MNDvRDx0RtUF5moD/Xss
n4jQBRqTn+oo1zMTeKHHdbOjTu9n00wcWOX+kJtoVi1x4ZR5myFLQlUgytLagGmylOXm+w25tMFM
xPtvYPTWFHxnIL4HhJ++NHy1PzOchv9gaJLAj8DrIyMnATWPhscgxwbBB+IP0ONGB2ayRAF1MarD
SFEab2onQ5ACThGYCRAqQwmAr0dn6ePfmErRz78HRJBXxicUxDJ/A007mtz1dW72qpM1tlHv6S8b
lhVp+Z3HhWNsSCkZeQbVFbKxP5fbbBvk3AekXdnwCTS85B2pD5lU14jZqn2ezt+rfLEoZq0aXZEz
Gutog6lv8Udf3nKJX07VnXUbgllCQxpnnnBjO0IKmaCpPnlBkVk6vTNMRSrQUxvucNqAYP0VeO+g
rlW/GieuP+BGoPNuvZOXW8YEZ6KX8AEZfW/FhBGwPlorQ4s+0GA5iCGxsmaZkJuKBnnX+MSOANQO
pFLYLHKh34k6FzlMF9JZ4C8HNdpgCNirK9kdR4wsWsh/1TRetBMeIRn5FH2o/9MSI5dBeEgvBArH
H5yikALQOdv35O48sIDDrMI74I07wPV+932uqhDvgqdOyzc2rLwVkbJgXSIpcMGEiGqrNcbI/I9E
eCzSBGAGqlGinWLE8T9k/FMlsUdp7Bt826VD3k2HCfChcqYVfHSEyKYHpEODMVeJgZapi9+1TYW4
A6RR6+3kGHfDMhoAPjWYRbcj2Awa1aBdKtOvExLZ/ZRWRuvS6e3wpdCLKx3ppFLnfeQ4oYY6jA+C
V7+aIFxJqyQ7wIHlnBzrr6Xz5qGGbN2Owq47BJ67OlA+P5KbUAnFSq4pXKR5Ee4BgcPWJTw+ERMG
DAmkllQBfBklms0Ke8Xnh4AN7mdT5D0n4eAJ0a9e/WqFA1yZmcr8NyLiTBPi02vN/4wLMLC9dt+s
OE4lyQmcXCAwGtyasuiD/gGR8SIam3UlpaNm8oJwz7HbTxBplEGGU08wypqBJlWPMDYKfMpPFuzq
MqtZsnlR5q58dwFKFgeIg0dCf0fs7TEPLVrMcyOLGQnxy+zGUSYZqamKLowf8+3vJGRDGW2ft2Bz
ZS1Ok8LB1YJX4gQ/gIB1vTQUAigu6B9dy2l/M4hZHdvxxOfm9GyD+WWw9CUHPe6173MwlShOdnnn
dfV5x9I2tqjDjoHxO1GPrPggVwojaNOSuBua+lGCUETaeMLcvFlomR4F+mAXig2kIlxsqst+7c2Y
/QnXdVvP5m9UxsmzWrMLZrD10OXmIa3Hs4F6HfvlNzE6doaVVfTKSyJv2+NjG+gtQjwy4RrWGV2q
FEm0A+k5ekQGAGxnnDkPeHaCnlm4UsqW1N6bg/NC0SF7g6sj8u8Wk3ezkUwXcfAjIiWveK0oKDEC
KC9r19TRfQ1puVSENZUZpY8gU7aGC4KvdfmehKb9bWACsNXFVaW/9iAi5EiS8xdIh6ZbmsxBnQlu
m9MRTkrZKat+46NdSFfgmbPdG+HAm4YisYlrH80+2VEVus136ExQIkS3NkCzTms6qVeYz8OGupvF
5Zn1YMpxt+7ckKsM8+XftaWVtCtgcTfBk6fvnJOCM3K7P3mcYW/6VhxGnpNkhFAMvlSp2cWaJ9gx
e6bXwKeHSxmM47IWor1iudi5jCtkphF9Pah7pgmgtWssHU1ogu/mqiWTQ5/HeFWD1C7LkSFUxdve
fXREqXXyfHkgP/6VMdPXaon/3FSz5cbkaXl5eB2sjEg8c7g+1CVSy7wwezr2molef4YHc6Lv+23B
TzgockhcGw8xchucidT+h/rDS3sjinkSE5+s7pCCcfI6ElG1+gOkK2zGuhjFwllDN2/8pxvcEOSr
cvmlwkNsAR4/3whqFL0fI7iXIX01A1hfMn/RniKy0TpWzB64JM8LT9vXAH6A9LJS8bTVA+Vb4HHc
690fe1j9FmfEEd8RpxHBfzldVP5dfb874wh303b7P6BgQk03kOQfbNCde1AaXJ9/R7tF3HBrFJ00
vPmvWxi2Vhy3cX+eYthCzMJhuCNc+Jvy1az5gxMZar+991PmwoPgl8jQ0eeQ7dYIC8SFa1hlmb4G
6yOQ4NA9NllWut5pNCHuE/GBj5XDvn6nvUGUxApqYI4wlF1DjlRaRKPK5OBeREawkcyNLZs8i4bu
u/bjZSx/ZaTF5joJeOvGDbcwJeqoMPoh6gz4Zomlw8lc6Zg7am5c7v2SbjAgGNihPlPS5NM2Sdvx
qsgknsR9/00F/vUK4MWmS70FjS5Z6+x5aff/Q+/S/S/rvtBYxv236kIFx5Npcg7djP44pW4iFElU
V3Z1RT2XK+39dLj6UDew7QZNowGDXiziaZXwoA3t6ti30UeW6LdoaS3vDWXr95Zm2vJQiR0hMMth
P/elvEdLggfu6itYiuZ/yb3deZuONnA7mucLzgsV3jGl67G3C1JpzFzEBxbECOYHt9EgALX/AIhK
PtUKVaXQ+W6t2urTppj1ftHyYaz3tUqqrdJcDtAKhT4UVDBd+yj8JsT2ioAg5/1dpvnYuCA+g57b
KKKMZhmnOs9+s9kdnkHR9Ogp1PjSEqnQ19AY8Hzhmf7IaRENa2yW3rFsDqZMvvpj6mqW5MXsD3Hi
BOBYrsQpsQNh9u/c9ss/FhRDFP3EbWB8O056E5PaP4y7VI06WWwyw7vV0DR+ETveiDovlbtSzLOI
yFihksJYeWTLoaS5mIKaj3houfKm38o/RppWFvxvUmxSfFVdiTIrPZXJkppMygw/WH7Gdxyw4spw
06Q/VI6POhypsogVrIUGy6Pk0bA7n98oQxq/O8WHIen80OZ5Aia3FR8MAUL+xUgOaQml9oqpO2VN
9j8sSy20VnyXiWZ8FxaiLLm8Q2NEWKA9hhhyJeg3MmUizD8dgn1imXerd59QDjJdgoT8aroujaQ7
JTz41np/fxJ992iWeEL7why+CbePiYqb/L++sqE3B+dg3xXVGzEuvj1MbKRMMKbGsVD2ei/okwCr
+et1LeEVnPDuX8dGz41ol9PKPj1/J88C2Rfe1F02i6oLDr4E14JiHs/Obo40BJmJGPGZ3YmZJEul
+gqXf8bb3KRxYbRDxscNgDsyQbEFWG4vOtq2exzuXgEVTDe1dapMQuPwoh6yDowZhFu6CEA42pSc
M4rU6I07UctqJkrSLUJkR2N4jG6ak6H7vh7Ffdho4QNWa0KfMCRXEnEAvDlKD0JWm3qebzGP/ySI
Ft5SrQiMoYfPEjeLz5SI2+2EGOAlyKB8APflIalFfIbuUOEfkvCXV/0CYEJ5p+cks6WUzqR2bGkN
/FxWvK4Y+P/Sg3p7/EpyIYGRCtyPV6ldLAyndzrVBGbDn6fSjU7zi/TlbfuNF4U6840p9H8+OtDy
BtOyVOoIclsBKiMUAFpJXlAXDOiQ2UFrY9RvBadiN4GpTKmMLcYm8T6Cwofe83x5KGrsHyMRMFGV
4JDhwjRq6jmBMmQC7Uf/V/wpzT9lMoNu8ycnp3b8CPlkzrH3JQWGznlKRamcwLnI5DOgmM3+NF7L
oVxrVNcL9ToWa320djFC1ImDzLehzTCu6nzXWz6pzmd2tcPTPXfSemiCieWG6HnyFV/6bogL3k1X
gjWSwoovKMRxgzcyEvFeHTG2a3784DV7nvi/CAZ7/vDDW8/ZT62aBmLqFXLNEW17zA8ljtJv60UP
hOBLtck9aWjNFg/D3Xfq9VoL7WaSGoONaq6C2nf727m7s9ol4USbcHLZwhIgbuzTcY0wHQoJWT8r
kT4/XLbA3WPLF7QLVXdqLpWMzw2HNKYXyRSD/nv9sRnFU/9lQ8ItC573XZGYz01CHGVbwXsmGvm1
WJWXk33TvGO399aeg80aKnQ1JqRfL1babBzInZhxVULBzSwpejIir7bJP/Ts1/fjBV4JiBhpERUW
KL1UaLiCc58Q7g/Lvt1SuXg6MaYDyWskNRuH53baaNWbBdqJMmPxz6u/edbn1fHOqcQtegqVCEhd
qWMP1XZjNJJwLeV5FMPvGm4KAAvDGifO2X9GB2AgdmLmPcnAuNxpuEuNOtOJu3pgPo4YjDWWoUtq
SYkaIPQEKGAEbi16im2j8kz6eljApWhlKzuQMSLt7no1NWnTxaXY28frXn7MO84jXoQEQlJ/4YiQ
mwLwixnHKotTFVPu85V3ija0DCiQAD9nYixNY0FcniyLHoCSpSYp+uz4nz95kdIHLDGZ+9Vm75SW
a0v1rkwx3XeEwTxd+TCyP+sbjMhxgpMJ9u9+yC+YrIQeWZFusG0+5phHmi2tNqGAyB9WHBnaTc00
HXPSfbAeTgUqvAOBRaPP8RgShDqj2+tJjioUGuVKfVIp8THDNvJJLQB1Rm1TMenTPL2Gj23xFiJf
c81b0rT1s1JCe/wYBlBxTkZRm/nY8blrf+x3ugeTF1AZOiV5IxNQZ0J658b3zouMymEshBlVtEnC
vvg7W9CEfraTf9X1aIBlim+rxGitM4LqHDB6JDoFqA1/qnUcEm1Dq8/6JQPuL8aqImz+k3wYd1Hx
soYEHyoqA6/SkrFKpQOt25PCrdVqjrZ3rf8Cs6v373tET0jkLpa6Nfpie0fwtd4v8kOwbPHy0nNB
paiS6eutdGufs+PWWr5pZjhhBoyJfQPVqCmE4mnCTrA/mAVHIvTEhHbwptbitGvM8+9XHPfFQSp9
54BcFfAUJ3pJkjMPvz/lY4a+cs630J+XfMPTQa9v4MeVxQeJFJnaMzpHVejbDvuejQsQxoaM+eb9
meS+yAuaFsS0bT0njO86jJ98hyN2yccyQC4cirGugKoOAiLEBKIfWayZqZB8TRFV2vj1ULVV2ICB
mfVqlrdVuAO1kv+BA7dxGUXqf4iNmjkWLLhrKkfveorF+mj+XgHTKxk/jgjGH9DiSZYjfCOUXTm4
Ovr5gGK8oJzTsRFdX4r992QTOhSzHhM+ldQqtEqBusfV64DOS678RsTwBi4JJav7zuDf3MymomQ3
xMQRNUrr9Mk/gcaXuf8J+j/8zEaij9P1YPSaOxT1wXjGspm2ip4OisTjcLmeDDBfn48q70MPbZDf
LE2VCCGsTJn3EKG7gd2dxkr0Xr5eBtlykGxzx3nf95aolIWLiFbXtHDk91s+av/a4EcF1T97Vy1Z
zLfJK+FSCqgVc1mneMkkZw27LlBEMWpVXTbLxuazmGEupbkVkix2cZN9LVekw65hVXstu0ubk96K
Ttk8iKtftG1gC8LdHCkEOW1UO6g9SgysTEbyUVlEfenysxD+O9p5GJjXj2e4WcWoORtRohT9tK+/
+UvIla7ZoiZ3zeyFaIrV+jhvKYH1EEMtQ10gky0H8sf5WKWKDlSIHkurMhHxmHdAaYMWShfhmAS0
G+ktIhhGQvJ9EcEvRvKT7acCDuNc9hBY8QNMMKy0Dxl0+ZKGr8d53d0CV43QiBn1cXdrOWZVytNU
ngoUaO1myr1T1qskwziOPoteUOipfcVZSPFMXzI+Eu8F0hH7sTd+Cex96SxJPYGbHuuA0hWFmez0
JSLBhbhRTTL3VhN9wdjly/QpeyQf+m2kHXQnAtkdiwHPziEk8in61odXs4zB6zxEkVSdkqaeQ1vN
2fOvHlKgnXA06J4Kh1p5oMqwrglAO5pI7lgCIHlLRgLL7LK9qrokg3DAA7x+0n4sLE2Jp1Oc6Lac
KTyuvDg5Cy5h4nyc5wexES/a5Glu9An+7dYGjDCqiS6InX1wDO4wxqefQMTlDyiRVehtlu8YL7Mj
DTy3QLO4vHnPDJrjFa9YtJgBCU99yKIaQAR/Gg0PMiNWnwzHVTQcKXfql9vqrEB/+eFQESnSTbA+
Q09Cj4spEGZ1O6sdnTge3nwXo7q8T7IpNAANptbnzQcA2Yb71ClDP/NIhER+tGFHb4JAm+B+83Fh
xUZAck0FYrgke2h58258/mHZSlxuPSDIGonyvBUzXBL6Yur8HVzk9rPjFYpZP0uqhyqkIoDO6Ld6
JR+1I0xgi+U3I7fAKa7KZwpFuYJBZZhFfqAoqIkiuGHe+LnX+yjxGXw278VzyydtzKgb5GZRwjBZ
kO8X4DLwIkFnJXdNTae9jKAb42O+Q8sZdvnLiFV/tAC1Nwy3R7QKy29pMNNFMPvFHibJplVd5+uj
av44/Vv9Rg0Mp5uDAbLDhK68s0OPPF+6GhFmmZkZ2XNY3zsZTmdd+wK0cupTtPOMdmVyXlLgpR/T
Wh3OA+YKWkRcGg3leoCLlYKIFVoiZPFaIbo7Tu2OPKF2zT3hBOYlScmdUDlZomMOGNU9tZ7F+ZLm
ZK8NjVLvOmDYfYXPozqcKC1tkjKtYtGbFHWLrXbHugRUXeZM7FiSYvrf0+rAP75QLTZ/4ljf9d8Y
TRNCHcuZoAY/aRzhBgYs8sITSIhWRJ4NjFcSRDYuTBEYAiM07QCniHwBUi7Fk/UjBz09Da8+RQ1m
FtgKHfewmNoKnnXkPvF6BblOWUiRQuW9NRh5P1YFUoZp8LWWMMWGDUEG8brRre2CE7vxkBl5fcng
ypxzT29VGxOg0zh0NpghxmQSq9+iD2ihBFO3UBeM98RMdqCXoP6jEkxUAXtr4bN32pB9Ruxq9Aaz
c7H8DhYpuhy4SPvsEhpdniqZTjyw1hfhUhs4v+dIvnWopd+clL/okzLq49dHJa+rgG8sITiIlnQD
ij0IjXbfoU95wtMf8Cyeea16H2DqJE6rfFK4SY5Xtbi1Elrwi4t5OcHJw4EgpA4m5mKrx2Sgr/eh
f+7o9iILdE6tfWIcgJLJPBE5V+3mHV3u//9YDJHihYrlxdMBwCSVGN5DcXZOAcxWQy1z46l0iqi1
TzpWWetFHzvygprjkVHPQhoyiX2AFaXZwgSsm93UaDCj794UbookMdhveoqZUyWQYdTnFSnROKwy
mRfBGDinv1nQD4YkrN/S50f5U6Fao4aiTEzeLmktwosVqLuwUq+VYFE5s7UhaB14U46f5UHCGoUu
4pmVb3OIuFNKwO4/klXxtKyzu6vJCswdZ7UAO5oqTc3kAjq4Ay1s+iMN/Xa4Lw8zuiyPiWNnQPoV
fxWXhrZsvDpGMWMH/ng5CU+T56xT71RttbP10cwxkplnyPgWuoqQm3vB9PpcuSq170EjdmqtOrHy
MpYSi+rkJGulGX5XgIatoJ+m/scNm3MkWR+87QLigEnvxelx5BYQjRVzZ+SODS5kr8RhmiwOx4yS
XqrgUWrUCIT4fBOjgAZncebpqFxrIfwGb1zTNupJ0TdMDGZMZRAbaSyhvXxZZMeXqXOGkmr7xPtR
WJohx8z+Ez7oA8yJEzoS6oA1TMfFTxaqJ+/mHEfGZHDHvSTAEmgxD5F41AKgZRrcEHegY55pT1NM
WeCFGiZSswjBgxSmq/O3h9vNet6CDCa2mWsWQ8bXUkdBP0v8fFDnocVP9JZGRg3GTRFvbSy0k8ZB
aWVejgT5kL3Q4fV9EMOOM/riCUWs9CkgMie0H0akzrcUpCncWeQmPRon9jnGocAz7n80S+sir6VS
AJIW0iMyUVZdHCK8vyb1FydVI0P3XL6Y8ew4EplJTL6Vh/hTUyjlB+Ins+7b2PlI5fNYc6l/E0Kh
/NLaZcxiAYL4yvtAZezH2UbrfQ9+a5Bk1OoVOJ83zoGhLs39xPRCex6siNw2DNEb6zWF9TRhiw48
cLLUsK6I+xv9fqvd5B4DefZ8SVH3iuVnxY4yUk4xR8nvp8xjBNJlQnT8CBnVOTNxIwW3kXweoYt/
3kAxQG9kxHVaq8CTkZGAQJyFB8RXk5WWiY9t6qwNzYllEcEsBuE4orrFzP2cwu9+cf4jdhJKVJ4j
KyM68Vl9NgSUTB+7Km1TnXZQNNXrMF/d8io7Ie+NGJy0X5tgb+XZSp2+/Nw9qeYYmlGVizef17Q5
pRVjPKT0lFKAWQAWycOySMJh40w87/C/BeG71Qm8ZOIfZ+TL4xMqehIoirDyKCEx8jJPq185C3Mk
Vp9VO9XUX/01vieKy2ZWd4sDizRBgoMhzPm0gZq428+y7M6Un2bd3IVCEhh7gI+l1lZ5SO8vucyG
lTXFdNjvF58RP8pEuA1Vf5o8PiDbQqA3nmaX0UUQavBNMXx9GhlpsLzd3/8yXpSsNME/u+r48Nof
s5dfyBV0EXO+2EXN1sk9u/DUEAU3uazmkomMtID/OuUhl5SCSM0gA5ZZ3c37kH/7ZjsAZDgxYsek
VkjxhgLXeMBCLZqypFyciLRtnKGLsziCo6XnUFOLetpiyD+etZ7YsG7jcH0U9p7NDAjtEV9aF7ng
N8GRH6JH/NcUsbm6AIo5XBmRisU5N2h7eDKzkXp2yZWp4lva9nZTZ1au5DeGqzCaQz0UZaQKSX8q
5ENiczjf0v69VCkg4HSyuKJGQYNJ300Aupvo86y6lIropE33/KSX6XF7svpH4/zntHuvHAIZDAl7
m4cnqXx3t+N5cFvbv5D2SzsrKL1NAFDOP6BtoHNj9zMpR2C4KAmnHfrrGc9PfE4a9K54Hu7X0yWH
/5gyEYtBrIhomh1aSxxgbalbHLDswI10VEsHKc4l0089UUGoXNKPeZIKvfmPoQl5KbZG1UOfS3MD
7EyKoae7K0c+czx9WemI8b1Njf/5bpNpkZEEqpYy0t78KSlDms+1RtmyekDlyOYVwf3f48dcp6HR
BgSNdzQMjFaaUBi7sApz77aYdd4nGQ0adCJuszTBEqXKfGiPb/VocalWJjLdweJtXoC87YpmG7pS
u0m79qIaiqTaiywdjDc0fgUv1340ZV0acvts4k7BKCph1JTt0A+oxAR5gaaYhAkuMzdGXdSXJW5w
G78HS+3lZq06Bd4+cVahEVyePH1llN3liamRDpPI8ni/JkIUpROKtteIjC1mv0LPu70TcgHE95AA
zl+TSopmmkpHR5P+jd6LfJa69oucNxPoLkVjScwpRLhNwbRrmYtfCqGsZ4+Y39gjlhGfbYZQPFC/
iLi+wjnBf1+x3qk9Ijqzoljx8L8Gq6iu/BsMWnTIkfDrwDXQJVvDAfdVauxpnWtW7oYuktRcmjaz
ssN4Ji0oNRbrZbSTIWJBcdEFU9lE/4aqzbWX0+d6QPjhMugcHrOqJWGWMFSV8giImyzXsR+UP+Fy
v6B8SSC5nyyNGuL1sNWzA0OomhxtWgBp+kDTz3gkOYfWhAlFyyOifavby0YvSJOsRTCvojWkDU9B
WVghxqDSmajgMQbUnUpOjTJVPeajb8n6LQn1lCic910WiGmPPh2vgo80woDyXWZUg8S8iBYl6nP3
/ALzMFHMUDsueHkUjaw0JiCIHb8t94qLUOk0Cp5rwnOTaeOHNYDMNUkPb7CObRPZ/WJwu+ksumfK
KEb6I54O/f3Z0ylG8yyqg23U1LIFxdqF8ihPMXhxv1VhAG8pyefJ+5JmSqinVLyBoZfzPuRLMjSR
uosYBWj2uiQ0qYoKOO7FtZtm01jLAIAoumIJcVJlKIl8/AvSK47UrglaXpBNpBUhnKBsJS9/GjmK
PHGVr1dBFLbYSRSySbzQdfVLEVhmQRsxcHWMrbHASE70C+DA0nDmGaq4Y1TIf6zeIK8lNGTAV2O1
t1LUv/SJTesF8FQ1+E5oaO4HnjvxRj/82BLJvTVCiRepZdqse/a1Dfib0eTnW2JtuY+mMLw0A2eC
bXYtjZXBozXP1WA2pFdADxxqvbMvso/836vkOegLgJGLXGch6Z0YpByOQFzDcKQeEXV7f3qZQzVY
rXBWlLCw6dzfHF/IgNGm0cunZ+Z4d55jOAdkKih3g/fjQgbU0hglswtNLIsTZdskhXfpAuDiXT7y
HNXB+w4QRfj+Izpca2yougPFMNWRexyqXjZZyFcpQK/1GNQZ1w2CiZsp9laGnDjGxr0Mg21btDBc
TeKulHz5mmtyISAkJ0xSDhPdru67lA3JI+/+VTMRJGwZv9wv9nBESxgnNYeP0WaYt0oeywWWa5b2
uP1AURfQp5vGZg0UhWNBtOAgzwXqs3qaQgorLwQHZJJyOBDRDH36QjY2mSmc9Qy4kriC69r+ib2n
Y3JO8V8bCM82YJA+Kv7Vkpqe5FYAclvpWhWld+zW87m88U52lMeihwG5ZLEsUWS437h2DgXnbkln
UrvCbN3Bhcaw3VyQhVnBaq6g68iolUoRspk5b7/KkiY6UDEAwdg2JgBngWmM/0tn5KcdC1p17+wP
E2Y2XYXxSnDQTGorgOxBhm6jaTg7nZHIbTbxev3h+Io3ZY7QFj7MkzeLreV71dX9+cBGmu0xhvJi
88PZYGll5u0hSOUQF54D92qmCcGF0jFo765tdcxW8J/uzbR3jqR07W5FcSJbad3p0MG2/3V6wENI
XOvZQuyTDZUy90IkGroSYV1S24grFltT6kPOt4wMGSlf0u0LJFMgT0SGKAx79bf67W/+keFirG9I
mo2qTDOgaS8EhCRquA/8S+8HH7Zi0QP8Kc6GyPdrIG0EdSy39Eopj/eKyQbm8YuStvfi1zrKJw/k
//9CO1GPePb+McH1G/boGDn4kc58PGF8vIENZX3fZKC4uOH3broEgiF4mveo6sV4VWKgXPx4g0J/
mWm00+HLqG4nWzJXba2uu0KjG665CSt6jLEYZ9dk+zJuCzvya9clv0bpVXMcNP/GM3n/D7lQnC8Y
ogjoU/bbZJKFPNB4nMDb9yoRSYJLxZzykdJpt7DVbxwDdSQMfSLoMLmITD2X2aMqrJ5X3LBA5dhX
1WlD/+hyDkGV5E3Gsbov8FeekidevEJRx1A/OGLNEn6QkF0Cg0UuoOUg88+MydUbVvBv+PUoSx4q
6oThwlHZ9EvyJWsShdHUtPZ05iKWjKyLeWauAV0AHDNlQvkL2Fuoql7PrZJ+odjQ92xasECXHeyh
zaeRpu2Gzx78FKW+Hl57watmt3e4wtj8iwot+BgJFhugLcQltJc+ppGYUTpBxm9aL+pIG4S/YwCq
F7lx6/ot/HR/hv5PQG8NhZPu7AaIjOEC/Nv8mQxfOChFgiCYxMlA9plrrL6tigihPDNx/xh5TRqJ
/qiok2y1bm20CVk9ov9baSdQOb4SsYjRW/39bCTiW/4d/GFtzsLPq5zA9dwfgOocazMAltHER8ad
Wbc9uL3djkDbeYEuia+iIde/hBUO8vJGejZgFjMILxSJic1gD0qdDavlHGVk3ddf60CUxf31E2uD
xNFpgk7oFKJXH96yA3Vx5ot6CQdMaReLisfG8TE5acMDtePiC4NJwPNf8m8dfnSVbYdy2+/IjDLK
IY4ST7HeCkUm+bJezgX1gQQ40Dvaa88vYCqsOSTkk4L4QM57rgrRYEu7Bj50DW3DKPbi19KhlP4D
31MQJEE90XGYGynkrtqNPzlYqkR30NhPqODe9hikHY7f1MQQ08f45CXh8IAM8u8n6Kv2xyaqx0nh
CKLW272Ha5zGowOaMSZe3mAEgiyfp1JdpgTaxroTyJjRI2uUglcYb5qpH/TIKS64Rt/U5hu4wUTv
vvUC3TvFYhLfhjBBAU+vK1vcO2QyzYghB5kI/UdxzPMUenD+C2AgiL89bInieqw2ih4/LlTE3JFV
f9kIWXEj1tcQX68Aw3yr3pk5IKZuIzH6Ioa5kJKwY6ZxLZlfmdWUjpecyOXfsxAW5xS1BqJHK1zn
Sv6G37BkKfd0L7Ls9lRYMjY7LRuxt76tQelTxP/uoQasaQYsTtk+cNpNN/XQgX/ygDLySgYdwytT
Nb4v3H8DX2h0NmIFydUUweq4JfvUojyrRP0lgVXMRNRB6Dkghf+F1QBa54/lK+OEq1uLtv+xzQt3
9edYUqbasl19wF66qc3P4P8wEhbs8UAIMTuUH5k0gUhCXI7NPRyj9/MRseRmw4BPv/RlE2Q9ntda
0oNKZvIWU1cOBNqN4k4EJqkRRlLsmZJl4Gau5XHPM03QMkF3rP6Zh+GNEuqboRD1bzevo2rLM0WD
DcS4r6EZOT9sLcCMO5ccAIPxhrOahaIOQGg3v8IfpZXOMUI+PaWohnDQPnNXBTfGAFhfpi6IbTMh
vqOJAZGpTBjCj+0Zvlz5DVnT+rN9Dr2o/jpBNmxmFPqX63M2Mcx9keSNLr0c5fuIqOfazFBW50Dy
5lh0iWR4Rx4sGwxwIB0hYPKm2WDwuW9obcdzs/RQj4YQkRm4WvFQZ6KwB9MOTw+yXDIqyoWKQ/93
QT4zkUcc0LhRcFSQWV1f7B/cySp7YGHFEdij/HL+gBbWpIy02yW822WgLi0CoQn5LWja5BGSIyyn
R//VycOLamW1rgCIxpgzOXijcvCzLCjdQYX9jNk8KXHr1HPxF/SYqCEVGzX5L9QpUaGSo4QimLW7
66+ZY/aPSyosxU8LER28INKO5X83fNq3uT+h6EkUTBbO6tizt+uMW6EgQ9H0oe0xh9dGkGupnTPF
w2KuQx41GfX7XJlm+wHtvky8W1D6tpzWx4WO0TT6Az/G0+YF8PywqP6OAsaPb/U/I3E0wDNi5dX8
hgIMbZa+sVFy63R7nEp+OuU+B/SdgVA7PYdd+UfbnyaVxkHO/yJy0ahNw8XDE3SmhqUVVOIFNAIH
PiVnSmAYGznNORoKlg2RIH1DE7wQkckIY6ChYhymg24R33bOdk24e3ZhjhGfgxnDNvlf3gG27BJO
zroxmoZbBBsDJa6YdADniRXHr02TC4FCXmxR5d8bO9kx7bffLnXi8+Bdf5E1dxX2sXOqBk+1lAuQ
unlRYJ+egfgy52ovgpum2fjLJmEhCExYo10mnQN7p/fKqdzIN6YpNJHyLUpgFo3hjC8gKwTmmzmm
gjXTpJka/wr0OGFKWYjPekKov++zPq+Aw+E9ZMdjDLDV7tgoDJZEK+Qkalvphx+2lCWJygyzorUs
yVIxfiJbaSzbSHIRs7ptmwC7EavYL/G3yusuvhS7UuU3XBWsxazqB/Js9MN21TRigKAQ/HCm8VWJ
Lom2ZmsDewExlTWdPNzjvH92lj7xu4htsw/zmgh+5c3bmowkJR5PrKTtNipyH+grx/XTRF7Zf3fM
EkgOJfsGKpOaCy3BRimS2HTWkN6qLPEYX3ClW7XnQK/vAqpNzE9ZAthQMS8epO9EYgl0uppkG1JM
bfhmI5GfrAQaSGJOazDZPprsOFE7OQ3GtBv5y7Hpu3ZKxWO2fXCsK4Zv1SLmxljUzk9uSUslAzGS
x1N6rLwiORdYkMVQw6xIlsvz+ykv3n5mR1oHTUlRLiFeqe54ndoWqcjQkTgvcSYCdJsV+Eg8VV8M
AJ6pHjiMkPTpChmD5s11zM5h8yV80IuuSAPyuTV60kGevfDoPec8C2attvzXwMMZBiLKMekC1TB2
QVhp/xpAxpK0taEolagOzDiF54AvJQMJMYqi9fz+ImYkBd12410CbhO+rE+8E8YItXZm+JaF8Akl
wmxowedaZz0wi+ZXCdZDgP+nCVDcADk0etty3UbtQZBRt6EpJChtfLJYu1Yk1qlCvwdWEVX5MGvE
Vj9kkN4+vRL8H8fIXVVqPigEc//tAGV2fj7Pdzz0vqG3a7cJFLWcZ7coB/XkUdqCBgBqozx0YrfW
bjxce0hV67cCIZ6XOYap8RGEMdfiQraEoNsKGX9HDgKc/9EFP4L5plZZS4qdPZhqY2emMxzAsdbU
I0lTkk/W5t1H1Lgba8EjsqBssmRfs7ax6uNRLvAq/eDQc336hRRCk4DWw49/pjJxM+AMqmT2d+fJ
21YtrZg/lzjKSFuiQ1HYtYSKoNTKj2xxMpc6L/6e9iN8eXQuwEZxXF78Ky/qxeXDcSDVFQsq6y87
5PUX86UJEaxO0xTAWlXdp5FAq3OTtvWyFqH2E1gFtwRuAPeTAvfLVlfprssFXT+eY/2X2l8OaRt0
xE1dS/pjPICWG6hzrQBFJNk/F9BakeduWuf2JmFUk43Cx4ILfJjMfnRYI59h2yt5DYnvswowVIeK
RickFDZHKoKP3U+EU4WHsVKW6ptevb68fpo8y0IshylgkiLwGuCelEv+nvGtNzfNCv1mvcaVC4cE
gOLLG+/YbeJDILYEzx9cC15mJKKiZ9pUq7wnT8zorwY/Bn1JdDNXz+CyvIHtaNtn9FkwJPh101wf
eN5dHuoMRr725veRbMz3Xlgqlqmaw1SCDdZMrbEWn7ErypuUAezlA8oAVPvDbGt8X/1l5BOGT1cm
x+/0J8f9O4HqsBm3KzaKtOYaVtuv8+vN99BQhYtNVWnZ9CIlil+yakeKqnjnS3CiP/CS3fi11Sk+
g8Od/Q5ak5lZpMHwLUSJnEud/Lk5E0wWtm6NlSCwxdnBiDfhCh5FmPxh8HUTsyM+hvAOW1O6s6TX
02evq/q1bwUJbLSpUD5kyqmORQFfAy7FD9zT4WOZ2b1eKNCvSvSI4f6nzgXu90pQ+YbPOZ2C6giC
GdRcWCRVun3IhuaYZLG0k54PHCaUDRXS+mZ1+Mt8LMbt8Mwp0omhBAz/sgOB5C0F5oiWP53ObiW5
J+w3htYxA8uFyUYhKxwpzy5WKZy/6FL8bmdZ10ZqExB8kLrZCyGCbM0rrIx57VNC6gC1/wTwNnG6
GJQdsjvC2oEYXmAidzpSPNWkDjricAdhB/b2jriSEyveF7DOrgBZTe3/ZgLxFWe6byrYxAYqzxD4
Q1O8y6MzK3mEPjdoTb5gGSff2x5qGr1nHzWmW6jydeVltZ2IXZElxee3hvk73al8P2CHsgGmUDZu
7TXAfhb5vK2l7FuTQomSYVMGGKkV2q3CbVaN3F9cJCnas+tSHWJUh3XoB7b7tCKxrmf0ttB+hW2E
nxmY7u5UgsZ79hRwEUtQ85K+oNAUJ4mIdHlZhaUt1S1bvOIZcc3vNJMG03UOY3r90ZWJ9LT2PUgU
+LFmkKBABOBzmpl4MVpfGup9tpRqP92bVMZeRiEmDAAXIyCZuP7Ck+XU4d2Qkaf4KeNKLK3FVj+H
ckPFwcBPMm7PkykaMQIyav0KTuC0O/zvJ1Gka7nrlZx+/VqD/i03vEqOsnSRxAeDYxTFd415/Igt
8ZH4mmrOdp5YT2Ce57h0iYC2sR7OzZFxXF4UhLp6k19mWG89ZvzFpotLvhTn77YG8WWh/C9K01uq
bDOvZJLN3HahWggk5dkhUc8f2hDDSx9KDUoCVBcxbNh/Gi/bmCGDC2bYHqyflRAltK+jtcRXOzvn
E4DXWbSYklu2pjky7YaxEaYyUzKn4+TjrrrjfCX2zpbEVdMBBuF0vmNkkf/VGoIiSLMs8ikXm1TW
ksz+t/SnoGZKetknCVeV+8m6xeRNr7lddqzhE5VVY5lfT85rJiw7aPR8AxQIUrcXcEcTwrCarhDt
Zekcn2IsamzTLqr8w3g83i5ZIXnnyNwOS1KKkf//WLAJg+wIq6JZ66wFIsIvkh7gibWoiUuAkC/Z
jODXDFV/WOYM2ezHj2kxJKpUodLPYW8ndC2EebIwnQD5MosPTBYJqucjcRCZXI2k2WWaACbA2za6
82P2GaqRlSDzAmt2JRIN82afznOOrgjO1R0f8g0lt7dDysDXcWcs9lERd0FHgwukpZrAMBp0EL4z
WGtGM/Mqm8aFG4xK8baYts3O1MRRNj9xbYwofE2c0KELy5hzO0wwymUANS+8N4sSqZyZ8IObf6LM
7fA4DbQp4qRP8DzUvqN71QiGvhzmfzbtnR181dC3zUO1ZeFm4rVvqUxG3uex7YATejAaPZEyZS72
kLxeJP2IcfozyV/W3L2w2bdkXnFHD0AYVKEwzI0SWMWCvX+hBDnychZrm/8f/eSY7vGTc7Sx2dYF
DmYDvXYwP0VOm7kNPBmDbwrL0L+MGPOLt7V72vqQOPXYCphIiw3ux/HGSF3yder2XtwiNIy5gQXV
8EHXU7bVk+pnYx8Sc7n/SQaXGcwxIp0Xnxb4ABxF2vWVq9J17Zrw1cgjSu2TjB/LPGRbRuCfwR0l
NLVa5mcI8CYfXr37MKsfNLxpJ3RWi6r+sq+DuM83z8VvZ0WvEdmE3u6Qt4n2R8iMvN/hOU9b0I9J
tx39En9lM4RZvZWJcSSeNFFXayrfiMEA07Yhz3GB5nUSJjBqeNou/UeU8Jrtd5yiyI0xPrwuUG3g
01OLr0tNgdBGu9HRlJT80SJ2Apkwi+OclflAJLOaB3oHLP5s0jUOUxDrt9v94LFIYd9Ef12JhgwF
c1U1CvWPDx0eKNG1bmKpfx874q0d7P5OIOAkSk0e+vQKcWtTcy3iAnqz0xHLx4WM/ZF/fGCZutdL
BN8wt9f/4kTZQFwFFSz2HTAaW2iWIPr/buv35lXAJms99iXaWeBCoWWEbe0j+n1GNJw2WvlhTY95
Fg1jWuuNz02wHya/5a+3Z4jagJNsCQ7cxiWt/OR7djU+CTrbaJhQw3jw5QlSHEPcnPyiVqqsYmhA
IVU6ydcngAtDhANFRTzAhaMkH2bzbQ3fvMH3Y6yV9dERmptl53XhXgu/B0aV6b8c1JsBhKsPVsEd
m2wN8Y+40ImTircRUX97MCLiHWj1eqMRwLnaXbNhJgmZ7g8ThRdni/ent4xoh+UUQbdfpaFZnKqS
LQ61hE/9mUduQJOE+PAWiTowxrPmmyXwV+Vh1JzYPQlffwTNaCNvLUoJwB9O097GzMX+PzRy/Hw2
XUq9eHdmJ/RCs4Wu1oGNouWXNfRU26mG8mtlr3rs8vVGb2SORTNcRy/sV+RzY9dNhDXVPvghQg62
lMVBfOjBflhq7ysjtGYj/0ne6SJl4GY+CgHpB0rsMBYY0rCcaOzQk7CPJ3b0CKSlfBcmen5Z7GaV
cOJHSwVyfx3LjFC588xXo3Ky6+SCkRIe3/6sDxhOENW1Znybn68lBOJqdOr4EWonEpDro5MPHusX
6Tb3fNwmnfpXJXNElIgdX2+xbcshMxoZ/nmBECxruGsea9UwuGfDbW3ZmjoKoBqB/mKo3IrMcgpS
JJLdUdLEqENtekIl/PBn9wtWMvhyq7Q5O7Zyp0gXqUagioGnHk83WpZJzny1BjKvCg3oTtP9HrK2
hTDHlqlG/Nm4WgAp/HoX6iRvA7+Wc6oGErByR0ZvJq1bORYPfXUHBdoXleNoDEy9P5AGwAteAOuU
ci6fXbzubuJxTNUsv26m6++ITghpgSaSRWXalddBLxybx41Az8dt5xAFqcdJOBRAWdz5/uo5sAcL
7LtOgoZGUF0CL7gzdD+KabP25V600Vn/xwynuoJdsT6uXBIyWbsgp6JpLty0eMSbP9QJWPqcLOmy
QBqwoYoe9bYw1rBX0i8yH+2AcvXPBWl3Vwdyhha46N5+mAe5caHmlxITurDWc2btglvbyYqzd8bq
p6fPF610taL9QKMpfglCsy6a0Af/W7c+icq72L7PJc13fk6RpYuI1AUgRLczpnBs7v1idIKDUYyp
jUhH9e35wacwxsIdUu4xwgHuQhrsMIV2tJqdh+joiUjNgulHHWFifHXCUBj6qpR5IHbFi3sFpoPU
XDPfKGl1TQJWMAurMpmb/7yBQZy9LiEJIX/3Gx19s0ZQM6t+NC4mJe0/SlDDlUSgbVBHqDBBd4PL
kf3g1FHLpRI9G1ajLgZdrOzA0WdDLTumN/y53RX1eVRX+Q67Wj4RFC00UREcEJt6aKQJSvTn/HoU
AEfu7H3+XW4AxYNEmG8Bi6sarDAeO4k4qp5BQfsh0t5o6ZiK6Q4eEtrkG9ijNo4FLCvJ6Ltf0bbw
G2P5ozJdGXEQOBlaciqEd4hkrtkzUV4UrJ3VtVLyEHwcLIaIKv9vkqu29aoubFAe9NptiexLIypt
PE7bLxefm3FO8dHYgbWBrfSE7l4uicJtbUR54gJTpG6Ylo8wASrLtXR5jhFWe0/vKtaqBkKUD0ZU
l2w1Cz/CMpAAyWa6fNxzo+klMHoZoyhDKpNUIaYA9VW/3yqGEI/PSAGil6Hp3k51gf/hw4AoLLfx
0pS1GVd01tzcXHorKSC3vyV3YYYr1nNa4xWajeQArBi+mNMSXGmFeSPJi9mWVxg5BP4wWbRDatzN
AkgMiwB4LyyH4Hj/pR1QH+4PcxeQG/3qDE7ewkiWFic0Qt++mApOzm2OFuXVc88Auuiafyj3e2yx
AZSnI0IlboydoL630FEnEitaOBWvTnmmAJgHcYxV06herYYkyCldB26x64ctJO9+PgxZ3izk+yDH
pZZOjd9aH0CtxNayloDjYicRBBiPsfpBY0KxbHEunG7npKgBEqWCO+0P6IhG0qq5hmRHCY3cNOXY
5497e1/u7T4sdlTI3+cBwJ2b8FDCsPNY1f7ql7++bXIrRx8ad1LQslETNJBm39Z/9bv5b6kLi1yD
KQcy2EOZSrNOX02nD7L1XcMdSchVb2R/KHsC7pgv2jKBIWklweNtsSkkIqgu8Lrrb+hZdzRA2Rtg
eyZmIhCQJuGzUHEXG9h1T071NZ4fcirMdHzsasj/mUg5FZq53ahho0cHmUZskjK6x5Nw2JExEMTL
Zu3TnA7+1oIEUQQlDn+s5dM19ddifyzSK1O0tlqQF6pdnjJS1pIJ54bAUsrFbHm+HURosen0rIE5
x0uEhRMBCg5QEMCTUnds9lN7hMH6urttlz23mNM/mfSpUw5MtBXaHSZUiWM0eWY1DvUetF+gth1V
9PmmJDwW8h3C2lp9Uyc6CjfE5LrUgmlYLu/ImAwu1v/5mhCb18MCW9akGrOxDPVH85eyY+zUp/0X
+TCvf0fLnUreC9s/rzoscAvusNJP+kGFQIiApuM8x8BnYqe55y9NhKvCMtBn9fTw/3W8u23KlysW
2HBCYROWIQuablK667NmR43tyNwYAY6rR1w26uD7uy2ffH8elRSHtkxWxaeOkKM3QfcWGk53sw4G
9RM+6Liv5CkBUBuZSBXvekFMCyrf0+5k7mf5p1S4cvZhdUeacxu3/1EN7SQnazT/VVgWhjXgaikG
bAQIDefRD/oUIodMo+cTw/u5f+0qI7xEtLbo7RdQUY+zoCNr/TCeYbleVirk/MKQeN5Oiu+I11T/
cO0JnZHY27kZX7ZIdy6C0BKD/Z8o7xFf7Ef9cpHJDibzUrCsyjJ/cjeORlJf0ptHvyxWUQ8Etx59
DexHgYpqNYJdUmsSebIhb23pHIM7nYC0VNfdI2HAe1cF4V0u+AqE2Z5wMIBge3lY6bzGsdJwRX1k
/GcA5AGglt2yGrYDKEdsCoNgMLmwxNn2GxWriQpUO9Y6avO/2ULEe1NQXUoD3rym/0Vbwoeb2ddJ
kvfFc4vj1GfKIzJii8DMJOo+pmC4cBiCWTL95WyfNXrZwhEW09+7dpKJ9fAIlWaOfOOE/YR1v81c
eytT3Bs4P8+1bsLkhwo3CTDoSDmiOPQOAoweyKiMKFNJ/sfD62ds1U0K0nA9lgPEwnZkQbGzv/nU
rWT6BWZ54Ul9Zg411FmHxyZ7UksMSGuPi8LknOx0sMaxhaoFJSm2QU5pdTjZtxz0Lm1iK8jhzn1r
xJRzHuetoiqVgBLD6zMNrvJSMAA34WrfAJhMVFebcztioj5Y431ymSfX+lFfWkFYEOtxLK0YgZ87
ndwtMBbtYB1FkmnETCmhJJFt+NwImzqz38Mc0wWiGDlTmr74YUE8K55RqK2YWrYpZr3LT7zmke7r
edzUfGdDYgo27oqqHQ5MZuiGHS6/txa2mQgjiZWJIWQxoWE+zbdCaGewbmOzoOuwHymZi51UwmNc
43S3742fwQZrrL7RcAVhiWFK5uXRsn+Egyj5x+BMrXj9FL3x3B++jWSZI/cTY07tHjTtQxBDQzA2
MaAe/nMW8PbTmoLwnMXciaDYd14N20mgitYxWsvHDNwnpnpnuUvPTKF1KEcnFejgETt3O6jz/l3N
6ogQrZySBW/2g2/bjD9c5KXPV1Mtu6jGYElK1egENjwfHa6FV1GWTGTDHfZcGoUY8YEaGdzXkE5Y
OTCzyFS0CLwn+jmFNYrMigUkclabdoSYw7QtdWbgd3Qk5AGnrTK0nXvPMv1aCdKaAhnv5CYz0H9/
nhtFb7XZoHRRbyEJLQdHsrY34RcTBYQJpbv6SClqjZ3hqLlNPSPHrRWELuwYCRHcRhxLC9mVZbIs
osncKNa5CG6iyd/efV18DSxMujOKP7ZqCq1TG+jQRZgObJQxoAkAxuJ5zIaPyD5wRMF2qS2sJYe/
lAdI78FCVK5QS+UwsickK104NIRbjwRSTC30I5ykQuqvuR+5iPONVvg8oQxspA5GgYsu5BLt9xGp
hwfQZO9hYFhp52An/eZVfURZWWF6u6Vrmh0soCxCoWXBR8yam1djPUCJWez0RWreaTpilrXa+3ih
l/ZQj5f6tG4gPzTkRdA+kx/kwCR1ooP6AA/7skczcTgHud9hRud65yWaC/Wj/7Cyi3As6ingWFiH
7q+h0XN5Rv5aHJhKOBs5qBjsobXz8o/jQCNdvkd1KX85GEJd3qqKaBrs4oMqkBYTcVYENhG8Qble
ueVcEJ30WI7TLsAzBozKZS4Bd4mCwWP5rOzADGdCDCOOpXj8pEVuK5sG2pWZ6QGV9s/DSv5RP5Kb
uEEwhM7j3Tbtka5YVGO6Tq1QWP8ET8yQz8AwLtZij2xTQA5nhFi+2GFXPwlDknz9qiBhkJtEJH6w
yVz+DXT3QM+k60Ir7jEwfYz+hvP6h5trCi5BVVlNxsa36P1E7IvqzZAN40uIM56V/zl5EUf+wmkM
wXkZGMhK+x2xTSaNb8eRtlMSRxpI3W0VE/2gOBF41ZU5l5sk0MgneakWGZ5kzJ/SJtilEdy6bIwX
LFBehM2hG/j83cZBhQQ+qfPp1+k20QSLzIoVDSMEXdf6T165grPCsabkOibFbHajShxjgky6j9XO
mgrFWksLNIwmLXmyFC0EO+lkwBBTMQbtXJFkPKXNzEqIFMYpkg1NdHNWxsR7o34RXhw+P1qkgJO5
YYarmsAns7rfTRNklEa8XZsR/mmt5acd02C/mkB7GBhCpN2zA5MbIvB6hCXHjculB5TCMW1vkIMq
TjcKl1c5jzX1BW7/nqImG9MJq8LjZnpAE5XqP6ZN/HTWCugR+N9MCnabbVNi6EUdFnj3diOm5xWw
5Os1lXvwEaETTIFbm70Y5mcGdIQFrjtklWHqbZGhnmUcRaxqy89Zyy+ZAIecskbGizq1G9B3f+Ci
IKqPF0/JjTiVqAhFSJgpkadW1wtwwY7ph8AvmNuaBneDA0g+9dOUOSEovJSchLtD31iJdffrGFPG
7R94LjrX/95oYUjvG0jSIabW8JKhH26WU3pr92lcDjMK3teWIyO4R5caAl4uVrzys0tHeDMyA8L3
ULmG1IMMggfE+eEIwPidpJpV9v3oxLatRuSsbFnY36gyIla6DJ1jSiIppp8IwsBhEDBwwIdoG4kB
HM4RZEv0oZ3ACUqPQFM1dI+GY8TM24MVmMrErypEH4ETo9xPGiu+N06OEC0l/9tmC5ubXr8BEmJg
06SSp1PcXQGpiQrJ0wtDsdhPbLhjkrJpt1AZ+w03ZP92ZbfnD18Sqbnvkg5ASDuQHcEc6mx8IkBI
LVlVNXHiJ0q5aorL68mDla1wM3UldV06vyOONkRIOVDBgbqZejSCcZKI31EA/lgPejfxAVf8tH5x
dGfvwE2cBSsJg3ks2BERAz7W2uDhNDpooVDjK676o6+e2wC3vZ83HDdXWwxOPDeQVlKl8Y8Ll3X/
8LwusCv5BFmHJAu7aSUyZzdCqXJXcvwzUnMuJV8Fg/Q+244ZdIe/mFrPK7c6x+7JFElOl2m/BaCe
uJV3GAS2OuP5bq2pSlk9/efF0f4lyxQkf9YStp/aWETYumGTD8BOn0V9fir4aNHygoiN3a/tjIY3
ybNiXNKCJ2VtsRgLPtb4J8PAO5TdXLpKXiXRbJXi/HBUHPQfKcPQ/6jLx1aCYC58rj8sqIZOep07
V38+3KRt2hHdJuPNZxV7onWHWyanBCsgDprKyAmT3ZboFIUimGvNmxycIj4ExIQ+BmvMKe4bt+Z3
OR+taN3GNRS6Lq40EZbYPADW4wL6ZvLdwZKL7W9trfs8m2TilIFTC0IlSBo1/bxwEN9VRJCPb5TJ
UfPlys4pMGM1KUplLMdhSVtDK4uHRytToN/WHx0VEEUhbp9XhfS68eLxIc6BvJFqfTUwAk/6AKq+
FnnGvONULw+srj8xkmwS5KxNDB4lHtizfEv9g3gIrPo/YEFqF+GWUeodXB1unpb3bL3Av+b/WDSt
qbxH4TYulyxPg3hVsbkLD+Au4NsHmWIVpbFtFMefe0g9uc34oC/6rNwtM28EgWvYB/ng1cO1eJNQ
cOvLtLFzdPqbR6GHK+y+HDA0XLlGS53I4MbKE2QWoznSpZo0CfbLilHl8F4yOyR5WpScVlwTCOrf
Wr1f7pFHsX3B5DTrZYwtZRqEeZ4i+dlKlFknS7Z5DeP1iXDNHSHK4E/VxNGuUGTDyHHltdY2iC3y
e0985BgH8nzj+SC6PVvmD/+2kNQ8dIOnAodxHusUitmgyI5Oex+ntjCC/LI3xwQW0MDTYw6panvB
IPYHuwqdiEiN4pmv6myOpauPC0Ep3J2Vr3ao3F/+2tJLG+Ve/hQRJUxjELKNhQcefinLUcjCaS6m
A0NaPgZnSHxC59DrrInNJwmDeArYcBjIk/M2q/MKB+hpCLjCQ/pFvvwseJbQpRSaWQOfdVxvvIab
qcWp0eTFnU9sCh5iRWJ1hE6LHHp0yhDJ3bGxGXcwhCxG6wcEN2W0D4fQiyr0Ixc+CHaUINFsYgfX
pqjkffuzt4gk+sD3R15rDX6PB/ms+YXqGf6co9akK6GH37ucszb9Jxltl8ejBh9ue5Tq6AcmM0uZ
N+NYfvdWlB6xUowUDxs7Gyz0z+s/ddwJsRpIJllhV+efvBf+Kwy61PENe1ngFf3TA14WqIaT7Yav
Neo2qaaWfRx6IPLcUUSDtrU3KJhPXQwuK8uN9YKkToOL5D604T5Vi0oiHpSDxmxJzB1/1WXDIp5e
L0NrR1DzdRhD81AluAsZzOOfrjzZKw5Bd7QyPz1xVhHHfnNXJr3NLrBg/Gq7PwEeZlRTq6sW3jhO
inlQjPcASCj7TK5Nc9vSLWjLBdAVwsHvohXnLBFD3gUwc3oGyc3xrcoOedsRrAswADNuD+UpsQXx
4P3PM6jP9yGRSRQSXcS+l+G1hXpef+QE8uXqDp927GUAzOXWpF2GoVy3mx2sQlns7U+jfdnQK90q
qstRGxtzwvKubAKSBskq0b5lxScyfGh0omXn+Hgt/Mymu6swzf6T3I4yUrxHQXDX6J8UeWWGoMZR
Td6klDkhvtCQxKRlzrBRvDU8gXMzHzxiF33EaJSJz++bvR2FpEWH5q7DIKIQWFouEuu0EpI/n2rX
+Ur+W1SAPXXG+Kzy9feGYSV6aoWhPjcTE3F20JLdl9h+OfapvILY+R46BuDYhOlTcUA2v3qlTSIm
RS9ZTrRWkFVXzmzShB02xg4X20bYvAg9To4aAn/W7ca9tHhCibGuyfTl25cJ4Dza44oZVs3ExuJM
72ZWdcIPPvuxZ4VOXZVQX9GSQTIIuvtNGHA52bECN+vAAWfWou1CUCarDhC+pLV+C8L7+TroO4St
SqY8rUS8xY3XgHDmOsKj5z+xyS5TjO1Rbqn4ScuWd1Cw/hPjjIpHc3qMTebERPoE4j1m4ddhBmp+
fqDldAHaEbJcyGT05C0DK3sj+E4MzN6Nufp7BcbacDgE2xawFNrBZxXSQrv4SfokPMvcHeALVjSn
CdlqhJCkG+Xe4EbugWCbXrEzi62isjRvzYQjN03Ep47jJp4kI2WPvyDxgy5WWgukc+m7EBnwafKU
Q0l6uGwU20N0gFg8iI6JzP5az0nRpbLQX/gKjQwiQ91bb4eHpyoVXtiwB8BoUNXZUbYdN7AanfIX
4P6ZkFoW0P2NFo+lOVQhqcF/HeSakUa0USz5ISlkxH21cD2BES6vv99orosfJZ82jD/5z7eYVKd1
vqWtJAm7bDlV2m+ykbkWBcx3T5rhYrY3VoAhDqT3uQof1S6PhBbyWqcwF67wLHIZJKALs2yM1iTH
8XGU6+r/lsLYFXjTpvXEtWONcP/cLf8CRLpIls7jf3UJtbiCG894kO0LCzzy5C3kaY3i866r6ZmY
qg179Wn/mq50pKOGb9WB5NF6MkLjSvDGiOmuwgiq+StQXB2iQaDpLUP07rKG3MyFrSwSNSGvJGKZ
He4u+MUWTvmOhRaQyg/RKIbrifDWdMenNgaMjX5LdGLaw7Nkz5kZgfmGOUPw8wJfiG9bMwNM/6zq
5kQBksOV504CChwqPtt5NZdUBskOC5hb88jETAt6KwuCoNLvSCi1e/hM15NVrLSK5l6t+bkbsibY
kDfDoibKy6jvaTUoosud3oBXYNhjA1x4f6+/qXBFkIq2VGmMjwA49WXZaZusB9e1w7SCEICHIuxZ
aLkkr4d/xMRVe+aTnkaQawZRiwhB7q1O79GtmQ/5X1Gjli4zUu/2/06m4ngXq5YmEoya1PNnJvsE
MERdg6Ds3RL1GQGQIlI0BccKZf2G0WfNfdhg6MIZ4qeP7PwVzWefo3OgNjDmnLx/wzcmnbkxVQWQ
gFrEmKH1BqFvJOV6XMlo5at5a9s2KOZ4sjp2+cuT2oLDhpWP2INnr1bkGbkHpIcVSRqe5FuY9SOH
FqqjA9bdNuTDcD6LehbCK2n6gVDZfZQb8PoOGNxHJHWslqgZ1x6JAWco3KaHXvqwa7DBeZyAe8zq
ey/qkFXfYRRmmdjE0HEb24lt6Pn19jsT+FrMWl8cA4zpYuU8f0CKrRfRAte8QTa1s2caTgAOa7On
064fW+MW2Q/XN8kAWox7jOo+H69tVuODLx1Vxsa7Pd28B1tJI+M/agExlqy5Y80GApbJ0HQJnMoM
TT2PAbiIZC7hUvvK7Q3yFnnL7ARHmLegYgE8ojte2kHbX3c8/bSEM2gK29fUq+Fl2CoIxA14KA1l
pTCzd0NhBF8EijZP+jUGYk+4gqvtAWL8/pCK+XmyABM3fJ2Bu4q+B+2Ten3b55ZbPU1LWajvX2v0
XmsEFwyLUV0QDoS5oj42uY170BjMYwMha9lq/vsifyohQtRvQ+4mqW8WlE5IF9HULBrqAUfERhwt
werG3WQ/pcTfsVeI/sdefpdFTkIj10ioHfkE8PdpdijVv+mP4zaTO5/jPvsd4z6BADYDYzGw3GBb
wSZCzBw0NVskEUuVx94XR3xjvjvyntOy8cKeEDkD5h6M11EjrcRTpT2E9qJGFVp3CW0kv2SqR17z
bR4tJZ9HH0+xrZAfykpgej3bY44gnARO126SdCRD3vUFN2zIl4gTUGleSgXK0XZrIrzmkASem92a
GcgI+aTJojqV5LlzBelyOseNPeAmqr23EkI42Nh0R2Od3Nb5bZoUHFOPtu+fYJHHN3ebK1yqyPLN
xs6jTx0ilv3XrrZe0ZOmQgf+hRFp3l8rmizmGiat27OPH9Hp4yGYJdIrxjMRWPJo72l2+R31Z1aq
EGQbu0XIRrOTOU9D+ytVDME5Ghp/SJa37ie8EVdCMJCWy7dNIqSeIHMfO1rkoi7A/2XB9mP4yxMS
Tc+YPwM9gDkOz4GXZ3/2cvxxBJ95A7ZotA6Uw7FWEX9nv3fmMk97k18cZ+O5J60uklsGtA2kmqin
gzVbeIjutwZM5almbWMlIOdFdWcK44+dKEs/8ucQo6nlmiRQPPPlhmElnljgs2GyCzGaHxp8z/4s
Y6zCZ7mOwtzFoSxC1pOEU5U3JUtg68Hx4M9/TndF59fQilg0Eguw6VyA0YDSrl+geMJQP6YMGWuP
ba1DEeFP1moowAwEdj3YiC2pACtS5+XX+SonNX12wj8YWDRj4caKu+uz2GXVHkkUxrVEpyW3IKjy
sb1W7GHD+5+7R+aQ51uRx0YnM236gnWiZBTiFwPb66qK24HdMPtF0kzpV4eg5p9f5pZsNdVe71cq
NtKJv2Ex9Wl0t9BEkA/G4ZZIfMddhps7r6LU+JomGVjHKdNpsViZhgqRLzpDplW2t/DbjjpllKPt
OAkTfI35AznglqR6JQG7vX17qmHJG0YWvvEShAx1rsol+z87dbhffqk2wcLDrwWFnrCPzl/QUu2b
0uS3tXY+ahwBTNJHXj584KfJSrlTKjFkyJJWPL4c/r2dbtvJqCmmBMdQo8kgTfUoOm5DAcmUGV0v
y9+Xz9OQWlRg04VOu5p9ZN91NFIlAa5sz2tKo+m1knan64FD0N79wXFEkypOnUn37DDzxrulhDcc
y6AFMLmBPjiktbNhxOrGKgiZH9C4a+iPXfFc1McOsUuPj5GkEK///yvjOqfsB0EogHhUHCNhhLat
U9sEMyjpCzZn/pjNcQf30OJRjC8CHuYaIZGm5IRDnF14wM/ihnQnKcr7o0zgt02OShub0eXr37iT
uwDniBdg14N5wnK8VSZ5spNKJXRo2iM4tzp2EtIow8eu2/WXM/hovLpqIsdPybClGXEpxcpU94ZY
oLQkqFhL/fPUwFoScx54jx4LJEHyCwQaLXWo1S2wHQPHRr5wbzmqAxbXlTn8YeVwZ2rraKOBAJV3
ON1NNZ+i61JaFPoDmRad4D5vOIWqfQAjOo76n9M1lkMYsSrvNRegL6fOIoqvmKFg126OJno/uLXV
mXxOfGqDtEEk/slWwcTFLK66UouHh/vhFgQu+hJB2zdZHzVX70KRbiibYAko4irX4W1AbJy6K8YA
Ln/vnxadRS7H1vX72UYqtNjZHrO5IpLV6UgkVxIG+AO4RWYr5Av2wroeqyc96HPcwE6WTUmE9nUW
bBEBYlnKdYPuIVf6Fj0in5SRn4Hz+9P52bWwdbwd4J/9ZKpLSjyQKVOoNaWT9mYfr8msfk8cru7O
+FomsnIxPBJB+qb4MCKxGu1IlxjzGSRbqipefiNB/dVoOXZTOK/DPHC6sYc0YyfwhM2C7Jm1kIRt
z4HzRfvDit1vFWA70ueMMefxdfOaUGAYYMfc7o1ePyvYjLeXgzoF08TkhCIfp8VYxvO1hpQ+laxI
ah63sc7FaWwID7hrvv/SDjgChP7YtHrgaBt3scwf0uQOnLcZ4dw5k6CENHnuip9O/McaLz+pxM/V
c3XsB48wxxR1afxFM/4MVPrSgy37LKz2Qeuyj5lUeJ8kpbv5eiajZ6ktlD1zR12mK/K5gIkDhHMb
qKsai32FWYXCW8T3hLnoYy7Xg5inje60itMm9yZxaVj3hWAx8hT/XODxCKTzolNk7nPmhKhNcCDi
dAXpS5hAYBYkUApdo4iqIuR7Fz74986p9OcRsyzPfgJ5DjRZ4KDE0e+6uyu9IY3rgbSosxAqMz6N
frHbNQqH/njGpGYarfxycOlj/FYrgw0rb688+z0X7nP96DVT1DHQYmC2ZxfuopDN9hMPrQ9mlHIV
8YcHmftBUfdJcyTIX0gQb6Gqdo1+mOTWdd2ZErw5STwlX9yOj6xP5zIEUZFtFJJ5kHQhoP6MVF/H
1UCyTNScOJ/Y2oE0IsQt5t2CWDrBsXZAi5oNV+g/cOs3/9YsOcZqr8EFoVlw2+/f3HmUD/LaFiTs
HI2s2SCzlOocbJZp3FKaePLDfFp4RfLQNPFbDR5xgkreJ4KWQyk51i7Cx9HJ4izF+5gnTAU/5/N3
Lnui3zwjMeyX92hw5gfaHn7RP+xXjU4WjWntJtlt6lKa5/5hMteczfLQvPi3/ByjFVDxdKmI1+yB
oWpo4AYCajI96WQ7GHx4VGzIkAC5i7DCwU6I9gPjyw8VDNz4/uG9bxDuNyvAMbvlV4XEaq4yW0iD
Jf57gtPKrCKGxLXogqIn5lT2sxIY7/tC0dxRwPoWoeMo7lqzfMPonQzdTCaU/7VymUCEuvwmsn2t
ZrISNhOgGEk5tjsM1Jq5CBTc1qB1t6sn+vGSyv0L/VQDq9HDMQyMWNeXeVubqIOM6UHTVofT46Y/
s4guJjTWFyIP1S3SB3dz9PwaLRA6lyj2s4YXHC7boyk8fHEtKcPP+sapDM8Y9N5FY4GN2M7JbHpq
1SPtKFyWfQs6WpIPZ8n/rYXleAS4tWzpC9AhHYwWWoEldZKkAknCmw/NtEkRfP47syY9ppAwIyoE
1cwFL25l4bJd4jlNR3Begt3KIj4nSzbTz7vOsTO6fgE1KP9T1HsFntPbHghIqjOLwJ4306S5Ke8h
3WhOls+ZAdURiriGNpM41UGIHa0WHiwweWoaSJRoVeG4XhZU5Un/1y8E/JHsWQGqFldCZD+fPedM
jIhEU2mohQGUkJnSGAcqVEW/Tk7SQo/A5fD5Qz5Nrr4Z60pqYZj4e4zbKUtFhVOuU3S2xU2lGcFB
p0kwuKgJjaNnDJjRKImCw1hReIX3sYvrKlviaOAtg6me4eNogqyHWceoupcsRLfZM63QLWcxZNAY
HsexynmZukl3aHAizvtPiWhchNVvXru7cAxg2fNIzIKiSupq5nvhwmDNwaAql/04m3IP3v3bQUpf
zJper5NnxwyQf408sxZS6WBUbKOTM/nXfBJZMegr2YMwFr1QfNMjLaKboUMmn6sJZ31Q1mk50uia
Diuqs7Hh8XqjtqSOROUja/NI/gl2d62VhGrvssTzagYlqGsJ5VmPO+BJq0JC9g7ujvZZAMiqaIvE
segd2f9QY1tApew/EEIaDQimdQ6BDV137eNTNTzII6kwJQI2C4fdMEgxXGiVYGKQtuOXRfOo4q6d
lmUB0YDVt8E8+ECgj1yPWiaBnEUPqKxxyd5eN69HxyTFnKEsGcWCo4uVpnwP0g9wxUCG+eeeY+tL
c+0XRIQjVlo0pmz4IgDCUTAkbhkTR3awcOhZAGHD6aPfyXtgFdZ0aX7u/Ou9gqXAqhcQNQxvU+dY
te99rHUS+JQSzLYjhsl78czzg5ivMKKYELgCCBcywZmcI/UHuqBMe3X65e+izAl26PSHo0ZKTvka
gro50jd9pK0boCUGTaGLVOv8q9eiyVyGVV/9hox0PhPTUxSXDrNZfTeuuVmxfkBTjO4uINjlECdz
mdFsxFRWuLIwoeyem4oQdTIp9npEpY6Z8GdjG0qO1gtgi6iXjmTZFqoP2tR9FKhSrvedKZX3v2KB
IJHI9KzWCkxKewW4B60Acnuzd3/Rm8DjsLJ2N2HTcfmO6m4fsT+gfnQudoB+GnAE94PR2WYDahGc
hmq9rfistuCvzE68tTrf226J1DqD5LWRTHUtNo/wr+grP8cZVib5aE4lLwe+yNAey9uXrCKNY17a
bnyc+lPNScLWPM47d2e/Qvmr2AQzALfg8nrp0X/Sb5Men7qjCjZkcAv+jLHzrLpHVpZguXejvkQ/
AbdrtB9hvwcOIBywLVg8CUJcCpFuad38NMAs4edI7PkqQEVNavFDO3DkPnhnRPeQCFfDbMKVMGtk
HIFOPD+0VTOnIr44KL1Fqe5i1RNryWN0ytCXQp7UrmSzpgaNU8cOi8Zc0w8qQlQ4TtCBcwqaINrB
WdpBoJuwMvTFNlISlkzvYrgDXxEemsuiNfixZH7ngXoGFCDa7aBqt1fD6e/yicO60A4cEdHpVGPm
APNqtECxW4dUdc0mwX7TT/7Cjq9MH2dllIhf3w76Oi7B+3StfALcwjUKE8QzCj4M3bgwjqY1G0bV
jOKCW21bE/f9U04pF5Di83ljvjNOjh/gg62IkaW8MRXhj44pIuORzUdxJMDJKKK/FYYHaxAsn+Tg
IFFf8ZIv3Dimcbd0roRPRs7KCO157rkuMv5b1ka2VsQ4Xl/eCKOqVfSK9atR2XvFivQSLGNZeG50
BW7lPYqe2jt8jcsyUsPAhfPtxBC7+wOObpsgoXKWWfpMoVaq2Kk3lqfJu2S64YsrcB4E/ACj7IN7
BijxWZyhwGffksKFFDnhQ4FXvcMODupLsKt/dfsnRtoYPBhqfZ3r8ycsLfbyVvbCxjyRmbGx6Y1l
Ryyw5NoaDu+FuVp+N7JLoVvFqihEDM/51dkL56KSDbNKkJPfDW5HBbe1Osl+bGIyyLs9/FETO1Lg
eqyrYNUqO0bJI7qCPUqOMQuVoQp3IWFV9V217I8/UHISk69neYmAsluPas4xxO16CbASYNzlScXT
vTtJY42HViqIyHWGccU4Sw7CCnpEK9xEsG8BYUmtnsHbfYieryi9q7odJYa1zAXfz8/4yDttR+y9
+SVVhtPV0IpWNz33Z/SjJi6em8LflTNfcLGU2exsivqkgmuZUyWjLncyZNVG8o84jeeVZbFrSuOK
qsmdu204F68EDIx+8pOqs2LdrfF/Vo9tNdnJLJVE+Na7wjF0dLysTOtBieI+q+iVGlX50sGWSTqE
hXAPwzwOPsKiXyLm2IURvT/V8Z1dOEdpILFhCHfQcooKcuL9OU3GNRrGtha9283RQ435Ru/v6API
Ii59P2sDf1oJm1oDkxIqmBAa0hvGMOf49hdOinGtlnfsQFesgg52+G3dt1/jJD5oVcq00MURhY5Q
alrSkwP4Oz3HXYUgwZu/72B1TYyRumudgy8gKZW0vU6IHhXFbQRDf7qyt0aRCqd9XEu8oHfHvbw6
6lp2jPRth2Kc8g3yJW+x1mIhuKnDBfKL73nlPY5UDQi5TJoUefe4pJ6IksyOYRONVXwVLtZ2ca1f
aXAXJOaOK0XtMx2Phaf8MnaN0PTrj89YX5NmwbrHtMkX9CnOMILIeCM/qkbig8fFE8yzeoY3KhLk
ytgioj7RMacycpWhRRdWlhL2wtn+VUPw20pcbOQx6KDTvIIWkw+Iiu/57xd8wiYDs0qpkFfWA/bH
uyYOWJr3XhBHV1CjOjBenrq7wGdCsog4EreM+JVkPhDaxzvoDGNp30+b60jib75xC0SgZnpDlkum
JeXWjw/IuPtrxdZWiqPdsSU7m5zwEnOHYMntCYFsOlRZxQ4K86NZIsXmeYei595TSD7/8PYGHVbu
NZ6yjoFK24q2aho1QlY5U4RBOLOlh1CQPmOqrPzpV4ML3O72GyzBkb2KjT637uyZDFAD+Nz/bInM
/vy1LLZZKYVgfX+xftkpd4CqAChepYAMTJqE3HMJiOVB0Yp6e2VYhjMjLiITWypSBp13Xj9KetwD
K359VBTPbezah10OjMZc6hPk/5xpSyso+2mwNmsKug981J8xLWjKn2SyPO7rygKM5iDRae6QCWQ7
H89iezy3IzAIgLqgzGCXrsyNryaL549KUGkspGfidF2KojfnCKnkeFDg88hYpdYvdCW7qL33Uf0V
6Ed/Fp3Uk7xcaB6lX2KWvpNX84LLdq1sbdVBJ1L1wLI11/JcMPqQ+srfcf/TfUv6XSRYjS5ndSMp
9RRjAjMg1RFoSEnfBwZ2siuPS46wHnSTm4kHqjRjj9DtoCppjVWG3ErQml1KkvyygZzmLoC/l/0e
jl+/N/J3RqXFG51ihJjJHD7KxKtwiIVKqW5OFV+t1BBOXiMg282C+qkVYjTvAb4Pg551gwFvEVkY
jmLJCmKLieFbcF3hWwbin65imKTL/zyGlAf7MIsMZ+KR7Aqj5yrK1YAQVIACZVF/MbpsQyPjWZlu
RXsucgN9K7nByNh1jEnWYgHbBzZ7JeQ/PFC/p+mOoX/4b45vmDVUUKv47nvxvj1zhhhXC7detDXA
75EbNHfquwUdAWYz2bTKrQ5PyG4g0Luoe/K7e2vdZI8GPK/U3pKrK3aPgaazrcPOjljD0tb/XBWS
sUahui3G/Lvkes7a3HnJkDZuj+ew8YoSROVzQQlJdElpoqkgx04NtPoOfEDzrPA0lM3Tv5mp0HUz
VNCk3cRAEe2wxjXNjSrlX0XFmVsQ56WsZ9HzR9Xka3GIKurg9DmtTBPjf6sDYu9iTN53hQNR1uhH
djcMK+SHt5AYRXDBBE3hyEsfyY3H9g5Z8fouSpKn1oc9tWUuCAIMS7WHWnB9FyxBEm0JDVjVApe7
uJS+niY/RsZNxQJbdBjtgv3mdg6CMK3tsWgZQtSsYe4x40EOljZLOuJkP1O+dzKXatrnOLBtiAi1
N9V6xSc+TZyhGlANw8cIeU8vY4xk/YQbnf/1+YMDgPdYQfi+tmjcU4XqEwTkXnA3DYRJw4EOnx46
ImcKFCE14gnB3AsBnqjd5OlGgPRDNDEmm7tGWDIf9WPvLisGkiEW1YD+XGzSW6UbBcxMm8iYjYyD
QX+wxRlo9AIrWOT1dfsjN55DsIpTlk+pB7Wr5DLPb7AZnO9dtvy9V3BCJXGaKbiL+xC+u+UtOpzr
Lgd9tHBunyRMZkDrhynD8/Nx8EpIAe5KmyGgfAAZLnkZK/Tng3ZbOC3DAAAe0UVY7E65mBbctwqT
mp1V3MeyzNEBrTx/V0RiVuZhLzh3TOMvuqvt22k5PeJW7O5AyByA2l+77m101aul4SZHYbkQX4d6
9Mzl7LE52f66ks1CH2oH2OfKxQRm7+SQbmnq2YWmSQczgMRg42r8G34G/JplzYk0UsHC5MfM8eU2
Wrk9CUptlDHCYGAdf/M+jvYj3HJ4ijgLLkqWEsx3Kz+c+7BSKNzY6G+4Q68Jc13/zL12/m6WsTfy
N1BGTOkvKN6wo99e0R3GUyUVCmaVQVNDTObB0Ay1mU2hNRsSRXBwOfIfyaz7IYGWOewzlgv053br
UymVVuFv+jK2HHwhcfH0W7nVLCd0RklH7zX4ODjmFqJyWgk4F7wohwPbLpMBYfyeWob9DWiLQso4
FcCXcJySMpb99jb4guXECikHBx4u+xO3MXZgD7Ye5g+NNdY5MthhMgDWgCI6iwfNpPvVWQABgcfy
NYkXZO+IlRE3a+A6XUSF13Z57287gOceErOk7xHdT/viNiZSddk2rgbwJKxMxxhlYcBmf9NMhXM0
hghFfRHSGlbM6dmc/IgO1wPX/mYhi6nHQAfkn0J6eZQEvrYuRrk8Aba4FysCvAezAlimgXAV2jt5
p060DwHvlMAVXPg5U8WAqOsaqvp4mAZfCzER7SVGTlAg1dIXUZ3ESQoYLfN61K6nFVzagD1XndUF
VUHkR2dRjf3WE57po9zv6gsOpmz8V2tip/jkTVY7evnwFkc2vc+kYlqvcKrWpHJmxX23CPrMjOUq
sOaUUhkXTVj//uvbxG5f1sVvAkb0bwNgS3q9HUnOC2FBhWzn5WuBJGu+MYEWYEyWPXldEreZ5/mQ
izET3qSbcXfvm3+FzkeMFd3q037/40AhgPjoZRtycxJ+raHVfk6+hrXXe5+sDa4PuNQS+fWBe6f6
jm6QxTWqzSeScJCBYTneAcynbSMfSxvN8brYW/9zbjkTvpP/H6ryKxKhto0SmCQLMSJarnCKYWW+
bWGmktEKW6qdsJsurWCTZnxk/H0/FG/YB+VL1NZZXPsS2NFjeo05fUdpJEqqE/fJYQ4wGQ8JSgTu
s1aLzHlhpZgocymUtRtNY5J8OFD0i3WS070K1d3X7GK4hYIA82lJYJPBFVtDiB1lKTXyD/y3wXIC
J6NNu+9VWkF9aPU1t8QaBNsItfq6l81cSVtP+zzThU/aaSnfoAwRWmmYxGm5JYDfrEQ0uPhwWPzk
mE84tkZGienXFY3KuDeTDBqESRDfRkfW64ORzUcao60AzjF3gXnUO7F7NDDvMZqwu515gSElREPt
yscou+cfzYGGy6wdCJsTn6F+22pBV7X4AHOD1LT4GIJHK7zR1UsX4eg5W5Vhr9tSYVj0xh/gRfMg
DkdUtjLi9xQ1kTqptGdtEgqOtNenSklDzaeRr+tgDjKw4aR1tUW5OpZAyIylk7ZB
`protect end_protected
