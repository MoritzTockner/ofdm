-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Le+bgd+JAjZ5/FTlR1N3NobE45SFjo2SvFH2krDv6emV1YAjqSaDA7pKABSmoXP0TRtvnB+euEAY
tX7kX4gJSPWh0LImEpwt8X8DvDauL4q8LkVZB6G74YZlSMWZbFFQqr7fjkQ+avzpkZ38jEM2W5RZ
drf8iX2FAwZ6FJ5gn1y5jyqKrhtoTl9qaUTQIgg9UIt4D6aIVatpsre3UcMd9qS+em1PafDWBsJs
ZvKhDSA3tu1WVUOjg7+AWZQ2RbiBH5KrdaXrt/Azf4HdJEPBcz7kFfX+koexvgLQN9wFNZ+hWAcy
d5U8EahHd4QabWekJY6sSYYJNHnteBGHLtmUGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
OmXicsJr/YA1wF2NfeXcWjwj4u9hNiMeLFwysCvsM4x6SOm1VPqTtPpM+yV9DaJnFSGUEkmvjqMK
Ii61H82/EgLDpEdkA91MGCI7ao8vCCnfPB5T3nMZyr1/UkSNOg/yLJOFFV9S7NOQNEOa+gmmuY68
43MYW91QreCyrfC17cfkReNGIWvGvG8pZ1wXoYSt6gPu1HwXuorLKFA0PA16hUWCkFQeqkuWbXA1
piJ0DM9/qS2X0R6SAbpHyXFLWo9o8TQoAT/GyX5Agr54x0mGWSJnkkF5DFgplvmf54QOHypCgaBy
xIN4eQocVyuFGns11b1R6Bu7Bt9mKHbjI1nySg+cF9JDtvD4X2GKIMHseLkh6zWnQKspm+mLB87y
6kBVmoMUbUvgHBhimnIxyfAdkFMCQ9jmykel8qVzCZ0WKM5vSm2uLn832FxPx1FTyCZspcBMnzDv
AUV783fxg4pu3Pn99o/Dl7A6mjCIO+MfeTu+8PqLW7ZDoB4FUsYGgFGzmFzPbZcHZzlLoz3bvtDA
g7PtiywdNFdEeZ/jdlFoWyYaEFiDc/h/yHhH1uiNXIjuCYz1BDqdVb4w8RhrQWq4BDXWckdX2zb0
vET9VMVYiBhwnx5T5obJ9eMNzDoHzjTSGWr6bCM7JervusJe2QrFBOrXxYJmbQsYz7UgKP0hHYra
Z4bGoRckxBej85Zc0dBKLb5Mj+eG2Nn3dt00Qx73qdGf1FL/qdHAP854rG/50DwQZ1zHNB95Puq5
lI/CU4KTzuOfeQmgvkJ74X/6HVH9UiWlxa5bv16RzQblM1807qi+isaM/2Pptfr3Sjk5r8dyP2vJ
cnU1zCnEHlZS+9XvOrqcv/ssUqpVJqtYRzcNTbFGny7yszlpazE33a0ly8HlExRnLRNsP0IhWoZu
JIq33cdfYFvZvKmQ0jum2EXWHK3Wb0LSXWc8/XjuiEhcXyjZfTcohQBGVbZjy/j2CWUcPfsmnWXi
iJoqKyImKU8dKqKIVdRCOh+TRWifNiJJ07aFDxXAtKmSYryUJC+F//TXHNwl9p7bqv5j2kMVz9Up
//HRE+t3HVXz/oxiVl1qMqwnd7M9TwU8tLcD9bJ+zPjvm9j9U2s5xCD6SMYGJY0JEOklNuHvikex
NLmdsIn7yRdxmKWPsz0ksGwCNRFv3n9mT+VZq9VBxJ/+6OiTEXbM6VZImF5ccdyGoJsoS8Q7feia
gkCb+UYUp5zWuIbA+oDAjeR2pyoLN5LBh6pm8XxnRPr9dFCu5NNBq9yq9WRls4QMZi78Q94jev7W
M6mkOnocJ7yRCTWeGENL95vMaUExt1IRm5y0+fVwPZw8E9K1KqYIpojPoSlUjsu1oj5OZbU1vUb6
Q3iD2PPuzHDdiV1uT+w+m4GUBnXVCqfLSWXp2s2/kyOGI7HOU2WIulRmItkFo0DHMbdUftRti4h4
36kdot1nps+wZSH3N+VE0RCwyjVh0BM/oQXgN1vlU9L1ihMr5iH0Z9AzxbQSgHyP7ycMcvDTR7w0
JZ1ws7qa67jb6PAiMnrZLSEmvuwE97pltJw6bLoEIXW+eEpj0WJvpc5TUg8dw1jU9TWnVGd1Y5VN
mx0o3sU6w7UGoqt4sTXn2NjdcpM0ZyjEapOh9gBpbCTmCa+NRWhHVD+MHIkupSEO1zYaQ1SRUYry
bR9V2jcBmI/i9CDIbjcK3b15Fir+35mrLUjIhXXnVZ9EIdFdh67xqer3FFdOSOpBU6smXX0v5Hf3
st0lyIIoMWJRc+gn48rBO5pbeE4G1IWLhK5lEHrAqD7+3xeHuqn9LC0y3YwWVIqG3j5X8wwEdRq+
wNm87qkhOVLxyVEEh31yf9eQ86nU6ZVPFkdL+cDp+ll5tE6ptSHbt5XVkajwhhqrZcjRbjnyykC2
thiaPweGjZW5JERfhqtNDeaIEV8L5OzQFuRfCQP7vw55bjYCaXy6pdBBCvi9rRwzCi/v9A69Rolr
BLchIeTCk8T/Yq5SiyZw7iLoHgpgW9AWWWtkgYGBtW+xgrtgOfSozmkUVoRk9/gxaU5lvqlN7Oyc
gL2pIUNi0IJ/MyAd5sk7Tlo4G+Tz7rCzh9z0ogKigop1LNMCtJrMoy58WwoyD5K838b5lNd9wsFr
yPkIl1DLBo1+D6zxslG/iB0nMcfo7lFdNSFrLBlUB/+85cED1MfRyR0mdZg7QtruOlMa55kgPZg5
p8y2kvLJGLEbaaoFaXvhvCHUzaCQl9x+qIY2MHseBf1QuARjUndAZoVFj1lCihvhfCM6YroioXOB
WE2Hc4iqVA0f4/HtYq61db6wqMNwO89ww9VALaKbijjirjcJEMbDZb2WzPHBcY6YbIEKk4r/BMjO
Acq1au9DMWnbe2aIBkeVADpuFP+KCvLjc954saTdNoH6mjUeIZH7zXQq6RI3bdNG75Z1pTvHtIrc
KN7BDg7Jjymro9lJjaCqtpPQJ9wKE63UUBw9akyzLe3RJWyzgo0BLjIzrmiWuNq0Pc0Q3UC4Yf7Q
kgN+eL27x5eOagWyMdUC/nlKLh1sLAciG3qiTQxUVxvYOSBqJQbjo0N7ICQHlrpiShhVbElOIxzV
HA2xBEt1uCtieLGwbyLFRU62RzCyrklSffZeZkLO+vylhrFls43p5e7qC/ybsf/ZmXinrXma4xfF
LlSclUx58r5EWfB4T03lt+6xK44+NKRKKEniKKbqiAAEOBrfmKNM9xtn1GlEByNNrcz0QXp92vzp
mp3GmPCOB51qe2yWb3OwOtjrRnkTwdDphjJHnbGPKI7aWXNo3Nt5SmTa9cdnWfEKblqWZvbAt1JP
kzLLQMhAXVPOvS3d40EPK7/PzX941dPFAcnQrv9box2cw23K03UGwz3qE/euQq1TwR8mYYSHxtkw
RKNjPwWvm9qU0Y3Vz1GDM2og7KWfvlUkrtODUWS81T8ng7bCMLtDBAr5YJSC5fWaoz18QEqrDJED
WKuENipwzn242CxW20bNeRAD77uWZkvDfuNyLsmYgV6Ozl5Xzwa9wGm7TLsoEqMwKO6ZD3rqIIfz
1Xu8Ek70HAdI78w9sub5qVHUhxvU2pChE5X1Wh1T1KrVX1felr/RzTa44XK0Yg2IoJ0MeJzusXMA
/QmoCA8TNLizqBRdtEcvhWcz+qDSI5MvSz3WUYjWtCGV3vGWXW5CPbb9XqqdWrYl9RXxy30W0TC7
kQ7KPe6Do9a6M7tXNSlRMxByYtEKXpdAcxKtSkD3p/6Kchu/Wa7ylXv7Z0GKUZtAkjbOVKnRCBs8
OzP1/vNMZNEcekK4cmenMVXTkMuiyE2chYf+mD1qqSpmInm12gRrIcY32Ng4GB0FNXStd/qRLzOe
uxO3JKOHnaA7TqiAv/SCIThNnGYjwlTxYr10JkYxx5TOmAq/otcU/9qrt5Txv52D6DE/NnCvoELJ
E98thSWze5+KKPAGTgWqUBsU5vhGAub5ffeAzYkeKxfrRINg5kK60vHkS2pxQ3jrpQXfidB5oZQV
V2+H52VDk24ZFeIXaNjeeb9PfDIFz1uIr53LrO5aCp+QTbpq8+z8PKOJHhXH+vVD96eEkxieodod
LXUEo8PgMfRsKRYaiuXWeD9uPEObis1IsyUQrAFceCn+fffxLldgd9zmtE6J6pEKJzUsoEnrZS1v
ty889nwdIAlPM86ITv77YMtJO9iJF/7l3uOJsUM3Tk8X1ow+2z5mevkZGHz8/E4dsR4TcjXr25bz
Xmck0XqZ37DdsgPyHySPk3oeelDIYY+hvucDCeHQ9kYtHc3xMB979zeB1s/7ilMMiVyUec6GSf12
4IPfbywLowcKLYxfFeLcTc8Ky8FjZ6emAdi6eGJu/NRJfQyAo10wuUA0Sm+o/rjBsUcJ1gflVOk/
98h/j83kX1QgQPa2nyIXNY2ezXMbUM9NVtCzt9n7wfp/jR5aTdphPrnwPQtAR9H8E7XYz2coPphw
966js/2BnJfhQsAYKPW3aoBpo49dmDlZ4Vb1ZVGwm/FkXKmxLHVz+bf/7FavkYW4jRFGD7kQ0v3L
dZrjlBYK3CSqh93/pze7d64WTOvRt2UnKxRBqdQTd/pGWsgFwBl2rnxiyp5ml4j1kmCIbqYkF/5Z
YSdMawOkA3qgrUBpv44gbsSlwZErvAql6oJZdkd0DOkOrz4CFD83qyoWD+BghknqTJEnKUTXQk+1
UuDzLAqD8zHrRKaTVkyfl5EXDIBF4E2Orstb/18EoDNOqXL8rJyUFyEQca/GTz7blYt67rLKVaih
GSB+9fOEKrAI7LDez//HEdjPZkqXa+bVcnttkr5L59303NzkulAYcpXirnH8NFo7EjVs1Kq2aVj1
/euHQU2DOZlkBHal0+9LoCKfdJr1BSYZ8AIAgDBzJ7YWYbIxXhav/nE0VRrpLFZHgxX5KbZHQq0W
uSMtAPMC9tb1QR7ZsCoaKrgmAdjOpHPCgttzI5ggrUNiLDPWlijy8Tthvt9HaxFxvmxo4WO2TpuS
tXoJHKJQJ+yB0CN1+7Dvw6rfgE7an1zzgLfA3VDu0T4p+PS8guL42Dr+yfHS7cCq0DOSuLG8MNbx
TxC95BKdtMp1H7skwFvl09mPP1D36DemcRiWTJmrckhu6S1+QelKlOdhDSvE3xDC7wK8rTaHk3dQ
jMTcRBMLEjbk0BZdfWruO+XSsDVljBZRTNvagYiF5W73xyb5aAXNb+UMR06V3Z2bUm1TYfx9Jsb9
yijrOBXX6pRWkasVNdwxTzgWbXrd2/Oh/rIGsBXNI4dmwNDTjD72jsQEtVEJmtOrxh3mp2Dyy+uz
NS9khpNkN/VjPNjbvOeheZNpUv8c9lAYCCrRZUsJWbDJ1rJPFioQ96WRafsy9lYJJmbWQYWMC6sC
Ge7pRk4TzeT7XyFsa/MOUSSbPIKpvjXOPOIyt0Z0VJFxHpU9X04Nq3hk+jIxFoj8gmhw/L1DWArZ
W2+cUS/SI+kkZuHQYMZNA6EnrwWkwURk7wHBd63FeI9EPwNw1A8V6/ysb+mtzIFM/ZS0wNM4dgYp
NAXeL3S+WG7itBEhUxERO0cXepAy6Ejmjct4UBJQXiqb2qPPXm7MOR71npY/eHSEPR8RvICmU+VY
eL5ZxQHeNrk3zCsXV3ir0aZsTnj7Q9b8yonCZtFjpX7dTWzU4xJfYClWK+1JkIAFzj5sEKVvlUgT
hRUmcVblCFh93t1LiIoXyeBfSyTQHiNLg0S3PigrqfNj1O3JNs3qlp5S5AYV2XsKgWOA9zgpDJ/a
neOA5blJ4vZn2ySdFxQIPJqxi01VWSIq1m9xO+95ohjNir7fzwJcMSyiqUGBqsh2NdlAq050O19Z
7pf40lxhhnTgqmYjzns+n5h0Jwb2hAgcrkD0rmUq4hnQ2fk8M+kWWyUc1P+AnKYYly7pPioxRFe+
WhrBilDWI+yuvvnSFZ/QcwhT+5jfV/CzLyzBml6YMJiMn40hDxfDskP0bUKcikDKg4tLwWgEHSZR
K/L2jhM689jWpNeugFBYcsWQQjC29zlT0Kd9CjA2yhPlQoSDzuYDzYE7+SpiWNTfUQ+/Gb5ndQhd
u7bOYI4Ev8XJfzWUegrzbUT2AKBP1h6QCN1nP98Iwt3EyjFYLuQeFpcUjIl3mDlI78KTbKFB+aY+
ay98KR0cwhvGjmRMhxc5o4eWBCJq7t02ErJdtGVIFrpe0/1AhZHPSWQLcfqU7VgRA9KKKzyX15e/
RuGgX4gnu8HNLCzUPz8miY4jao0pbsyidGQ3ViO2u73lAe1ozX2Evc6lfLvLga6W7MaRMq89oviQ
y0XxuxvOZGIROxsA5gp4RbkRHz9XYzPCj+t1jhWIpOVXl3JSGyKmO4MPggBtXrDAMPkFLY3SoIpk
aVwv8CPqef540iqtWtRiwbb7ViZZPtAfV1gbvPisuTQZYfztHvDGncGPSGhQ2ncRIw1GbHxrdF6v
x7+Jmtu839ClPVvEJuqq25RJWFU1PTH0SaVTGR61n7GiwnxW879/RpCKd8kFSxHjle0UUb3xqb//
r70FOh81x2s2KwVtgnwRWwUBF21XJnrOXJuyoT/4SjSfCoYmckaeimV4PXumWxNIBQkUVEIiSHsT
ppbWV9yT7X8ZYd0LEk/pFPdf6zOKU5pIYMmFsF22q/+S4Or4HuQNi6hO64xj+XJaNpIFKsk8sGVt
sbeawypLsOv9y5ld3wSdkH6RaPt5bMeVtyLkCK1s1M1rXnPl1/RRmDqUv+4L+xFo+cwrAN6RV6EO
T1e5VUubup4rHWt93WnP//6WiQysewuoS55pNGL2E9ExtAKOgC27LRtU/PNdRQa+tvQo/0s0I+9R
KyahnCydo6i0U6QSBuzL21R7AHfn5teEYSr3oKfo1e2LFmVmJCC1OfLRZvcLzDsZZyxYuDGnWscg
Gq/fy1157Os54EuF/IB65VaJ2zJ8RF6CiIvQXazSPeYOJXlqKqhqvivEMkWnal/kS5tThFcAWXoy
i8FrWDrdrVioj4ZUEMJoIylRwb6R6pg8U32UpU9xRE7SHcB0Ak0M6lM77GZPuCNzxHem94XI6ypj
G5/bd1BKw/jKLPMyh0HXf69joBEydOlA/+LpwtoKa7A2O0OYftkzE8v43mZzHbAHDh2Xwp6rmKVj
Rx4EELiqY4hzPKImrsHlxWMpvQKVmzix5zzdic00zBZteuoJZvMRedyV7+IOm+3l7e5KCROPK6yb
ZQHXZNBREfvrzC1/U5CwanSQMMKSasJSNK1xuxHU26ITf4kLO9TOOeveHhKswpJNK7M7Bm7MdnL9
75EjYmx0YO2foqRGFhan+LfdJca93G3pXX8bSUFkQRDjhWpimPv817h0zCCmUfl4orJlmZrr1M64
DtdbZD2pPwq3JEELDRCM7pk7CEZVTwKZrAt6kH+cOfCB+tNGHWVgtj/mgn5zpIqpd5Gwde6K4iYf
b11KHI/wkJd9ObosEjh/U1XwhC1paaKOJItE8pTPc13dRoOSqT7GblC2l/65IoLRK3jsYlRrHGBR
OM9d+iRmi6dviOjL9cvV4lIYW9miOYh4eCxGzFiHG+0nRXzG8HlprLHP9gN6op1uMiudDlfrVBwy
Z0sjmioJWMJabtYxRwSyvCFmjQBQpmZYl2MY8GHecpG9XGm4ogdDLU0r2fQK+4DOjN9qF28fTIuY
mBLsP5YUP1lfifeH/xdmpJU/dpYh+s2a9RZ+QC6PP2xrglUAfMEHgRPYz28ZK0CUipnwr7Bhxmsl
xYPsj1q9lsuj4EF8xJS7lKd4hfEjNVvXcMsFWTg06H/r9wI5QCW7if3Yvbm8BRzceKpJJ17lloWP
zU2NzANCG3k55RHIL0MBvboD8ASNsSHB7bp2gMFisjuS27rV+b2+XpOkvlwQl/dIOSt/M6wHWunk
wJBRu/oYOP4FNKO27dkgl1olQuB4zHbAzHEFdGlJ9iCKfsN6qU6efZsLdqrLU/WHXA1qpmgEk/tF
EEaiUBRkXG7uNNjffJaWS3fBrkA1/l8hfK9KVbc8Amh4Dg9LKEZjm+fnjgsQRyJfwuDv2Nq/t+jv
OUiYCl9hHj0DfE8lRjFa0mzO6n5Xx0Z7WJ7J1LRceG8bP9jJ5FmqMngIcuHO54q0uoiNEtZfgIvb
aTVEnDsVQ/hX8El/HGrkKZPG6u6FufV030pN2S/HjWWxwXuvSKSIaQcy+3Zsk7+0tGnEh/gXersu
P9C8rB7Hwgf8mM6r90941ysm8DK1KXZSC7mCp9mD0wRrGxVXBu4x4nVQYAknLmbtNMs+j1Qfjm8y
6oynkX3IhF9TZqgjW1eWfnwbmz8SY69R/MgqF8gW8q1PFLQgPQyoWgP5pSUWXGaBbRe6hEIONBmm
CxqSilE2YVX1sU0osmZnXw9FrYmr7z6OMyU5mcWogMZKS6yiE0sj3WzhXohC1VuiV7lGGqYo73UI
idneV9ozfx7IiWpPG/1BoXhrBWBxVzoxODDDRz6YyTh+a5dRerH8PClO7K2SeGELKU4G246Ux/4A
X94EyrR1c8eZk1pLzDGoIOpYUChE8C3RKob8mrvEaG8oISEt4d9OGbLgVDpBJFdBYrAdAiU6m+3s
uo2QAU6wQApyJBEjgq1zkdAoLxnKlplb0z3BpkDwe9hGuA1XISW7sAW4/vgR/xgsMT0ep4tS7Swc
ue589WBjm5KdivrM+sqVasJQmZ3cgGBeFor6ijVR7af+QChaqqOP7U8K4i2XppqCak3M6FtQodeI
Iq7trvmQjVgBcSx/TsUPNrkweakt5bGW8MTGpNH66Uxp7xdstvNuhiMUIw5M0QTzIp65rZvhqalj
YJnEOLiF5a2Z2wTqqBV87ozjwo6uvfpodrutWqlx8BsE4MNS70CT/5ZmZ2hT55oSaXZZUJ+7W5zY
Cc00tfGfTeUCFSm+pQlmHogX54ywkhgeOo5yPm+Xws9vgpSx2RDej8JXYKPP3Cg2hOuUd4D9LAst
n9GlixiMHVjQUH3d5QfMsv2CWGKjLiSuqmkKlcDI+O1pXHE2dI0gwIKC16TCEH3hMyjrucoXazRq
nTNfNsJA9BeMEyXe1oeNbHfugL4aXzaUXYwTg0GlmhcVTFR/pXbMe9ogRvq7MmQEbWWNDR7vxiHi
k+tHgXxMTnGihJbey6otUuPOXyuBfkaemT/AMoxsD5UpxkwahoQAELDIPZGPcJwVMimQm3L0CMyc
qKvH6SrxNcobnnwZjCyr5AK0vsh9w7tvcAz4eTflpym22RJspMDi86/DwyIFECvPzqlbLwiLZr7L
nJBlTrl9iDQIHKQTgOvdlkdAvvch58KaNcgghgVDlv4OIB8lMjTMkefk8jjBj3LIVJUWWKBxzG+f
YFYsz1Pp8TCG+et+orTS199Kt3XZXCCcCDw4m8AILcUNNmm+mQYja7rVPwyt2hfza2/RjOHkpJwW
XLWQTssdG55zTMH5swF+BG38uJjf1QU7eTQv+IXpwZTBDsEGKiPCRE6n38cDQXjYOkNReoLvtbFS
zzb0WKFy9Gfyb2RszmRf7hsZkmL26rBNTWYVGlJoQzQU4Pc8NHYWPknK/YpHJ9FnQGoFuZ2XVu4r
XTonQKCIUA443S89uu9X2FLfQSYSHVJsmvKxyh0lMBhisuhUbYuN4IdM7xqcjVWhfZg1vPCJgQ/A
6oXnw1yQ48g7LF+ndA+COse8uu5N8P8krK7fWNpSTMMJP0UAndcvaJDYggsdIfcui7m0aFPMLEiR
sAxs6c0TBddyKrE96G3DBi4HHB5jwNhyycL9pM/KZznS8Z3jLpJ244be3RirCgNPOLHtgyyzHIfv
P/l+QPSsxGXS/V5/MaLT9WkhF8TLFdox1ixd+l+5XeASgb1anPxE1zkCUUGEPst8E/YwOFge8N7h
5SmcMi8j33vzXdRwgN0TEhRAZxCWf6htol7iEwnwmmQPgd6EUaAHsuhQz6ENAlZZx1IfyLhrsNwR
hXKoMrrC9rMAJ+Ve99YfVERi4DKV/ALWkc+OopVfZZvc5j1Jt520yADtRwTKfJuudTHSqkX676u3
6kq2lTN+HD8SRuMlavrYute7btV+D0krP7iFI3Gg9onXf+xKoL9VBgCTvMGB746GvK8Cv2JLvrnV
lQaPgGB/UQlRGHQymMsTpeFnEESIOdjUevoPmLw6GqlpsHWhkZv0pUjYwlWhr87yVKQUnZVdqYel
5fzG+vExOTXXIGxEMDnpVcB8v8Dw001COGIAJvXzAkfr5D46iKNZhBWTgeevJS1iNH98wrN4p8cN
9Y3flrQnQOO1jJtEzxAqhJRk8WvMYVfNOHRUVL4l7cKjLVk7Pa3wPsQlouxylu0vQGWkVtPt39XK
QoDyfbfSWB+koPTVlW5iDDcIVygtYQjpvOGEYKOpC8q5KmMdIZ/nLDPoSQXz1+AgpQ7SCZLCDJhc
PlkYo7HIj7MRCABnSrGqqTNSvuiX+2ICPcze9qzQod4VCHUXS1mPKPJMtlYmBp6L1vTnDbenWXPz
JXUxTQ1D0iD7E5jhMHnOoQb9oyCU8j5D1OoeJJVQRPEGMvDARQshKsHPvfmXv4xQZ8/AwXniILxh
6fj1fJ++vq1ZAovP9F5Twsybbto6C3PScf3qiAc+HHAr5iNAcqL/99D9V2XN7bAqpu3eb5cv1Zw5
Ed3zzEvjHSUqY47Ey8GUNnKTOoL6ciGR6a3kQa00dM8WWI95HxGoq62sN+VE7YxAJRSXC8LUGrbP
WZkPY1k0wOgaGNFab7vprmgF2JcHmrhMtvzyjPLFuxUz/BzbQ3UcjxDbMHS44LVg3RcNSQOkBeFT
F3owOS0UehTS2LaYI5vrDFKO0DnoWvibnvF9siYmNcH6buXqYUes3GjuDy3i0c6ZM4QHlN5VNEW9
L3oNqQYOnBEj+urLSrZ7PbPT1HnQekaYHjRRUxPfEeG5o/aL8Irv/r+8vyfBFSYIGjNXU3mTRXKH
tmvBQ3u06J3OjOYdtEPENBiX1Gwbo58MfcPsvykVLWEbqYLL4sQoBKTDHOUtD82MlAc8ypczw86t
xmN/UDoZVrwHFGhE6UqPKRsNDk5AUhuoeq3JKg0Pq7QlqrCYV8xoxMWTObimn2yUncQw8cwtZHZ6
hoJEAjYCsrjLNWUIPAxHqGSJyjc1rNg8WLDU3orG1bSO0RPJI1L6405vE1yf2oYfGqO7jNY5NOUr
U0Nw7r1KGh65KhkI5ktYn1TdGX8djPlzFTWGIw7ONxnCvO9KkK+87wVXPsM3cmhrFRmLp4D8707a
KK2SXoXTLfAtyfaYY9rMCCKY6yQz49yXZKcxOZvsz93/lkCs3pqR8uPemGaxA3woEUftXTYqdsQv
mhponAytm+1UgfKACTHVTWAQVvPpI0CORPxyf8C/VFjQsBvtQnTAS1TG0kZlU7vMKIEUWD8VGh1w
xYKB8xX7sASaSotUbuqZ4fdAloA5RDltU45w7W1irzJ1oGehDY22cYeiF02LR3AMqJQVIhdF1o5x
AgwofSsx/5QR/ZnFESvv+mCLgTOiYkUCTwNOAThTfjPZRzxCnh/GLLX2FcrKPjFOzSD9cC4FVDLE
fegk6SoRanSr1IpkWpVRflRUEkLRdxgBUWFP2U3S7Iy6n2EpYZeCOKvS86itQgGttRxuluFU2OXd
jEEAluzN2o1GsontI0VS0YSWaarJloRIZvjgJ0PzLYeK551pAcQwNCDjD4AtZ7HzA2rxgKOGeK/Z
lPQeYFOD5rouzUjU17e4pnWLDTnYOyVFGx+rHqpBwhFemVmYkwcKPYtiluI+FokSlS9rmYP//nyG
VGkBUrOZGSEkjGa3PAS+6P7R5H4Qmxw637z2PpzCPvtnJVWr1TUdFfldfTLrh7JSTOubhYvxc4aO
xtHRtiZMg60dXzvxBF95/Wv7D7DZaamcpIEA+Ur4aDIzpvbGtoYp68vB5UhjTgt7cylJIKEaarfP
9HBQ/qQZWD7pnDDOa49VA4jc6JKOnd5A98PFRxHhJrOMLeSaBXfPcOe9IRfGeskGXls6oeNfO7/5
7F3v5ziyFOtqusWHJ6dTkSthp9KwTEA+E04MilEjrqQ22QQQZ2dfqP7qHz/LFU/ek/tFAbfDR6eU
gnzTjoVHkTEmsf10aR/yKobRtN7MYc/4KYaBHtFP3d85poDPAOTwXlNJdFvTI9Lx/0kLTkO27XsY
8tB5XRmtoTAcvif2H+6P9h6HtqYAnW+bbg9HDkW/soli0C6+HmGzgSt0iFG/kqlJ8XQPOL/r8Mr0
6wZ5ElvPTg2/53yDRsZ/JYzFbynEfnVaTSq+NlEYLF0tmRHwMFZtAxSYF/RlCu3iRtYstF6oVIPt
Y3yoQBUZxqS5KLrlFYTnbXAfoVGAZwwLZ0ynrTErJkZB/Bk6iw4EomCwPi82AiLpElWUDbsbG3QX
ufYz5Fn0cPo4cmhF05VKqR+wHL68Wwv+hrxNKTVpwdCrzbCpn3K9q9inXhBap5SjPCtBCiGfYkv9
1/I5yZdKqne+baGJB/Qzg5dG6DPBe+z4La3izP5RUWwwIm9FVQuY4YxNu6SN2nKH18crMaRAtz7l
G11SoVwq8do2XV93Fp/xcEWuKEyOIlSat3Ct8WRlYr96YNInD51e6qRtx1T28wuqpNmGATSW5qZd
oZgwUrJZGOLQvpyXsz+9W8tbA4kjgXaDzA7koyEb+U50zbIyPNoW506yJSaS2TIR6j3V3kE25cWL
9lK0j5OJZMA5AT+sJoVrexqI2P+lXbqFrEyeSKCqkYbZwPRXoYjxWLvZbFDv0mWrCODIS4SXUxQg
9T70QCZen3BxBksYtng+DsBF+3WWPttqu7BJ9Z/NiDuwVA4Qt5fifY0vcxojMr/KsWPud1iYMlpe
i0nEqV6p1hR8sLWuQnm2uJBWFpil2FLNJK52uAZYeHGKpw2gPW3CpKZ/Chg8UEi4IAt39nI/O9LS
cR0NbG940QwkTe6pzssoFU7dSttYAvnQ0RIVOgUlF7GTdCaeXpqZTsNMxoGE8SxAnn7pMKBbX6TJ
KCaAgDIdwEenmgCY+kwsJXC/d0smFejmFEmPCJrIKil9IwNBlKIzmB0Jck59/Z4vLMGvX3LYj3Vi
qoYSbdAF7jU2Ev+OHahkJZL7HKXd2EGFUD/FZHngC0Ze2GwDGcydWXJws+/i/4Hs67iWd/KIQHFC
So9FLRh6JDRnMYaOga969+QdzZ/VhQYe21TcxToaJsUvHeNZqyfbafdxA7SyjlOjyqTl2/qXobI+
SqYliJxM5bFdAsHkw2Mbe5WrXuPVLVxJ9tzeokVp8EDmxfH6DgFzkQ5jCnN/vIZwkhuomqF42G4D
BYRU6ZB01HjNixMZZOkMBF0Ntbs/yimBtRPVFvBcf7xO98jBLFRMxmvyYYclTMf9fcnN8xvOrBAp
AqCzqLUZ2reXPi6qH2fpp3PphuRFI5T/3qmt2VPo3HHzUHOyPmvX/2WHzQGL4JnMQcthAHD/if/B
06KIRlDzIqKco6PhaifWqftvI+Jd/ItyYbUYzYoB9AHAhESBqmnz4H4Ev9cWzbNz0mUBSDieKsMV
SAvqlcjwEy7PMylb3s6ar9YmtWL2iiAbe48tbvdAkfihAVXSAIhZoy9nEBTGew8Xjphe3dWu10cY
mVMxOyuzxZdJkS+k+mH7LYE5lGCrYH0J6OMi2a9FBRFcdRnq0kIjTgesGaUqvAhuY2/t47hzp0fJ
U0TvyjwUnHLSmhKccS22A5zxZ46J5GttpanaKcuyZyWdC5rKeco+/9NvM8glNpBG/kS0G4eXdJ3f
mPMMpsOdzohVlqU9I+Q7Zkkk4AnLf1jFgEP7Scvx0oytxoPZ3dZBX/cghmVyteInvIXvjx/CTL6W
YXrQmRouacKsLnAZ7rHEhnjXh/untk1zTiZ2tiKo+mu5Go2ge6DMNPS+ZCZPxU780He2QPX+v7Hn
zxkGuAtB+usqLao4dmzCT4drZMeR0lopTiJdGTS7W9y25koxdJwD0+GNZSBgflOfTF3PD8YaGLqW
hKR07k0fwbTaBWdXy6CwBx7FMjJX9c7ejG0MLIreyJsQHmiGSHEbj1epnCEb80z6CZRdOEVh9Nsi
YGnb5Cs2m96OMTO4Bq2E+a8Ixs1uOYmBw+GvKYbGQt4AVh8bdvFZle+EGPvlR2JBUXDvzz9iohcm
9j60seC0AVpLtV/Xpv4D6YuPs5nmF8AgzNQ9xGy61uifziRj3++WZCz8ddLlWuwFwHDj6Q2fOBPr
p+7gYtmmT89JeGieRZhU0aNAT/zP9XDHM7Sb/zEfqXrmbtyZsxEX4XYi0OyQWAQB2nf4Ro/sP8c1
PrXSN5BIz5VZhrHRi6bECpinndVkJ9bWOUnYr14xCK8AZ0v1Cyil6PtwAr6h510Cfjc5HlC1lu13
sNW73GjxzxHeIvCZHxbNdQkayTznPS/fDKuK76Ls+H9xOKIViZPuv1Kjj7euB7a05jtzapufed2r
jPvmsMkui2RlkzHk3z3YnGz7DmchQn/VtDVGbW6n4gszZbla8GzmQ6IITGChSyLQ5S6mrCVHA8Xg
VR8AkIRMyr6Vpy4G39mrQFK6SXsVLsytogQ99JYISylTSwB0vUkESK1u/vkpM+n6CS9/7sHeP67l
64psmeEWbliR7rRrGCeAEHt+tW/CPuVntlkzqA/PgsZp+KRmSoDIdU4NVoO/rrG5xAN5GGJGi5IJ
R7DeeYJ65bZy221aXCgW7YKG+QvfKxBeNd4s6k/XC1Ylw2Ygn2rzlNLDRKbHhVvLRWD3JWS9tYpw
VBDLtWDRDTYVcCZQmObc2+BooNib+aewUScdAlHhNzB1T6Xn2oEHKDecS9TWw2BRJqEgBHwHgSBl
UHnmSDhZaHxuQAkuJEg2GlbMR0v6mLMvRlviUJnr9a+q4zZcbwW5Zk1iEUG5HxhPArg6rU24bYeS
9BNK2hn6MOaUTW4T22dHUBepcZTXN7al/9GZeyl4C7/OowsVeuqEzsKx5kHqem/WFKnNUmD29Ngi
JrmDUwFFrRYGNBpArk2NSG8FMhlhheL7IG7sYRvQQMM8SF1jUOzGf7vu3DR14Ez6KIhUaiFGHWea
gNWihSf5fLKJ+wjjoywJ6NhMjq21m4Nmfnfuhu+JlaEFA17rw30p7U3aq3m30OVsDYof0UKxH8pJ
5oE2IqNTD0lz1BYsFV766AA0YTxCn/muky2DN5T+9h6CWvLVR0ZWCS6lm9EFQ7GUqVwX9nJGbRiw
ks5/fURbIGTbSMkVbW7N0Pf5rfls1aAeJrRoB0ufYDzke4MOYted3FzQ3Kg+XrmkSp3XoGuHHy/9
33uHZjlQEP5F3uHRbyaXipAOtftFMIjRwtav5YTW2XXXKVbHprRoE1UMMTnnAqexnAxkd3vzglFL
ddPfno/FNUrGgT9Yej54ILMigLmBLVr8U6K79md/tQ390YqWy74meJaaYO29oI4dxjdU+9OlCuh/
zlnH6wWRcpafH9twh6SAxQnceBOPrjVWN7ZAc2brSOz/Z82SriRl5Tnp9fOancOOfTX9U8amXvhP
3WzbaHeCKPCz7WIGYYKUvu3F9EgtbA3RSOvQy7EdW84DOG5/kAIlYr+pCiZ4ICm6Y8aWoyoOZqwR
9iSxTG9gM5/BY0LgC6nw5TrFvcXumSoDDxGuOxktQaC110/WmEoa0Z5RIjzRfnM9ODlu8y3lcRjx
DQl5F1tQ1lc1jO1eHFRhKzd6zwDZUerxoPYs4DBwRoLCtGMTqcAphUVJdrLGZWF6n7DmM/XUdm8G
Ky36NsAqw5KSttXBeEYX6ih4hVmXxH34WV/PDePwcyM2voVhdWqey3mNh52uw2pYmHynJaFLNKOx
n5PFZS2CIHYHe7Nz/eiJZBYkJSUC6uipPiU5kODd4izA0YS6CouvrlaMeXG3AAyxrRTw5zAxB6Yq
2kG1SOIbTI+dEI8fikpzs8X4Xrzb87c2QU9WHPJyLcxlyRwdwoEhRPPcL+K6WaYZfTorPB6VQXKT
Kg5ewm4N+e6dvsbIpReA2VhRynddXPF4b6s+igD4+XdGebYxFrADzdJzJoxwcQqQT1QPLC5N8oQV
v2wrMLyg1mdaYNCLyjMy3SVNlnyepfsmcR9GzAcHwj0zKPC/PPNLyz+sc9ts9Qb+L0mCXNVvugHq
AgWSZFm+07Nr+HX8ynTWhlDrNLzkgBjxtDtluQO108RZElsQvUdNUkHoNlYSZvbTF5RFKjIzpau3
3DkW79cvVxm+W+F4lBM6KHeQ4c2bAJCkY+ExpA7X2PxkGMKOET820TL2jU41auAZTtxIjkEVwjpA
CZ8fP4dUEBgfWXdXK5Y6bzO6MDsVEcp0n4EmWaalSmAlkxhr74TsLV5wSc3Dag5XKXYEXFWy7jMn
rV+vxzzGTyYOE2DOhBgUFCd/svSMTNDwsYc7/MRVm29zTq2tMo7bAnEGIIL/Oqb5gMQV4hCzh/zz
vn3eHNYGYFmVcn9KTFTWiUHl59rLHMmOzZbIexVLfO2GaUjFuC6NedRgFIdk2b18MaBCFo2uSgCB
4GWtMMtx3BwutuB+jMJtg0y0yUHKjEGUTfDctcLCDshzVtNSeV4tQL6LqYPAd/0L/KfBPls66zC0
u8wwlBQBuXZ/nRm2vZ5dt0Z7u7IuQyievRGtkSZzG5Nhb1GYMzR5njsCThZBRmF+YAus8NxD6uU+
2UATQWSSEHpjWM0kHiI40gbyHF+k2Rg8GJB6RUqDcWzct5fqWUW+8bqHz3mQSdaHPWXa9AsXObG8
98FoXcS3SyeD8tdf5if4cJYt8jmYiuABrv+FWw5L2fNUgwEs2QYOtjdzAZmHl16/iv2JV+zx1wJ0
GgadhqczPVb65vJ6BSdRa/m4ks/TKGpKiTrHKZOchYFDOh/1WSWi+o+vaoW+x/vFddyewi47b3yf
17fWZYgKPN8jj84jSTLF/gLeRCt/qfJE5JPFC8khE4e/mIL1bD4Yif+QK3KMSWhA1Pke1SOrqLBj
/IEd9V41UHFctFHX19YqD9g66dnogBbV3W7sbY2LlPDI8cHDYqD+WBgpp/e/yUXs7j+WDWsTiECX
pKV/Jj7mGE+dl/GcspcxCfkSaK4QsJJ5D81NJbgUC03VE28lPdyjah2UOCHR4aIbQ6gTDtJaE8TX
i6SrH6w9vFkH1xV0pdFqsjeUL4ZW1d3NjSXeLwUhzRTMIcCXE1Zc+cJbiZUSuF/A+Dljuw9prR1G
3+Vlfj05dwQA/pCWuMdjAOgV9bGjRGb0kkN6ZIL4owIfxyQdX2Kmtf5HoOwVK7Wecm93td0iGUD9
dg2lU/9tOdiPZipgmhRSRW9k3eI9dt1empINbBfwlicAh82+/9+q0xBJT5LNcV5Pu9ExFkJMgJZY
aS8qk+7Py5u58hbPsSGc6KAS18KA0I7UXCBRuL9jpe/lsk1dyJj6i2uxkH0/yZxHEGLJUKtLTh9e
X89md/YKtUEMumiOjypExTwUyY4CJmEiAK9/Iq8i8qtPsmNZH/erpLTeO81IlHaR+Ft2MlzuZpsa
CE65m4xYmVeOU80d3CXdDip3sWh2NOr1K0Sg/DnWXj+/2LCIojjzGRR/NQXfpDrBKA/n8sqpS+rD
x0G6Jpu6Yg2GSRB5AfM7DHggcbpFH7V4KLiGt7bp6X5c7t9yUbQ8MNCKAuj/X0+1l+YR577IaPCX
HVSomGVgoNSuC37PJJG/tFDRnt790B6rCf6F9PcdmXFoO4D/GDNK6eROQae7tDzhz8OF1W02XIo+
kAOPXHaYm0LmhwAuj3B68wYAooqVVMkCYCFDos8TDOOZndrPxQKhtrHk/6YZQdHZUMvjIIc05vd2
7GnvJFs/FjAJZw5wtOsSteE4kWw9TueC0NgzgtfcWnUXzvG+YxYQnSlBGIqvLhLAgm172jyOqOjJ
GGbaXedKDfu3zDhqqFJkmI6WgG7d1LxRRek7kZPtXclsMMeYALFpSBwt4HD8Gv46NZo6VbBpyYHK
Gwpa6tWPHCFNCSbUgKwxSgVgSOmot/oLkSoiJksOuupfAB5kzEn3cyhhDnKmddvqDxYXJWl6deJS
ueKo/Zq2OUrUt5SGgTT7+jbnuiw7sK9Nd/M+HzH2yudzLIsHY4zyIirODyb04kG9TE1NuO5LFZ/u
pxWCbPc4rl5hDvd8jY6+cqpZcSbPUEPWAcan80XROU+8bGqUDv9E9TG/0Gu3SpnoPrKEk+8XXp4w
RjiHf509H7MwCLHoZvUvv7DnVdPUwyeHgi3/HEP1habxh8C0HAa+UuYsiqF23CeMUhGHBdNCjm3t
Oo+co3hYd4Ym4gfA4fMtRFnhW2FKRJ/NY2kTmqdu71UzRRy9UXNg8Bjl1TGEOk00/rbOE6hipRM8
F8PWCYlbSeRN9J2YWtuXa3efRBiZEMlbLqrtGM3DMG9XHKOdaSVUmXlkzV8W8NznSQvDJpydKFIp
T86UBCInVEX/JLGVC6pxSS2RgFualJxVQe4T8lJWsQkbHS+qVjfszXGGDxt/ER86cJGUBOrvq1Pj
vhzcxMus+Z1kUVck8cv5Iyqt+WAgnJoxEUk+QRc3HEC1KmzFoAdk1bzOqwFOW2rvlCM8uzezFmP2
0A2n7IefOxpMsi/0aah0wU+601eUCL+6x6uIN4++Fdc/mlTRbA9clnN784kIG7u3hyL21aQn5kIN
fNWfWzMnNmoQ1ow3llOD01zAdPX2ge9bs5gDjAwoMfLruI++2UJWhKWmkDOoS50riNOlbP9HSs2t
BTDDGxVn1VaotaQr9AAqTO2XHLBrcwW4Dvl5V5eGGc2J0lYtCNIjy8pYCkTfWGDvS44NCsEA+0ce
p5YcVaJdvi9adLs3llXMO191TpYTKIb0ouC01WQi15P8B/nfPI3r8VSxy8kwHfJxzGkC+Abi/ZVH
mJlmMbf50WRn2rBGKiEfCagDi9SXDLAx3e1+gjXJcSoksWz9PtGxAUFl/a+xfK8TRTHSAs2gQx0z
1DvcT4NLndbUStEQKepN8Ztw03ULsZCE4O8Aro4K2Sgp+2U4I6xOvjcDTL05+uXYQlfFpUAXz4Ru
JGFDOU3KI5FBTg7Qn7VlXuCXXGT0IKkYoDYDbFzmCrJQHyxFXnDqFKGtzHg7h7Z3J7mobJtfmRne
ATPe7uiMEnpga6Sex9zNLxsNQcZO7dk2DWMxizI3+/k5EMQ9CLwgdLlbHZqmfOwvU+lpBhnTxtag
FlrbPsuWi9XS0RMEmP6dPpk9S5TQCOMQNVKOVXKFXdKZE9OHedQFKnYOubnmEOQIWM25sSzaaOBe
xgYHdRLUXqRxpCEbfEQS/5IudDGcagVZOROcHV+zvz/5zu9ow1oneE19+Z5ICzIZSVCPwCFC3vkq
vdPndL64SSSUfG5iRZjxaUodsn3t6mHnXPxUOYb/r2CP+6Hba36aD05cQOYt/eZeqMQJrymp3dSH
94WOOrEu5ezjB5ejymUj13hdXAU2P/6DQpDBHEKgcMooYYZAMxhnYON3E3Z3xKTqeNmk5OnIOp8Q
ePo3XMw7BPV4Tj2NnqhLW8t7R+3WKx7smn7YOz31e0Qq8kDOq4nGM4HCxEFv2kznBR4BIgDhh6mx
J64hexhlUwnUNd7l43niZWu6+opW1yJEtWvRC3VVhpkhpiGrmV51lQA6CEuTo6GNQqdxpEkPWNJ3
UE+aKmBGX1UGlnWztq0OuN7zKbYMTzQuX8n5Wz1UsD3+2/fHVk1I3f+zzDyVdrSIvH1OJZC3YF7R
zYfbxKZl5GILYzh7CyhXYtxv80zqbRwKnBcf3PQ9UeNCrMBZ+RGFurpgFgJSbGhhmkdkpyklJ39M
Z1iJ9biu0AALfXULe6+IGB1WlMK72D/RuGoY4tPMge4KzQPtiZeiDUswU6e2+31vZRVmjFsbphaP
KPDUINF762HLuV1XdJJfFKKn4W7HDBOC0dID1CBY2vXrQxCI36d6lsX8koIKoZVBie3+wBzd6WVN
q+4gSE70ZCvcCsGG6aY9+mvLBLzbvkKR9/2x6cDHI92gKrL/44aAJoqg8DPwOS0cuHdd4UTyQxcR
XrH/8pgDHE0ds/zxUOjwrMuuicrGYzSZ0W0t6vIQFNly27ITcc8nQJbtabxrVMcTq5754VAsqVR4
ARurYnzD6b6MXj8plw85lYy03Q0vGuLHEBsipEhAbIFrW1WHEie7ROAOaPVUIHkWEKfx1KYsz7sg
5RgkHM0cALrJJg9kjEh9VEQ/FalKXBjfKlZRtsbOj65QUswkrzMUUkg3EvjQUm6bh35nS+mtd3Yp
LzySyEY5Z74h90coA8aTapiDlnKncCAItU1XUc/E7nPuDRj0FnzzaVPYjZwqQ7WT7EZFvg67ulxK
ctbLqdwxF2E91DN4Ds0A0GwqwgB1ENFU2irccEFOoqnNMVeRBCZHqx0VkvhC8f8wighVHcmzdEuZ
35mcJPbxRdUIb9MPXxbks1jW1HuLeLYtTU/V6pBAOQHATFJXmSTQ0xeE2xLgfelf89Zm9fq500lB
sW71CBJxX0Yt1GUJGhQy6rg8SOerK9uHpd1vF9HDZE+hTq4L/t+xt2KKj74vUmbfxvsk/7tUWWry
/zeX2X7sRP7wJfKX9NQ8pipq/T+w9XGO77MYhL6S1sr12SD74Eon9qAVWR7q0Z3kLFn49dtHKmuD
F8f9zEmc9AbvfOrEcEiVy350/ICUUjFVcoD6V0DtrCzDOAHpbNtigxU6QUQwVkwyFpLd1apJozpt
hu5BZ4K6SgslZgY65qzxKpxUdH1g1b7TVbRLxdr5XL2JvUDXojhvdML4bNYoTCoCljhMRuF8tAKS
+MHBxeJVuDoYrW0cHfZwYmMnKkprZHqOoxFg6gEEEPqmEJxmjAzAto39BdCg+qv4RTB3258hp3L1
O/vc2dZ++karHaDXHPSIep4aTqrYs29BwxI8IzBZSKhQQFQtftI65DfIzrPs4QdQquBNYAuNyn7m
7IUukVg822AqAki/e3RxgGaHaBbDpXjKglFeG4jKr6OU4A6PStc9L3zvgBWP4FIY2ubRnCAPvzpM
DaGx5I/R+vB/DAXWx61RZLqw3HvV6D8Bluxr/GTflZW6mfIESaP6Ca3j15KVnr0ZGok2CTDCvAps
ioAVd4mUrNV61a74oGZwfuDOoe8GHBtHbnGAhSBUiVXyRKD+3sVtoASbembU5B58lU2HqUHpnEP6
akMeV5Od0ei3mrnmpVqyt2Z9ZiPYE7XL6R3hfHBxBHXAYF5vBVG7MviAPUhvvjDLeGLxonEEFk3G
P0lnPYny2bV8X1i9j8leIeG1dX1cJwAb2QHUEaqRJynWuO2AdJ0yv1tCHIhtJaTycA7zTdRGaZIq
BOwd6nMFUsA9yBq0J9eusOdBK7veKpzD9HGBpB9SOaO2UgI3dwgVl8B6xM9uQADAeVDNaJ+4oXk1
g1Ja18G/AhLjQOV6PLAmu72eL0UR/npOP3aZbHvKdWkYAK0TlS8c1aBVU4LsUlpN3fk2H8KSFeyj
wPgLX/LewYh6lIUH0bPPmkZLh+lMEYMsg0B6ckTg0OijkYyFvfmlJTHst7XItkb6olqoQT/aKXpj
Kx3/2htFAKnRZhxfErChCX1XFPA7X4x6qB9c6IFppc76aLWFVgPwzmKid/56v3kJJN0ewjZnzlan
qDlIIO+beRuM2d7seqd78S43y3lGzdjclVx2do3xi1/u4WGn7tnoZUs0Oud4PveyoENRwhtv+nkI
dTxuWicQWGMWUirGTVmKzcoAdkFGAOLoXFzNoeHIpNkn2Y9ou+TCz1xPQWEIQ6xRp2aiG1kNucfo
dG1+i3ueLA7GBTkxwcoTWD0lTa/s87I2Qx2CSZBHbi3xURqkKPX2yZ6elnJiavSeI88+jLdT5F3m
4Jj7o1hdIq5/4cvfV06Z+kuw8OdVggHMqZNaGuiQtXtQFVy8F8gPO+q+LB4xzYzKRSia14ZEKHga
zfoDyYv9vBI9cOqq7c7o9BXYgovvKnkrbngx2qlAeHRC6fzxHSCQhYFzR7EMgPfjlu3Ss1WpDZ7r
/MqpT+NvHcnE0iX9qnvHmRJS1jrJlHNKRGbJQZ586N5p1F7WiW9CeFIIghItP0TSFNHoDUfszuq+
r03M117VG0VN32LMB6sFdov8o55TJchPAdYdXhrH/rSKex3roa0GBy6zdk1M/JrR8FXsIhLdwNN9
LrtyNTH2BglCaia45fGkTk1DbPrLK2ORVAFUXNhr2oGH2TvbCkDI7fKDu0fTIR6xoFAeWOaJ3z3w
FzYfn2sCsUtc6znA/RRm2mFiGzjM5hSXl/meNPEZGZ02ieDWa7DdWNlY3nJY5w8T/0z1wydwPQu5
EvmqldMcGRlgadKpizgbq1w1UsjMBB+3yw0tJr2Gmw+qT4mHDl4JXR67aOCMoCGYWq0AvOF8ZV/p
2116t+7fE2O5RqaX5/0iuoa+zHH204m0W9/5ZmkKfC4rUXnxcrsMMRhkkrZaQ3r1ku2p4OCmahSH
TYol08stcmYKklTUWx308V7kQXP/OJ11/LGLWrMsJ/wfjezcSwJ8dtrss9wq8vzZKfs6JId9VmRz
FPNL2YmXpAQIgIDOcdzwyYO2ShTsfbuA7bjgAufrCwlef7EFWka1cgUn5qMex6CmrP35GNzDrrlz
/S25Ld9e6wMg+TDZZB4j7z7iplnLADn11Jk7D48wWfUT4cdNeBifcTiQTTjPx0nJ5wZYFGRHaXA3
3eDbqXdYltQr6hXFaoyCWDpg4JH4hspnzoKxTfFoos8/gVIBOmA8cb2tVOpLJap55aC8fUkcuQwx
pmVHj4+dVaQNieYQMO4aHgX0cR7JyJDKm8JrNMI9wi40gjMqeJZh4/YKHoxDOKB2kezTup2G/2UI
1GCjqhrNRSURUd2AUAQsFOuLntm9Oy+KxRSkLbEx2SDGvZbflBXVqznTE+LWKNDV/mVIqimHI2p4
OoyoubJWylLQdEBIj3xEXbuFX8TR8dovAb4l6AuDPUcKLDXvJ2Z95RJZcpgwV7WvukiZufcP8HNv
+lUvx1gE2jM4dmGZ1FD7ny0cRr35eY/sXgmdkRbZP3mYoLCkJjecSzGkz0eBiDZVdXXC6eDlZZ2S
Q3hJPi5ALDfG3pj6VbBQB97S0Si3JDRFGIc83q7CXRAtnEDOvI0eb+0kIkVJ2ttcBEvNxxFg2F1V
noVk4A19aTnNOrP0ABfgFVTQ8VarN83v8rTVJwpEb/NdTSKBOopfR0EdC8w8QvuSWKv9edUuwZtt
XT8PoRN7BdoVE+l8/iPikZB+GhbvY9EOMHiQDuJqaFMN71zmbyVRNz4/gWh3m/i8YzOR+fHyrEN6
i1ahUaoftnwCegIfnKJczFKHXLprlcVzfPf97tulpNHQ5J6fkA+GMXUWX/pW05DpxsGqpYVXpgHm
/0mgVntBEmN6iEydFMEaU+bIvtYo0w2Y5se9TldtVbzz2Zbmo+r8nUvELLdlpQAi247Yrpofltfk
IkTt4kEECYAwTkmV/d3ljngjuq3VSq4KK9oX9ZBZgU9FjNxye2kDVJqdziBDUA4jiSGBjQvfKKpJ
6tK1Iy5sKzLMwKYLuJmqrJNN268wlxxkLsZA03AQqitZf3DQ5bTLXiBrGQwsLV4ixPjJgzp5yIN3
k1P8X5dfl48f1lT6AAsgKUYoAmagYcYYzbN0tSUWSNgCVaC26madTzGZirud/aRY5F1rMH+KQBHm
mL3ohRwT+wJE5H2z96Ad6JbHoFd6f8k3Zx7mh1KQ42+IVAvgeKu0bfWqYbnHwAswBa8xZHSBP02F
eYno9V3fA68h1JtSI9XbJDb70rOA2dVCgFKL9jNZk5QkXDfC6gCYc7ZhnQ4tbseZWa0LyTYnT+xi
gsn2QEweaALMc60EQ01ixYJZLi0MS7XaqHHcNvjHCzqbe3nh5tQCNWhf27676Drde0tX88NJuBMi
C6dGpzulj9HxeAdlwpzMaSPEu/q8ftj31QcAznIXX4ftBz1fbemmtDqON5q7GYORFp+oMzGXwOnz
QvTYNakcA9p3uzewrkMVTjqWNUYRfSkJMgnQmnLTaUkQMPdmbz/JLwFcACBZxZsCZfJyILREh9lw
QHV5xX6fwdPiaKQiOuukxiqlUXWVBjAZ8gdiiJ0W6HrU0nFkh581ReofDzZ+YoK26LyygNMfAmeW
PBKiT0Db9YGnOeOTdzVK2MQVi+FhN7Af7Hvp/jdQI46+YW3Zuw0saOzTxgs0kQqeoWNZIKEi8hcn
DMJmDHwFGwA+lO27K2JPPySYASmkr+nIrwcB53HmNgkKV9GhbF7u2FKrcnYcYJN4X9ovV5aQbMtX
o4QYnC1EV1fk1Q3DUyqYbuWv2SlInMfQ5CzVwP03mUV1ZeQ++ilVbZZkwf34APOUMQsdVU/DoEi2
e812kplJjBr16mspndjD2TlhYHBxwhn5t+o8v1iXS6/LZ+/6oxcPXBKEPGtE1gAjxJ38ZunzJX86
wHJ/LPhOgi0fHQyB0BL48pJNNv3w3xaKWVdsHNevyXV0kVU42me+igBRMNOhZthy96w4Ng0xEa/P
X5rASzsqy+jYgbOZxKlpTSBPPJUTynBBP23WZa6lHCXoZfivbLyzbNVQnIQfcXAcTqpZWmV94rkO
/yq5S05vNynVWDWYdQOuoZsR/okVPSCjTnnGgHcAZuEzoZnAPKWxNc3i9XqHlKwN89Hw7qIYDkrs
+cOR1u6KJFYGJqJEQE6hhCGGGW2RAA4dAFPl68Gdmnyxx8iVGDw/KQYSc7wdWlTtqK7OIHkcmprB
rwd1YF8eRSztWPIFgHI7w83hWMWPXP0EU0dNA8yYH5IUyvsdDlJOTyJ0OssY03OXzXDAUYxtWb8s
2sDwGjklI+ng6cVeMfi9vEeYHu/TL4FMUmdP76wcM1jPHkqJEMl5XAjU6XOBKtYj0Gvf6NOvk+/b
29cBqEoxFyfDpsVkRONmzWk4Y+lQrs8dQ3r6i7yplHkSu0VpLEJyAawrJsRP6uo27FdO3rZ1BLbi
8gvEv+xcjeQ1GoOFp+T7LjeecosP5z4XdRC0ldEdGRk8tSvhEJ4v79HZo9cwm410FEyKwycwbA48
zAxAKbib6jIviqkEYSR1QvGu7+vAZPPP5wIw2If1GGKaHtiav1jf6RF6izmThIiyhJgZYyKMvP7Q
ImSIowX/PQMBbA3/3QjHF4ObIujSq9xOKxPMoTn+Veskkb2n7riuRw7SbD3JHYTnBtHBm6/AsxT3
A1RbzMgicx88axNhvDh6ogoXXerlOBCz11tViNJ/Fbrjs/ADvDWX8/5voNTuKJNd6pO+U8kVSyVP
LPdEZLj9T1IQag6BoPEF+lYios21PaTvnSlmGct6ruR9o8Bs+Hptlcu6XfypS2wHp2DLrHxSQrc7
O8cW1yGgRCf2bx0ubyeHCKJVlcPWrIDfjgTA9T6MQiVmF9jVBMgMn5dZvMyS/C47ULWV34TYrUP1
LqVvZF3WKNZkzS/P59LTJJrYv91bSaZcdXOpM1k7vIw8CqIHch8/xV0pw0PejgllO/rjD6YcGeUd
AJEzqOfuuQZczWUjI4Zv/5ef0D3Poa6I7MO+No7GvtCczf3CzqHQ1OznlazhW3UfYcSAHtsmd/Pi
mxevw4RzOLvfNxVhdxTo9a3PJciuwiWSVOAHkq5PgZ+VVdrfwFnQPx1mSulUf4Qh3CvGJf69qlvK
xBN47zzbvB6BrAIQkdUl6qPGzQ8x6rLgg3UgtdSNB2+sWvuNugviZlcG1cJ1Pg7OYjW4MRLyuwkX
2374hSm4xokEsIzJaXJ4G2iuc2P100QYFM/aEV9lunP7VlW+8xtfAMR/6s5D8U8jjdka/UXSE32n
JKaWuVTrZIWGiwoAP9tQehndWDxPYk6RIkro2e/SllQ/U3Zpi2Cgzxs+MWpAQWHr3rMv22bFBMi7
3G4u+rlZYigeTGzmOoZm7E6hkQwGDSrwkpzyISOZ1cUVmyO8uD1z7I0/WdqGCUPZS1u+E00hXxeQ
5ZTU07oV3wMsjgFxsG+RqQoBGKgctko49tlVK5mKrnfxgkrbPV8rKyoQogHwKrRfsIxKdKDgP6Ux
ipi92mPtKdKtyjbBqZuAO9gE+YPPe1M5PrOuJwryLemTJbKq7brSjU6BSZ8BAU8Qy4qUmsyFrhYv
AfGM6UadbMb7wbjJPl+JkkEIUToeU5cp/2jsMnCzGP/hph+hkIiJxf9RntCFqMVVZ9jipI92xuUq
1g40CdFm1V+OLXuXZLsJ6k8lg5UL/2miAk1iwyKta0kcc1PuB9EwqKdiqVeWFd9YaEc5aTIL62d2
3a6BKhP/7KmJ8nj1RibHNWP/hTWRR19/a74shtw3W5w6GNd9BLRuwJfnUnfHKXfeRvOIs3UIvAYT
JMfTS1b0AQHOx6Ttvb6IaoWE8f65hT8aeVcBefK5OW3y3tamVDmFIfsEFyT7O64Zxdxsc5Er2eBG
FvuYWVnEv7J6bOBNhKnUnZOx14ApxK1dTu0fdnWmGOQlNvB94TzR+APXU45amBcbNMtzeSK8S9QY
spSj/Z5M62D2VmL1MLFeP1xwdOP5sHBSzyvBdFJjj/whSvbMq86L31dViFeBx8/UAreKpUvq117w
qK6OL+H3TSKjy8PheVCElvBzm4xNNSMlNVHEEgsuJEGl70aS1hfqL5hLPUW8uOX5kNJATFeWRb++
0VTCUlcYk9LKBRRT/qoBh9kpUdBy6QMENvUUDgrSONkRX73UnFbCId/B8LL8cYPXawwdxeOVgWIP
MTfe/vNK9+uvAvlDIgUtEh/feF2aQewB+Qg5+Ih4iv0MljJPvFvwpunLQjlRtgJPMQUL1UueuHzT
+Jl5B0MkvKLZT3aQyBDfF0M7v97BPIuPswEZ8i2Z38aRxZsCLlKuosWddvGnLfhPusLbh3YO/QcB
4Zfiul2vl9vdzDgjSbs3s4H0mJZw7ZOLKe1nzB+AeoCi+Buch07BdY4DhO80qiLM1uC4t1oq/U+h
K5ePtmc469CD4uiKcVsrgxRfa8KbAZrJ4t6qMTqZSWI3WP4rxSDedXyvaFJDxfWVEARiyzq7d66V
wsOh319gUk5Die1OfIfV7apP3dV19uENVUmL/LcpbBHgInqjpLVy6InsntCXDC0cHaJRoZG8bZo5
BmlOsa3rZwNJ7gx4+Lie+OxjcdWWmQy9btKVbHDMsozC8JYSVcdb+XueG3qyvKeqwRx/fp7a0/li
Qn4fIobbtfiUujf2Bx7/2mi0zEI6/b0czsKGIKwv3nR/+qzzDBgQZtZFpinXwjCUIDkFcdMcyTbj
eZ5ke+HyKPogecP9Sn2RZ0b31m1nO6j3JvXwHxy/htGxNJky8quCPrHuS8B65k47BjlXkaOU0NjI
bOnjjHA+K2diX/99IAdTGrPxvLIEGESA2VAMmQX4byM8S2MH0kxP8JgPthcRnQu1207NRKmcoyos
JqNmIflHbyNgpyUN++WmIE3FWiOQZQfi9+oJ8xLJPN5lUtLaRMWk9zM004rsuHCfPFsWtSDyDGXu
bQAbECjAA1J5Sn0JCUYbSFryUhnAb0wGFv098iZD4ovzxRWzGgoU40b259gxS+8fovfCg1dbm9HS
LuzhL4nsBRdyahcKjJaj0Vht40ZAE4CD46a0khCZR1HycDYl/f1YJrgRN6uJY0vnrl6W4RpZ1FQU
URmgWN6Po762sd+f7FX2TjYWis4ZL7ILnibTM08q1R6QLPLsI6N/+hths4QO4DgAQQ4F4YV+p1LX
oDaIULKcYVOIEhf6eVgq7AZNERpRUEq6NhRCrnQSZ3Fa4a8KqbuvLgg4Hh+DSCi16vzRRiNRaZXP
ER1OBQOL4zPPGd6F/M2zrXdgeJG8haCnLFELvm520qL5Jw3FQJdY1pjs43tAmM7ntPH3ce+PqEMu
q+N1noBq0Ou3W40GxpTjFE4l7RAzA3CLIxchhdNA7cwITmHs0PU3ziCYN+qNzpHpmct/OWxDS5sB
JqVbpWyR4RkhMQaICgxy9sYykKzCoyqu1nTNN9dYy9iOaTkddHq5xhLE7yTdh5gCzYpKa5GVcWoy
1E2SQjzZRv77xbgRKu6sAm33tqlrVMNham8evUgwxNZssroSuFFgVHBFamxdwMNCakvmTxhFseA6
Gl8YVFdOgYRlYgl5XIMf/q/keIfeVmdB4hKETl/2qpmBH2B+DlkUxDyy5PJ1IHiGEOFcCM+86Z/p
WzlpMRErOrtd+mU8SZQXsWCALbuDIBqeeexCB0iGfJaJXEvrTcKeWLn9vhaZLrpxybUAuU/rrGQS
abOXFNDbbAbnwRch9MJ+tx6tLNd4Gvhcj0AdfgRlIm1heLS6B30GRu7rP2QkaUAqTtOP+odghqQp
DMTHwVY+DlmCKwVcsSB93sxz4KU4sFtXoacCqHSIrNpiZ37hFkbZuMix7ExFweaPg03+a2YGmnSn
4m6d2iu3tzRkxZUd4Z4OSqoFXimWB9rgssruJEQ2thTtxUkoSiVLXFsHm5Al8gesevbkwJ9YqPUJ
mdv/PWYCs51RLmzvSgJxEtojxYpAnfqtEFdrJM6xPpZ3YWA7BwwJaKGpsu+MUCbcYOO/j66SMi3q
vHTVQfM5cqGC77L8NDlzY3/exPjEXvrlTzVP7OXDYH5IovmyDwBg+0KfYKgY2YYnZKopvjuiJhX4
DSnstYtjNsuF6aSnJxVlxOK8QnG2z5P0pqRbKNnhLbcyc9UCYCKj50vcEQNXlMTFedEQgHaT1SB7
SWbBse8CE6y0GGxCaQNwSIMLDG/IFMhhslDjgH1UsAgOgTASAlkvzMv86FrtzoJ9kjqdli9u2Ttn
4Xqew623OkhphMTkWFsTcXd5aAT/uEc0hGsphcLUWkcWpUJQ2oaN6esGH6tVeDaxII5J57McoHQ9
qjMn6r00l0B0Eii9phsDS4O6DeM9tTI1jD0SLsP8rdqH9dNYxWho3KZZBaRJOjj8/kSUwoBhLA8P
hfDTTLRjgbEkw7dSEtGe8Yqb7ELU+vv+Hoyy+zAZOMZf8DQ1Umk5SIaGkLs5S2h5RorKpvOIuhQs
Ao7ePmlUtniExvNyXXtTiDTSK72+Mf5GfZCeA3dkTcBaYkDiqe5CfZrnbRm/cAvcrOfeenX10Q4R
ICvrzLzaaXM9mm+Eane/768yPn7a6QtQWheNNvgJBuIcuFiOpA0k+BEK7pVaLHk3ANlDbkmlNmjp
mkpzmnvj2/gs8Ad/VRF+gyEvgJFgVoc1//a8HOEwdA+NLpoPc9IGdn1iZ8tbPfyPzmiE9WoAo1gX
WpTWhGeJfwFywDZdAGtBOj16b8gb4s5/xo2w2vKnc1t8jjnoyFIdUREZcVN5UfYr7rwzUufytNGM
67YCFOKjIHkV8Kpr/JfYrZZewyYRZ6uaYFMlDd9pUXk5GkwDILTwWKq3Mk6xnNkNX6W3RYRuQcAa
Dx+zXk6df4OXY640VdnXqFgK41qWTjZs5OP+3K2exMavkm3VcjRQp3AUTdIz4N34RTiPIcdJOOpF
j2gI5ETpc5CVpAAJIcw9jQcknvT+nuTJQMp70o0kGWI+04kg2jYUGp7LWYjoqk4yWCcHX2WV1tri
zk4m6wTEMEk3yy13o4SWEh/HkGaUUgYhlLwU8pWVGlDKwIABSE4merXjVXmZLpORUiU/jBpCuYuq
ImRUKdxEoXq/s0q2CJBcxaBW8omeUJraVelYv7Jf6idmk0l4HRX6VyVjyMEx//znPJD/P0bS1E5i
alP2EmwRiHGux7qnfTWvzSiSxIV0/UBCDPjNWK7HWg6nsTISoDdBl88NLxVwlYSR71SdiifUJ9vy
F1Be3BHiFRsxNH9iX0dN1KMzcimmPPpYqdo/E0aIByPg6dljCwEmCtjoA91FTlzv/yA78yW/W8N4
0+V2wFZTgkVJrY2YDTnK9I3kkb+qYGymXvprfepzKEoJXZzYN4WufWP+wscSEYm3PxUhT4dzczLD
ExyNVn24eLIVYAaKhLlXTYtMizcG71JiYT/q9+ZAvwebHAmGRa5lFzsW1Ea6TeCGqi/0yb1LxcdU
oGKSDGDUzn25QZIrPeAJJErrALMHP1ubC49wwgokOG0LETUyulygkzpC/kl9GyGJA1l2dBUHCcVY
f/BknakIF+JYfn9H47a1y15xPpwvFpJFV/JjPKEt92rpyfdSG22qkbATNyZihRmFBdiNzrZIdbRn
nG2rz2ijwqrHp78EsWrVrXMnEycXVDVoxzUXKZYLu+ePSc8fJRwXdtjUbGfLdb8YmBMC5ge5QYwi
Xrb5lyIUUPrpDoci8Fvkh0uhat+0A4JI+dZwtOvzFFO6JO6LMFmt8UP233slnqJEAHsxW/j2bJ/A
EQkkX89YeWSx/XTbA8rxRfLXkzopktyMJobWpHp1OtkfErSQALKwRcD+Eyfd/QgFl3YE9C4UBjvP
vEmHFE/V21/ym6mtiMwU41YVRO+PFdlwoQ4HQ2NrB5XYDqhREuUGuUCFK2BRsLxsE5tlyZ923Rtj
wuH61000K5+f79+DXbgfSFOenw3xKFBflcWTo+klKoGQFKmddexPGw+HWgbzHhi6lLeBnhG3+3aP
jQN6HdAjON9f7fXPGTd2CCU70w7q9m9fbULk56J0ShAbxQPebjl+RlFMEmI/JEaWAVFW9uB3e+Ad
TRoyinfu0+SGU4r+ra2qE4thIvlOtJktlCOHTyaC2SyFtT/nqCao8/MhEMqKoMpflwjyuA07HjES
agwZjif6BUpjKqhmNGYB0seoPTXLj0++ZU/oIdc+4WYPhdgEIxsUfQAyBfuV8tvwCmHdq1K1C7fq
bjrTy5v2isr+9NG1jyaucxS8A1zux+vv0y0hpDKUxFMOtTf6KHi9kQOUABwv/MCAJ4emyXuePzmk
deBosRkHlKuu2zzTNNKovFgqUA8xtOV75rPgwtZmSvviHIb9nA37FxoexaJ/dpIX/ynzY7sd5tW+
lpCnRelmIEwKzNpVsw0BBOieguINVhPgxLs0JHhMbBklFbbNDcPyxIPBhSvUkZvbTXyFE/PvMsSP
NXYE3tVuLkpEJmM990sCUdR0dH1o23eYNr6/TQjTTRp0qAYR04uPkrZQjUlN+GLh0aFCugQNdh+p
UBSUD3o1jt5hiVFgZZU6QauBc2XZ8Wyn7KvBQG3JXnL8wgpmSTAETKBSOOc+9gXEPm2oET6JEaed
Waoin5wnMDiXRPUV3kJ8cUYHKbAZWENvPSHKp3ble4cViv2Bpz2gWt6InQ71/Nzwy1l3x5rSu5of
mANjqxgoKNWdYib/0YFQFhrileDRM6ZdoGSlhAoibguYQlecGOVsIQz7oAdtyYYq6LTkv4OcOsPJ
r9GFErKZUyEtVru0CRo0zjAEXlTzMwIF7oghei1kS+8tOAsGLv4jHAY/tqJ2qzRpaqEhUTEQyKmy
3AAa4UCckn9UTSJVzKU8b2Hj2Zl6Gm71TUGSApJsb2xGx2l1sEcVrOYl2DRN2lrdWIXGF5tkDrux
h/YTFMT67HXA2LKYbZH2UAo4ZSLWnRaZP9yBcmSmSIXNkNnyyVUDiLlzxMS1yzDbQhmiseqVlRNa
qR1bocktdrIGvMzpZiwujma49u/DLNOsocquxLfDxKQ/A+8krEzFZ39Ti0vDRuUbTawSRsjJVrup
/Hw5QoxltSwR6wuQ0tLZB8gZedRDeKUfXczdHcnY2p/Dhn7Jr1Qm8mhE4A0bmqpLkP1C7X1S6rHF
BBJdTS/HLSv9HtDi5Krxn1e+Y8kEOGgl94TyUfBgiZdfM3VzFldleyu5ivcAbAnxThVTXuLQHlHq
pk4/FaGXrdxHVWR/yohufdGmonFjz+eumfiGxu1Uk3wXP13y9yCVJhiVluX6npI8v7zPYG5zt9fB
l06kROok676DIpZYu8xb6eKAP2WA3kEqMYLo1WmfwwLDTIsAiPXyPjSXCADcUD20QBZ1JC04+1QC
Dl7xPxD2C7QPBiNIr25bKCwI2nqH6ZSqQ+FMksH/AFaUZxEg8vGvf2RR4qo6tHuIJoQwFCoxcNRY
m7gmG0M+wJKS0g0pVA5x4XQe9C8YSdRdru2twyjyjQO7ba0UpxuxkfNTpRam+oK5xYlq3B7KaBV4
kH9idL0y+EBW2RzTeenBvsTcrrht9Ia4aVb7eV3q3AK0QdWpK5/zKyKVgmGl+J1yr1g7YBGJdfse
jfmLMOevXdBPAPBoRnMJctcL6hBA9VjGzTDI4y3C49fo1r5wJiyBq9jhPgcagzvZJzKm6CXbjyQ/
xBlRpU8RDRE2NejLmdwVdK2qPGnxQGfTiNCBV6Yi46EAJJJgsJt08g2wwrrNmNIUiV22sNEPxmPp
FDhDSUo+qfeeiTnzxYSG/C9loDixfscODJU36MTIv/eHrjV83gREkrNEl0OcB1sH5VuZNu8p8TBN
AguzLl/EHjTmEJm37Wg3O8cTGqg5/qjWmdVrlrW6i5vFc7FEHroIbO270vVU6fdzJy2HCq7thfwn
qqOuIIcpQ8kKngAzKe/4LdeuF6MmXqLdLX2VQ3v2SxoL2cL5lYd4ZSq3IEgsHoksHOTGqbA326JX
EGf53C907jKxGJnM9K8/zifVIE9N1G6dAtzPFYj3uvbIdgnY3148uR94BatQiFMKnwHpHUJVXQmE
dd+QwepbSQPRRkA1VCsb60lWGvlht/LMM9RxdmGY6NA8p8ROqmh9K4EpL//ouYKa+h78RiaeL0Td
hgyrK0EvUNiPweyM8EiBQLUJBnj1nfaMadQJZFQhTW+UvRh1ktrH7yIzoYLK3062UwRL1h+n6K2g
DI86tSC8kCHexgxq3Eid9sH0XMeynAtNwt9kf2/VWKZl1U/aSQqJ6uen34gnxFAYkz6etjBw5Aj4
rwd78mUTUehZxC1inCRirlvHmAzPgocOctO83rjIrQW0Vrzyz0FN30AvugrTru85SNxO8ldFiQv4
dUl/iwWAV1gQoc7iK6hutRZyUdxAfCvxaIyvoRbWRowfMVT0E3uV1yd8DGfc/R/eIjPljUm4CpnU
co/sq7uLuBnmMUICLZPXPzR+eRcebPacLlru9n/pTJ5JAryq6GKQ3qh8wQKzQGOngCs1BlStHcab
CGnSA7fjlprmjZIpEYtqGFqy+69ho/MV+9Z6eg7J8Po986RiG9+0qc+JiQzmNndQSvPw6s4PC1Px
jN8YhWVVH8H6d4eArlIeQDCtWFJTLZ+XqFVY2PVph3G9TiEz4opchhAZH3Z3Gl8QzReZcHIT5OLA
zb9OC2R/vWjFsMGDYtuk6zgKOFQ07/dqmqAdTfJ4Fwc8+bHcVCSipacP6FoVHs6q5Eme4snHgJyq
o5IzqcjslofLwjqDnpaZFQH9zvtfAPP+TeOU3JAKfqAEyYl2/crPH9b636QAqNdtUtmKqrGo2Fv8
7aO+OcJkjGncShtUK68sytaasefd2OXtma3Zi7VsH15XINioMDoDODF/YSiwa7bhzJJr0BypiJwY
KY1Wu7H2w70hYK3BM1yhXpZNTfQgrr3dGUDrZQFXBnTBhhZoenEElvjT4IpktIDqEh1R2R4vTwV+
+Z5xyRgbUA3jHcFZxnt3lKM+6NjR4ZT1gef19IS+mZ+J3b+eseh/2qQ0DZwcVtSWLajBKcmbaFaD
9slkT/ut8oZ68I/HYL8vx7n3c+7N8pywVsYacEGv4vsdjbl7ySN3ei2Ow1TGy9QE7yF4/IeuKdy9
JO0olzNpvrbMJ7XTAnD2/IsHu/kN3U5AK3Y7zzy3ioUDffg4fW237w3PmLPPowWSxE609+Stewvk
kj2XvYUTrTm44tpGwpxlHieiJJTKuj6EYursCZOBqy+YyxUqgv8TbLXRv+Qvdc4NDx93ELJ1cOvc
WftvNYH3DpYdW79IsUj0oPY0Ep0GxfAALOQZp2ULSdXGRfrTfGaQ72B/XiGsS9zifXdM0RkR91R1
DSrTqeGm1bF75LJJmWoK7KLeP+O4pZlg1dYuA7qMxIv55vnD65qGAnyIABgyokp7LlRnBlaTRd8m
E3NipzP6NbGTAN0e8vc96dn3xGJV6lz5eGlMWf+V8PJ9ZMlWt40aCGq7dJ7uaiQjd3g1W8fKSDuc
dLF2qL/gh6fC/sBnco9a4USP/gMTndhbfXq/DDHsyLlKKjHrhJS351Fv8IZw6lNYbzg/1W6yNtYr
yzB3NyW0JvZaTJ5H3iHModAh+G8pG7VVIlF+4kJRSsevI+wBolReWz8H+9phz/YULJShfic3fkEM
L8i8p9wdN6jyw/18OI6opCiY5NRXXilNDzRYnmDptRlN4wGDcl3ZWG0UXd6RnixgfOikJ6tlQU0Q
/s4y1LpahYlUoPE8XCgadrfnzVia/M/dAc5Wdk3wBpj471pVpAT12M55WvbLp3inAyXodTMtgudb
CwdpXUWkxgKEa0hM1eq8lRoDVRPk6RLIjnKjtOOgTrgX1S5kcg6O4fwMExxplgEeBD+cDe7i2Sgf
A92Z5fjUm7Jl4fedw+2JpL0hZQx7D94iNDFtLIXtShAoJcxkZyB5c2kQDdFDpCDolO5yD0O4CLOy
wyIV7JNzOJdDcI9hw3qVx+nYwDxJv8D1wTLktU3PGjPX5sTK4HL4k463/KAYQt9B5oAaI0GQVkLn
axhBYh/ak3g5OE/hkVnJuc0k8hAsvnAjBWDeX9GPmPJWVOz/SJNzUZJQV8vG+rTlbl8ibdgNHr8h
+B2j+rX7tf+D5/P+ECDRcixWSUtnCQl0xQmkBNXWWm6rsNfPvQZylqtVviOkpwN5Bb+7WvTYlOyP
FB5MMf/cX6ZkobpP2g7itw8drgiEZzoRNq6+tpjAAICbAn2tBhs/Q8JgRKxNDNgMONlQrQvT31tq
9FKpo4Z1xA9f9aoEhjsxQOaV1Ou6+rVwzjZY0GNgBiuZBh5/i+NJeKm8ae7DhN4448qZjOCJJXbi
SFcg+ru5gixvTJkNbzYg8Zsw5vbLxkVacTkpNRU/h9qF9a2MRg0XKvnSKZ64fw1LCJ4upRqJbXmg
El+tIVFo1Y90gE28qquCEyBDjpcLqcUccHBsItzgAHThvNaUWzG9XZwWICo+5I6jbZ9UB/iZnWg/
5NIGlfAqE+JMJsTmuxJKGjk0V6VJvUuS40sb79rQ+6XvGNSBvlSaA0Mh7AQU4OynbJ40MOsy/Tox
/X/KhYPih2IFxMy2sG7tPnzaI9i9A1OqTw82y2TNapyaqUpQRSZRCPa6MEg7JT1gjJAEcv1q49yT
GhaICmP/HyUWCA4unm9yYo95DH5qKP3xuKDDbykXhTRkRkV6Ftdrl/YKYeAK4LHSRvnCqRfUxhOk
2Ooq07utfHbdUmL0PC3RxMWusS/JGVGFL7Go9b83d6ZDpsZ12PCg5oxUSb/nKfWEHCo49iZjBVD2
6Fe1ljDxrlFCasB6OVUW1jcWjfCUsclKuCkcIU2QYpuuq+2mZwbwsFGu8l0dtUxSTAJxLByhxdnT
y7s+jJN0fUFTARECrawuAwvJWrzyxQXmJWPo0C494UVX3BS0qj0sEf+VQArOozmI2d7QDiLxE4Ux
ZN+EDw55Ixt2c0DTgR9mLVfJJpqjcTQkAjgRpOJMEYgNFWIz5BbZakCVJ8p5ngHraWhWVMb0mjWC
UdJHGr2hcIYIb50UNbELueI8dHk8kbd4yJgS5+yB8LAB5nYmA9FP7/qOtXSZy5jQPUV9jKLsgtki
JyONqIvm34iXPerznKWYPZUWoB/dmP7iP3i8TWY3mxX6fReQ72WkQ1lZtQW0gvzjUb+sbxb4DPAw
6SYzuZWB462kI/ABlLcdY+RpsZphG2G+s5dfMjq7X9KxUyXkRfpssWVykmx8b7BGSjX/OXUGwcaU
CfpRPqqAFhrUXNCQvBNxKkzl2WxztfODW3i9XzXY5XIgyUTioyco/vPP0VBTtJeRJ1KEpRgRVhq7
yVIzzE+Nwrr8AINx6k2j1Pc4UGuuBnpVsItnGntETmHl/+QWHLRUENkUtthA2RQYlZB0yyrvkOMV
LBaTFnrfnedfFdMu0JxsaB/Wlkk3f0mQ3QlDByKjCUA4LJvle9ays1lqWe1+r3cneHrsez/aka1e
Pr5uzSlgaiVK8Vn80RrWce89gUd5/XQtESch7u0vTNr9tdKgbSCxCkdqtKstyKGJ4721YJBDghhR
Gr2OuAZCV3bsoZ4fvSANTVbTMfq13HLlj0zqWYkKpMXDFr7fCIySAib1Jvtgsjjx78LIVOrrPXzS
BJfvN+TSh6653v94hNDkiA9UDwlfsQtJcfF6oZyhEZAea2Fu3rX4OhSXsO8zDZloC2hwBx6OprBz
Wgi2Vp8RdqzTkAtUqTaWf8xEOEuiSSWGq1yg3vLgf22nbN9/qrv+Ps1Lxqqq4yArp901s2UXEQ35
iM37xn4eX6bsDvt5+5zKTEwUPYIcpOhyb5nm/qif7R9LKtO1YwGUAEqhditoAQdqH4ojxfEc+OXA
xNpp/8s/a1cIRtJLKLldItPWuu9JB5BUBbuRTZcOMxva4Zo5ewPLNtyoYP9zwAwVI/qYAvIg49Vo
zEbyr/hr+NI9Kk/VJvzEzQTZyfQXM/CF9KrxOcMnV6AEVb56jPgUW5koJ6Hk+EK0yHJD6Y/JDhEs
b27+DTpXptvdkMYSj993uF2nO1eV9GKZtrGCevgx+B9b7ktid7VRlWN1KvxSHO7XTinbzXPdiuD6
4gHTE7bljF32+rIy5MyTi53lp671gkL2ILwX2U5yL6fCBH8UB34x+BraNEZl6TiosVjjNwJPT4FW
N7KBccRxXEur1mHyPM61bavU9vyRDoG1w194CxcboMPdMZAng2YMtGchHskXH8qEqTD6GmkzhAwX
+BCFSiXkHqzj8J/rRFHRoJVMQ71siDW9HwE67Z1fWVKBBswqcDUOds3hhUjaUBbe8TYD6EXnzxzn
CUJGd+CQw9g0WL2tZ4yJI9rULgvA7offOFasFrD0oxJJEf6T4itqBJS0HostWk24ZRaeW2c1+r0P
euZpuAi488/8dEU9T99jfeMynEw3+UW5wG7m8NOkp64AKKjeTHOHc35FcR3BmcScbkvLL5calDoZ
7aC7gU7pSr+5nHLvoPF0YjaY2vegVzAl3UmKvyvhnjL/IZot4bpGDL+x8/c8z5INyOvAIQIlVgWc
Oi4FcKaaJnkRXKTcpgpa8yvJyi5LGQGfRxf96n0ulo0yTie2Vpd5WpS92WLZhhZPXORAQ7vquhnf
DVuVfJEXPVtUorhKu3qvwFmeTDswjYNaGaHQLLCuO4i0e9sxgyDsUYI+UDT6zr52JM6C5HyzIh3B
nU/mLO4ARQ6igfPOs4wJgFgraLVghB54EXno97zoiF55cgzH/QkKLqgum5jAsqfoT9dU0wYscj8e
zBRR4uv3kBxakKHhoeY1N1QWMk1PJZdAY082YM4wBWdilmFvyfYRYkjo4IPJ2r5wIOh1/4SpYFfv
OyDHYS2dlQLFuA+q0z4aOmNzJQLK/q4KB24MJvEOhaypBWJRUmV9chR9HthX2LHIF7pppLRUy+rF
8KzGXq3W0KshMFdrKqGAkNt/E7Q1oVq9NihAaqjzDHEeuR5uh+5vXxwm/rCgSyP/QOfswCiSpJp5
Ng5DLORTa9ThwHuEXLYyGDHqLyOS+KN9BpyZFUU14X3XPB+OPE84tsWqxEbABydhjTfyO+/Oaf3S
qJTiRk4a322oVfdgJ0BFQgMC+jYI7AXT2Z9LF1fsKEXNtFYyX88Q3etixvusKJlf1SMxBluTo6hh
t0J9qm2Fu9cW0lbxgY4LbkGWGlgUc18d1a4S1a6ykWBrX2B39L+3hLx8Dm38B9Z+J/V6v8rv+Tuq
gBjmbk+LT59OfW/8mhJnBErrqxMRp+liKaA6T+1JYgUkLh21VY3EEBvQe74rczyCSeIDpbNHGZtY
wDSU+hkG8c7Vt9z1jhQPm6HVQctHh9mbD+ifefvmYWj0a/Uic4str8aNKXWVZQFmptIcpgCIF71m
zr55RJg7oZQMp+LRUi9ufoqNn2yg0MpSb5yLGR/ectQievLt2wzog2+XUErdTn/UlAuderyp43jz
d92Zt8AW1KXwV3UI0B3/ENfp7HhyDL+us63jAkbawFA7Y4SMY3KyKaH5UhZbHY7FTNIVb5Ai82+o
ZE8lKykuMiythrxD7IgZUQC3SZwGLW2Z8Emz8OhAbssr1//3XHQDx65sqPOPvF/kVNx+dj7bLo4E
/uBu4Oowp/oJ71IDQrEUpH58pqImaYocbriuLDATpXLA52DRc7Irahun3UhC8tOSmg5RIOuLv2vx
KcUBLLeuPeiH57ySFifjWMpn0Q4KRooMzwtBLXlyX0J3oDojQZNcSrwSc3/QSaBZvt7E+ktkVTwp
P4KsjsGySwxFBkLqU9K/VYoYNITyddd3dT0Ypjr21l36lgCokQdzzetebhqZIekpGl/gE7apLHFj
EmW/LBpr8S9CTtL2gv0/dV66fGGqy5LpHK8Fr2e0BTtuYPGhyacF7lK5CqE5pIkP3Z16Fwol31i9
gDKnoqhZn4OYZ8WajhkdhKNZsBnjDQJfxM/BmEpLHtOq99F8fI1aPCxbqphAXlGh4ltOqMGmGQiy
IO+kMjSJY6EGBZ8LzcxnOZ4XRxLdmW2CD0aZb7SoHyxswso7uGh7JWhq4CVqaHYy9ErOAHzElxbD
213Y0kmP/PBZE0W/wwAh7lOy7SIbBHpWfdaXJMGtxkYxFBeaPGnHn54sfgchHCHvBU1BZpVPnA6c
0Sw4enCT9vnf4unbXA0cN2NGbUi8xHXoTsmDrRrdUcJsi66GDpT1z4kziKagyXR1PfOK/zc4B/A3
DzRnwY7+RO3RqJVgV1NTKCG30ccTkvYwZlj9vf+/yjQcr4jZGP2iGsz98sUJ+r0x72YVdrURF6A2
MuffW5Ajh35N1PbTaFRC2xVTt3BJLMVQdx8F50NNK91mJJ2aznqBSPEh5eZjUoMUCl++DPkisYaz
LHq05qUIkDNPIiWCm1ByDvubLFW90H2+TuTRi6cwNMZQi+NiRBbwhIo4/1z2w9HPLgkabFLSAsV2
qnt1jvrTuzpEeNOk9FNP93ilLSyCtS58sUX9R82mjyflLd5L54Ji78xRWeRh+8Jn0XStMswaLbgw
TMP7btfa4fOYfvPfFZl6QnGgPNhpD70VyP9RjXN4AoFmSpz6zpvpEG+Nb/u4KCVW7v9sNyF31v/B
n+bj2IDMwRf1Q625OSzu427o6QObuwY9rOSXj+QhQrwtmjZr4IES2IqVobkthzKnxL+9IovhgIks
52GmTohY68iIAgr0i3HyUDeBiCHQ1IErLh2HQn8WwqV70V2JmO0+XViQ0uSxT8gRp4WmwqHnRg85
fRZbJYP9vArMUqmWLPuJ8FnuNgzPJpCeZvK0Boq5ThBfQsQJPT3hZVCcQxFRoeBBo9+DzhuSIpu+
9Pzx4rPC4RGp3iEzQaxunqS60SD4QGx6Q4nxeex1OLp3kfWxukJP/9ovvF4N+0+PX399uDTgiKKS
b7dluVFCcVlD/5ps7SJ3UDR56RmIPXmlT2e7IhQCoZjgZsFnErYO9QyKssvYT4rbHxNRvWN3tCj8
NsVLsEwRiYbjlhX399VPxT4+u157UW3RV9Yp25JQVp4dqZp4Rp4wxVebWhrhbpfbzFNsQvdp1fgd
gcEvjROlGlaR8HqLiSrwYiGaMeLtObdNNrqi1ND+SI5Ntkxny22xzypSu05iaCeWzbGzZf8J4U+7
+rgk9FA+/8QRIcJptvBucr/VQo9BAw4L/p8GSxaWS/rPYwTIMZekVxiZJNwYAwURQ/zIwC1ZIE7p
38bMHDYRypHHjwdFfNHXJXkzk+AlKx9lo7sy5WC2bRrv7PnVEg7+NJfmArLhcoJ2XDJzOeGFdk60
A72TqVhguMCN19Yq50wA10rsAZhWgo0++vTSCBntlqfzK+o++AWcuGUFjr7Hug4IsN519qmugiv8
y+bSPO0NDJtLWvFaF2HK9BOkzMALKtaQAnBG5oYz/1fO4DUbs3YrYzGHXgTebeAfW17lbGr2yq/r
jLeUJsjEah/metxY1/ueDLEHyUyRCy885vbAmbonhzUngcfjxhkeAu3b0mBIAOd4z0YoWgbqSvfl
GmmKT+JmNwFYB0FufITPUcTbPOi5CKm/hOOPnrl8YLZzv7MYD9ev9t6h0Mbyedbhu8g4Ji/F3dMX
NK/UZDY1PbBjLxcpqY2qVVcO6EKMoWwuwt0XBxSk1TvzJPBoUqCsGb73/USRL/w+zkAPOHOSfRRD
3qF781R5ctAD6vZ7N1omZdgm9VY69fpafg+d2qeLwHO+ClmvppFJ+Ca5UBe12p1sZuUiT37obKQS
OOL6WpHtSHV+wQEu3t+0TU69i4aEyiTniURqKYEWDVEpGfPYGK9fFAsexPSQrN4zsKVEMxNomL4J
FnjUTdtl5rE8Tumcz2ZxtRPLDsweEpC4td4ClSrLlq3bDgEZDZ7hCr2ROkbaXKuevH/Lex60aChV
17fSZeHEXQTOm9qU0dw8umRiYNHTwtZ3edJzcjL5Xotac2nqnOxSLdD7d/B7iClyJnLqXB2U6Yr0
9mgQiYi5JRHLj1MW/nL7GuN3SmZb7mNIcWeP40DGZugYcTbYiyRZOz+Q3kdqfgujAyG4VMRVht5N
rH89E6QIJYGhxepTT6yKKyO3heZND530TK3fkNlQhOKHLSceqiIX3XBCyI5ChuYH2K5mGvh4TooT
SeQEfTnyfbi3eAQlZ930/RkNptvM8nrgkehhO8kjZokZXQUM27DJTmcji9Z6KRDZBLjs0nQCFVxh
6rQlrqqIVJBNsu8Ai/+V7D357Gf7pXYEjTMj3Qd2wJJhGgJOc5cgLyOLyBlkY+f1xGgMsVQ7/qFV
NSJdCLJKC2jJm4bQ5fh3PC4EMlinoNKwOs+KRIuT9koDm737zOhrW6mMM8yOVOce/zLNh4PB1el3
0eTm6a4UhXd+vAFerFoDOF07jI8Yshdo8fRF5q9t0VOUpqJtHL+v84J5pzxyNiMmxYkjiWm0pcBQ
QUDwn7mgTaYhX9HYV1uNsWfw+ru6GeB9cRSK5UympwVRKgXaduIJql2x2zJcdR/kvrkh1ln3uEtv
chz3D3DWP2Y6+6G0OqpQRiQkbeTiF8gO6yTsZ1IzCsYr1vIJ4BLnd3HDhEaKRUW3EMqJeTsFU9dz
nrRsebLFoVXm/mg4evW3uV8xG6fqw3fhqYCrSmKX1eOM7tiY2iwguP5ZHBUTCeUuGXxUTX/IeFh6
KYioBMgQYqJZdV+Mx+M1zDAXOQH5VH8Vi/UuPALW1nrlLqPyxjwjHtGGsgZr9UdmcFkC6qq5hhsI
zeAXYowIEnQr6rqryvhfAmCJnt7vr45mEPdSYHUh/mO6ptYzQ6PigIAyrEyFKbr0S8dvH+YboawN
I61lG1uhHzsSYaITz3r5GqxxKiXD8O4R87EJUBZmuUQXejNgWaR5jzvHyiVxYgRMyee3pb5Wi0EY
4aany7RBC0+h5lZ+ovdQHLOW+vFTIBabvnFBXTLAN3S7eSu4Rwn+Hkv+FMiI2NwyMPrUgjidpd5J
k7eAMhIDaTYcEDSFnyxMRBPusgAtuKxXZXu6TxJc7XKE6BQ4A2EW0HYJaw1pP5DZiRXujM1qYHZ9
BZydffybUzjLrnjxGeb7IFP/TGI/fVYC4nT3j1CqMEYNRue9gHBZiIbzb4as2/N1hmjTGjGV3VDe
WM2kOSqPux9sZvuAaehFxC1/C8DGQBB+wcJcI6iCXX7TW014MAMRZMVRoF7oV5sBANUaItGMSwnK
Evs8gG0AHapu0Fzy/RQitggyf0E1jeGTsqqjHwZ64WJrffSTFAp4s2wKoPxa5q3AChNEOr9lVccj
mBRfLK7WEjKTHeAn+rRBMWYNfgtdIGI9ejpnhJskftRSzznLXju68dmaL512W41VzqJrQwFt1I/j
jvUqbZiJFKl+yWaE3ZF/9gjSKUWr3yOsNXM/K3jTcJPidUUPmzp4wLknlc9CUR1G3DSYNx5Dp5GF
5Z4HP4+PW9OjCBuvf8jcfsk2axL0vaxuIgcuoUA46cIoeMTvjgfWcWziEnSqUVfUd/RIh35+/HmI
vzamizKv8DFbZPgeXFVQf/pssWLd7tnfERP25+dtZeMY9/bXHXPoHBOZYz+2g3+tn9BJ/r8Ti0pW
9BMh7PTImD1K2mDmlS9Ig5RiDy/mxCoQuogm6+nFmTQe5ZZCx+tSEf3gGoVEr38FpIBBbx6Yn3aL
bv7XEm5/ySbEUCtvjyMT4XYqTePn+Rs40ti4IEl5SaYMjJTo6/WQQJrihqwYFFBGd7OD4QWO3UEZ
tsYfXfUFp5U59fb/Ir1NRTWO5obstlluCQl1OLGwLrOqrQNQa7pAMZTsjMx2WwXTzZP5c6yjF1wW
xORsan7qOeWItKFjmUU/IRfsmJNptA299FgPntZLsrztQF7cik118SBhEzi17yjmg6teudF07GqD
gecyhQWkJ5ncTVXlJ6R8ksTkMO/gk+PPX2gaM4qS0fPWQIRrpyRLdXgHxrWSkRko9OjWLGD1rslo
jSEaf1PS3XQT2lYmLGTQX4JCVVLj5v2HYDUJUY38ki8vhGd/bJZ/IkBqUKtl6J3nuErZehCnVHDw
+QFCMRW8ICwoTLv+ZMmz4GX76eABopxg5Pieo3OXALuB0ucezlvR/zBvtVsSOhbgRgMgFOMPOWAm
5SFL38nvk/G/YTvjH3uWTCL/+z1ppjE94zQqQvvsw7/vCudLGuragBaiCGTMOrPv3LN52IOArl1j
kKH6pUWGxR7HJkmwpSJmoqqNElmPu1dueBN7DKtVVQl1L/+ntPeqR7MDuTdMrgN/Njefvqc5mmjr
Ytx+ww4DqC3MUv/yRXqnT9YmqZdOZNuGah7N0vrw4xAaubPtKp1uzzjaP4lMEHP3l/GnNFLBMNJc
G3RuDJllEXfXZco3yYby0ci9bLmZ/fHs9dMTj7DkxAELTzH4d5sKKcxkcXz4wxH4E1FmPGijT2tj
qzH+JAAMSGcKPlbV7VeTMr6tNblXs6NxCKPlbiKZCncC8KGYmh74nJnG64zI9IryKA9F0ir9Mxnj
ALZr2h1MdRi2XkaSPbS5WaeAwMZbMoartnPC1D/V17miyp/qeJBVRRWOQ2D3BZJWtdBrqOi9HJNW
n+WEEIeshwCBYQwsJf5Lkh/4cA4xH6yXPWNPwIJTE2lL1ZPMIqNUOEuD29hu9YOzlf4Y9gAwQIYk
IHLfLYi1Vvdew+vlUTY8AeRVOLdfPAsvWz28GRZ5KvYuueClWtszfbpYvUfBn2zZYpPtpej+0/Ml
xlbzgFbMjYn8nxCmKooumBOQFcmj4O6PaJ0kWKGlkWjkGWlteymVQ6lpXdUhWKPIeT2lnwQq5nXQ
snUncc8Wao1SNTrrZDxidEVYpC3XI6sEh26dJzc/tI8CoBR+B/rUsv6auU3mc2CTbVTMstbhHWy+
qcelXA8C9znBBvhpkHdvK13LPwxXQBfi5bvVM2rmliqrFHp2VmheRRzmo6+tiZOFqdT1yrK5KyQv
PglJkcV3qiSN4Wk9yqLnbSu0OYf3pgQevEgA6Mr6b14Jcxo3HtHYKWQP7rovSSKJ+Vj2e4lJg1PF
mKN0kJdyohF+aJA9HABLnU1jYyMzBEzxcyfOeNP4gcN41EEPMDRmGsn8pW2ObPdQpl22FJbjRyzU
940y6XEwnyotxEVwg/iUOxiiFQp1VHj9iW7tbbfX06MOmcFV2PWwrqRb6oHcGK+fFvO41qQiBxtG
tZI/LnjQLNwoxxpLKXEf6lr2BkZU6bnUTWnqzD/Wj8q+n2DHIi7Xw6HPMu1pODp/YRg28qDT4wC9
ovBbophyu750Zcx4Uu9K5Gqmrkqc1rkqXmhxJFY4UF4ireq/HdHtvlN0jHWsWjGZRNVt7XJSOYdP
yC1mLid2Kj63DhkkZdLyI/5tyH+Z1nxuC9cgYfppCWLKkpFy4DHzQRdT1Xthk0wZBpkfiqZJUfnI
mxwjwrR5vYWioUfUIELxMXdRyo4VRt/AMvU8BuF3BLgM6hCBSS4lD6YQcqJ6BlO3imPHdvh8lau0
Dz1dJdZLSMJ5TfnNFSjt8u8xyg2MPVOEKt3VoKFJhgt78lZT32w9d0hQi1TIomx/44/WDIX8e80H
Xq6LFWGAtqDXRaaSOy1roQnh06QUFGOGUJGXjh36D0mlRYSAAIAfBpaGcQdAPzy3pXIgJVsD1gEL
+tUpdyhTetis/3AQSK8FN2yh6Y9nu87hjB4hUbMZTGAnrU1UKTk0lPFvO4W+xS3fM6w3RTTDkNkr
RWG2sJaDGmLuC6CgxPPNgJsZhuynu1EesMaEpazNSZQpLl3xEW9DKLGvc/LXKMnMDpx0xzDptuSG
QXQK1TLkTeOf9uOevS+UIJn29Lqe+GmTGU1OawlBBlYwPx7YCw2hFV+pXUMeDY4v2yRQIHY0RZTo
xQocGVgS37Yvwop6it3rmjEXsXK/cZ2f3KTCG7HL3si65L973sV303b/VGGNM2fFa0MJYzCEdewz
WasimtPDxS0pKiWLLMopE98K83flLzr5cDXc7VF5me9jpxi1UaBoLiFr3Dqtv3/mivNreAhvTJbA
21Trb8jO/fWE0xMDW5LbD+SJTMDoS1dZrI+HQdQa1I1pS3rA6D4F62rQlJZZOEyQ6Hkna3D3Y1Ys
75ouZnVpYQMQPjT77UGq6VJuMk8D7OREg/bM9mIjphV539Jn9W6ys9BWiEk5d5xJeZ0bEaLrHQzu
zD9bqtekvP6xIDQY7QrZgUV9uI96J11a1+Vuf2UZhgPy+pI2h73s7d9m053mazHCpH8JtpBEKLlI
uwBvlrucSJQqiQb0jrj37kv3eQa0+a04f6WQbfDPmconKYZ1I61bkkcmxZvA1OPagfQVmeWfnDBp
KfSknXj7lVBMc0PnIVvThUhnRhQXsUWu0v/sBijTxEZBopgg1tBIq6U5nhuV5yP6sfck9Gt8Kc4F
pFjfichq3Au/P6WB8adFBvE1lKwbbY37pJ7j2dpuOBAocDoyRwDESQqLCRiRStHAdeN0YuChCZQh
rFqnzKdHRiuNBXqF1PoMxkPO0tqcaMgoIUxdFnXuXIMHhefVQif59Z6ecbTePxhASkrhW5AmkhZx
LvKvo9SIGqGVhii15Waq76bSPjl+OySE3/WyLU7DmoRDWWvFIYMvK1mIP1e2/4AKXilw7DUVZ1un
hRLRV6SSF/gX2E06RjHVqOnoD9D/0bsClOASU07VrsJafh69+A6wqmuJGca3iOSPHlfgwpkRUhOZ
O/znJfnI0NP2CSf7mopCDCNdGBnIk6JxPZlDG9H1wqGDyYRfQ5cnxEoma0/jSdYckHEL4Wgyz9K2
kD3C9jmOE/7AnJS/6SZpbUZsb23xht3i6G9518zHuiHK9fG0/dpUJDMNnqWIe1h+wZpc6i9xKUDi
3sN1uFH4STu1RSv3jr6T+P4nBvtjtAOSpJodYRZgGdiS3g6fYEUxGtxKYVISvGTird3Mo6KXESVw
ojKbVPgCiqFDi05M7ad0ckvUYiUv0CPYgJEYKOBOIQ2a+PuDHlcwqT3v8LmFhv4hRJvrPR14SVSC
jDsGUR52APMOeEWczjE4jQdR6/t/1tMZzt086wfLxXas1cks3yFUt3C7NSCfpdcFNHxvI5xhjhQC
PNNmvUq66gvy1Cw+27X5DmSp57yOpCBSi0cizBSWrWDO5+k0Bt0k89a26wvq4n6g+MLMGV89XL/4
I5HYo8d/eSBHYIuiGUf79O8GD7SqXdW+nuUgoaLkkUKQ4RJKVrH9u6GQCd93GXBGCKNEnm3tu8o6
sK1d5jHspH6ThIzbktsxnEpmFKVMY1g67GzbHl9Z5gjCmN2BVmftm2TKIZpqxsWqH1SMV+lo+mgg
pcag6rlfmcrKBH2nT11tSNrcBXgWj96Kp0O5xjS9FSZ/3Bc+RbWU7kxSfixq37mPauJ+N8B4ffEp
iRVCfQQMunZhfkJkrq/EkhZnWUvsWwdxAveOrv5I8UHKiBZF/b5jpmOEK7hcqDT2tGGepoIxRq3P
R0C3D/jDs2Re8rNspA8DEErk5FtWggOfYZSDHeDrh/s8H3QQY2etzmpRcMcz7/Qv9lOd8BLSS1OX
3l92VB1PW6hPm4kEgzCtjSgdFsfSWUvCv635JPwCt1prLu08s7E9wjRUWK6vXlpF1o7owlx+DJtj
bc2Kbzic+p+61Xy7os4d03DfJi7WOy42lThAOqLYjB7nSL8JTIQJ1XiLVQAHY+tdpbDsx08Uv4tN
JnYhk0tDl4Fbry9VrwkhHEErvGqyELvbRa3Rk+/zsNnj4pe5e7qFC50bUrmKlkcuzPJXJ++MKz4W
+pcEEQP4XyMq56c5//pxkX0IWV7VrDg641O7e3u9BktqIQKKUUPlb7/Vbeo9S5rJdKnMYyk/sobh
tdupCf5114C5i5miLrK9VSOpU85pTyZiH1mFa8XjiPbrQ2DQUklJfE25uDJHk3JyXZmjkFHB/gkk
FPHTQ54Rtf97U8AnxQZ7YRBidrtMCaom+UXO3LLfYkA+6Q/9MWAmk36dw8aJwY2H4us6Lo6QPHLp
ufOuSUYc973zmJM9tBoeM4FSI5AlU9m8xxmOvSFhcN+9XaF8jbd05hWpRl06Xk5So/JlI5ucpcdG
+gzui8uURNDmSRX2111qOFeZlld9IvDLFuKYBzerJlZtvpzR7A/JHyZD2xpYgZjoRpym6bCJeCwV
/f9etLQeWjEtFhrnfjkaIU0bBY1P+b9/xRJ2AppC0lnfkKUfZ9l0O9JQdkBnQlNJItfXH4yROsMa
U/or15U9hyv934uzKtlfgVYLyRLxe5NTZjWLZVmLMdBHven9vx2V+WS19GQ+tEkU+cfxgaC0vj7D
7nnALneJwwYzipQ7hQjzzpI9p7zAYN0ruTczV87PH0ozl3fB9k432xGY+fpvfhqxeChqtRnK/U6B
37ichiPPnvNV3pULJffRwAIaMXeebe/nXrqL3eAli67zPOeUQZ8g2a0P+I8BJn4eGNOY7D3b0I7E
zDq6D03wxM7VtupEyByaFZSfn7luZwv5ns1DsUG6EBiXX94/7h6UvRCqxnfQclEqoRA0fqGO9ajW
08g3oUuBKiZKkvzLlbpHWnTz2tmVl2X+f7rRjVd2nSip8uXnUHBmJMTF/ZN2wi3iQgEE7jPPDJ0I
8sz2mPW3g5vynftp3ADfeolqjOvzYv0AxRUTbZb97Xo9SMzR69vNzk408jqMp4m85gUxDTUAOg3T
L0unQgF2rV8EGVXulw6wcS8YpI3Tf7NgiYTuOVNcavdjnLWE6EahG4nYQAWu7Vc8t/zJ+GAx+KK9
7CrwAN5h3B9r1m3195JRWRfxjUQkvxZlvv1UoaDdF6le2jSgvC8SC0Lx9wDPxSUtMrUdwF9877Um
YAXPeNOLbTl2GVLT2lCrRapkfTBCwVWLOs0XilNJUOnBgHd2JgzKcL9VPE726IGkMAbah7T9MVJG
4kBpiW97/0xEm2T29WVyXaeo1tBpdhi7O7hC3s4P4fpCHH94xlidC5HO6ln5kXivnatA4HVn/vHk
cIhEtxXt7Gin7EgFMCjkMp2wJ8INfpJ9H1tfA1bXQ04xz4gD6V13HhRM2JhuKScYq/wD9fM+CZg3
B/T0vnSTfe30KQ98Q3vOX6qQk/y11pdfns5xcUMCPAe3HOQ9SZVHKkmliNj2CONKrO9Qxxpoh77J
NbNSfTbr62rvtp0fKJVhydBoCt6FoqrYCBmiAEXu9tEl679slmqPMJst72XbazbfqfUQNzKbs5D5
aEGaqQBAhmBeeSY/DzLKULr+1+AbJDF2qfnXoTFaof2/+92GcUQuemHv2lYnhryedFQTBV8FIYHJ
gH1yvo9R3oiCsdghoyult8cN/90xGIGSPvmDncit+kfDEKQ5zjaU42THGss5UVysuyn4o2URm07P
zzbuPZ2VvXZGqlMz25BmNBlZ49G88E2XCsaF/wb5ZBHs2LDH4la9IzibZ/3tVqgQzNv1oDbhN5ZA
z3cP/tXs1/DcZcoW6wipLcXaOgO9ivvY0w7fiNAaASBbEQ7R95dDyzF42iKjohDKQ8p04rxxp5q1
oy9PsFCK3Cl5tvGRYfUOyf44sb/OO+5IVj2VarntyXcwz1cJEMNwAAC8qU2FggAXnvEjYmOoMKOA
WdzT1ijoI3J8SfMJnh6BqjL5eErM02u5mlcmXufCxM6KDJMjpXgb6rqdd9lPQ3Z1tf3Bl5VSFUOy
4QoSbJ26jRNhO1l7RiNk15j00EZ5kODz/r/TzoOT5wVRqE9tdgd7vsMb0ovpoVFlko0pg/OLZ8gH
QXxV6hltml4zMglQQ4iVpNnx6hf6P1xnll35aJgbcqX1vTGY07NLmoFcz3Xoi8Oe2j4nc8/roxYY
4ekrvT0eeQ7KtQ0aYinBMEI+9R92x5KCfIRKP89iTLtSS3hXUOzOvFDpvjrl1isOhj2M3/jfJc6E
Uu8HhWDagMLSMgMdmCLXl1ir9sJoSNLVjsG6y8Y7638FyevS1YaGRn8g0TfodDy04XT8p+XDideL
RFSQvcpwSEq5eiV81kg7jkOstiyKBop+RVGObpDnRt36eBQ9bZjSZrZnd9REsD5BtiVci0CuNlAW
laJgdh653J1vxWDdAkmSowtTNGETbwSo5/ZFW1l4wQ7OHL1wzDF+lvN+3sq7cPhTSxwS/dxf01gt
cW+zwtXnGZTAsQ1uX2Hb2ryv5IW7nqPU/xnygz++VhA6rs++EkpQ3Nark/cmwE/myou2q8Bg0YqA
dcfePxG+pxHfCYWddQ9hjKGZNIpX1PyT53sKMmUDbgQSY2Ym/ASHbTexPonn4QkdC1uIi4HgKRXy
HMhvn9F7exeyYfYfkxZySxPpfHIpA8NLkEYTeq1R+asP8qcMZphN4GGyPBD4I1tmo8qEkMY9rWDV
8fvfXOlPCjceqtDfoqLLmjzwS/DwNd10s36kN9OhsUx3ax3PLK+a8UJGH1M7XIy9qEqO/KpMVl7P
elPtnDH61WarLBK3tHjhWbVUw1Y7JO/5/BgnUUnymMeIgbvpnD8nY/pFqHhUzox8bTCFJ7iEj/7/
gNoMF0MNdr0jSOTNyPPJyzLB3iGfyMBtOP/CdIX+6H71Zzsqx2jx+oBZyD0jHjy1sTIV4wvhMbez
MPGVxeF0Aynn9pj8q640UcLZX/+xmhyd9USv9WKHwLTBZA1REqeT1FcbWSt3snVjuHP4zy6eZ2Gq
49WNQnx1MP+eBsuxLitq/hpNiAGhXp4Gg4cWwIlsB+JCOaPCA2i8fyP8VhGuS6oQyyOsNkIuMagx
bcpuzApgXtFffzMzw8f+B4eWUuR0gnxbAs5AVomNlvmHeZecQgDwKvKi1E0jl5UXiYIIYKDhxAJL
t1Fokg6YtQ+HkjZ3e5Yk3qnLrsm5HRokySlpoyo5ybaydd6ZV/DkAn6ex7v0UsakbNjYAGLaEcDu
A6sZ3/oVQ0xGobxlG8DzLduuAs7UBAHkchmcXASIOGXv8WiMM+HUROIb311usfdbybRwutga68vA
uwlRrYeSFEk1Mf/Wv8tWQOYoUPTW52loLA3v+Cfjdi2cH18AZkmedfN5MzFTSQsSy1tX9dzUEZe8
+vmY6+MOzHPbzoeqUdVVG7GBBdk9sBb/CHi398oJXxI8WmSE+3mN3gz52OoJi1S9Jl3/RktaEbxz
BWii+LldQs0CWjV6GX9NuLdDnvdg2+getyHPVPEJBBz2cm5ofWxdMLGsIrdTytf3ubDdiyrjHmks
lG9Llu0RpCt/XV5qDywkvAtthVuEV2+2SfZoUKJaLjpoSAG216hgAtJsKGSSEx+Dm85E6uOFTNhx
ipe4XqaSsCGajNTDjJXKvVWBEdiDf5ybYcnaNkrxuLHWMSEfmG+TK9DNpBBaXz2m6RvTs5mCAwFu
2spQNJNxZPGlkhRBqmhMdahrbnGQHRoTYWvW3sTou4x28DG2TlH7diB2rFlxtPfRpw3qzOLyT6ey
OZlP4vGhTBKoJpWm4+duIJXtO/JCkM0Z/7lv4NNsbAVlMRGE6yigzK+otXVXtcHZaoSD8mfgBIRx
MCrz/Pyjj0bsQDGqRxxtwaj+FN/u01esNpbIWkFu4QFjyTCgkMFME1F0OgWVcDQD5KHurx3QLJ4c
yWjPHbbbGRhz6yO5WyMi27EBsHTx8a3nqAQIjsvbclqV5iE7V+yuP7tbekdbzARtN0KTUjbtrrrW
3gIBYRGAQ7VsWP9qi2bzmRzNlgvw+7MsUVxcdYrjaCw5jpG6IydyzZLdVKArf8mzQBEGOaaNpk7Z
s6KONcszQz/gJTLk9I9WNWy1pNLZV5edI+BxuEyre4RMCvZuL1vbfIgvhT5v9Jw3EYT27EClOIVU
SUoPLlK1jyWTcPb0sX0QBYppgQ0WJ4iZ2ZPCezlfgD66GcP0EKIIkhw28yf0+v29EcwTZDTjMspP
n+izG4qEZ4vnzoU9CeKzqu7wPpDm/bBYQsl3k7CJ+kzoAIy6hspxchVI4kahoCDifEQuv4vwJ7Xe
ZtHqOBH+Sd+WwMvNZgLoSlmvka8jnBS7arFTrHK87UWq/JaPacf6RX8Dui/Guhy2/NQv4QM64kM3
vlYJNT2w494GZ5RpgQ7+WaHJY+UyOSab/mkQ5jLpSXTiC3Q1hH/975wKrTy3JLQwj7g7fyNH1R6s
o9PvgUwhDsyhTeXL4VvhrBFJcFU5SN7+SIJXYpefEDrSXRs9dzKoM6TVgFHwRxW1IiNoKmhuC1n5
Vr2CYvhLuN5he7oNKqlB5m4Vk6rd35J5q24GdKvL4ibDDF6DRTWi6uKCTk/UXTwvOEiL/dFNLh7A
2sG6DN8Oe5OvjqmJrnaeK9nM6ofIxQOkPHJ5Sgnz8MyyY+U2LEv9X5MFvM6QG+8re+WorIBPdAlA
LNyYPp6us7LgQnDuYHND0fDMcMzUoy+Bb0sZn7knkuqa+7dExwDPyUY7ImhgUZ/Rxcvgcd1QN9Wi
7qPDc13g09xg+g3m15y+0ZdMK3AsXikeNVdutJxTtxz5X3fnZwOfYn+jHR9pKTeQX36RMROaC5Ej
DmqbUd3vhxXwM7w5jIw1s0GDCXMcVloKikGeD5ZJzct4MsAUi0iST1NHFxtWMCgrTAkXZAi5zmc1
aHq00uu1nVFKbYM4gUaE9kahYWHUbjnJ5MsebypfKJxLGpSKzMTkFY4Up8sByMrpQbHo19+pEnpr
eoYl+Q6C+lKfCabVRyajXUf0VNF5go6XYT9Oq7WooQoFSeJ7HLKoopMXM//qVXLR77IlK5MW2wyY
zOAxc8er/OGO7WXcKJhajtkg10xgUKS7az+NLuhZhfIbWy1boF22sEHyL5JLbSzX9oQcNQo0wWjU
byODj2hOZnlLvos2LQRCcXbU2YFsvpMrXkY9c1t9j9f4zw8A8SkiKXYT18S8vDahh/4mJyrrqc/j
NlU+1gI4YPLEKgLiIksLRQOdSepBOsRmuPJIcIiONIh56bDj8woQeCkVOdsmNoZlObmRTH8mB/dt
fb21CPk8lSDDTkPA4nCrRmTgGVKEyGcX0ZnaZU36ydmei99DBOh3bc51lGStKjPnU4O+B67f2nL5
m74NVT5+K0W5RnyJ079xEGmb4wy3BFHiX85xpFvh+6gS0tRsGv/UlfxhkAJY+DXPaYPfpn+fPnLu
Ra9CBeZ152zTUQAKCfYAgCbIBUjLOM6ww51makerOahPbN6btPMtT+KGtb/9NgFGuHsrm5BYkceb
TXZBd4kRYktgwR2Qn45qeZ/F0qsxtXZ3KIY6VB9nbpcYYRtgiJy4KCuoosfyt0Y1D4CfZSg5ZLYU
NnE1r39JZcEOcfRevxRnLwrRK2BTyH2hfLiTopna7A39bLEvRvZxoiSaix62zgrem67QKkpbkpZQ
0VoRjFa9uHb28mZ3m7DZI1tae4nysNaErjSd3Ew9esAKGo7RUNKcHA8L94oGm4qB95sM0JXyP/PA
wqHbAEsp33Z2uiaEw4N33jsIEkrpxk4XB0b2+JJaG4bpY5m5wmqH2PTTldRotkuFVm9OPvieYAbs
03yqPIeApCSnBu0LVvt8351uPqUZoW6qFvbaBMAqgESow82Reval/eBRdn0P8YhArk68eIhM4D3/
uD6970dViCnv7MmhiTZF/S7pB6/cfGboGU68THtd+jOHwIRUidNbPXgJkH0cEtMjLrlWV6Cs5sxI
zwSAkAv/HQEkmYkrHYJ/vTH8irjBGPca/i4I8wVTCNqd4yVgdUpBCb6W/2EyrmPRRV9jW0xXUKiS
A/CXRnGzff5EoT5y58Po0uiRVhK26g5zqp9tt30dC9E4rOuxEYNZWiyswf+oTZnV4LfOmouW9e9V
N3d8dO5GDU15vTVIhH03+NTSMFsXy/YDHCQdNvqVMB4dDS/AFyvB7vT7MRLd5xkq5RNRMQ1YVDaD
0uYDJUMlKw4bbq04EehSTLf1glcXjIgs5Q6JCmeyLhCxuHjVcPSUPXcqPF8qaXi6ulOkBMN7RA7C
PzSlFj4evUvpjI1i4oTo4wvgpuZMPICVwica619SLlbIvdJwYeEvoIfDcum3LzymjXEY3/eo4ZeC
Ckh0tG1N9/2ZjH9NKsZp+ji+nNLxv/jNm78t/nVe/Iym7NVkKS9235YHDjwZjTksJCOccKULgsjA
S6cYqooGydNYNdb5uCMtRL+rDlNwZVvVGNUNH/LeMfBwSVoO62JKv3A0GIGpCJGrIymic0/9hM+a
znRvtlM6fXmX5nOCv53JH4QmHJSL5YGlvz6zg0tbdTCB5Ogf27xbc1KTXgXKc8JmJumyvCFXK7vk
TI0SCLYtRvxfmzHMwJYC+vb7cJfqp/F9bSw2Z3h5t4lnqCqsOBpWcIyUAjqy0ZzKZ54pAPbhao7k
+rQkN6Kdl6Rk2o+YrGPYIpVNAwHoy0eAleo+Tt1Wvqg4Gr759Q/GBpEu4aNjqA7+u2vK0F4yzLDc
3zCYpZHoBWiSPhNLZt/OvNbFqfYYdZ4qrihn2gdD3zewIQoBLW9YnCCvfBOScCjKX/sMJmBri7Qa
QG/AFaI5sVNx3uNgRqrQ6jb4/34x2UvfTj6DNkO/0x0Abz34c9E3vej0sZ2YbDX8JqdEF7L9fUU7
WdcEx6fwFgiP7FTj2GEAAwf7faWN0mXCINtp+K80chmLVJCRw2T9+IgCjSyHMItU+T8mrIH77f51
SLF+EZzkdM0t67aOApghhdHuF0RWJh9A9FA1l5Da9jJpBtHYAzdIlkfHaz3LqeNHBx8x8AN/oM+r
+3iIyTxC56alzii+43wxB4xoReWpCe81N6z1OKeeF+wqWS51wFGEgaj/qXPuDj4TrhVtNne5eWkh
7FMWT4MZghr8KJsU805sfx6dsetDaEeYx/2ROczNH4ZKApEwYotdv+mlCvMJwhSiEN6uq21EtULV
j7A0rmlzT8sT8RMZpOjFK7f583yUNyqavm2mweSBEORRAkSlCc0nAAUAw/jNfngiJPZt3rZS1Rsj
+hNYKlNUcitIFlEINdEwoIiStKvP7kjUJdyqgyXo1+aCx97GPZ3UH7J4TMGIFEmltlR089CZv/gi
vjSVPbXImUmsYILjVvYars2BShY+Tmw29/y3lNaqyV9f2yMLu0zrFngXjFAY/qfDBuEOUko0rHm4
JGMG3t9u3/7snhAiQLt99bAeikiRgePddd3zOxI0NqE1andLPkCcAn9K7+8/OfTp43OxoaMtkf38
7XA4CPDqSgVuAcRM5DooLE7ADh8nPMh65J38JDPBz5MOzSFdoJKbY3J5ct8hwUIowaNsHShtMmUP
fXKU2yQse1KI57aI5DXAjpZZGwBhyOcrm7W403brJS1IS4ctjaeGLBuONar82c1pj7093kUvbdBE
YadXFDDt0Dl88g75E9qo9nByh5gZXHWrJjXIkDYXz4/smzOt/HXxID8XXXObHOgwgFohzxipaJbk
IbmhtxyO2RkvR4e2jQWzHcmsOuN9v+fZwZg9n3HjCzldZ9eCc+Y5mV5g9GKi2hHvyCLnaEidaqqH
P7qHs0USZK1A25c8uhdWsus1UHEVAx8NUmsowzmsEKp6uslQaOqe3ioYxSIYilaXHGi6BCAOi7QG
SAXv2vAMY54qMcTS1aKL0/mfUiR8b4MVI/vBIfcFLypvAAds810X4DU5aFX+RIo6rKHQaCO4Bvub
qAlr2tLgC1KctghJ37ECG3DmaWRB3VTHviVHGPebNsmnMnGIymN4Tf98q0gmdQa9/m2Ep01G9dIL
KoYCOIWIasRiMLYF5TswUjctbfTUeFdpZDRPjAGmI160FaTnKvdnMXn2w1MZ1TshdFqrvpI2EfRC
DKIUMlVlKjBuIyPy1b5VYiJSZjERFJfEzfY2AONv/+KZwANT3TMk5sK1wG3akNFgTTnvAfDFe1Go
VjTtU6+2eYkM7a4adGv6zyo6zX6/6RZCjzKE+hTQ6+4ZqX83QojClNjhXcRxXVvJFkwwU2JqXfIf
3GXIkrdfiWEFmlG4ReyZC3RVC5l6xpOJhItLIwZPIHAgy3WeoHeMI51Ym+B9YUYoY/1pKCbRSc3/
BoclgtRFuhb9u8uLj03NSvqhUyW/hugQcHg5nb8rfKLbRLx9IkYKW1PoeC9U5WCmcCtrNh371CvV
fK8bJs6H9zehsjzZdmZaDVdv2szl5Dlnt9Y5JVA9sQpvJyM0hzi86E1taWK6+eZrPqhb+T5FPB8y
f49HbFmQRsWIJQM5LyF9opYXilsttJDtXl50MJ/5nJ9fzRPmWZIk+9kuw1Gr0LvRBE8szy9DIqyd
4YXIj9EDV1mLNoT7ooxpM+rRCrjoIrhWVLyIOgqzR4pWUko9PntS/vocjW3tOfhwUg1h5a/k/pb3
3PvYunXi+2MukXEJ3FSnxgqJK7/EkdiV9O5jLSO5OFY0PN0FK/MPpzXpwzGgkX+wdK8lhFmjePF1
h1qgJn41m16rEcAr1l3f/OOy3x6NWN8EAhWVshEvHU0dpkGJ67JXj37DdZdmhAEE6A6mS9m2jqUk
8zwIzj6fawLF0SGiJEAWsN0wfweQrvZrE2SgVrt0CyRC0cC8GfWmwNg3sk/P1jsoyyREBmTQeZGl
Kbo34i57wl9tdTorBMnlBZAdH+fBXcfgaJTlZoS3OfbJZmoTnnjrBh1838pH/gItL1NDZkHNGn1w
T0IWvUnfUd/OIXbvXF4y/5xXuKJo+S96NdFC2GvS4y0VD1qdXcv32Wgy7XfSkbwoyvF+Q55V/Hgo
OaDsEydUmXdeasO0Y7CEHjgf1AfzTcPqyMqRnAUJvQxb/JPpHfi/31HAprHnuQD3k3mzg8ikDJmv
yAz0mK3y4v45H82Fjk6KaPVsz1wq4hmWEkFP47ecbdlGINUsJdZs//K/z1UCo3Ss4Yy53AdRVbC5
17pEjz2ApeDUA6QutS+zpssMqlzQRk/Hnx2jQX89jMPKnK0xnGdjBAfTrnA8NhThLLobkQ2qLodU
CyS0VaA5XD2O+K62bMd6McjrCPioCMAdV06flWFWkxoO3TH6GAEQFQ0RtYdqNhgpBf4id2Z4MvWv
UkDPDCexrR7kQWymMDeOGI8l/PauogA0Df1pYHIhdOFK4fb58i/B2Nqe2ZB1iDe3HkkVYIKnKFpV
CeeRGimuaVtvco30CSnBj3I+yjTkmP1VJv24b3mB+Ms8kGAxP4Wazg6SaueM98ydMYVFjd6bJg7X
EteLj0p6Ir5oAYCSVW83bPCSwkOZiFKyO24FOBjPh+cfsehM7QkCB17SS7zDeE+9EEnZl5Y+V83l
KHgCmdCBzRJDEBL76S8oZjVLvTDkNySZmAkdI6hEOspRU2IfBBDp8vHNJBWcw96e2HuQYnR6Oaem
iRlYAEugsh+0M/c2JXe/0W9EfvTb1/MBSVbptIf+pFTOGi4sCkm7CF2BT/hWYCoxwkfBxCL3wuiz
OCKaOA29eLRgpqwYJsd9d8P217bC7QuyQ0IT5YQaPz9RR45Kn94iIx2U2S0n77YSXYDwcAXarzXx
YNYHtwArKnskqJKX4rx3LRag4+y8Aunilc5BO1/rNFKP6aBf7iWDEhOwYFDZcMloFpYYCJaPkbjt
koQP5CgwdMuHuGg7MmZLyXQlEVpcljkUgDJSEEVfO7erOWcGUi2N0OjJgR0hvHo3Dfa1q1m4hxkV
Y0jgVtbHJdzugZ8l5lZKAnmZADRXV3fb72KAyClpSH87n01//owvcFgK+3FMfxfZNZ+WkHDCs8+Q
4DL/qehLyNrLuqXxxmweMWEUBDBi09NutUrs6Jw6KvPHJVPzdnZGKWYjbx9KWaFBzjn553WjHyps
4XN8uR6/ZIH2TQczJEMqe2vp4DotDLRGEgjK81kpaq+oLYYexPWm0VjK2a1CviW9MrmvtLDpnAQO
NCgnt4d6xgmIhb+GAKOgXoWSWZdofu1FVTV/vvSZ+zssne1B9SK0hgxBo7gKm1EEKDuu77Da/fBX
IFFy659qYKaZPtBAA+Du1V2gz7yQGzTnFDxXpHIb2vGmEFX2vkwj3CAxQ0YXmZutMXbRzwrlWzq5
qlK6Ql2ufcEPWvBsviicYfbi1C76B1z+TgoqJ/Z/X9gdiOrcoyzm+gu/YZ36XUPdfBIDyiLlTYCp
W1d07gJ+LOyyTsrWBAnrRr6eZRQeqG6x4dT5n+FMbv2wtytPFB2cmeLGiKZ0BUIQ1y9geguGKaMP
9XcoA0aYniPlPByBu0piRHjy28KsqSLPnb8e2T7nSXA8DGR3JQzekiKA7ReHwV8h5rbNIIohW8jp
K5KtvhNMYp0Xio3HDI+vSms5/i0LjwKVfzWmrCPkxG/+8LEPjtWoNeXHj5TAtOm4j2BIdkRoRTH6
pEiYu27KxV8eu20ReXNAAqrEGa7YD0OGP6heY7kTXNHML38Blo40c9i9lucYhXIf5j7hBVVdbkwK
bKibIMBa8j/xTa6Cg8Q9au9rQmTQMQhYZ2pwFgMjMrrdCdNG3pr8MtzmWJQJUuxShE+q1N0gYsuY
wnFX936dTfCj+AHJmeQIJyK5+RJFSkIq7dAC4QUG9oAirf6Mt+Rw1asa+4PrUcet0dNLW1IUGr0S
YV1CJ9ltrd74zGiEJF5NvyEKr+yUnsewxCp63rToBbQh0K0flmTkDTpYhsMsZ7mqFddihx0yC6v+
y7yVPfiy8UnBBSAWh/iNUB55Qo5qisCzOxKsd8bP2cz+AnX7I/2fREvuwj26XKex7BGEi5WSH+dR
O/ySZiAr93plcL2vZa8/a/VIVy/xWdLfCsJswWrwAJ3QUJ5TDNA2skE4sJykmlTyWTjVXdkaHrga
fe1JNGoHh+1BI7FnV919SL79xjtynycYXBJvIiAbdhFVV9/VbPlwd1H5EMyyTD79Zy5Otoz+gI0s
UyU6fuenFgtRiGafEc+L8yJPkg7AUI3m9k8sH2dr3CRCkOmIEIT7IEc2+pyC05IkGFuJA1x5ngw0
kmwRXy3cUAwOEoteDf8qd2P3Zz+w/7kKLmO/wxw+rgZ0/BBogXoynPmzaV/wrS3H+/DHbqX5Msqw
xlnlLma9Zx0l2cO2gYfnagM+fOG9m9yEnpno4wwCN51eGdbYkynyi6ob9dN+i2KybTlmLmSu2q6R
344qYejuAIUXLHFKS4P+rT5W3WrNVdrCAHJg2H7qY7GUBPY/lEwSldCAIyrWRka0TCimG2gGgDSN
yZug3f7cX5cFuK45ls8I/WMk/12TYz7IFZBr2KBAyAiak9wVej80aA50pjlf/LSpKFS3/UNH/mcs
KA+hIPEfWWjMFSlcDlT+bYz9GMNYxqiRj2ZqLoWYUbwvVWX5k35MH395qp4Gl5yFN+9NOVmb5tkv
SoIp54C6vPuR4OG0WLv0A4KS6TK4zfzE+ybsJU+RRg24lJ+kYDhJ1IzFJN6FmQzGove9JkTyoHDv
L8PJWguLAPyoGadIjv518Agqn50Q9srOsWBUEbg60Ge/Z6e1ILbbMceTMqp5X6kFkvXnmP4EUZeC
/dQPTZq59DtDlh/7ldrZUdLc0fFDUuLpWOOTs3Ca7W1y20JrPgpUC+zuQzC3skxqbxCD/z/QRgKO
/ms/ro87As1XVZ+nri9pI7IkzeYDiFDzaSE9qTpdy1GUl5olfs57n5MHThEXYyQmBhOYhd9Q9QJC
eqArCkdWzP2OtJprfUJ0sg4eO4rHnBdDWI5dW7TihCgwGgqK8ajYVKJkk7q8Kj+F83lyWMFnZaEh
J+TQNzU7aLQ+ZPNTx9HwbS8nUFMbPeVkIDRIvut4HdLMF0D+jELZJo7hcH5pNiPkdozBEdDS0u9P
IgyRe8xA9HdPLgdASdf7FYXbRcKFYElTbJzZ/NOikH8y+LX/gpeWDjxRxJahwC2yw31nIlJ/LtKV
SDeNtGkazyNCpxUiNSecorzkus2JADJkYXj0r6Of5feCi6AA6ACkBgVJbwf1tKACQt8oWpigNIgQ
WB0JTxjajEuv7biM0AScof5lBGQZkK7CXUSsI/u4d1FsYteOobh4AmjLp/0OG9tx8vweUHVsKPgc
5cO8JJw2VN+8awGr0SwhK9N7u3QYpiPgEJXN+5iXgy0g9h0kAWekKtJUHW6ePzboTEP8iayprsW2
KZ0Zh3hWbJcGHseQ8JYMQ9ZNHGk2Xj0RtUHs4caO17HXABtHJjWu8U0iHPz/cLOsSw5I47RyQejc
7SkTqcXrV9trE600MyinyIGDA88KUkA31GmpiSBlqhtrwrFyZm6WzoYHPItogkl9Lxapx58//15S
r96BEN8MJaf+KhQSd4pOGuwbiVBakOnu3nckLHKOC3Qdy+vZ3pHvyB4/RJyNouMTYHjIBgGJe4+z
tUOTIgl3f1e5p4rYyWr4w0anKXu+eL6TUvBQkUR8D2/TkvcWcIaExyvQnTuqTfB+P2TkkmUIFlZ2
9I1p2itsvwnz/tt0GNzo+fMsA+YXZD4oIvKWHdEMreKz7A8t4p7zAEJO1puHN/QOe9vF0HSMdiQ/
e9n//t2iGYvuZLSBrdNf8OL+k5dRKEkQzqYXpkvsY2dvE4yEQ0+tn2nGQbTfrOuotbCNs7OACD8h
yPCMV7oZM1qEEVhnljJWoegguKuWJuc7i6grD94XXPdn/HR+bHru7LZRBaQ93JGViU/AjfEX0xe+
yG6HTkOcD7Pez6B7qoxW47zm8hfNjaE8bh+84cG0Ebh5tWSvQXc1wFYQXjasSKhSN9UkzN3tJdkU
0H2bON8KFSd8AJ/yuvzeJmDZKcRSI8L7c7mvqh3Pq1Jev6q65unpW2vrapR+GAGWKWgxq7E/hwHd
03fpUWN/4ZTuKlCBhx1IboYBuypR81yin2xikADD94oRMWfEWRkLmW8wFi69JvABQKyXjssSH1jE
+L8I7uCd9y7sEu+7I1WgCYboSThAQ4wgciMgwfEGc99IcsTLr30fSEO2oGd0CL211RdJhapwtjcA
rEgJgScMnme6+cNp8aRra2wPHawQZDIgNJ6CA6S60LfFcBB3bfwzaLTStGrXusOVcTtYnBdmv+Rk
YT9Mwo3fF7pMVwuAfm4rITiUCA9en2oXMUI1XzbpUAmmGnqbVC73IOjUWukyHswCf+duyg0LBVfY
XWWdRzWbUDNZNtE5LI6XJJFiCHS4vVM/i7bzHmpCSNik7dZYb1MxS24jE2anRHA7nmFS/mh5+kB8
jf1uVEWtRe1je+Aq17vYmpTJ3KKYn+Xpoei98C6002qKPp437L98f2xs0pKe1t8LJ/YYxAcEv45G
Kcaj/SKD69aF7wHZmnWKC/jkoqTsvHBHueafhvvf5DwNGRSsneOaXl/CtZRY+zMwcUJsFqIaggpX
OJbMRnW4Vjk8EGmkj++XfY3l7M0Kfo0wZA1OzacYbFT7SPvvkb8rfE2BqxzKUDkfJ60/PnqfUSPY
bdBB27XpCTUCGhRDHvp/rgZCCdb2UEEAX3o4hNclCoist0Hme1Ge9tYRhWsfLoH4CTMdw8yO/aIP
+9yfVk0emB2FQ89XD6FYhLg6vMqGZU72l3l3gyRJ0Enqv2yJKiX5t7vFAuT8Yo5hFSLpNJ6QHjYx
+3/UaGNxMVEhTZOy/XyGtmLmkQvOvjgMWypBHRAWUcDOyqld+uf5H0JARo1n4cz0Elvknt5PvGcV
R9xOWbnMBrj4Qp4QRijGmufkvrMZL5NJGTellMubUvBryflXtQIMujlXdPDdZvp0iXcqaQJF/nYD
X1IrJFWrMYcISthbdHl2ClijYjHqQPv+hjD8DYzC4ivc3D3SzanivlWbHosc5j5LK8OB1iHBlrT2
lmVcx5t7Stena20MyjT4J6J0cGPzX7foUkosmOYhcFQQPFyOj90HWMfQ/TRBiyOgkOXM/80EvIkl
2wFOMYl8p7QssfJfkT5tqfN1GFVabpXza83LE/afawQw+HzT2bgbnF9sSLl8FBt5/4ENhOerYhv4
v6S96435AMpTb2iQaKLtG3X8DffKWk8Px6GHM6tIOZoQG/i1Hspq8DlI4X12vZP+3X9DdOCdCSI5
TBjRMNdfN86VmePFfzITQHmhrwOc+JNPNtt6dnvGmmlWSa6WH4NyfhEVAMc19HZdfSNJWH7IKzcq
jIIQZOOLZl9wvGDX0y0YLQveD9rdqeztNW439WCV0qQMi0OqDURv5CwOD5XXmXGUXeWeSxlccBkm
qZ41qbpSZM6VvrY7/GgXSYu3cBvKncufRgGYAM4wdpwa3UyqClNm4pPmHNmAaepovSuty4St+9Ty
xfbowXv5BkgZazC8dVqVIOchRsJyOiOCNo7yO5VJkwuzvkcG/qC1jo5G1DEOZPiJaZmVflK7G0PN
IYcAKKFVTpcALKQfvETaDBSotRToM2fszJv1d4mjKXtEP5CBnh6ymw3MlH1Ex5cgEOGmBXrjuYmv
AghixkqgVNrVcrswKmcMJZ3RTiYh/RQkYuhPUsRAmgqsoxdGB/u2HCqG/OE/34M5jUU19adKUDFc
8n9kkT+qMxQOqnWP8CnKj9O8b7F5Qsx8UsY+xceoYfXcnVXh2UQm/8trPBY/SXnxwm+DQpHtfvxn
ofP9Le5EJXVQfSKqXZIPBmPRDT/gz8pfhTtuvzxheQl1hHMdCvz4Aq4FgRwwOvAdpJvzHdeY/tUe
bKJ3EGFlce888zAgQRaAwZqZGPLNn8Ve7ldWdPALvA3bCwIDZgdOsyPbE8O3T9OCP7A95X9VssmC
ehv23aOUehU1+9rcnqmzFMS0FIF/uA+Aa08buomHtuYS11iYlmATJwGpEvnbGWaZ+sftmxLw9Ycn
5+tMAXWk8s8552/rXmMCbHvD2Zi1LR1yjxbadcdKaFVB/ku/25naq2qjJykGxI4heJwvQkCtvSuy
8wURYrS2sITQsDNC02uZFe5lanMm0VjXHD9GG22DtVx/P/NAYb1hKgWm1e4sfjkqlPxiaN+WIUnS
ppC5qGtQf+rFPlle5TqlRTe1uq4+uHSbzy47/2EtZ3toGOwsx0zHID2hWwoRCx233g8K4MLRY6IL
/PNF557cMH1JmiWi9/yQXDgglHFnEK3yHYCEMf7ZunXyjPDBETrG6Yfe+tjZwa0kX1t2yuopupyz
4RgFSLhW62sSUZVu7gfZNEXpBYwdkPt9U9NTi9dhrrLTLZXNg5Vfr79sMXaejCU9JseUxmCIE4zL
PNVFyHXSSO+QP+bYGAyjawXIVoHsUhGVPlCM9F3MrXr9KcLJnp2aVJpfaC7E2ZlQ4R+YUs26TGeq
jN1GndZM0SZUIFLzoRxW7SKyLYevdpeOmiERR5N6ARjZdDma06Lb9opx0SUeYf4hovJxP70TGBrQ
GeZNF+Ko0aUv6wB61URgbQ4PaNGHYFGCDSUqFuOwsXpSRlA2nq/BGhitTm8AYggOgJAGHdw9dZy9
oq/3ruCz6StuPAYo65mQ8bC5B4psH53UQAUeG77PO1g7Y9WZWqGrr19QSlIQw+CFJ79YUlbw5FGy
Q903DKJaKSV8MWEio6gT1fRFCFLsV+Nq56VaXxJ10xDOMTq9kh0duslN+91NfZrO3T+XWW3/PBsJ
XE2UBqCkCSeOJytP5IcismvfGlQk9mfwZSbvhwwrVCxeQsb7tixi0WIDKAmydVRPB++udqPFozum
NnPn4w+3O9CeEDYo74WAD7nsf+5Q1BwGg5viOIlVpzPEHyPUhFduZMQPqk2Ri8wZioJUz/y/dixc
sdDo6B1Mgg+d2tcS5mJLVOzr4yuEcjFG7K9slRX+Ti88H0yCLVd4cX86q3ExN3ehvekjIwX+1PRK
kf7Q72cCvZO5+gRzMe8Wrpl61l3+tBVO44NwdAk36Wc8rCjqfOFdm0RHebPu95CMtAuDodRz27rd
9pjkTpU4Tr5qm4Qns5eza5TDXCWFgzlc142FI9HyF7uWYCJf8OQw0w0ZgMTTGd67mGSyPLVF8PdP
7Hg6EDLF39eaTeqAjH91Gz8W9L7r18P9KucuQzQoKRa6yXxQ9cQxtrKE5aCwUIeQRBNWdSg6aAS9
WP4liFHwPkPwsQVE32PJd/zrDFkRugs/TazUNmuXrBwkQxdgWN76Ufbjcd8mi8C4VVNrZMBVU4wU
DllgPrpwrvvoOj/YSQ6gW99x8dFe9PJGrxFRgynvefpgLR0z8RZRteZGi576Klt7b/PmXwGu4Eds
5/t9K8sHTcZTou2VzUkqg7Qm91NjqPAn8QOYgtVaOoFp7WYiiUBUZ91/gxjQXzZzNRTBBMg/NJN+
njgfbHcxwzpObI9yMtALhBOXViVl+/p5PwuVSv2vSlHZZNfl9Wyjg5bZF0smuF74QoMIVtUgO3yy
i2Rth7FJLKZHtLYtgDWZDrI+arssKIfggMcUNOp7NlzFNDSUMwN+gml26Si5QGD+HSHjBXnswYOO
pPJvvKB1aFZTrvJlqGx/YtVwGlb1SaP44Dv83IhSotdr/wAzFxLrvQlWIw3sk6Hsb9RL5mMssJgs
/+H0D4EnbF5UU+Mz8MwMVIJRUsCQIYgXR5Ize1taKRa34lML7oNkBiHlofpyMvhf7J+b/assW3PF
HB8fjdMSHGR2Qch5+CHJ1aCpbyBDfRZRk4zrFO4smpGSJhm7dVzKgGHAzD/4wlqBg15s3rwJuNZb
ZXkZDA3hSIu9YIdWTkMDTw8Y2M33NMh8AU76BKqfD741WvNCQyLUBeH9nOeT8D/XxJ9cmMzxKw8H
ahCG4vTw7O4Z28VLPpP8A138t4+LsXWYkVPlV9YIMKFF9y6/Xgdu2OkipJmrrc1Ah3G5N0jR09ZA
m3QqKn9jv7LWw9SL8+ZZD4j/2q2tWis1pfCy+qsudaTnVvUhD7Y50cuHDuJNuSTYbZnGykUu2RpK
EMEqa0vIHpD2kaYSPIMXy5bv1yKCgXUmbsFc6rOViec9Oz35BW1w56kVHRMilgEXYryKGRo8IqKS
UagkzQajIClFD3D+MA0gkER3BLeYeKsZyWfZJOFNFJc2K8V/VWJBRYYYELqlpaJa59ISaO7F6Q7U
sJgcvR0Hqsb5WXan+InK3B1AN1qhFV+rB009IW6dei3cgYmSi8NF6va88urNTHUTVtUm+2BYErWs
liQjjNkj+no9gkZvfDE28/A+4pBlQbZChZ2tLA2/tliaOgs3jNwXjnUGE4Afr5zeN76lqknsHODI
N0fZKYh7vVQ41RY7xmJkMkKM9XrPuylRUgJHNCRzBhSjCXFyXeTTWfvH0+QNdwEIxBHwwC57o9KN
00/u/cb545PTd62HzHmB+i9rqIP4auekRMJ52pfXPDA4GpEE6AdBucSedF6hQpBUdhfRVFEinm+o
HMYYk6sEV8GPYoRRu1OFmUpYZJkFm700mb4dUtCm9N8+Lar51q7k7k/7e6v70wEFd6sB0SA8cVr3
ga0xhgM4HniwuVDBKQqu9WRCF8XCureZP8aWXxqDO3qExmUqGLWOQ8EUyNsWp/X90rI2FF93H3Nz
MLw1YNh6CbdEMClsSgAtz2SPe2BETyVe2BJ/qHIZ08xTWvn0y7cTgUBuiRSPlah8zEFUuOLWFOu8
9Im5wzwoSz8W5kTwYLLvpRMj/H9iSAxE4mT7a/+px9Jyn6jdmmeY+T4cmDQbwncY3LrLpJ3pjHCE
CvlQVLrVqNbJ2Mv9vGsjdXMxzqxVFzvF2kIxkYnGGVIxW1/d3a7SDNjp7yg41TeZeBVAXA61F8Ja
2KweYC5C30KDDfPnoMEvH1eTbJESX6lgI5uhsqltlYI7Q89uNcMa2O8/z18XRNnHkOhdMbu1kre/
DTkhwUjfKw0brCW5daPuyEq50F2GllqZJfMPM9PHBGqctFtpfwYniw0YhRAnE6sG63pg5D8WPnmN
M732T/hPPf9jtEQVEnuf+3kjTtGLMMsvuRpAU8ylyMWiP6n5YTkBCwxZ561QJdBNtitnrCfdrOBF
9Img8hlq/UdMHRFGu+1XHedaUbKMTMACgOLqaoD46UAYdxo9mooSLiZxWpqmvrvH0Twt+Rk0iVsq
GVpZbUxFjspBuWSIzX6sIofYAKI7AqwJSqRJv8W088MCI75DJ3FzpciJfYs9r9fz8Aoza1g6UnFW
Be8RFbtNSk3IrN1fRtohwlBdLyEE8CZJIh6O768GtcvCH3u56gHTqkUkhotnrP3f9YJrvcg+Z2LP
rpkQGvyNrbb6KVv1hABC+gsMM0/BBqoE7Q86BdgxIpnb658GtTTINc6b67u5zscR5qGxH8RtmcIn
fsN4CUgStcb6rPT2AGJneOF0/O+LoHTZkR1qFtnwN64rPL+lFIJHuZCsSZ+KwoOS23HF27JG2S9c
shs//1e0PgjXhIz/k5NPP+t6qOGIoJXiHmuZPcLwCvZbw11/j9z0Y2Zl69eR8T1ZwIK2G8EQxHFj
4/Zm2qPhXrtpOLd5VyItrFd4F1OfKL2d5+0HSP/obMYP/pxRNYHmqvYXoZhTr7pxNG4DHIurTuk4
6r2A61MSWTbgmvDie3B1xwgLFQcSGROHxDdm7WEozKIkvpVpwJ1tHlbyOOL0VXGV38pRC0G0x2S0
fjGn7qZv4ZF+WcxxP5jcURtf+Us/wtxFrpBB0H/I9DThiiEDa2AXAJt7aGpDEpIS5HvKEVJ6k47t
izsARvSQaHLhN25q2sO+73ppZ5aDKMWYo9AtRkc89KJoddCZ8o8dtN6uYAX6P+bZbJTUoO+WZeGT
ziMVCb0gP6ZGK5TFGjgt4PPnXwGREsJ2EivA/JZnXUJelkjWQ/KqDlh75UUeP92FaRUQvrTsFEnh
EzApPQhkVG48hV9VEDZbJiyJrJuZwAbPonz8DMw5oywdbYUpsNI9LGlVSpsYmA8NMAwDzgmcGJku
nvn0p4FbzLDBfC0Zqm0i+SGV1DWc3BVWo74W8pqlINqQy5F2ZWgE1hgtIm7idZsxyCdpVXxAeT94
U4vYq7InLwp4k9pDzOnV+mjFSBbCVi1qS6E4NkvpNUGuDlHQZUNRjxOgZNB66oDvyxH502N+Dkn2
RN8bcUukV4yVrB9rWSaLEa/Xsy0MXz3ry4iQcdpd+50VPv8npmLyn/tlVIdWzWPgWwd49Xg9b8sm
2v0Zt2DP+cVkQvD76IF0mDggwxj320mmnbqVci37mpTj61X2isK4VAGHU2AtEWJTK1NZIaRomRxu
oZ7e3S1CuOUl/+qjosLvFWvsr5yCSOPl5Sa1RXqUpVTb340SwRRllVrrRxYHmFrQZZzo/k8bA5gV
4QMOf1OwpXR1YJ/qF0GSIwB2ueW046k4AwJJjAVZbCT3S7+3WzClmaCczXOvTESruI18/ko+m787
wlce/OKqLm1Nkgc/iasRyq+Ja34wfqFrQOiLSGLvD2LnAp/jdY4z02k18DbHPXNadlGf2cv+XGqg
5tQgD84nG1Ftkonxv7BF0fyCmTFVPwRR6lEbpETlQNBLuVPU0SYddBh9uYYZraAN7SBQI5ONesD4
VQz+2po9GKOoqP9jTm+XcY0WECrEihjlDbo1yeMyfIjsG7gxWFWZbV9EM8pnntxdWO5M+5u394Iv
yt8MUGQl3NOoINjjPIk41V5aY2KingG5uSCgc6hqOXtX64gbWWqsrn33NUV3YtZpmlMI9LCkPR8Y
+tdGJ+dN6JAH4Gb2/euoTuX0BQi7HHFeEA6wmoN79CAXjrbRJfiuRihcrjHfpmx6OZUspHq3nkGX
n/t9AL8orTKaHPg2YKElGTLTEX7X9xVEFar1uK2+dGsAcj7yhBO1k/4c/A6ZQ9Z++xsjAQApx02Z
BfGURGXeeYx81VHteif3o83IYvKaDubJ14llaVrGsAJSsL6hryuWdstA5ZAooPErc2Q/NsY95Vf9
6sK65JgPG4vN86wRNLWVQJ1wMNXKtgMG2/UEUuXQJLSHC3Vr2PjHzFhcdBGxe+7z/GT4Scp1FUU0
/15uH8/0CFTX0E6u1EWR3d1ZfReNHN5jhlu3a7plSoubRwa/3+ggKuBCeeu0gup5CQ0aR0My3Onk
jP7DYsV4XxfOhaSPYoCoEi2be6PpuiuZck/21pprbt3Efr638Cf9SFZD5x+nz7efK/IrtNWSqnSy
hQrDpp5RIkFc25KrIvLVBPqSC2YtOhPNujIn7vuBKCZYRih5ESnPTUMvAYrOS1dmQSgheEO73Zz7
VA0aw420AYEehbneYJTnqZKKOxTONfHPNEIEC90LIW6om8QO480EWuiuqkLBa88QTetn6Y3eHGyV
Uh53B00VjunX7rktYDnwCH5S/U8AVrOyCk9kTtlUpRhjiGVckeGMBwjpRNNytLKWbn7lxfCFB4bz
AnSnHP9ng4NOicV2FcnOu7769eq0H5QvqnDDzoPe3p/x/sJtE+Om5ssl0UoBP7IJDD+XiCXXK+Of
d10eYh6er8MZdTOuqf7QKMxDVNJfhrEb0mzPQxZTn49Vw7yaxIUmYg67gOLWawWWGQ3bNLlf57vV
rSApk6B+GPDCJ1dq2izg0l4GIEUo75pXWPlXa5qhmH2NFtGb3OtX/1EFY+CS0N3ER1JDB2/emHg5
eaF8IanYIHy1yhLRUN3AJFhVy5N5k9gEBtjOat/+ipBp1HM9ZcTh0Amh/Vxgiz7VbUFZtI8os/66
AQlI+tPpwCl4ecSpQZEmOIdSbnJmHl2ItMaE4kqY/qg+QDRzEm+xAiXfkkqDBxn4ybXDve6h83Gq
oC5E2tdL5T3jZ0rGo9lo9lD1utS/7/QngJ23Jt3Hurg5pPWvhgHrycH4ZmrgjOBDMRt3CcM4mHez
aVDs/vsG4eMGev2zl3DjAoU7DHlAQ5NkCjE8Xo1F05GJajFrvdzUl2hWPjCc7SAeiUsKb6+6gi8v
dLlRNAayCXnYn0cq0jMDAYvAwWoh08HrDb/boeam+nid/dyrvv2UlbOjGkVY1oojWi+nuYSLGKf+
6h2lUXeYuAvzVD+JVzMNkBDK6QWdCSHeFftL3YfQX5XLQpRs16cSJqd7A2jGZiECbSXOyjY5qPMT
EPFDHYr4ovVoru//iRPVCDZosahL9zxt5m8xGb72X0ZSssEimygFGFYa/Uu8LJcEvs6sOFYMsRy+
EkoF1I9krPPpI/UmwOzve7cv4s4kvgCWACv9Nv1qrM54ozu5ZgwQ2oDDt/pRLbVRdCj9mbBZjPcx
Chr3MHbsG1OxmaibgkLosFW0zrx1k99vLhtrCDLg8WOYZBZ4ThSp19Za2oDa8L3X7PWRF8g8X7bS
bxXZGl7khWuA41bbkoJwEK5SuNLgNiKkHhe0LmJ+mbvZ+qSw4q0cAVbnXG4bMXghgysZ0q8oTpZJ
bJca3TfJDhX6L8cWJ2AniKZWAt3VZ72kl7zbKCx/3C0irMjHp9BfoB0KKXVyyK6QlmumQID3+Saf
gRHbIwc9Cdd6Wvd2wh3LXZVmm/tJybGQ8CL/ymp9Nkytx7ukyFPeONyETbUg92Fa5qxi1TipqFRP
IY6C3AGtIwDfoReEsYf3ApIQ0mx/Uc579tLUOfViFp/b8OcwgRjrp7xspN5n6KxlH/L5Up2nwru3
hS8ZCQSXaCQWvyvu7VijXAOdY2ADdfFfYPvQXht4x9nfrSnmakUPjCfGnjw1FMqd9prwLAcNZFMY
hhF5QC6Mc9ptEC2Osw2P189K7GhcRi+m03fndjdzMdteRo7EFBsFaNXCnOSLKtCGlHZoVRX4QiTB
39Oq4K00R06d14PjhlCPeSeu9ZrAM5r1VBkjUtmAPGV9q2kkpEZL1n6u9hMe78B+5dtZsSXZx1Fg
pACFm62UVv0dAZl/chcIYhh1eHA9LpDyMq4N5mwoHnktlzmYTKA73lCTC61SQnW4TFTiRng1Si8J
p70ri4n1WFaXJuuUqoQo0NQ4yb5OlNua/AwJEyJESo8k0S1/QYQ3VHl1nb3KBRsSPeFgUraBCP/X
pQNilpxE0iFLF1zQMxn2pnYve+ey8rXGEviB206Nro/1PSZm+Fdw2tk8qQ/8dcsTrsBkBdKPaWLT
FQFB11yw83JCqNlz/eQH/OFuIeifuuQnFHFhD/LbsUFbMIBEg1nn+1/rswDWkUkSuYOAdo1dDBiC
qrN1kODsnArizs+jLEZGRuPHr/A+5p4frE+tTjkj/HyF5FiSYWWYMK96LpwLy4WjR+daHYfowGUR
Qt3f8ILmN0iOAsM/KHAWFWE5Y1rQ+rVO+Py2t+42BpOsZDN7u6f1B/1El8W2IXZEQnbG9abQrXTv
EFYE4fMad0M+Z6Jil6vr3umBTdIDrCwIVY9dDtO2p7h/VYkYb8jZvKQD4RGw4X4aUvDysVq5uear
09XWXVOdbZ6C413j9XbhTBWI5UcDSwAehGOLZGL7j1F0qSiLOj3FDd1i18mVThCemUaMF0/73V8P
sO/NPjZSRDQWyz5D1nzvFEltpPyGoRr+EeJ7eH4h6E6VSUrajPz9100pFT2QKZFvXGKuBAewzNX9
mO79K1/kQkpcDHbOWb66KmfE16QeiCeeSudqe9wV+ZAsXSTAImxamLPPI9Lukk0MCrAmhzFB3ePv
xfIG34X979x8E3TE9NuFB1EjMUl+ZGzsgS44YyAY77c9vb73oHiyjbIXJyywmvceZoKhO7r1sg7C
Wla2FmcXIJLb+2wwEPCmuqfRGp+BkGaNSRBye6NDALI5a7Wl7QBAIp66qZEjAtqjwGg0pNOiCdUy
MLhQGJPeCm8Sbzs7qLXhDDzof6JwvZI/R2h2bXb8gTgOwAxyIX4H61FMjuFRCaPgepfb7BpcSSpr
B5EVXq3hgS8OoL69PYIPrjsTkeQ82XDfMvFp01+wrgvJUGB+gV3dmVjdw3H0G2KQFHSIRVGR5WiB
PG1FEDdGe2rRnef7QAXkitjyI3oQQy3/Tm/SWM4FrXVY7fGSrV/sXxfMqw4bC3o8nkhh0/8xPtyA
IiLzZqb7vk3dEBzR2XvKC1fyDrIgmCOf2x/PpnUCm24fvHj608UKRYqDvgsdramu/7wvjOmxCo8m
n6i4XYkNGjuhbe0p97sg+NT3ljdjSbjiZrSkD1wNIHtc+8v7+0NS/VgbIBykWEysJalnk5vb7Dv8
JK0h913S+Ot9QlTjNxa5fDDYxgfFRD92F4qak4TMQNdz68f5Ntd2oR3ytU0nc6ThMwK4wXQP6107
GKOPuEplePaNKxntpFI3KtPvE/+evH8U9DmmZR/1MYexCqJBh6QkMai/3U0a3/SDGqTgo4gu7P7N
UcQFSz9Iq32V1kzTLD6tb+BbDwDZ+H56wTBFUNLbCt6wCZN2Iq0KyY3vSaSpEw2ILAqV4/H3LvKP
8Ba03Fj2/teIf5aDJ5gAHRwSA1hBoihDFpdmmoKiRhXxPIkxZfQj4z5G8Kc4e0gGYwRMnyYYmip9
p1RRZGvEO2VJuBl7nb4I8/fivYvo8k+ZQvp1uyw6vF9LKcdrj6mP/cggL863BNDlknJ1Qqc3Oy/n
0JUAT4KXy96rozAQMuwDIyKrOJ8KcOUaOR3grHBmURElwj4Pbh08eQqwhyHcIZBWYG4oxbVS1zN1
//UZJcEEnZtTeoaP+3xIVl3eVQRtHssnb9ogxMHL3khugRyRMXUG90eYdHeY3c7Au8n/O00ohgEf
bPt/z6XIQ2SCKzgMBAIaCXISSb8eHUk7mhgKVYFblD83uasVojAPIMjBfmGHiU/mz7xJ94UsPXrv
2G437mVKhyuqqZs81HIF6V4gVdjmt6QYV+ykE6WMwNcAzZG6xtpWlTyQzKmPQX3oLSUyQ7NLdNTW
TU4gY2soHdSK/O7vnaNtgeJONalHT6i/SIQFd7QyTGH7LxTIMNXrZ5rXAN4k4QhfOOG8juw3bb8G
FezLvGdlitfXCAl8s1CzuRBhf1Vt+w+bF2j3VAiqw2HA3qqbe9NwEhN3rBvR3jr61ZoKRtgGL7A7
B4qLSCdNaOkk4RBJkzHdfUSdyKPBJY5TMPkctg9OgqqsLeGN/IOgAFbpiem7qS3ZujejuEo17Eee
dipolmN9maJyL5l9eJidDgxZg2NxZNb3VawVHh61AX0TXTxySRh0M6kVp/S5MGQE0cCToRL5RTiN
FEnP/D/i1o/cz6n3B470+iJwk90DWO8UCfPKmbBYXhjoLXnTcWSdaH53gnOib1AsR11abflFmaTI
C727RTFTrhCDusYMeUMFp0CGQ5l9dCv2kwv5tPc1UZafn6KAXsdnaNmQcV0u/TyIYul6tZN5nOXW
g6UJFX0SMeNWOyvX/4psb593+IOOW+OSRtoG0gNalt45uDsfDn+hCPrlWfO/E+s2Lble95N8NL4o
U2z/QCIu0+PQjbhSfGgEtOhGUrN79UlWipnt/7J8wbRQd3xzcOZdQw8VeUznCOVJaeKTHF2sf4mc
AtSsi+yymPr0XOfdQj1/az2tP2Encm4GZm6qDh9UtN9YCzCPDwVTxWIO80bajzr2yZWGNwhsVn/C
MtxHmLhlg/SC6gZxNcptd9LCor/JoXCc+2yz/EHphURSP+lZNdEq86tkOCO/HdtgUF+H6Ah1J4sY
ak2c6Zzu9+lPYH/Rt+5bOb5nKI2tXI2n5MwzmbZpaj9cKAIgHbkDbeN5dZ3loTS+8gJMN6WZWMxc
LEhEVKwS5yOThJ57khBFht4QYXenZN7HK+0GuRGPZTt1i5dxKxyEafguAcOKfSsKYrO2gbSf95ag
Of8ImzKQUfvuQgFvngH9COneQsbLu1afpfNEsYDTeB3/6IAHOxfCgqf7ndRX295p5o4l+L2k7eUB
5ZcUPeqIChoKxJ8i8QJdtBSdUcN8FG124AA36DBHg5669h+3AjguA+wZt2+mfoZOE301zcpcQI/9
f33Qy97WIsMu4PhJh/b3wHErYIjqixRcy9k4Fxz6lZHDYnaTKmVn9a6zcmPW5hcFbGESBPGCtBFU
ZFgvXEkh27YWJxPo7wicn/T9dUKczHt2gx+XYPnDGSiX4M1xaijVhY/Vd8xpT0dGu++x8fQ/ld1n
633rrhSAwOIN70hvmIal1BOh4lfqg80urxIdKpOePczedKa/e4Tjo/u8/lc+0mWoUAemTgr6ZRd/
+qMdmYBhsblX4yf+lLP6krDOeyZLW+uPSfVmrtO5k0UKaYUQz0PFKMnsYCI0+FxiQBa/bZrIdnI/
oU1wKFmfSKBxAw+/7pwtU3jE8PBxiqlHB3vrO6RjWoZ3CrGJGx+dg5YbWxJ7Xum+I2al9dzsjWYY
3Nl8DplKQx1k0in6ioajEsbWVhaMbhxXOxyPRxkLtF4/oYNb9xhziF643C4pulo7dgmSBJbGwdU3
HXTjAI1eCkG6TO1wI8btnicVZl20jZsro0b3uG1brIWshUJk/gPfj5tNz38O3fgU0q/wlJUKn/0C
VYrDB3+YRN3uwg8Fd/MVmdXt3+30OuJMeq+j3dPFKoe3Q0ISjXRYDyaDQvp60VigFdyhXU72Dhsb
Z0GObOvZv0vdeiatfxObgMI+vv3zEvyCbApWduf2muWW2RS9hto2hySXwZHiolM2Z0f2kEO87k6v
yiXZGvrZ39KgHT7ZeLKUTRvYinEYXozZzzjHOJdUO+k5Z3UlgXZZQc0a77TONf2aorCkd4nb49F8
H/3FAELSB8lJd/SXy8uQprcYYBgVspJ74Sb6elmJ3Dysi+H6AgmSvULta8FuN1TLkiALhqkgdh6D
NrQSxQTB0ctMeC29+f2CXiBuJD76bWst5/w9youV0pvTuYRqf1dbEfuG5gkwVLiJIOqB4aehI8R4
q0R9dJwr5BWPs3chZPGGDQ51sV8Je/G61IyW/GayU9zuqTI6ZvgCC3B1xaI5IZPkWUJ/NaiktOhy
0Zpyjhy2K0WTlS6yyxbI3+ReY0s3m+2Jv+pN4+1fMR3GEp7WZmyF+iM+V0JQdxg/YFeiNCSbEtlS
5AHHkIpK4meVfUIHz8ud2+enxMGH9yainUigNU62CzvDt3+FTR7MY3Z91UdFIuFZNVvfOib8GYBR
qgs7MKwhMlv7E6GnnRaxW5mn9ewh3ZpDiiPxMyTHZH/vNAtJORmhBEJRsXwbcvF94IOqNGF4U7y4
erdg93LUycmJXVtA/pWSEDD9RxytltN6Ew/mLRlXOlWGs8uEb6eF+OjJJpx45XKJgeDL3OtrjULh
37VOKcKoXuWZMaHEnVFOL6rIvHElGkDK1VE4mwh+rR31U5FH2MPuNiteb+upT2tiev6FvBnoQENP
ftC/yO5vuZeEr45l0WN0TtJtkqgbdHhf7IAIgvvNOawkjgk7U0fswtFQTUW6oqwN00z55Z42eSQT
sx/9iNXm2gfGcyLa34PTIAt/+6Hs2nSBX2dGEYbTGzK1Xl6FgWSKmD5fJ1ZX1MnZgQS3bCuPwpv+
ayXZb6JwCR8BGgK4sAKv27aYFHD5i9V1WzPmu6HpSMxfPpBgPCBWc6efcgmVagikGl0lUZ3XJKVo
yJdOjr6N+Wqy+axQwgOzJQf6g4DIpIcDRm1mbobbWZT1aChVgiKcs+1VgvIb4j5Fuw92j+kREwrp
J+eoExuj4QqtbHXOlUjQSuZSx2azWVwkXb8FGC4tkvIVPqrPFO3NQxnBh/s1I4uzXgNRLIYV6WpZ
RpIBlXaAMKzpPdXASltGW/ZG71aoXRdhipy/JJ0wmWKZTR1y/6NRb8t5mQDUnTTJ2SEBVlYT5vx/
6lIJOzXmYlccuhw3I7C3LVSFFdmlmfWkhM2bxox1o3ZbffofQadvDTkKSTIZ6ncnENj7dLf7uMhH
BCVuCV33GPjRYTMb+8IBF9PNo8sWnkTJmKTJ7TZ/7AfOd1Mx7hlJqZj+avPpIw0N+lw42oy2g+pf
klPt6hqjZ3hcTe9yhX2ADtFQ/M8YfceWRgVpJR4DMzycN+dlzIF203Bw9AGUmJGJroLJq+BE/gko
n5kc/X5FCgkVB99U23Cse37Hh6FCuoJJFXALx4Q1cazcIPNqmrlD869Buvrs6f0jJogT8WLwRD77
KdKVt+Wp6poIJyBNNIGoZdb5sIWGXDakvYikrYdOzb+3Q2fYow/A0pYAi0prFQB9LXa18FJ4VDnu
uXlzyJWREYF6+hU9tzMFzyLLrwneA5RdeoNMNLlpgdkOXNYg9jzRGCxcBJpuxwFSY2sXAtTU2MHF
5t3V8Djv90GX+nZ25aK18T6NlXTQVNrOb5OX56UxUGYQrPe0JFWCHO6zLbaFzTFRQoCziU+ihXC1
rKpRjZn29Bf3h9jkMI82oAJKfy1eDMPjPsnBgiHHEoIjvoAZCehcIcIC8/oCUQilPg7GDyUbaIPg
wIvZ2EF5N7AlliFaYgBzixnIsg9jOkziLoFzOo6zHcUYjk86FTt87D8nTIJ5Lv2mLixd6KfVJlsW
9Z5+Mtnr/IFHq0eKwV4OtvgMqJGkVWem9Oem5LtWKIPKGT71aGaOM8ke2/fw8OspOqK1bVAZJVsZ
y9A8QjV0UU1UVcFRmRzN3N80n8FRPnUOXixaGGvdOWNC5sQJAHUhVyzcKdhso3QlCALV8in53y07
O37/f2ktMkK9SnU5sbrADPUg1jCnjdvsP7DW6ZP6JIyfE7qEHpfWluL2Yoeee7m84e6QWEEBepY6
zaxGT3nI0KcI7jrNxm+aN0qEn6ySlEtKWu5MvWvFgu1AGVwlhk0fDLHeKOZ2Q7IJjw5YbsbjdQ+U
vbe2CHQzVcvs5AVaexOYtPIROdCNyRBN6+UjDTvIzg7izFD6adQgqN85sFcK5TeXL3WE787QTMl+
3ok+1CfYPR1fb/3+hcA6aWow4f6Pna2sfJrLtcFJtHSuUiTDi2YPFn1M5fh6NvdELDw11EvnMx35
SJUzaWiBvkZFwT4oBAxRzaTZY8Ze1pB93SnmQV2VhVQltuR0lvE7UemfrLrH7zlMpoP3sNQfUoqu
w/hZqwdsOJUBDvMVTeOuYUhLcgfG592MwYC7BXqfJitftuu+Zs4RUYPrvSXuLbwts+dKeoF4SU7t
4fAgBZ2wFDAvL/iy29ldpm/NN+m+KTmHDnFHu++ZMtHTtBXpRDI3W/7xwuHET+w4yUvM+RCVCPlP
Tpq36Rwn5YJk2uC0+KKLOKnKriyXP6T1vNvqyfEtFgddXCXNL4cK6nZKX65FDbS8HmQftvfqsHdc
uNhfYADJ5nLoPLgVAyAabMNTrkBy+3H59qZ6i1eYBEKigDYEMZl1vjOndbkx4hqZCZUyZKTQB4MG
subKA1xirM4CLI8me1ZtjtYKXkeWyqDTLrFVYD52g53XIvtZFv2ZTnEq0H+5bHaOEEyat9JFMLt+
+SoRvjXzoBwUQvXYoCi7zvxRJ4aKQ1KjzrWDd8srj/nhheIu4ebLWcpGOalFaOaXu3v7mzJn8jOX
sOn5LrQvbBoGGEZcZ5kLwX1KSQ1IXMfmw3YL56FLNQ9Mhiymp6Djk/+fOCqJUF67u6BaEISzWOr6
6S6E9mfG5Lj0X4NKFnBLCvsDEO5LB0z7y0b8HxvL9NBiJRN7eJnI2F+Hh9nZC1V5jbIkArSZuoex
UDTw6nyWn3C8o46mZ9ZI+U26EJgYp7WbO/4XO2eWR9IY4sKVR5spK4exCHHR2xBiDkORxFS42u5n
7qfT6GZLLVkdn2YCnT/5B8IIEpN7WtDko8ikRMZt7ft1ylg69U/yaX+d0PIgn4N2rL4IO8QN8EVx
osKXj35VKJc1f1JFQ6kOymFqA855H54I1jav8Zl/87V4/1e4Ts7rlCB3QTLouJS7mfj4vlf0JwLm
BEw+CgC7IvYnl2RJvLJpw/pl62XFvAhJvf9M7rLiEgFQBKdolRuP+M560PWly1APuYGD8AsTnP3u
U22tfywSE3yy3NdvEB0SgyUBzEJzQPtzZToQ3qTTOF1xk6dDS6Sc9YDvte8g4NPh7a0KiJ/v5jK2
jJ9bQ/vY2Tup9CFZpmNwtpm81RX+ZGFt6uv/33PiwjKHiIhZXrg9k10PygGDKR2ebTgmMi7Y1i+h
PnPDFbfrMHAHIUe0mgoWgHNhF7dzPSdgyNdkT8kVyafXt+TMUxQoFV2rZ3xMB1AlUlAhgutFGVbY
Hln2ECOHT1ywb1Xl8KVAiZV6JDiRcbSLnqiQQ2+BPuCl1peZ4e7AiXhnwOF1eBdw2PmFX/EfIchh
ElMf5CHAx3/Euxc8wlqKDGbx5NivncOcGmJOeATeNO6L9flhHemPWxtVUKwA2/J1Rv30y45zN+T3
MajmEkfGwr6D54nVf8kXx/4pq8M8+S1MwZEREWqiR8ZJO6VHMwgoWzzxwzV4YPEfmcQTqCjh87SB
kmlHsFM7+wQAohO5VyNj47vlQuH2eKKMcfigib8SF5/qhtCcmGiWhQSbyOsK0LKyfT5GHSKZHPia
EXTTPDUEvyuyIX5KQTxsJtXY/CMNucF92D/HTdcPTUCA28g9XwcePdYNyQu0t9022+lOpnExVDm2
V/2SymO7H3KO4Q5eYCypCF7S5o8vMzHgaZW6tv+6YjvPJqm5QnRe2x8wtvYn+ene+jQSa66GutIH
tvISp9nWmoBP5HCjN94kXKC2PrlW/dHk2iA8hRuha0YcshwnUn+5or/KgjkYrCfCT/v5u3pr1OP0
k1V4Pmu8tmVDqXK1cfA9hyFUtUXzF+CMyKcjMuPqj1bCY6NrIEHbDdjIXPwyNzzEltnnhZZTqABD
UoDUSESfRksKXKcMS/jHJIuwBk2V1cqRBmreAIl7avhZ8JCiQI6FnrT5zZGTaBpHnNzHzec9yzt1
/yl/Rnv70L1qESGIYIPAPjZWAjs2ntwwYSR6vKhYSt48LwiiH0CtR0mVSmQnB68ODuwTRSVu5q3v
DG7yZNWQYLLOd7jbW4bwFOjIypuHgOtMzKPWvotnY8yp8PAERgVd+2roERltzq1JuHISyaEj+eRs
Qoq/Mu5TwU9bUq6KRnTRaIVu7ZRp0E7ShLUqMccSRklAiP0GK2h/404rbv4Nlk9KFzDtcODzesLg
koszt73uphdZWB+cqcCejSvlUoyVf3wDXLTxCxnovDlww87CJhoaMygU+OfLEJxN7+HipHCpmQMb
z7WtJAYvoii7MiOFjvEodL1xJ50BhxqaLnVJiEje+MtP7hJBjvGeOIvdb16crGVjUEy7G7bN7dfs
vOI9E7tNXXqb0IorcH0lf+rN8VGldPW2BkW1P3Ll9ZQGmimcsjOIGruyaef/oWpwRzCpueWpzBtB
ndGEhoHRnkXGcPFc3YxuIiP/pKDvmCSczQNAR765d46uXWPuDHFopujcJFWqtlemQNQS9H8gnoxm
Wh/koI4h/BqfRDqlb6nJ1sLEDpokEuaSYkOj94oy5nRXGgDIpYiXd+/7ntE7MnVMIPbCcnm1mlwe
B3Vcv6jP7GQJyxdV/1e80G82sen66mF9DL26rhqUsGpO0Iy/wSnjIgDVLSYET8xtTQUqjESuYd9t
Z231aQYrq3l9DqItZ7+EQgmgCLURkhN2GLf42XY95G81oy7lJbdMj2YiSzmkFqDsYjEZtWOZ23xG
7r/MzYFURppLkSqTNTkYYoF4ubKtmeOL10GOX1fWZJLnvsTQ1VCFtvhTsERF2dRRTQIp6N+Ro5Xh
ppl0XD4Z3W2Wugdn2cdKrJVXc69mstIY+ai3VTJ93Ndd7BmiMwPkzSN/ebj2FI+gVnGWzG1yQbXu
+cjvfV3hRNGLMXI7L/6EoqNLPTtTVIvn4FO7Z3AilUTpCcDBhY4rVz3vMRq5Aiz2pvgTZVaMKY0m
3DhTWD77u0gBUgzvSc8BIz67gIrmYu8tgoaDpE7/7IMKGhf2iGTBxE2tl5fZOTCUBaLrJNyxtfqr
x76lxh29ePiUkeI3PGU1gzCCDr+d/RsbNCMlACdyAHQ5TY5mzQniZFDXiyPSQJzZS+3gBAG8aPjy
CKLvmrLkf+2E78mNh6K17c8qysLQQ2mBrOEs6PDknlOseYi37AuTjW5EEMJP1EN7vU9zSWdVF8bv
FMrO7NEtM/XDxdvWKuXL8k/UXamUNQUoHHOBGXWpQsopuOK26Z4E+/VmXp2KGjgnWUXXIKeiLS/O
CCHM4FlmqeNbU/hTOZ+0vz/D9x7kXXGY8PpyBkT3qqGoT4pXqrJCclMqAYLeXTi1IydUyp8ixZGk
ljlV4dedza8oQu7/C/AAsK98UkfubSz8Js6pTx78Y6pIzi2lrk7TgdyX7DcG9mcaO1X8bycuFYES
IK9kkrRuosOtanAm12kIezaq8CLXs/BGOu20tLd1S5agTH4GWioRk9Rlg1M8ouNje9gnLxvquW5h
e2eYFzjablz/3BcG51UCJN0amzXT2Cr2SwQWevZgJSV3A6w+Lf8/vENMC1f0QFmeJuMQURhrIUNv
aSY/ZgYivF4CcBQGwVuSbYM6kooYr1c99KpOdLQ/u2hqL6oQbaZ9GM2lr5Dne2s/JWXF2vxK8/z+
3RiQSHgR8miAhiBHmo8SccM9nr94cVo6k0nOOk82uVpMJTsbw0mfU89YPbZtShXxSiQJHzttPf+2
OgdaDAVCaPkRF0qI+Po/Nr4Z6oZReF8vWDeSLS2a3x6CpkqxMKlkJW6Xr6K2nsL8cUGFByhQ3NRp
RYBeSR2KzUS6upGuvWoPCpxEXMqwefx6LnbvIlS6lcVCXoTspn9f7ZAJDDPPpLOtjmoqLNV4XCln
hM5C2Ah6PvUk4yv69Mo8xsAnPbavW5KBlJ06oA0hhkm2/hVj7UeBD/3hepRQzpaUPwHPJhFyQQIw
3yTyO0VhU8GEGUqvvUGsVU5ARhNzal3lI8HRchG08kMYgor/u98NwSpo+/3gD4bS72MDawpDj0ye
Tv5IjkfOwF956IEnMyTGm4PdSC5fDcVg1ofQKMo0AYsFJwewZ4HsrEuHnNB4Nk0XJnzh1+be9kk4
APKytzt6BrK7iP891YTgLWtbFyfxT4S2jjFHpqUMC+lQgLjkz7k10nmwMbk8LDyy8Xp2wg+jkPa+
w4M+l5LWiRYnQb5ghhEWS8XRi26He1mURozHqtz+J6kPOybVZ290Ft3c1JqmJs4I7eGNE+faxaCP
ik4rSNGlAeavy+MMTLjkHKRNeZK0uIZ5FaN9Gig5djpqRWLa+jCY5tiEG2DiBPG8fPnykwrYZsYX
SMLeoEA+KlLb12/dL4vwL2PBbta2Nc+vl52FbR0fuqdjSjwqFROWtxD5woSkoMKCalayvxIUTxNP
FO7bhA7mojR8Vl5k0L6byRBvkRNX1jR+OSLf+6FZ0hltgNtndcYNSz7LKBZbNvvICh35pbH9wO4A
vfEWxx15kmbZSU1enLc9xkDjDbw9vt9/fO7UgzCDGRPEWzhEdipFfJ8WDqJvv/ebVhnH/1ircW/Z
hGI7RzR72rxC6q1PuVj/47TrRsBu59gsxZG/95kG86Itf9BJCFnjNrACW1GTDVYEJPjoCcOP/fsA
7EpiwodUUeDuVw7YkPqQ7/MmYzZV/BKHpjUFc/3HPAHpqN8xPeOenlPDc8bjbfHymNi5Ri2D275T
pyuTecl8GRXiO2UOsf6Un6u/Bg67XpQC2w70SJsVE+N3tBOVrbXxUDumYhYmQHFm0NeKi8+d7IlH
mSm29we8SRryIIGKUdZeNmXaeZ+0nwSECcL0qg6h4me9g6zNjBDp6N5OkBRAE0wZ/7id2Id/WLL/
kG/baLBkxXJ37f2BqLGbOj6kHgDoMIdW9dVI9A195GJUhva2w68rYzyJz7F5/vCKHpX4nuHgxlTm
Ou4d27F3ZYx8guP5JjWOZhsmHOU8MO0yAuQ1YkSxGTqMtTp4WI8qbRCk8cyJWIFLudE4++t7zW62
GqG9/aQQush1+MfFwKqDgL+/uEUJZdfNnj2yDAQpwUwF+y32GMYAv1zgY4rNfdYl9/ecljHApR8G
wNsF3DAIZbUI2fVgfacP8e+O5kxIV1JRP6vjiCN1MTjopxV4lDgbOo05N1rtNJmNtJ35S2dIolgW
LOUuv5sH6Pvi57rtHEV8VDj9BhSlMR/37Uc5Kwjnwk6ItUvjTqE8M+fBZs1XIkkAC0CRYFCp2vY0
3NJgMzoWrLVpAilhg/aUiRjKjmP0FEtGKKmIiKnSv2UIKiE9HYOL5xrvDFvb0p1Q0HnEqXh6Jq+a
/elLSBNItHgDzrRjUIbLHSujmikip9bmJ8/ZGI9WL2Kkd5c33EOc6DXejeng7RdNm91Nz3z8ira3
UNsIcyfSxOwBr9RvnSAqjrdmUZmdC1LeNZourE6ABTHZhBHZn+X27yFm3L8/TIbX/y9VcD/2IhL+
679xoIyVXJELDX6KMvmOll/uY1MoF2WVG+vdLAB6mLVTFDbpNcQ/CEvxMuhNHXnozC8C8EuCiWX1
O/qg2n0W2y5oymRL4qA2XIf39FrwrfayjkHUSnMzMuvu3dKO6WONJaYnIeqlnLvUDauC2tJS02F4
LzPHNdlmmqccQ5dNScjxKD8UaSy5pRHAnZH2R0EY2J2sd9gfG12iuqVL7DiJ/aLXET1DJ495COz7
Sw5N7AIccCUGrNX2yv6VQ4/yqyWWwhnKPwX4nkAnXWTZYPP+gK2Jybb7tcqIoa6Q2we+67hbj0v6
lT/N3bgQ0ay9WL4g30KM1tpj5u55ggu+a4sWkUInh3FzdlMvlnzMtbFaGWeRpjQg1UnhHuXeVUQg
Ljui8yUyCud3BT68urEwNyfhYUzUU+SGTCGOjlVIMgyJ9R3mrfmBpr+efJIygKMYnoNbwj12TAAL
MradnK35Wdtaw0OigzZWk3n3NNT6Lw8A1+8w4HUPGg3fKDTeGaP55aZDnv0fV2BjYBJZ6yv+Kssa
KI6Eu5YmGLvGNZbtDEnHFSA3cuutJy1ueDmCeL8fN4af62Hn+iNPypQu2rJU0PTjjWNcDrQPYmpZ
qpK5gtH96BVB9BCDitZyXC89WFN+TFqRv1wB4w35Tcz7KVB46QjCslLlw8Q9MSkwiTpVWAZTEEag
84gURMchBsiHGdKzij0eCEnTzH8TaUFyTYhoQpqYS8whXDkMw5qT2f9FF7jJu459wnnhOP0I79zw
V1kN7W0DwkxSPC35l8/3WWko4xMERZcwBvy50eDbcjW/IvECjMnEqTF1aQchzhox2iVYlW6Cgzuo
SuHh+gb7MBY16IFpP/xooEYJaxgpWhWxUHEBnNydmlTQ3meW9Gr8CbzP4p115a5YubWuSD3AT7qQ
1ucHqlo2jMxRtBsWGI4DOTseuTy01VHjkpTQ+2eZJq/Cszy3wdBRPQ8FCI/6hNaxiTgiOzx81C8/
YWAug1A6nADOljM5WSuHeiOg4SuEsreG2Su6kakfaNyFvarKWFZg2cSmx7d4+EDuP+MjqWo3ffQr
5icoXSVL05nQ9gpXlMAcPpLCJeyca9OnjT3jZCuaCKX2q2YSD+491PIps0NZFdCQHwPvcHvC7fwG
FjpfLba9o1j8XI1zeBV6RQKnai3l5lnjMYSYq3l9/bRchDDZK4qHlihABOgeN4wf2U83ppvXpEiM
7c3tr+3naqhDeBiCzMVmAbAGB1DjaTl/3evZyO6pN1vpqdYyJ9BCKC4sr45rf1VBR6LPe1f5DFCQ
7PM4kTQGUfxNxiWAoaBJ6dM4st9jckkA5amy66m8XdAg8McVK2ZDj0sI5C4tzZdbr5uY/7xZ6ffE
d/k7OU2XSuFxGhIbjm6/RKRCaEPE1t8gtr5RNYYky7ZQx35J3hDib5RSrsOp0v8GMg1UWHF2Z3eq
tFKFnuR4A/mo5GSh5WFhH3fLcnj1TzSqGDhdaKFliAUmYt/RsCqwjos/6OWgkQtUq8YfSaHL8jEC
2OzYHI6vB+MA9AvfQMsjSKyA6z9lobQ42vezBQiCrQ5wt951DLjgfbMlSzsD4lb0er8H3mXXKUwN
4sGD0BbDlMR55PcrtpSz2y4FkokjAVQ5Qj6r2kLSWvaUjriZImnQGLfITsH0RBJIfmDVFRhGcCnz
biFcZWM8a68rfQanUHYJ2owgPz0bXQfrSL38dKoDTuj2EvyVfyVwfLB/49JDL5rpqqsATmZRz/Mu
XqnsDchpb8ahQls3w5MEoB+Jb5wEnQSbTCZgmfkME+4BYM0AslMQl2IuErWj4HM5dkmnd8KkzcDp
l4cvDUWMqrYvWzzopnWxiS3+sgv9EEdNK6QtnYIv4yg0uSodif6V3zQIopf1nDOw6iQ2Qr0z9h01
2sn4bcuenfROanMMVBTkTe7b9AV0t+Te+mlv5Mj+StV/XQ95pNKHp4d9/gjnDEZNGzkmLHlSunXy
1D0lTsFPEEl6PFMOXtF7I+e1TxWiprBXE3gM/Li9nA2WLBPsPCbagn0OarszhXC5ZSlU5NJGiCjK
kNjpE6M6A4lpHKt6OliSM2O8Fs5gCrI475NifIwmcoPYn8+7+YpmVgayuFQov+70bTk4GsrEvByf
LJtel87uEb2bliUMIEvf2SmGMuPnjts+lcCu9f9htpdNsnPL111TP2u6NNavHpLgbMMnT7PtEdnw
Tv9SsVIwnZndOef80uBTFjPciOjqMbzm/FAqBsC0wfU9Cg3LtHoE6coVxmKkBYdED3BNV3nHOj2q
kA61UWK1U4Z5RXXAQmn4A1YDFOn5nYsZZhXrYRPLKji5eN0VX7GclC2vjuU8VraNnvsX1JRMed8H
tcuQzdk0HwtoYqrO9128++TnI8Gj433xZro6FHDudE0oCrHNqDf0MGhpa9WP+DpENSOnREf98YMu
YuYOy1cyTxakRa1SnpP1nI3buj0sb8/UO7aTOSr1e9B9zAw/7rOD97jj9wXLtjKJ+JPW18qzFaRI
JmUVe4+A1t6/yBdD+NxUaLZDwCYrXsKtuw6j04e0tM3ETc0mdas+oMhbZuL+6ahhtN31C2H2Lj51
pd1ohFJC6Z0Ye3raAZgcd80alzxMk/Ui8smMou3QOsF82tNQCG0ajBtTghjuR7Ig1+gopBDv5T60
Ny0xe/4pMiM7UQ5xsF6gmrEj2rNd5+lWPLSYjTKkS4IE7Bu2NVAeRFAnYsFHv2GBQwlvk0kJehP1
bgyKnE0rBFDN7HUTPqV0x9E1JilV/+omvgI3ji7qIzTKlFBg/mbFrSUDrU2ZNHFKbW1EShP/vR/5
S77KHak08vhAWQzhWhHCZdyCdhYNYegK7dEbC4V6TDcBglgl07TmcCrtzbfRIwYoFCJUkPyXWkgy
TGBzpyzazPgX0LKAEI8wng+vRdHRG0OlD+SaewKkIrPCeMatLatnTrbSOrvVLx6NAJDC9W/TnJpG
fqxT4m+kwdlniBilbndhXN/19zFEfL9UM7bDKPvHqUPNAh4UYPGYX4jH0rJv363lLY9kpUJe9dB9
eHzSnlWcMBAfwQfOfBpfcEiXFXDDI8lfiX+IcwHS2wfiU5wFicnGApj2qSEch8LNEDfRw6/+BTRe
9GHkHyzArf6GxFwJGoiCYdXzNjR8EGGpf8bmEa+++n5K1z/tTfa+TWt/1ZBGjybjXS8RxKPa4JOu
400Q6Ai1h6SZ6vStASnSvxzxc88v+pHHix6KP/VW3ZB/bn2AmJSIDbEwRwgwKwS1DwQLLh881Dal
LDmAYxjugLbikY9Tzoiq48ZEW5l1vZ7aqkxh8zfOg5wwbRaDkrbLlT9Kxn9YPo3cr9LPHQdRCf8l
XHpUvvQg3+sX7TXtH95pBy9bMPt7qlAKA1FrvRy4k4d+wSrW+O0diTIPTeL3+uLN4eZ+68AxkQOC
pbm9ZDup31ieTF6k5FetMPTDmAp0uMEbcu2D9flB2+4uJG9sd2aVaKfzrTKC7seDj0J9HquY92yT
+aiOg1SMpNTGidR0cjopG898IGWl/1iCNOhRmWVZPjYkTQtisYXGkBh0QFvhpx+Z2ZcjMgPRHyUU
cRaI+5HU/uvsDQ1OoSonVdRHMHNpRTVxfyYKXdVzU70pStw4nWKD+iTbr3suAsbatvhniFPR8GKY
sRNTL3q+W43feR/qu0ASFpUL/VT5vsO5uumFINZXYZAYjuo+yXbldf+a8uE8e9hL2415NnvhTUSR
Tud/mc2sgXjZsS7L3yBhagYQplK0v9DOpA01Kr/MrVLdaC8GVpSoAEzlRwcAWZ7WWoenJKzOGtA0
gvVPaW/we4xuX3qFGBsS62rwItY/CehmjzZwc64iuzYW7ZeHfUi98a0UmN94TLqS78n0kBCzvP4/
opRQaN1L8E20hVQjNWZMEAHI9NoyFBqbvGVXxAums5fLqyclOlJlxLl+FCCiDxywYDUTsi+XyFpi
P/rW7v+9WjKOUxH2pGBKRqnhMMHd4Pn595L2Tpsuj/vw8RDQ8t8KslKR3b3hmcywfL1jYUCtWAo1
oYDkXhTQ+MZ68ip6LxfvuZgVlPuVhPnH9xyg3X0Tz9WKMU26zoPji2cQosSKEsTWvB01nBhLXEcV
L5NLH+Mo1Z3WBmD/AQqW5Dfuc2Me9Wj91QvJ97GYzDmN46oU/c+d730kaLlsevxrlLawIUItfBZ4
24zGQZV4GLC1uqaobUVELmNKYkWX1DCj0hZ49FNzUQruI/yHnZ1WnUTlcI+EFqCOlCE+Y+fJaf7D
1pUD7BtpAbDnzSAsYZ3xiARJ45NiJrfs/xksLzdac1K6KCGw04eeRxz4nWSICNJsxF7kNFHExUtT
VUGR8yO0irQ4+q0v0/OZUjulus6oQMCJmoy2ZQtx+rt/lzPlUuiSlaHn8ZGQN3I9wRXQ0LmbFynP
fW65SO8cmHSpv+xxVyF0mtOl7Vvxz2XHP5wsTuKUaF+9GFU9cZ/vB0e8eYNQLczvRYBkEY0u49la
Rpmfw2oROEoQsbbi56DSLOeGU6Jf9sHeMPDCVIptcE1U5vyT1rnnR66D+/aKqjXpXPV/PVr3YOjf
64R/22KKI6xWHWSN+BpW5jLVYx4xvnzmqPZNDx7vMb70w0sGRDe4oP4Qv83vIPpUdm20HhwrqMMM
Nvh1tpAdXxGa/DaY3S0AS6lTy7CyZB8Vh+BKlxdAoi9EL4+H3k2BwLRXgCtcdIfeWbwLzVJU6Ql7
4sX/E5Qgf7KSbjg0kkqlMXEvscPmfhETML29xoqxLlCoD2hmiqIUHPNbGzvlvnygH27gCEHBijEn
jjaK3v6OBG0vV9YNG1rlqDXXx6DsvJwIcpeg8q3k7uZLXbIqNtUFrdzADk14GxlB7tM5nKMHmt4p
7SmSf2ZHrdu/h1ouvTObCLR7N9hkL5qX61aU6UtT0sfTraD3/R8EwljnugxWalfm/4lSJ9/Mh7Ph
MjyskVFUBtWKH+kcvdhEXKHrUaafjMqYhOzKGZV4uLnC57MUN4Cr+kvomp1rlH59/xTfjWObjUKq
DQeMzev6Us5MRHIeZFjaY4vAuOcUoL2vWIxCaaSQTm6Dal1fB4mTAztqoTlVbiBTL7vLaBgnPm2m
XccrkeSgXGgrieDyAMJ28CV9m19mHWArR8Q09BHpokj9kHKLM2DxTJWRUonAZrfsuIyjHhtmIg1F
rDjxvkFV65ofnImUuI7MzOBhUzaQyzaeg4n+SLRco6W9o0ZrgYAPk+v6xtoVBE6jSc1r+hmE282A
WgJ5jo9MJO+X00B+ayQa1FUI26PBL/HW6RvV9ZbHcKNs6wLHXugmXmnOk8kAsUO2JNVxzQpB0qEO
p7/I2s2OyQkaBQNi5qBWeU7+Jawjq6OUQHSSNd6zh1rnhLU86+tkDrwE/CyNdInf9CkqihN+DSH2
/g95FXjLN+Wc0OMOqaWb8Xb0jlj8dkvFy+SEZNt7XJumbfqv+UClnmBaNRcY1yXeM8ksPWxW3Z0p
NQMzt5JqwyFG8ezsnvaGrsrc9dOqEtqIeVRI6eO/vTilrR0zIH1JqYfhjnA07hvLzI3DEp8/Y5OY
smoiPW/AtrSJZe20ZStmYkadS327fa4yqXXZmvxSNX3VoFMa8AxCuw3Auj9xocsrfGSz7aKluD92
SU92pQXH2OrMmVTQQxCgVs6BuQPI/JNOaZ13ANZLBEPiP4TKhOtvbegaU8NLJkxVgOslw9MAPqUG
z5lYmDBBUYGjNJKk6ownh8lhpNvtRkmqJJNvu3US9RWBQRhCouUh8xAxmyqz11gI2A/n60HiVAub
hudxoORbQtZgB7ODwgPRBxQ6AjO5atewO8CFt95ic8MqRi20IKXOFi6xRvLK2hdkZTUK4lODSSJs
9lxAgYLtlcFGsujM67d3tAmvsI9Alj1TuJMCa7F5/3W4HVhGUaew+ZSO1u6ZkSyQ5VTnFPtmYH1P
EtTSSMHhvziVopwekS+SMI/mvR3DBO9rDdtM8P3gOk+/MT5iPVqZV2QrHJ++K8CIvU9qOq2BaRdo
9bZNpfM934KNxBlQOVmp11Faj1yzLuweaGS0u+DNNbHmtCgLlIqWs0Ro3mj51fneVJJMsIFwekaS
ZQuiSmdYCDxkEG9xyUCkbTHrNN+Jqqfnqw/6bp47YMKN28B3khC7BfRgxFTor2UTgCswhe67jW6m
DDwQmjeHHLhnae4U3cdl4z37wd6H8ZsMrAncftXeQFtnXbL9e3JEvSp/AwhzHGRHmfgJxxEO5Kpe
9+P/Y5esmcrjdTxLe5T7mzx+bIeP5Hhgoz1N+8hifUBcMaRW2l4MozddC6Dp/I17/XrlFmMTrZ4m
KL4slOZlgubeKrqQ/cJVnTD4XWWBErVaQb7KCIt1HSs3ajiE6lJ3Q43fmLK5NJRKPQ/FHoe0pXhj
7HkNiD3Jrzy0wSKsW8NhuJnE0jH8RBcUthYxyUeqys7Wbcfjr8hz42NsH0FlQAYyx3Br1Fb3HizL
kWcWCfxDyToxDnAcbtFCVIoZxNafpxApUhGQtG+d8qSE2T79my/t5uWfORQ3lK8BkqpKCjzIRggH
/+H8iSyAJQdFLFz7OgwWi77tNGQBUyCQ4DobaEZezr9PCD7969eND5ZmRnZoAB8lE/nl9hmRhexq
XAR8bSxC7Eow7183SHY9ChVb2L9/ezm0FuMidIw/T7Tefg4PF56BFyyieE2BNXzHT8rsn14hTMgC
nEDVdEHjYY7ECmWDklVjXtEGSAdyCAXkP8n4de/cYejYKuqAVIkrviPONfbMKiiygbZ4Uu0r+ulJ
4c1N0DnDw1IEZmqBK6PUpKn32jvz0kqIp/oGS5YMRjaMGpcaXE4xLlntb4ARaMims+dRUot5/XZe
Cu5su2kuNH1Lfs7MYuLNY8VqIJpFQxULL45ZyNOraFqarVPg+9OgKglbMLjrEsRflrKBTmJc4EVZ
00mBUpEGFLp8NcCAWDza4QIkp4fkIvCOQG+1u1zWi+vaw5r7QBi0nck8UIMAN610frrBlUKha+/U
Ly0OL6nRv9FgMymdBIJu4WgJ+2MGeWa6B0zBilGjjyM8kG7+usuTzT5tpA/nHGQ4irBwmydrViCY
tZ8nYIcX/Gci0ORcQXtT4Qk3cDWEKjg1Ll8lonL1mxFpnVNQV3KhqIqD0Gyb497p48IOh5Ns7Nk/
gaU2mJGFFhobarwxsIuiUMBKxlcX/7cB63l+dWVEESkMNYFd4uP6NlDRkmRIAXTwZ8+4V2xeG9rZ
CwwLg9dUZlTi5JgIVk2vcmkjX5kcFZ1OKb1Xsjjzujb/rkgse4t+VVaFAoNAWTy9RHBUWvXY+a7s
GH978igrf2jkfb//YphIxFnpc5r1pi+fi/3IEd1A6P070yZe/3pgI/vW1ybTGPkq4S8sccbBBISH
6PweMhguoFaQ+1I9MBB6CG9o+2l3zqjC6USzFiVPMsCdmrVf/7lDqHvMYKDMqw9D1E5OU4Xyuo6D
xobGXqos9MtnrmecbiNKnIC48iGKOqPhaub9M6VL2qzfY58EzR4tmqV3yERrrZKPilrj6YyDeaQC
vgcTdAkz76ManKb95KzqsR0u+2owklbdumQn1nCvYt+VEP9ryolW1wEq20qLqbJwNLZS8OoYfUOS
YpaqG0MyAK8D1kWKqr6gAu9UV4KDPAf7IZuOk9cW95aCa2cDrMkxSI4SwaIO8rFCldlsvGtH/HLR
m4qwxmg8zItkmNI/YM+ebxQBNWaRxbLBghrl8p5sgRVOHS1jm76aoEyB5DNIRQyL4KPTq7MwQC4q
NqGA9EHyoWpmxkHd13/N6ISfBiyjuspLYcEG3nGUpW7yomnVveuX1cwCvDIAAar+O1t4sJbDRAOT
8EslckhY2BlblcllDNtQ0oUxZecxgvKqFVtRXBXdppJTRQboWyp3K/naf0l4MS6AhvdF2z29O5kT
rbfnkC6ZbWpoKrni/oyUUjj9QmYMKjF8JDEQEbtfKT1YVtPw1PT5R3mjjsK3cUo/BVgPc7xT3GLM
R+o4YZAWvWLP6n9j4ULxZ0k0yNlpVn7zRkuFXkFUuhJqkTjVuG4nPlqWg7u1DBRtZOvptPwqD/Y7
hCOR18fbavM0NWmTETqgp0yaxTxGqUQ0MjcY2C09Vtdv8llCOpmbzB1nQEdxqE/82sr7+COXfDdW
uhjGKgIqGj+/Tl2cWqGIHA2RqYP+9saM7Tw8YogUMODwiV/ya2teoyNe5lqW8+EwrAR6ew1UXKZi
HGKxmAvOIAuVc4G4CcOZTgxWxzcd1MGXo8TD9myBUX+7cT4iU+Npncvaa4uYMLQ2rClawh176BIr
LcyCJ2onp4KlKl0EVAQJgr6+TMFHfZx64qQMXpKqbdektTrKp9cKi+A4HWv5I0XxuQKDCZMQGb0r
9KbNycm26BAntO36NyY45vX9R3cGQbwi8hWgaQEF5lGYQH1feom9doIN69LwbSqVZjC58eaDrcnE
FRfsLdoAVZsJNOZ2s5fk+IbqGrKL/hu1sin5YLStfnHz5y3EEZvbHne/enJgXK06fviC8BfZadX0
5bla1g1xPxiAwW19XJv6L55Y0HpXm1lMNSUGaaw07XVQFJuZJFrRfQlxs7KGbQ29CmBi7qZ7GHmS
bKzKpSedORt9X8Hyun5OY4Y6ODg2wpXcONtKlOecjp/s5E2RKO9bTPEhTZYozsgr0pem1KhTZoGM
hz3IOrEqlXVNQpGP1uRJ+0/uD2Yan846AtEEy84R1OaT1cm9+agEPUsZ2cPttsgP6uperLrlGOk+
HonA9Vrezry3TU7NF90JVJ7n9+n9bpz8r3aO0c/TipZch0zIEAC1XyrtyNtKpgq/IIa5yYJcwb/A
0pKEq3LgnRheSNXY0TfWAyVsxldmHW7BgjYRf37U939W+wqj/qZLVP3U4bYw+6Z3ByrE44nmnO+Z
dD5mcuudoMsBkl4W0v4wFepf9Z0IiCKHwzRTbTtmRm+DqDwVZp62GSF7O7TOC6K/UzcYiAB0HXmR
OlNS8NcbqDpqVrVBBEY9byv8kVH6VbDEwuKHFhH4FmXMcZl4Eji06cktXUrWnMU4nE+Vrfl1LqgG
KglFQrZnzcLQ7j7eg0/CvNkPBDDHaT9O/sB3HG0waZtC/rRIHYyBGsBDMuHwr7scWX6GbwQ2qGgG
AlmfiucZUCC0oLTUfF7QgpEl1GLJ4v6yx6O6loMGxvemQQnPFI9qVlFgViOKS/h2Iv3XbBkYSdGt
+hCOsq8N2X5RK4/v6Ha0P6+POPyfURVbaRNsdx6uGekPDT0QWaazjMVJNhQc0afRkHj7aoDpJJ5a
JuJwqZn45rDwz0xWGZicxWuvLC7X6cQkAuyjxrZeskLSPjlr55b9io7wh/8snlnU9dwu7Y9lVrPs
nW1c21ze4hoM4gIE/HVOCDyVWWtcnfGuC2rG7kc4UvUF2x0Z4Cdsho1/QJCRqJi25Yyhm4lZkHef
gUq4yw67nmgu0lD3JZ055WhkAzXyhtnYYudgRvCvE/5GgUBOW3+Hftt2hGRZhyIW6XLFSdZ9Pjf8
CLDM9uJjTtkpjJ09Qm7YJl719l+mE0SMSzraVLhStNaZF7qpHgEH9ZtIp6RA0uCVGKu+lgn3yAGO
bm8sohjKcXw+elfVDci4Ih+4b7dl2P0zQO3PlT8Xqixu0ih7XjrY7TSaJy7n+bigOfvPsUYq7M9N
XOP6jjNbmeKawpZjahd1FyDc3PVcEXkqChAEYSRyremMfavCLPhZdmbyjqjNYo9VnkWdnX5ncAoC
UXPuhgoZ6BE5P0UFhOKBxREL6EucvWYnkdWTbRXrFwnRvLw7cQfnm64xoNfe4f3epMFhLWElaUWr
xvKbiyGCw9iXy6yMdekzLuHnGA3WcpbDkaWVZ9t6FUVzyoy+0lXeQFOMNeCoABdR1Hd93vgTubh5
E4VkwA0UzVq4F5htsh4lleZCkexu4Fll13i1vRlKVFX3ohTntuKMlHph1i2FoxY89fJeVHOR4Gnw
ptX/6JNtposX6lofg0IDc5NAQimGuZYsN15V+vyhzOW4CI4rkE2dmSjrnuOE7MVLEadkWrs0lpzn
MiglbZrX0w36y03K270ckQgtqTZoC3YIvopzPjNKhvUmsoCjFX4V8zfFXRHyH3Dv5bdxsxgpM7Tn
nzHACsHBJQ5dzU6f5rJprPZz3/HV/AnZkKtAMp1SYiPVvzZWD2xwX9Em+DeYx7AdGlVu3HA9lXAQ
IK+C29alwX3bD+BwfPAazEV3/AiG5J/KyY30xDfFjGeWoczfCdbBJfBw6G4SakN67PwkeJMUAHHQ
ONIuXlscYzjNupBKW0Qb2yKFNtZ7gDz91o0EMcvaAfmPtrYusukNpjkEDlHyLDTCKOnlmHnWzuu1
pFqo3bEsHel0dbwdLBfFZijgBtnAQ1gxFOwpJEenpiikL+1LUeyovp/lUdcaP9mx7aiioHOFN7mG
lJnKDSstTD+0LyCES6OoA1NWGhGZ14hlCbn/8t1xXVkt1wMtsd9+MXk3Q8EAOnNh0sy8cinOMj87
zcrE3HwBBqmW2hG7hCl0f5TeFAcnFxqb5zAz+kYPe4CwG+3atiOtUBsPWuU7xmivwn3/bED2O3B2
newTlIJNBW7b5rBMpolvyLgvLOMzSY8uAL9jTS5K1vYQouhvdPRV6jMKp8lBYXAPAoNZwKFY/sJa
Emq7D/EtfbG3U0lc9k518KNbRJYSJrgP2+eLeTWzKih1luSFD4KzTNPUnW+pnVHHgGEN6I3zOawm
z4kZWoftFJfE2BZkIEjq8ejdaeRTFZ9l84P4edTtSK2AKk+AGz1JrHR4AxUN03w9lMvpVnRaILPw
Bvzh3AvYT0bk6VKlJwKHfF+SxoQ8D13EVCRNr+1aVcGU+KiG9pzDe3H4Mqw7+F0DC+0VzzYjDYtT
q6fOeEc/wI7ssDrTkCMB+v5bqI0kbaDy/ht7kqbRpNWPrPpsFQdFk5NXk0qHxtlMEso5kKaIXlBN
NwAM5Idvihgfvbzvxeqka33GjTZNOCpYW1gDyn/o/UC6nSlnmqcDb00l8o6RHMQE42PctzYJ4yZE
0pAbJVcLLYiCieQqJhfpLjJoV1T3cKoh3iFRESTpfkYA1Qg33yflGpxX5Aw/TAY4ebir7fL4URov
iHrS+OaxKDotmSpIRZGuMfsfNBA521KKZylLhWDm2ZfK4eHzEt6sHwSCt+pwTqDDtcuBkBzbpoQb
T+hdzp8CPgm7EbEobzTvaI4E8OiwUcDkcYQX5PeB5wNGpAOtPE0l+XqhG1MfT6Lli+iyCz8Lomsy
xV8dEEy8yUFBHrPs02nT8vNRbEIbqAPd1t17gLtkdOD9tinXnBJUtHR3lcNSEfn0QOP+h8OSJQdB
/gGDBYkaLoa6r4tFT9XMQ5dnBi8/OjIcK3JXyyx/tsoh1C6z62A3F3en8MGQhueRpu6zX2Ob53pA
XDNNWffaVsuVISlkpS1LAXIsrXSKJ5DIAgjvj6tPki9spwt7xM60Lj+LbWStGAE+clXxWfo+J/RO
Jmt02d/MBNpD8yq05VSZVrnqli5P6+xDZUb3o4T0nkE1nthssH+Fd1FRiCF+IuIxNS03jYwJ1yrJ
f6pNlKVWPnLq/NKBn2CbpRedhRiWX2T1IzC28JeY0Y8RHtaD61Jw1C5XFCX3O8i3eH2Q8JRsGsWB
3p9elUEFhFs5FLsZZEJEXnQwjsOA4g40wPEs38g/XCq30l/jiQg8DRd9acxIBlgQygvxZGSHzDud
WJHpKHTHaKNGzBTPAk8KQUgI293129AB5vusBsvUUpphqsMnGAau1IJ3K5jJPbubW0jEMN4dZC31
1lVvi1cSfLvLUmmxdARqOPgcQp8a55or6SsJJ/a2zNaKDyS+k3DK/eYUykr42UhLfOdEn9kzxFIS
ZMmwbkGbfQvh3noeHrinsdpe2HkZKNOb4govzQquv3hyAenUlTtc4YsnJpZJJSx/v3+b/8UoR8dn
E4T5XubqFq5rr9p4jL5i4yXh7GsZI0qfeRAnLtcEruMQiTLr3hAN2bWihLGQKHntPLSkavwB/Zs7
0Z2yaNgD4reR24Ezlu+pkjYUT/uSXQ8aY45Rh9CGP1WwQgxUHonR8uo5lCky7nMh5sR06UMon8BR
U8yZ0a84fxiXnbAF42lDRfnEnR7HJ1O3yQMJgHhH1FN7b8CVTxLG5eLkTeMMhfxfzyk6DYpPNOSO
4QU3faNjlddFf9Yb+gsVxps2CbQXuqjtBv5cpbctQfZR+h4TxTpCxxkY1eXZSELRyHAPcK1srWC0
0tLkdXiag11Ehf4M6xFTOHd+JSFiDzxvJRnGBKH6XO0qz1kvClHjOpjanUOWrOnPRRD1COaA6jH9
kHGrO8mmXXuPlg2++/IdDMvAKRFf2OY3cYoFH4n2dvB0JqxWlNxQTALpwtylntroBezl9BxSQl48
rjOL5ukvQJUpUXq0mxV9F1GoszU2ZSgBxHV1wgl2mDQrSnRZBeNF/aqxlIbfaUfpALY9EemmKsBa
S1uGqzu0o0ssOWHwx8xPMjsZBsa32nl1OiiO5K1uAazhM8WkHvY/XUKYFrZQ8AVKFbQ8YOHY60M9
FrVKCJcEcJZ3zKM6epYxSEahRuzeH8+xpS4QR34c/ZHxmgIzLJ/fq8G7y8VJzGMOIcM8ACTe62LW
tcdsAkRCsYcIkV/1fF50avgTRlmtQWSNRLxiu6SfbA399l9cxc3eJq2MvmZ8CfXwHV79Z3w1tns6
Y8DAllOKUDKtIm0ToJBr/07XsfVMtD6lcT3B3dRcTNs8RHZ+Mugw2/dMtAzIVGvxRv16YkTpTRH+
sPmK4iFX1aMr4zSBpucK4HKdULF7g7TpQ5EgqIkmpHB4I1D9uGlMAr5ttrJ10vi8MIesWnl0KxFY
0OMB59rfDiWvasoIAtIrrAFgBEtftBHu0drB/oN+nWU0CMiuu7W1dQ+BpQ2p3C/0S7PANFt8RByZ
ixyiH9zpY9w2cnTkbiXm4IFRrDZN2DXciHw66VTUOorh33bHFwTHK1qGX5vx7NxQTggcwsdamFv4
DPs3ocRzxhTjZxmTEBh/GFpISf1sSdUT+Mo6TT2sFrLRQmJauytTSbf6DXHqy37ohas3nbj/h6Sc
lLbJg1YH+lDOcLyeDJjCBr8fOhHOjXU39vVb6OpAiY4L2e7YgS+xaKGGxAAZGE3MjQhmXYtQuKeo
8CInVsKNcmCGJSsgbJPWYtc/TDgzmw/CKSBoX2kRWiyM61y2Sv+YW8GlMCEuQTUtsHP0A/9YMgoN
DzEksl4AosELCzhBh0JcUIcPq7W0vIPgz5YA/LhNg4/mG103YLGcEILyxrFJeeE3NsDqjd1UVf6B
HhEx4HsptXMlQbnhL52XCF8SGTgyORefil5f5ua9nNbAB2t7VxNquC1BZ7OlHvDXAvU2q3jBRyh7
CqJqApWrEuVnMQOAzhKUgQLngbxLPSu2GYuNtSbXh03De74i/AO+IXo4yL98VcIrxHXq1yseYKGv
H7Wbp85QlGUh1u0BvGH9pbVP3GBAfdlKCaNfaWSWidzOc1N+T5jwH7tTXkwsmYA8p5rhOpEMXF5N
ATm0srvcrDqmWPN81xxF0YWOLpjNfpeSj5XUevm5N0NJuqWedHiZgxXR9OKpI+jAJaG8XLGHkvv/
kt9FnATPM5NAWXvru0BUrcK0d2s2zmDrG8kJNxvVA/Y/FnCS1wvploGekPSUDG9Hsp6cLno/NUrb
Li+pS3x7HjsCnsXjGnZcqKSUhMOZYDhvGrb3YtUG5wWBoWCEkn+C1waQEhAeOXj9vNgTOAJ35fyQ
5bQXPfoFCXhR8SEl/a6UdydGTfEev8WbuIV/Qrd/3Lr2/6YHES/aJvQCnDe/kUL4oXqf0qLhRoo1
4Kzx4/3nCVpTqFM4xDvT04fWhCBb9X+4hkZriyVPnoTNfCEl6a7ZCMu95YkXhLYCavkP2dh/51tU
ewf/r1vspZSi/RlyT2BNvUVpKkOT0E/RulCWtGD/kdofnVkc+N4lk1/f0JCP4hGqm9ZVzfeOFY1C
A6UEmbC1B+xWaMY9CB/A7Hv9uxj4WdkU+sglBMDaSvSwai4jHxbJ497oAq79j6vNA2ki2H3pO54l
YAFPV4awSM9smKzriXSeyQCFdrNfXi/36LVpVIYK12mjABr44ZyRLHiWXFURyP6K/g2gB9t72Xbo
lV/ltDryaObVz2VOrWKmlMVGiUgh+juqnm4GzTBQbPlBjpzsmYs3kpcPvLqMBE8drNi/YaOSx7zD
C2OppGpRczNnuCevbyrVjp4oXuERzG0BDgC9byTJFpoFrg/+Wt0j9BuPSnql6WoMDfaoYvMQAG5Y
jQ8/Uip8ukEHn/MUorROh0V3gtg4PEziyIbvQzuofCJ1jjlN7Cs0Od2g0jwou7ZvlUsLGasNLt85
Wk+JkQQYsVYP3qty3KnCv1MoaMiDfHXLnd9dTU3pKCCY9gnAXS3vQQFdBsmxEzBjnVmWj7JEvqbF
P7jWu65W1R5aA1YDMATao0pxXCL2Dfuw0pV6UVypAgtschatxCj8vqpNg8Fn8WYfPCWMZXQvdBGR
Ft+KQKya6tyeeaVpsp/hteayPV3a4Iqf/eonD07o9vRTLZ0eZNB1LH+XwiWJOMgJ45qxAzsVu7pD
E2qust2lnokLzxHiuFb/IfSVG9Nr6OifizmASpYqCuTv54WP69RdnZvKXcsuc1xqao9f80wDb8+1
jHwk5JLqD77pGoVq2x9EZiKPrOOeC7TgWLLkJB3AaovwPXiDMLfhBZH55QcunOJ6R6oxZBdt2das
EztT6ONk1w8lRWdSmlUpHlzZylh79A6/8ygsfDTPDhfAkZt+9FOahZf+/aT3sSfiBs2l0FnBbwSK
rcVzwqye3IrM3Q95E17tJkKoD/2k63zhGuf7rWfnat8t9DCzq2arldXiBp7i9GEvaJDrm41oQRru
2EVWI2ky3r7K25rxAQ8Ox4xOp4sZaSQbPTJ8JAZjtAlJYRoL1HtRxkgnS8Q1+XeFpS3xzAp6Cm4f
bAo+APqRAz0uRKU4Y5W9iXls6PgxBKAAwOVidRFDK/lP55ekbSDPj0vdFzj8Rwn8O7D1q1dmEuhZ
YviYypKvXwLDRfbr/qts3JY1U5EA5Y0lnGrJfq+kmRzRrZ4xxYm0sCvbR6x3VLzAAs/PbkKbDf/f
oVKAl/JIRQKZPzwVg9Ve8SQA6AstXC3KPpRO1B0XTXv77vWu4iH3Nm3S3KBJ+cEB13jl8DgXndRN
2TWEC1KBLxTjAdGinfGE3uGhcvfYEFf2GepERmtNOYgpqz6o4SgbnxCGh4hYGiQFb1tVroHGOy5E
fRuD+NKsgT5KFb7RJCfG7F35XBsQUfIyWEgjP52hjXzJA/+UVNNjmJLaq1pBesEvhK3mNqh/Agx/
ctJ0QgmsHSY6ZiXVu468d/leJA530UnDTB3xkhJcsl5+ftAGGNocIuHLaSJzzYMcDcTglREn0bZY
Lx8G9TMyU+r1JSY36AvMRx23fIjWWPVjjgI8+fVomG8qarAW8NKguEIm7uWsFuP92kauzuaWPm9o
LRT3ZVs4ZiY/nj4g8xHkMuuxLo8+IUwTuN+DIMpD5wBli9XANrKPqc+Jwhszdh9844RFKI3mkdz7
6fGl5UsvVIE2Spb1YHOEj2JdXakcihWmgTKpH8fmg1kOdhIRcCwEtfG26YNjEpoiFDR0ROFn0x7A
CRNUTGDU8ePZlBxLLWM95ZF7rfH2HTqVp1raEjVXr10htPuNjdwknQN+tvEWbCta4uXduB7MCnIN
TK2EAuwbRDnK9YOlD9VQrj4Az3ajINhVlI9xBufpVth8g98AaEtBiHE37UboLIquHgpFT6BTXvgN
1RrUa3nAE3LYZCy7RlmJVGSH7VjKTE38d5KWM5+upnZpxj8j5LcrU1r8LgUx9NPC6lmPYwI5VLSh
wTR6sGgfARGfX+JSn0PEfLemKfb1HC2Z4x8wPv+3ieCXTOuRPtETZXgm7FeeiGsWE2pJY3lmELq9
tS7zZmr9DNBamXj+gS5k4jh4jzQoMIm1mgPTQSooCXu1rPdZKVt+SBj6gtqvKLPApv0cuRDSvH+Y
9C9q7Dl9tY3GvbBaZrwhyYzJ98rIn38wxWSEtuTxLod0J7cezZHOQpxsYw5K0jNxP8rRYklk74R5
uAZhdOU8BQTFAobbnOOY/2033ECpq5VXDRoEAOO65LE77heeRTSi6o3zFEX5C7rTa0LDjiihJKIe
vgOOaGm+zw3QLbVf8K7Sd+8HPBLDHhtqHknXrzx3seDxI7Au9yV4CgqS3oFF0roEHyBQytGr06Dg
lLuLVS3ETgNC7clVwtkfFE5LA/vLXDbjGFA9JAVbhMxfpdc2Tg8AjGoDsIsfgnFPcUqypTr6aVTe
8VsSWuahnOYhnm3idKLqcDeIQPcl63WwoMlvJCfMK/0Fp8eKLVntRRy+VaPsumaZTK1xcMcAlgaF
5mngqyc3h4YoKe1Zkg44+J2Ajxhx7ZECvRNo/s+PDjiLGKKoV2J3yidEnlIg8vbbk0T2AD4Mk3yS
dGupxkwmfSx/sQECYNN4/a+43Zhv1YWeWejbDB5bi8ZmFF+7A1nOd4Qz81c3gjt4OyFYtYWUnWSv
Y9VgjeH1ll/QLtSGpd0N6U+uqtehPirgFBTcX6x8hHbLczc7LBaBc+w/MdDSSlDuiumDi7TXadvp
ReBXE43xSQRdUZhNFk5tZTVXsc7RZvcZzln5aCnfwwKwHdEbotFmZYzl7uiGH2y6CJQrEfeorGWQ
BvoU39DtCD145m3+fZfQ53kyufsM63cneC5rBGSJpjD4umI2ibZg7TbfRN6VkHpoDNC+zrKcbfZD
sR/xA6WGXL+GeVdM2k73KfRuLpPJ0iMTlJSFhmOtPSNdOip8jz+jSrqOEh4kAEaabWTxqFAFMkVt
C9b4tzzIOc/ZzsQqDf+CXF0T65uL33dvZAIHQUrH2+/AhJ2LgfbYilrrGp9HAgB8RnuJONnEGLe1
D2aIyiSvfH5hNo/rv1825AS7aAvrFxizQF3rbCl+agh9ySYCQZ/u4H4cC9oeFCPqcnJ7N+8zFoVg
8oS3CmAnzGGiBBBGBlAPJ0MfiokIDvBV7waCmsLCyhIZ3MyaGSG0d5bWFh2eh4kCjVfwEox6pyoc
DOUbG3we6wFmiPNPGmXUYnD8zRzGdJFbnMU4FwbieeTxRQQaKig/FXTFEjk4+ykJYGbgPsLsVqVE
ISHzFwvpPuPW0UPT1jtsADTPydMhrj6Hqz52lislf3qNX20LaYsKAqQql2CDqMCSWuAsbSQrUmkP
r3Ivtngih/ldpDibMCd8I/snDrZw0aKtT5BIuCHEsz9Ixh+imxw7BvF3Tf5v6k3/X2SuhHxQNq81
msxFoBCIQ1nZVQuKNSsh2ZZlUGeHp8/9o2NxWqSX4Sy6ImfefxJDEcX/q7VNFhQN7+8wsc0Q+Wct
dM9gs8P4FiH257/DLBZlrz1fB9cNxqmkGHAO9ipr3pUx54uxh2ZKjcQz2KBbredvxzlGruHBNEp2
5cBe+1wNwMMHGaD/DxQwoK2vJFyao5YFEDhBPIIHW/eg6AXDYkDnDXCZcIDIprw1Ds4ffMP65Rh+
CJao/KgaWQ8dJT4I5e2NtrIbGDSvx7eCjUqfF2ZIvk9Pl2b4tMSRFUSdiMAw2ej6Z5//w42LbDRb
kVIQ3BACzDLbUJHvUTfg0HJt5reCFBoY249yFlHT8K/ZE/GtFLAyRk58HtNSt5dOOJ5IO4dLA2zR
3r9U7Q6MX/AgC+UaK2EWllW1GuERnBoNQOaA0MkM0oSphsCJC8iKwx0ZMUTwEGir643blwIAXFf7
ulX19scQ+bi65ercqe1nX8S570NxyIn3V8K7P7yDENmpSYmJNMCanwte3YkiaUcGN2+stGV+GmlJ
xJTobEXS7CSrh3t3suHWAdR68BxHBlSz3cK96O3lTF2QVIUZ4a1j7vuy7TkepQ0nFAcqENyLLTl/
axOZ9d/8teC9/jLAbbRrkZm39riqf78atiIfJ1+8WeXAWXWGeqjgZc8nHIWue09pl+Rnn7Bh3z8i
CIL/I3ELa5PY+FvH856j7W1BLkMFZLS7B0sTPNIVKcX/y/fQJRlwwEISx0XgzGB2NyYaoHbeUmhX
uvtcE3zyLV+iPldCWnzN3uJp5f776z1+QqCd93Q0baiHnutjyFxppEzOx+aGee7uYj02sQV1BsDq
dew9NwmJSDVIyYASZSWZ8rRBVb1l7l+Y5QpZ+3FEmAQ8FR6PCG7itdzN0S+IBnX+6R0o//LTrves
ORox5cUqnfpCoomxU5mEZNnnGX0Pr/GMroavYJ3SwGrH/QMV0bEPADlHv2odkqB1kLtHZSGM9C2S
2KZM3szsBtVBXhmFDkGDmGhqbojrxf3xYTS7xvAclWtLpPtP1JwsuIufPrLRnH95tBClDMpAuLsM
KUtqoO625LtKc8eDCJn6pMiAXv10X68OC9VqYT309ChWnqrTWrXITYB6xFQw7Ruya7SU5wlpzpRh
7jwZm8VTCoVYfZSRoFw6ztsr1EBZsA7e8TlLAKGZnbSo/jyOApYtgI0aZWILUW4QZpErnykj6GaS
zk9G5F4FeOH96dWHheUio1xTFJ6aBbYCfhHPgjOimr7PxEBudR1Y+mAfkDd7mZKL9tvKKqVjS0A/
K/cGteQk3oegPCVSQlE9PegJZkaV+xOTHD5TygBks9Xk0S23AKQr6ZOkrhNDjPnePEXtFeEpVuz8
4cYOAtmAFdZ5B6A32feYa/HEZe6cXzPmZ4FroY0sNb3wZhpnpW3MdbIY9C61eAQ/yF2z+/X7iiPH
ZZQA77DXIuSEJfIaUmtHVpGiDv8X4Xd3BSRrmpv+CLRKUY+sGbQOYCPzZkjIcUUMA+BsTDDqL6xy
U8EkbXFGVm0VU9XFWyOi1cmIjUSQy9TP2niLt9Ll27uL1EWKgaUXgYqOx80d7fXIblCp7H6LDnKD
z/JA+hK9C4M1Ybfj7EURPDg3UZ6g320o6WbwDaAIt/IZN9cDoZPT3TFpumfelrBJAyvI/UTKgzZw
KsKC3QMGhS+1rvJwh7vsqnDYiCNva6CbLqNXxWKRp2Z22Mlz4sNVifpynqO6HH2rkomcSJ0rVOw/
KyXcGPYeTcWEdI9vwatjYB2mo3sGAopRh/vtlAga3WpVmAw594NiCFmxJ+wkIYdeEo+jCsAaumwg
hZYobkIp7xHWIA/E7MZiiW87j9+JGHYgAybPxYBULTKYKOmU++LWYTwqk+1e2try5e+zzaBRIp09
V2iKmhVMlawscp7IvIIPSz9gtpplJ1BV6VfCT5KyLixprxVTttC7S86uvJTKDLA+0NU+JRWRnNqS
dCfvGuIahkhtWWVOwR5tXL3Qn7khKsAekRNH5+2vEZlh8dH+KS2ntS6fkIp5/Lp3sFBAXOXVYkbj
qI3rVMhDz0KcWR+J7s/XyDo3M3cZ1tT3wxz1zVbZfcHQKK0hgkjJOTePxn7GcevmwkxHfuwzYe67
kys3MrzBa0EbZc6j1+0AdgW+t1VKV23EfXp7iJCD0XmyWJJTJYuUp+B0JRDXZiGY//RWZywues+w
laaGVodJgRXO7+oDyVbqinbrSqtnAwgMnBUmYCCj3LwWWrX8h5GoE4SJmfiDwEWh47PCZxwZEtKT
H3hh79Zr/bzxTyBSx1gu4BKlLdcmbfC/wsC6WadAIc9XwPlnwpgqrZSktLivw7VLgW5Mkn96jFh+
GSVUyDRopkL4rQoidrFmoFAEZQDfdJZakb/zq4+9j1kkIZ2Ffn9Z57J5h8iJBokYkDIGrEm9TZPD
MpCQltTvTOMmGkJJrKTiNSJj3ODxHrnHI7ORr6UIY2+YQ0TKb4w/6nyU0VekZzED6EPXrlecvUx7
RTiIjjTX4lk0N6IljopFNF6dltIY2kVm9nr6/FZCf6uygybqgjtOi2C95YKRVTWs9yrHVNTFrRJA
iIvY/T2pOS7B1MBBbLgomOIQvg1wzbeBnvT3yc5fc91XQ1WkX2CMrNeMUNmnW2bkWhzf8SFUmeWz
pTIHpLHhxyJ0UakEy++Ujni7JOpc4WK4QI0OJFAoxJWB8wTalncGT/WH4Ofnyqm22xC63Hf1qt3l
yx+00n9XGI1RfoaF9xRSjLNsG9BpvFgf7iffQ8ZP32fXGhCChWG1lklWoZ0cSIkxNMo/VX7J41Bd
kaHLS+GhD+bVM5OD3fVDJ0SwO7R7OJcNhgOB1fWJ5BTZa+K/VOj2RBlIs4TbVT3vqj/PPAIq97qN
5i0emw+/Wg4a2Qz86cpwgYAP7RBTc9waTG5tX0VfDq0Ly91gIWYB9bl2I2pmG+GJ7EXX4jD+aEiW
tZsYX9uJvbQVyRn1HV1iSAK3puuX0RbJCyfsbbdrFtprE8qsCIIsozXB/43MfLXc/w/nbmjimiTX
gnaEUxlnP04p1GVDQZvTrpmqDJ/XZqMj1h033DFfqBykGgez7fQmziI/Y57dqCQAlA9iJyyU2Qxu
/ifY+iUtsqOgKtnmokkAMMYf9ka/y9LSe+8Ql0aI+NUeX2BQgkaJ/fLw5jdlrTcaJ0/U5doeMLYQ
rz/ZlZlYOeGicaQAz3rwQa8BuT8rwke/9hYth98Q6wu8xCg46pbQI5bdY58/yjqQheDM7d7XnZPa
7Mclm5RmD6C6QcESNoRcYac/hRdLAG3YJKQx+zq1s/24Ado/oQA0qc1/J0aSMu5GEZFXEqzg1c/I
KXrJOdne0jQ46F/egWjWZRPm9qzw62XMRdum1NlYSOYAEm/gaCZySZymXCdIlRFFFTOA8gXfBWpT
mnYOr9X3prgNIJEgkp3CO2JZZn2yz82s+h2ZuLlV7JXA7fIJxN3pzT2mDPg3fLrB4LY4T3NorV5R
PBC+AjeZOE8FfE8Grol004dtGLQVH1xKML0lcnQnW+aFaEWdhna8jmptz2icOJWFTcPWJ7Z503Cc
QvFCKuQpAh28ugR532uyyOpYXCpbocRR0lO8RrHEigRPb9ArRbKLhdO7nNMw9ZOW42tKplxX0BmV
wuSO451ja6OmQ2ks8u9kV3/GRKREArdWB7dHX2pUVQ8yRmISfvptBgxJJwE7BBwYz8gaPmBYaq4W
54dlsR4qLB1QSVHqhZHQw3ogku3/UbIa5eB7xrnJoBnrmZGgzKCNkIfY4yPN4lrDGL3b/mIzE10p
mMmffyuOPta1axFwsr2xEoKv1QRQByiH2L9Mb4dookvBt1LPmhISGkkrzWierKtR8GTFt6wPvRsj
kSleNCORRDJHWD7WB+uv16gjja5feT9TcuuV87XC6k/u0axBz/eny/FVSEv+w5Dpj4H61jKkYTie
DoOHSGw7+OMR0Z0YpBON/FTwiK4ZVwjpQG/9kRm+rhhhG/XRaE4oXO8n4Ulm9j0UYiUzRJmuRVQz
b3YuRqYahxd9EjK4k3+yCh6Jr0hb5j9OqyEED0LkCV0f8NRDkDAUMSselfQuAiRPO97ibGRUbRDP
m+w9tn4+JIsVlbmsNikkzbjv15qrkwFflrSjicXpE4TeYQ595C2FD5vrG1eJAZke4fr5J98665IX
3EFIVVdzQ8FhNjSDA+miE3XX1ALXwaSluz590eciNRTWbytJ795s6SSHJFewdod+5A4InkrT48pI
Ik0OpjE+uVMUPfBNtfWqWd7MuXHs7P9q5KZlbpSQZVRWnv6wMFqaOnBACREGU+OFhnJy0t3bu3Cg
Qyo9DMzt1uohSYdObYdO72uCtycwAM6LiptljfUcpNBFua0bxM3vj2UB7dAtcpih+TOFbbn3JCRW
M5t9dK2+5WHFhj9xWm9LPCkDRHP76BL/O7cMr3y80lw0PdC+tCIH3D6i3P5y7851Uc5lyZ72V+o4
eoZ0c/ynqkfjK3cwrHIc6vRxzork2ZAU4dOcCtssEtlGv2l4NbOwoQOaevbvqUPek+wctEJ/xCsJ
J+OrBQ3OfEyX8I2gIooiusLPagrPqfRayfqGjl1UB86zmFSDK+5vZy8NgDjefabI6SVeAJyMOBZY
Jvl0Gu6WlfqwlmmmNKqfYyNEIQYWQEzJVDfuyXPqULnD5DePgrfRqyQG2nYBKTzw2V2FiWmuIkUZ
0zwCDpV9j0aCBcr++sG441LEe2uS2V4ng9ucMMSNCyqKQo9BLjFrnTLr0dwk+/5BtuwtIQjNzz67
Z5h5jJQtmR4y9mlcZYF91bmY9cGDtj3KIwlgDClL6TKSFBZ605dxtZUT4Yrv6rAXs15LW65jJwpl
omTnk7016dP/J4dI29SzBdQbFd9WKJZfim1cEEdyBOzlCE3W4+HgZwfWSBfRuTFuupy+4CIqYDdV
FFNkFdQiqWpR+8rvzgAu9hPVyGjyYu5Tmfs1eTFZeuowoL3BX2M6KYRuPOlhb5l69Uo1kgRLv9ql
WzUNuUMX3q5labYJhJlc+AGto2+tmQaEY7fE6Tncw5gJGKORhjEmrFslJ+7Cb8lMsdcbIo3LMTfu
22z9aIv9o/71j4/9E9IibgIH7rvQmR5r2X3MSPkctPinyXO+hdOTTWHCseGXBFBY+57hwYhrsJ3o
EqEf7lt5zPPpVPOanZcy84anB/H4v7mz1EMNEvza/6WqgcllTHrAPhIdfshQ3AR+6Y+czrkWThVp
YZbuIa8vwwTjeUO/es2VJDv0JcuDLbfZSiB5uMPaxnJg+O+RhPboJ1Ul0/8x+U7GZ50CXGHfab5l
DDqR1mp8zTqfz0IRdxIb0Tn7CU5GY5MaLc672edJOK/8qdwGkj5l3Vav0Ua983mZ3gxufPsMZM1S
csnNZnwzq2Hd1ZcR+cUYIMCM6qtCQzxBsjIG68UZF0RXvmhbkVCLMWZBHpj5+faxPpzL0iAdYb71
VGYPekf92Afm7ALNR9LuBfBFr3D05VrX0UgkOZJcqdj2X/IhfvtGycYq2SwLRFWFaPpSfe6bZgZL
rtW61tHl0w3rZvukV5bbthgOOs3Uk/xDs9gNEyuemuj/GWietx6ItUDCmQRmRiBpsvggNWgGkenP
oZu4ymub0hFNwfuUTn2forgB7VXzvbLPynwK1PrvjfKFWvj/EnQ70yMbibUp4lec0sfL54hIRAwK
ACnwlI0W7TZdHV3rQs91kl/rLRwz2LgeEs5fXNdCpc9FSxXFF8jemHx2G165GbFLtZ5CAKB01B9Y
WpnCRJrtMxCPKgPioKgN2ZMMTc8K81KaZs8mZ5xONMQLLWFQISAmJy0IDyxtvVzqB97gI7MyESC8
ckLI5/HNMOCI3UpNz8B2QxSEXF/WrU3Nggpnyij/5WO34wn2pNYAsaSogOblf4Gd150/uVUvcQTG
OYVyh1sUdPCEBViiSocpYPIZJawBdLak/LfN8g87jsOzXmhbADvGx7gWzE/rD/9P8XVH4aNnFVrm
RNGXC/my/uecEFcZ+Flf/uRCsvK7ukYZMigEwSpEHANfnPoqDXP9C3povqhjjReXAKle7T92xMhl
NXQriowARpNp38D9mMuCrJARocQVxQV7pQSNefFTUw2pKv5C4OGJmzBPBUtRrwjjQESaIX5W3cby
BX+vSG2X+hfOnsu1hcAFY6NRAqxlrjvCUD5Ag/zBbIT02wjPWBHWRSpILs/eUGs5ZPHe9AValBpx
4xgrBeZQgeVvvKw+pjvrBtabJ82ZQYkuZC8QxlziTQL7X5tCZ1GabeO5Aa1PkbuKjPfFTSx62WT8
PSj7NTdigC2f8c7AySyc+ml5OeWRWV1xKgNX0kDs0rm1OP16WgjEXxqhNGXfvmTOUU1LPVZjKsja
KvWmgm2Du/LUoFnwOjH06Zm/TiG+GDinXwsWnaB03xRoYuyDlnwsB0F5HDFvvDX/fJ/sm2Mimi7C
76RMO5V/IcEktoRLN1g9LtTMeQeW3cO50khCUs17g4PPxzv832avyg46uIGeSjJi/DpCLIwQsqLn
dyOUwIy70iTTvcPc0f+/S2slItsABNjxG8/TOmEYKiwCdmH9+SKSE5FeRYjW2MCKh0Ra20isnZar
k3JSFvmKuJLWJ633gsrdkIp2XNFTaf4uGELWoyIdLnhAIJQkpHTETqHPq52nOFcSxih03DGOdyNz
ePZoHfDp7txokMMh3O978ZLZFit4dGe/wAHreUHktp0QqBSr2OxFxRpvGhgzIvV+J6YyOc79cicK
LkMsGZzi6soK1us2bjhJ0qr6/5j4uObFRQEzwIbgOv7j6aiPxnT1yH6WfmypOaM7/VldNR819bki
WFg4DYYqzyhdJHIwWUQ3epCYEAFsUDXF5FDLgPHInOoCJ72jVXwpQ/BpQwxpBBNORz6yau20SyZd
bsoGuOezIeq5IjseszP8ospkVS8UkAW75XGWevefGDsxf7oukbx2hWSvGqPafIirH2d/B4rOv1TS
/kgwVcYxDC9vS8sm3ZRaClIS79f2WXDAVG336VhLx7imbe8I3MhYFn4HdxF8ER8uZijJpaN1AniK
ENTbU5p9EXzx7mBWuYBtHB1/3+D4LCjKfUkkyvh6iF4ZxOvWJujH6wM+IFsJW0wqiq9Euc/skS2C
fw8kGOf66rKV2wNa+KcPn3qDCJDX/bdgFaQ4cJj2MQSknlNZOEgcqoxpA6FHA99iKtZ8B5uy5+pw
dbOCuJ2AuKtBMq1K6P057E7/66IEsMj9zLHvQNNsu/xNeVPhtoaRmyu5smUUpH2CG0+yB6OI/RTU
CzBArHXfoqAIGSQzeUSWmDK/A/YL3uqAM9wVNgbomCpH/oxFsvPpGC9a7oWpHXGg7KUsHMRUbHr5
W0Jr3/NRkIVZKyTVfKwQvrQCRkWYZkFUj9e7mvZs0OJgIEmkkkgYwRN7FSKrI6kBN4h+sXriNYCj
cOHI9kpRYl+RzB2mKIxLmZYvPGpqwyWwfT+iv3LfFPn19MwjBjDf7xswbb4yZxMJ5qQUGJfT0F7r
eDRoJzEg1sX21pZjApDlzkhufcc5YsHzhRq1pAah97VccZN43d2hUOrjTqUmrL6/o9goj2CCthGM
OgpIJnwBAH4JlRBxE7a/ravqpsW1PiDhggtJQZ9pWLappzyz9JKCSt/B1m8CjUSSudxJk0jOjEL0
Pp46ZBzN8rNM7AlnKd7fFRLKz9qYMjrB1E+c3mbVSRknnEHUzoiQOkBLRaIZF1Sl75UQEEJs6f2W
a1dYQuhzpPBaRtN0D/8sL0dYKcw/ZFXkCRFnU0T6irelA4VWmxTRYmsJ6GszftLt+Nyn34QHD6Vu
lc6LXsCcaxbtV7X69vGBBD1BzVbMRdV3rzaNTVXgQ3ScuzO6pOn+TBRAYA9jqaRjO65uCAEiIjP0
++fzLI/AKTBKbVN4LWvAezQCbdfUphZ/pEX71WH1tgwYARP+OYHmCietgCXcn+1GLcqlRJOgbVGB
aT8IXdpJWDCjS2llIvY71C1VfJJF6Zv6gXBoDXsu+rq3o2B2lLuO5QN9Y0NZrH59pvm0lAFuai4d
KSFsE1j/+2Ny6HU7lz67EprAe5TYAe/WSi1hByl3XyeGuKOLB8wpRm+KtyV/3P1ETV7Zypu6demq
LSbYhb57Ks2kJNrxbiKK2JCyKTGXzeqF0hYFzfYkdffxgJYHAil8dtw+msKOe+LnQpZPeh04kAdx
I9V15jmjNHsuSdSAYZXf9YwcSojWSxm1SuqftrKAmqUbBebgeSmK0OqJ+I9HMtvDskh4PtKbuOMF
E2EzBOOAhHgdJQOTDaHoc/oeMZKjKV2zsubCI+3Nz2MQ4HLiVhh3x9Q8lVV4PpYij+sdaBC5mTJx
P2YWUbWjfQDJ9eY8ZlK1G8MOON/X1ns3ITc1TQmDi4R4vlw7ER2XJc1lzIdrM+RY7/ROYD6yFHCF
CXVK++ngcD4I1iXzT86JC4eqAn2+P9TohXMiHwuyF5DTZNcqBnVo1Y6A/U31g1PDgQmSyUwJ1ytp
epdD64358ZHq9pVR6ReUf4YqM8SYB1Z043AXuhScCkV+a4hzoXZKpiojri/Xc5CAhSe8J4pOSDRD
1lHxaMtmRClFkj272aM0BoOd4+Hzu0kBH0pz/EWYdiH1Re9gOCdkcC60fL8zeR59b0pZQVo0Dt6w
zjo0op5n6V0di58s7Oi5AVc1LKSqGimBNjDkax3iYNPFSZSYuJ6pHw7AjtxYkg21iJCTELtpxY7J
Qtr8fEH3CBFaXJpjz2AVrQaYv2T1MuiMf2saJ8FRCgNUbQovoyPrC8xHinV5gSGbkeCVYPHl2Obh
UkDl/YA3JGucDJ4M9b5RK2t4lH6GUeYsN1kdqH+XKX4AWoW9dfXmUWGbdxq/crN7jKkDwDoLhB9P
4RAr/1GIj/4IA9OC9r5iZ8qrOn9H3fLlFCQtij+iQnqKy6zeYGEabXowX/MZWnxO8PmASk7gIw5E
+bU22AImaS0MmUPq62hYOfUbWVc7EdYCXfG0lJvECwNm+xwnMDiRNNXK7/lKSgw8RrYf8AQq4R5Q
Wp8ebfVPEt/OcJ4/MxhhUpIQQ+sN0WZy4mkr2j1OihbDkV2UMLI9NQoT8ZpkKqVYns7oZspDoGCG
jkYXw1YeHe2FrxyTW+9ugD4twzxTUQUbdzmnvVICsjZLRz0IOfMc8xWsBRsvBuG+VkRW8LMc8e+q
cOrXUHiD4fpQMNcfxXL3qznKXvE9QZkoxZ0sZKaT5RcpI/oOxfPKEnq1rRmO4njZydMbigUEVFom
tEw6OT/bKjLxAtYB9Abw9c3Xfa+dmORLoG0/Gv2hedkwJhBD6Lz2jJNBVh3dwosSSBQjmTjQuKe/
sqmtrR035HoaKJSeZ2ugioQhxf6CY2bVelSntf3HiYrFuoqpu/PE97QrqrI78b2Tqo+sVsdN9Xak
CICN5va/hZrg614/3MNERKidz6O3Ip65V+wg/kAPuHMrx5hu6WzTGmrqds2HUoNxDymvasm1+qaP
OMISuVGccRblY2O3gsRhs9rN/9o70HF4vvEtoPSxT7WXolz2PcrXtTPCrW17aftUZPlHWmqOF/mx
rwD48V0YHVCNvo1WetLKfhbWs3O2jN3OpRltJjoXM74SoMo0Zs3LWlOFU3j5oBjr7Zyb6+6j41uE
NSyPtfVjEfbUVjmdnjin3wEjhMPC/viDW5iATr0OJrjCIyEQKWG7njMi0zyCYgOhlYu4laX7GDpV
v7KMiVG2CotwfYV4OD4gYWT91W/Bz40VOcYLl6rx0GKGT97Jk73mqS3aozi1/oaMCISF8EFGXTHf
8yOq9ffIllmGNjjmpF4NqxeG0fXlnTlrHXU60OvkU12hgvLiabKVGiPVqCZ0afYeLcXHPj3X01Bp
SZtcGAcCSy6Sj3NtY1Bx7sNlYukva6LgpH6I2SzCLfSZuyfhh9shL1qMBF2+JaQxx+kMmIExhZnu
0L7VzMHMWG0bIDgcxhB58k9IfQMyXIYhGq1HLtFTNytwl+AFMy61sP9tBD62IQKKXfkXe07VHKle
uHT4OSFF+rNJ7AZMqQeLUv8dpGDBAsMcJ4kxsfglmyVwxiqXd5Hj5BSvulLVT2/02FcMmr2xAw0e
HAegsY/fpkjg093qGXXnltn8AC4UZIQftbst4tXDOFVa6l8wao8uKkfO6QoIjs30+CY1U8GeZnO2
Z8KPduW41cPuhGTRWMrzcdLwdQWCzyQ0DqeEQ+EvNqr6WzqVKsb8aBKH9IerUsMz+2e0ruK5Ag4q
PjqotE/3x+e0qQd6m3uCL21ZtK8qbRoB9XQGE4cyjgZrEm0lX42aHmZpKrN6lMJJWbs/hsNjc5FA
j3Nc3azMAywYUejksl+pRLI86wF4AIEyhEs/5nMClylEMoHC9dbnn8C8cI6Q3fJ5exc9jLKhAtkx
V5C3Aoyb+oM0Hu6SFqpyNNFK+kM1ULRBvyit13ajTIak2zW7My3eYoS5OMhNsSEnU67So02MivXV
Iiu6Aqpff66aJL6n7HGY51AspP7K1FkEoalmz2d3kDcdCzQiZBraTDJOtnfNgbmA8B+cWGyXiWfr
2DxZVMWA+NbgNKpoh57kcIzAe8dvHiRlEBeycvOKx/0QlLpfcTIoglTz5ftD2o4p1CXs8498DuSI
MNzBcFGvkSG3AM2GZTfUSae9lq4qDQoeu99Yc3+ic0BIKKLHhPTD9luiEOHemK4DVebqYW3/xM/9
ukTr9vM2UPARjVDx8eMYEsfmNBQXZyIRZpTt78BLJdONOYo2bF4UWjjF5YRBR2+BHXllV9OSX2CX
gOJLqou4hALyq7bUB/iOtxL1Z0q0YVn1hI1eFaewj7P+86sTjkj698NFeACRuJ+7bm7w7wFcFpJX
r4ToEFSxdezue1AQCmcY670wHe5Wnto9frBtYwwMdyIhMQI+9TH1r5j280hfv19G0zJfuqx93U6G
vsRtOjKMklpat0gcyBuPXHwoBYxvolTn07SH9+TbH5xOtN4+KNEH7JIKky2eb2WjiJFzeZ6dEpr9
NC66PYiCqKSjPPby2lwgjSFA79OL/hhWKgp/gQwWQuB/OMiIPbf9dd30rFL2xzYus82exbcoN6QI
BklDXJktQPB604Gd2/vxodboCc+tWzx5BSLPGxr9QEzne4TIrUSBGkFyuZZcWx2uYbLI5ORfUHJt
pjJvx48gBnIL2uO1+G6eIwu9jsYBF5sObWAzbxzITXZJCo9/F2TFunsGNths8xxhJLd3CpZFwG5K
hH5Gig9/nPTix/HR126S/gom/Z9J7gUyjzUvNuS15K5+wwupXleokCu8yaXgJyih6NywARcwfM+R
3WJIlRoD1mI45p5ILqkHnF6cO7YNQLK2HFcYVc8M3Ae3fMTMzVOLA+CDRt5XfKPQ9e43q4ReUlhT
0PpNt03dPx6Hs5Am3MPupqOXJ/bTWeVBNTjWA3p+kN10JZZ/WEcl6jlyO7sXqMHc6FH9DqtFSndp
aWO+4H5S5kQon/PVCW0KoEKVX1h6Sddey51O4Wl8gEOdKUxqEL5rjN6lCF3D7OuzLO71V3XJL3Pu
sEAOxUOBX7tjn0+XVLpCIC0HFaQVVhtGScaQWrG5l8tfRCXslEcdkCq72T+ytk2zulN7HBa5dtPC
bYNzInycvi4xSCF5gJlkfeWAEUngIiMYxWwQbRcV33ucLPhTwk7w8MhGWW/X8Ord9Sxc69PzgApA
bsNLv/QAggsb6+LTLSDej4nXxbnRTFuO+1N+kCap/uNDOcgyZvBFrQrDxRdxSHh/fVVtl2XhbUNE
GEwSPpt7OJiBBeMyZ9CbcDqvxqU3hoXx8WC1d+z6rNV+s6/SP0lRGy7APBlJkDBehBM9k+ce4gQa
cdoeRyZ4ORSMN6vQTg83Id4T8u/O7zBJpghQz6UutwLY8KoG5L8fJjkNjwMRF3jtzUXRDTRmJ6mv
EwwAh8Vd9CEQjhg5Rf7Uj/tkf34+/ahnlxXzANOgwkQRzckRrfpIhWSAzleVqZDkAT+u+9JAeB4r
3s9Qw3RXSu1GdmeKlY38SS8+C7IxspecJjBz/cZrhpuMDdo1K+M9caye4ii3Wice82UF54i2AJiB
46y5SCWVWBaJCpiP5CNeIQvV7Q7jfHk/Y97zoe8FoMSqF72ajz5C9rW6tQdEL9WfZnImmrQ21Df7
JrtnwHml7EkCnc4xgaoYq2wDbjsZkyfVhDdGeoZn9gEdoRLLOcelEX/5FXw99aRKJumDzZ1zd5++
HCE9++qIRgLSOZsC8tNJBW9GiGFr0MyBt9KV855D+LIQVMIRYyI7merX/tD6qSXZO12174BNXC4I
eDWEa6k9i0f+2GGs+XfYKjzrW/55Kz9qHvHFo8TunRmF0ci4nv9vSr4b813Lmyumn1zscsNly2Jn
+BbeYS8RTql66QXhaAlNwLnZaT07BRbRSfMg6ArVzaCP9C/J+FUauNXMsdoOj+wbuMqC2OE+S1hU
OR9jNFvWmENNCGcHKmFymC/7u5A+3rLWwGDiIPvohe1yNRGF/dTtZXWiaMsjmUjS6QBlJICt652Q
qaT9Tl1+MLncOS5scLNKfsrOQUGqvjed7j5WjR0CATdRk7u+PKaENq/bVpCj0q0dAkS3+eW7+B9k
rdp/JbqtYaPU/DhBNLczm2ivgUr1gL4xOL+oqPFNqufurAAI777t+EGrejkVORSmp/pW48ImcByS
p8mB9WQCveG8OIGt5UIDiNi8IW4sRlNZO5UWIdpsOL/Hd/9cB2KiSPYZ+01QlxeciRpMWx9mpNoe
3mF77Wr9IHzoOiTX75gZ5GrRwiDAp2qnBNVugsCk+5bAlkP167sQbwi/5EhSNG4ktJiKA2w7IqRZ
weJHQnfzPGV05toPWV5ADptrwMWrJB2sIDvylkrxuPNL4sMO9YMvuV4ZM1kHeI6OoZo27ohjb9gb
EyKUQ/ilMQpXQoJJsVLfKNFvbLexHljdgzNGYxAcXoOH6rtbZ9xPQpyxUjvwz4C9lJbYCzOt5GBu
wsS/Nm0TCXi45oC2lJ3gm6Ns9GrbmuW4PW98OJB16n2xT/zMVcSxbxbdqCs5ZhQsKs/NmuXN8Nn/
v/CuOVvujuA3q1taggxAilU4VywDBPGbPFQMQltu4mIPxRirlkzTSVf7FdbWA47dA9OZ/KgTqgwE
5zo1kZh2HjCb2iufDldJX0mjfLVkktx+fSPIaKATQtp1YyZiKxdBBxHEaLXBbhPe/FE7aSw0nW3s
ArtZ+LjrP83TXtUXxm3GSBOh2QaEVS8DkqOtltlR9xClb1bUd6aD8QEi/bCs3upt4QqgBgxJgnKM
1FFx8tLHx4riutjXMHtSLtLNoDME/wrPRzXSQlmYTPzYYPRxy5ftOaHA3L8vh2caSzg45mawUwc9
rJ9R3wieJmqN/54YHoVeT35aURok6z9DZ0muSjaRXUEjnpc7chdtrD5jwpQTxH+pqBCiDcGrn6Nx
/QIBENR80dF4yOMC28FDktYtuBrA8c8DuCqNENRap/WjsPBx4wqLeRp2fijlEyRDDhKGqm5WL2mc
mB5ya0PraAOPgqXKGtaelf8mt6KL8rkdygOK9tRHQWIlCOBUbuU+/Fr7flbjEDbcOPpciNz+zAwR
uROqLj49F1hQuVfXF4WmEqueuZbTiCZSiyoR27bvrcvZGQAKYjevtr34idTb55TfFbIncm8bmQca
yRzMEst1lOXGS+w87KriaiULKkI4lBH69tPnYwpPwycttyy771WeWjNU8o89oWpL0ESI0tn9ZUL1
E+OPVLCH/KFeo8ceB2COuh15kMcLkr9cbDgHMZQ+TZlYwXpjlRrheWbe19GX6vCJSvbw4rMKZ6V0
/YP1wEBf/VGBU45GRJAgDXXnmLXdwsm/iU77fwVAN3QoMmKIccQlGp+uBXVwx+1S09t5RV65M9Wh
X1P2Xtu1bvhIN7WQUIzWawNypW4voOwbt/AyGb+Xc1JXhHchwSLRY4suf5kQ1mwhsKF3twobDUx0
Y4fw9W5EoisneUoo7v3t4PEdNUigwUlWANfjFKWHcrGShp55fLIUMnV8lk++ig0qyjutgoVjLPCV
VYKuT5hX3tovIs9yuaamikOhExoos0wY7PW8A0wYeWSTLkDpuMB9YTFlgHF8ZxSNDQMyZpT5I74R
afwMIYuNBHiEFpkXXE0dwBeIPKblDJhQC6oeAvyUmZPmp3x/EcIJGPlO9F0l+5swPNFY7X0KRzRC
3q0Vbx9vBxZJ4nvNQGD+VS8xWCGG2CXgofiZzOO8eZYZYbJXAQDFNt9hbxWW36wMtuXpH3jeXUmD
36Vk4OfJGBVAyNk6csSI9fDKND9Wd+bFxKhtufwoIyEd2swvX8RedhjYpfz3k1qgtyEUsQrc5PZ7
58phhjWV7hfX706FQuRnqNWbA7rpVlEtomks2JVKGsDAosYncMfZRdE9UPwmBRiA1BlgckPiXawa
24oPHnvAXHPVR4j81c3NDDyD0dWXQNcuqpQqo7aBFlOt5acfk+S1Ur+2FOsO1Dv88Gq3o/qn11lA
gN44ZNHlxmD9FsYJrGeYXOKUWDq6PJX7ywyJ6CWpyWLK5m4vgRDQHQSdBDxWWYaNXNdVpJhYUI26
QtuN4dYvxUOPxqqUM5GcleHEbZR8qO4YOpeDDdLrjmz6zqa2LAxQCwrgSLx7baJSiMsBIqhZvMAU
tU0KyB3ND6RSbCoPOxO8/4lPm3W+ympmVOkV9nGU73cH4tSLO4xTv5Fe4tw/AAT5v0+msEESD8uC
GRTRVy1q0kkrGb96XjfJQQ+vd7qcpk4cSsWOV/IPNy16S60NJGp6BGXHbkUIOU3bk4m3C6reFDis
nlCmz848HYXSJAohJLIo7WrtAJ2LYOhb093SZPeeJ0tcUEOCGO+q6lUOqYJpE2YRlYQ+qKqrjGva
C82QgAE0wdt/GREDZtaG/u0wNsGwzVj7vVUUfYHh9wcMEJJrukriVFXPmnLQYkkxJxhAPTZ5xJGm
FvJpuWQTZnZVj9w5zKU2KAAdeKfvDGqqpZMQvJCGbCvQTaOe86iWSghLA3CWCx+FgEPwC4ofO5w1
lROyFrNbsvc2g9+s9v1WxEAiBitTbNeiXQsEWPMVNjC43INSPFO+Le3BSnmxfdfdhYYb1VLORWHK
/bVIisdTgMdmPjgC0rI1giRBwm9DvLF/QbKNSAtWD/KowkwLMeD15QcGbXfCuDUzzpWzXifjDffw
9Tj+8PlvtOzNkB/tOy9W1+aecrQcgTf/XD2EJCpJc6hqtitK5bhtYGtK2VciM+Ps45RFem4OooNz
nxqhoPGxsaTajzl3HHhOq+jvCRf4PgnKH2Fqqyc1620Tu78IMALgdqty2e4WTQTcf/2FqmOwBruu
5s3bNyOBqssFqq1XP1+lqWvpTJ+KsF7bFbKU7Oc0ZtxJbGqCmdBjbeAzygNWv8jR+RTZYpyC0noF
TjuK4J2DLS/cBQkbw9VHFYw5Ut1S4xWBrsVx9NSfxu+C7z0HzXX+0eCofGzSXex+kQa+7LDcc6VG
IEHT95qhAr4wPwNhc7jORn1cGZtekM+lueB9goo20aPZ8G8WJHMyfMNEwkkStks2R1LdAnBt617S
DqmHNjye6wZa3+eDAyTgRhVIEdv8rma6Mh/uqmNA7e+cUMECsgDSiX03DGZYzCQ7fWCMLqiYl2kC
WYoUgcW2fH4NWdEOt9NHfR6ZFF7jAIuntP6rI8TAo8DtxAOS/qY0NVR7jWEqejdkmHDbDK8jcv0c
73BnJ+kR5yAWdQJC50E9EieQKSEBi/X5c/8OcDgwaiVolHq5wl2j6L8oBqS5k8X7Zyr0EKU5Ezod
1dZ0i7Ra38A7kTMqEC3ZHoG7FvDIMyxNcN0XC6TdryajvUkTht02vIpnE2K4tLTT2l3RSukiIB3t
bwpKC4CvDmWP9hwLzq+qVlKPkL+/RlzdvfivpDKCpqH61kFARlgltPYLpasX/0lgHL5+Bjt+vvvh
t0hAU9ggVF47E4OdUR9OXPqyxWLir/IfCgnM9hj8Fd+eXkVv9TVqlPWEp0rDesooLZYsgp8bV3HQ
rkBEepSIf1ExnDm+MimiqoTAdcZ2QAnCQgS4DedVBbbX5SdbmJeWcKVK7NEatnZFVoDzuXoR748a
VWMa81CnUcCsy20vc1QRxzjBfgm+YJp2DRIBh3NBcCIRfa95VeF1VETzC97CgDM7W0uLvSlIGjid
/VhAwi14HsMDmfftk4noUES/IGFHfwNe23byQ6t4Ydy/ZpGtlkpbzXUyVVC4K/8IfYInkyDyOW1t
2o9foAsQEVQoe71TUzhv4Dfc4tWVnf17ScLY09UN3ReIBazOwaokLFzvD0yfO+2BWR/KEDu5ibMH
nlmYmPxZ5ZKZyuP648XxvQWbr1d0fXgPttksrE04s2ZKiIz3qsEftnvf5SBfEXSepcJ8uDXbQzhT
a7lFBdvfLam7m+jzNb4Z1ienBZ0y8xOzGvHPGM4ur4eaPHcal0IN5G3JIVY0ppzsEsEiZjnqRCS5
cAsOWlMiCQIQzs41SevV0pxprEnJGM03JW8nw94o5ROh8fDtjDI2DUZ4Q4ZBPKqXTohNZ24wa3HS
MV4vbjqi2NUuvLRutTO+ltF+n6wnfAxwUaJiY9kZEg4OKlrC3cehihsf1xhtg6IEXCAuJ8adM0DG
Q2dm//89EkxRNlPXhOyYROHHewh1atC34R0O/2x4dNsx7xFIlNXvrI0Ib0ie73vbPpMjZ4JZHE81
CaTjZMqaMAdWTbdT0NAYVGjlJVBlTxGzTurtr/QHvQZcVw++eKuAE5vyUsHrJiD0YqycoISSXQ1e
TWZyV4bKiDR3Wj06CL0tVZUqdX1V3ka+IcfvC7Wj5fReQMwfASjgXHlI2ojqUwQl31orV6IzxS1j
ybUxcvDZOiVteltltHCeQwmO3m2d3rpiu6yFN9He39Tr08mzNRGoL4c6oj3pz45Rr4ynfrwAoEgq
W15k6Y4HO3BDHKCDvmZucZUEhZYWQyFPp3nUAcCD+EMFRu4zKdCzdo1eaW9xQ/mnT6XBq+zy3+J9
0hDB+/gBTxllofudSclPig0sFU7LCXYfuHkeMPRtCOFtCk8/tE8Qi8nmKHjJS4QwbvKlIRPyV/KN
6pY5I8m87zasaG5kFp0PDuSVLwMM/ecvn/L5XbL6VTn6OSikb5SdWeqssdgvRlNSbwFHqno0zU5X
hqCfgWNf08VEKAigF6TgIUzMLgoOcouv6cCJ9fKEvOyP3cuRM6mMkRBlFZ3YXC2DQ1bqzxCmoFbE
MqOrGWrRuGg0ZEW3XV9bUtKm9WQirg9svY+HnAYH/Yc8czv6yedkDNespvX2gzkThXniErlUyNm3
0B3OyHjIpcSDVsnrL76UcVbF+WiesNYuaoSjj+e8xKZvYpWQ/RjUqswp/Mwps6fXcNFyUfeT0AKz
nBOMfY16z66nDf7dL3FIyhEP8vcNiBWBddiaR/I0jexNeUp1hZ2X5N8AhCznyxeNZ9PC2YzSSKJt
0YEHz681Vhdi3RbbrQuY3UlKBLh70edfm1PEq4Rr8EiqSKNSO0z5uth34FnpCmvmOAgNrhzjpSVv
fqHVgPkCNBnwAep1Qn2WBrGQRePAlAlVtrOkywVQCFHLRXnkfw3Sa3E9D7JQs3YGEj4vW5kIeK8b
UTPODQwNcdRKA9Z1uve+e8bzIOPblx3x76AGUEmNSZ7YlV6odc28oNbFz1Q0QjAnIVbzKBsplKOO
PZ18hrUrfiehLA5WTb1lmdDZ5FGRXE0uSdQUkY8ldeShKzuVrhZsinlB0nvPjO1S6dU3a8oJ+lVY
vY7JilEFVZGKmktnhgvVOJyPLhVR7SIaHgR68bSMIiOgRyhAJkk6dOsnhYEJ8WL4ZG/a1mV/mxQt
TK4bwjjkgy4JyplufACXUgzHKYZ/aNHgW1KDImL8fRmk4vl60j5Gdz1PDXNeTFTlYf13JPqJ+EKe
75Sh/kfAyEABJxswd0js1/5yOIv9qNpb8dwlspcs7+Tg3lJ/I6K2lAVjlnWIWHCl0220W3Z32+x9
RhwgEbIOgivqMwQ9zuK3I25lwJzjXCiIZy3DQ4H+Rxbsoy8bPcl76WHN1rgY4NsMGvyJweO7Ky/G
SwfLtah2vvsidoeOQ3jfl7M0d6vgDBJna6sNlxqD6a4RtpqkDKsrVS6mXbQakCXAS5f+0BlwhVAn
UicPhKSKqYqlXJsf9lpo01zBBTg6K0PQFVrAWyX923kZGIgKXroaSvNxHrDoo8PEDz94ESaW58Gm
erXBthIkx5aiXCAgS8+z8QBZc9lLJZhhEviTJDldCWOGqBRktICI3IOm4suTFus7vHOBlHyXzscF
Yd4H1TIFTzaaUZ3Tr9Jas7ixOHTb/0yc6amF6YnIo4GgOY7YclIWq4e69Tb1GbLAk14tReLqw0wN
+a+Sx8tSmRsVbkn4PwF47iSiyCtn+evjNRQZNU5a+worv/b4FDwcqj2J8/9l5k11lc4HrthDvM2Z
DMry/oEq3RSds4EbyKu3Gf4MdOe+i8xBiGHxNhwiU0Fc0U58EICMrvmqFHgD5ZMmNxv4v429V302
E4VyapOBLnXVpaanWsOKXJRR3QfZDVNETwRULlzqzhSro/C78Bczhn8Hvnil5lEDHqBva2GIQPcs
lyg45qNexZHpYC3k23E8idJ//IaJHXWcz4uGv1PGhCu777XhAiPrFowYDxl/K9In8SIGqL5hQhtU
S4XUOxeuikTSTpoDA2yxO3nOt2J/HE0FBsKq4goADgqeMFcR0eSfahZF+1/IgQYn6EW0Oy7j7l9t
SKhkqj4CwPNVJhmZrOTCy3YFvafEDZ2KlKwJ6C6OQhh2tKVJZpTndioOKiuGpHtiDY4BckJ0tNW3
F98idiOn1LVd+QWNPBQR0I9PzjxbvML0fKTB71LndF/3Q8NXilIsKFbnMFzMjE2UTnocm4d0DseY
GLbJeL9TUDCOUYGktIzrfv6ZqNQaw2V2m0KWv6VEyFWa/1Jr4wUU1tRn2slLcFNK9sx3O3VSRnDa
Bgk1Og8nE978Blmc8yE+Cc28o4GirMJgspc7RaCtkllixyMf478drDZghL0Cs/tNBnB98BuV3ZsV
LAVrFQJwkSEwJNo2N+07U+Szs4vU93HtOqyxIuTI4jgwRCoEAmfb0lcFtKJ5CWvU/w8bQV+1tF5E
PfwMRSi2itSnP5n7tiSLPwCZKiPQbwPA3ff2YpTBTR5bWwwsp8dgPGIxzB1fqar4UyXpZlrMfz4r
cojlGvi1J+kWvPZtZyaJia0q0gwBWQNeR43unJoxlCj6j6RZlv72uwYdXildFP23QW03u+Gzx5jc
DPium0Evm5/wEhpsJqHdXGb9fmByw/lRVoxDuctNbLEBQmEhneO844Tv/z7pyMW3926Z1DORJREV
eh1ZBnsHZqE8ql0zBAQlrLZbtluGEgtDgWzWB+0k+A8uZFDVkj8i2nKRGwkdznIoLqUpuoqEip8w
XXMPrARbYdBpnT+yc4MVHVclOOFFgAC775X8FT6F5bjO32ra/Xjj5MwkAGujzP2a9oqjG5CN1Ise
6GycLC54WgBbVqMtdLbW6vTymwmcdes+B9h2j8r0NfaZk8If5LpMK6m3j6XN6+QABByxxA/zGzkV
HduXvAsZxbryuk5XuJMPMm0CpB0qTzNnZWBeIPL93zLDSjJamjv3xWnsp/lr6DSfxUGXkr5322VG
3IhtwxufLB3FEwFTVSgUe2Cf6S6fR6D3yawxZWvC5cdFC77dv9t+LwyeZwFDH0k75NiPQR8Dq+9C
Vc3WtsMaUmbB1NhNOubxWe7/kcXNnffpikjnkA5a1uWzqpfNlVH3gil2KfnABubbdITcPjDsZ44m
7Lp//srUxqH8JqfMiu+9EGuRKLqpV5k/kFix0OvQq8keP3E9b5rljU88KHu1oOT6Wlhvb8oG2GJ9
yfPVYZtGBBQwsCGAUC4REmHxuAbABzaaBfCNdvC172fTcrgl2b3zOorzbFd6RwjTqyrYVBeFH/2+
A0QVjcUzb8TfDfgoLjzETJkW/jd+5xwdj8/imMSC5jYhXhn7pA0yMBSzRNv13/jAWFMQ+MI4nWRH
bDgl9BiElHvDA8AvrV/cUiQfmb6L2h4073gE4EhRm+mUGXyeQmPq0lyWVl6y546iJ0Qi4wl0nZZZ
53ZPvS4NE4RkRXGiQlQrpGS42QwsTdSwHTw0Ml6MEtsNxzmFc8MYm4cy5RAg02pzuxujGWaT0Tqr
f82NYKuWQ15xgfH3R2qwOUyhZ+qav/j/8IsORPOW9U4dQF4jIJBPs/q62n1A9oLo9hLXqnGiSajJ
g80Lc8rzk/WHLcfIebJIAVnaapqCTZbo67VTsDNyAeh+perjhwQmxjE/oBW1cF+vvR19BC8qNf9G
D8v+bzQwW0ue25jy5lGrmt0rz0s3G9dV+ExVgChmdcToWRyHuBDrFJ5HLRR4yMvof7o53MbF8WiW
vdrjbS1G7FXW3jMHX8OJaPoC/5c+Tn/AeMo7zzGtgvR7b9xmJKa+LcVwjSbygEirDUJtg8jizPk5
EjxKGliTxxFfK7zdHNR9mKDu8utaTSM9QNmyqk7rVMBPZ7AgON1omc1f2dtDR8OpQBXMryGqg5CX
KGLwhcAjdBUbN/N1JVLprxfowWo/hAWSkkgl5mMMfaz0JgPwAm4DwLpPjpvFrjK1x++UMdHcT9yz
teXTIiPdkT6dtIchqzkBsVrUuquUrvVkOmlJckkbCt7rcKqCEa6oBWKDxYYCQyLrwFlyTVjA0rXK
qD/MMICBWpHAWeDDAuJ5OmIrHsmnQcKDq/GKpE0wtyo2/T0tTnuaJ6mJ14rTW+CcFvzyfV8PgWLq
J/N/DTD20HXzDl9BCy15gtruSh3mhomMGycasFAXRZpfoZFLizYUz5Qs9TLcQ7m/A718Tw4xy6mA
rC5uH4Z6iprkjLHV5PN3dONKxH/AYSW+4S9nkSJv8KF1kw0XX0Kmyr48ny5UlDehTNueHR1dZdFI
fJCwwkUMRTsonUuc6Dexua6qLSlEzFvrfMkRqFnCbbjGQp7cY+N8/Yq7iOiLYBX1w1Hwv4k8S8Sj
Pd869QIWYjXgywmdi/2gC7VYXmgmXzXv+GPapf1y+9E8lEAJWqhUulthyVj57n3LZbTK3x8bY4UE
2kBw7zX/WXsPua1eX+c8JLYHDFE1nncUa9A49rMhHQM7lpkjaOQ93MyOaAbTLIfIPw+Nvb+H5Uim
X1NWxgGAzuczuE5jm+UA3lkK5Jffy7d+Fuwl4ifuyogoPnToEOIodzXcwI36tW1P26OTIy4tfWPa
5zLu0+GzLHJpqvhtHm7Pb3ftpwZC6YZVsCvEBkB/Udw/iZbEY4EeUilN1gU6BR2n6hjJ+ciIu5A/
Fc6rIuGuHRyM/FyxqC68YP3K+PFDOZBHnL7hqff50AdL6AQMy1//KhraEAGB5R74bxX1GaDhhNKP
IBr6jJEKIzhlirPu66x0W016nDpf2LXUxjuE/ds3jDzouWG93CnbiRjx8eHSJ2f5zA7C+7n1aIHZ
7S3qq0mLbXftiB+Q4ajlhP4vmk1l9sZBYfkhBWeezYEb/xMNSL+x9lEJLG2q9A9XLJHGL9VayAsP
YlfVHuwLtbMNi97atYJw1u5GDhNyre1uznMnoIPFUitAd1WngxbFSW9JQO/sVjUc9Hfbsda9op+9
2VYT6e+5rNlKYeYtT45ZiPxUABdrXqsxXj2jsDhl155mEWFU50Ky/IzJpb7rmj3h3jfHsPTEvDup
JyTLgO6ZcX9/jcaIjki1hXisK6wtYa7U3aYU5cCN6m2zHZmgYL1npmXCbxrtRqCoz5ZnGuPVB4Zc
4WqonP++IIXOyJMlBGg2gcq8erzgqmqoldYuieFXKaT1d0I6klYi5c9PVH70LoOPPFDGiX7FIKOk
05FF+L9kZzbwz6mINAj2VM9endEMwxOtCNZy0CM6KHGOnkc8NxmSYRFZ0xTJpC+FS2bqncKxljaF
ccPzUWchqxgHKOvfpP8G1EVlo3HOhj0EbMSGnmUQ9uwLFJzclde+l9s+ycVVgdf93LAkxL6n7rHC
boLPpBguDrH+UGdNM49vezqm9COl35FBvUXpLabj3UE4kgfQeRAsWXQkIfSHQjFQYmQ/D1+CcarQ
S2OVCIlu6c1Ef7vHIkMNBpu6/6py/tabfFSIXcUxz+tKp6N2TxJITYHd4TnhuiUO7az3jAh8k12U
zkolJ5Dh78Mt2vYMdKF//0K+kVLHcfRXojTFN3GCOBZOjVYFfH2+akGT3xa38yD7i/ne7IIbM4Op
VmElbvajWG/rgwlBerVQ62FlBiWqy0DF/6ZcnP3i0UN8iRJZB3894DweU/6kOiKi7E7hVc/y3Utx
a80WUe8hGJp9YaRIDYgu1PBZ3mpyoi66VlDZCCG6lElV5DPpzv3lo30QVb9U6Gs5yQqpjOT7Oaho
JO93VdWYIYPgegvBAKvodNnHMUC6M/d31T5OlMd43AKIFrvKkJkb7aq8bvOt+YnkySLnZ+lVeZ88
YCAAgtctJkEdlbyNgJ9BMM2hbPAgYZ02z83JnMSrlO5SF/gaCM2JVUOZU+xFmA4y+KTOTRAbChlg
iQ9aqNiUq5C5bcjxK4G/oqfGrt7Aoeset2hnx37TVDC6dixC3H4xpl6O8bM7RqE81Tto7gupCJOV
zBRknnA456VCMP5noqOoo1teUpz3DKbczoP8rdVEeXTEZgefbV6BcxxQ99/8Yxi8/dy4uHMrI3Nh
UAdg35AqbdFb840P8m2guJCh7YqEAw+JNxbmCOAS6uC1NOXfNGXdo7s6czV77SBDDORj2a/bu0XE
w5ZfV/5jCsleK1kXQnflIxQ6aM7NbgQ38JeOGuGYY8YonjsTNk0GUN99GCH0gaWyq/VjoReexYCX
iHMn81ZM1E8imn+TxmDy6b/Q853YETdMDE+GJYIenRdBtsXwqUt2yEbaxkRSObl0Kf1jJGtn/mLA
R9iFW8gx58DRKmKwtmRKujbytoCEb5IAVv/FYg9vT6BgCLqZ49Q4SweCGlbW/z0TvLoQV3e1jbvO
RkXJVAYpCwgePA8bGxlrWhzUMUuPrY5fNa1IROspRRWyRkQ2dLyTaZvWadj+VJrpuWgJwxu3+ei9
mJ4mhtXgTk+DSW+DWRQOtu8IkLAIxmKrQmfbywhL15zt7/bzF3jpOnlXlCDkt1dQ9NyLIE6XFsAd
6BdGoTXpWpzTSuytOyEkKKkY+A2PLMmRx89cVVil3bszOhIROZPQ4YU7zbPrHGMWUdAUngrPMMjz
Bvfj26IlcfA1R+wOyt9JBKWg9/Fc70R5bLQVjKWc+n+H/ftAUT7PQ3XOmwaoPpIoJ2kR0Os2x9QR
wABlu400nUEsejLuetLL3V0yvfqK19oHWAglT36aGuavHpIyc7Y2oCkjWgCNEM45nk6sACZ8bgYc
aBL+1XZn0G4rc16eIo+bkcWuIFBqno9TpHGiJhyfCRWNc/1kP2CRbejJ+K/Qi7fvUL9hzEkYzzQW
aDWhBwONXsplo04TzK4iJVjnebWocaAZdpPwrfc//Mr/pfAvMMqRMeLM5Q9EaQR/NmieN+025JAw
H/3AIigTPj78DhZlpr8WHVBWWy8KydUNgSd1pRVryxkqxs+10XxS1vVogdrQF6Fdz32VlMd4nBX3
xJp3QMVcHLKzqV5SkRNGioAh2OjxpWT9jeslfQRnbU962LN7dS+LrT5PV0k1A0CXyRIuPdO9BP7i
CFBeaUQrKY2brLSv76eaciDmqRpNjOOtYb7tzITf9/H9S5O14NkEAZz0QOVVRrzqZSpKY82xOx7Q
zelH/iRUinLP6dH0tx7f+GIs2Tbwa4rsO2kb/ZINMNqdmSOqAHlDXi9mK11aYMe7P+r2SZXnjYH0
am0q+C7uZR/jZpwM7zBrki+9d1d6Qbg9RU7oVOJOIhCGZrLkpbDIW16Xb7bJexvYdnQH0116/47r
HZ6qFZVT7j6TVueH3rY8SMqSgkS18cICIb7LTwc28vo+N72FQvPlgQFHnulyKvkm+GtLn+n5ZF2Y
QWc8bjcsn0U3jw0Qbr00FC8CsRWOqGtmgL7TEmdjxb58grVDKwufy88AUIZOCNVYoI3dBVfLD2TO
oTu0t0cG193x4UpK/63kS4FrgvRkv9xm3x1DPixFkhfvbeAmViueCqxFajNT9B8Kg5Z69w9zYb88
SakXZZEMYnhPgv0fjXHzqAx6V3IjhZFWKznwvg5WMut3KN8w6T+wbtdoo1zOXiGLdmImZ1Lm2gH1
DvHcEVoHtOTmMPcmcQNmeBg+xfGMQGxVCFMgusWiu2Ki2TPFHi6OAtE3Ts6eeeIAItqMi4t8lmnQ
Fxym2AS48lkjZLaI/x78vZqSdTTdHwefP+GQCFSEeAYcGjG5Je2qb4fIqcMfQrhvPmBPvAgVxQu0
N2YzMxDIVk+WgYrcNd8wRS3vJp/IquW9kB8yn1ZaKmpnW7cAKz+Bv8CEcSBnMSkr0x698JdqSu2B
cILrGlA/9nFRMXyuatzdNvSTf0skaOocxjNTKRb8YowbCnAN0ETIXzseWS88nhiLJBcS2Tt22d2W
eV/uus19Ctal1z4QaPUsJe87nJ2OOnDbtECSyrMiDjbdlWRBB0nwDwJG8keLv2qjTrwwPYxxwYtk
A8CuC5iLDmOHpdQAIZTEEWRcYoYO1zFZZQ5IKJjC116bqIHLmAkpdQKvc6ZYjnoWrfBphNk9BPxW
Z8ciPD7CNyRjlj3Ua50vGrnq0T/U34P9lKpJ7rX8H0tYb0qr2yt67ItNGKfZJnC71hd7fAWS8r2F
Nc3WASX3hKW9O5yY63UhXLLdMwIQ0JfXzuCD+mJf5z3G60VQE6VFHR0Z6lsz2/t5hGa5gD4rWvxW
Nven9nFgvMutTRo94GtyPqdmCI6UNw58ARcPCvwRGIxq++zW92yvt9qdsTxw/hWozPrqCDLkLtYU
80Y9EilBH3eH6HUnoUhwjIVfvfN5xyLicDvg0ioez1xwt7qussPxJ+MgljpgHvHhu6r73gKyKceD
jqy7EOwvbKHKWnXaCEcAE7ED0EzIT0SO/bbmBMiATj5NPqy60mU1d8oRwo51dVjkouRrLDTnjSds
wYjg+Lk4dsbrhf/ytUkNn2tlgcpdvFuviwbpt8nZxZoMF4ofkS0lExS/uUUD5qLGvPKGdgCmUYtd
e5uC5KQeyW26phwgbUYshF5ON7iYl7dY3jy9XqAJmi05BC1q5f4dXKOK5/Prz3R6OLqWvJplD2wJ
A2xqGqT7zfPbgaUhe6Xmbf+IlHrCquBf+hol/ZBm3yagZoKJ0boT+/gv0PLhbZeNBFkx8WeLB/zG
lzl/Z5KfPkA7Lw2N6N1BA1AjEsiejbpdqWHSBSjZZplIjiDDsX15CLFBRuHKqr0Jdx+gPKqL+022
uPUzBH5hSBqeHJZacYkkrEj+R2ZCleVO8hY5hzENoq9XXybn6++36jFSbUJN03SCQYp2juhiiRsM
0+7Ujs7wDxYSY3eXMQ7OpY0pnxjyDy4rx8WyYBvrgxTIWDS7UZRBF5UlTeD+n4Av82U+kU2X1qmG
EtmHRs8y86MjUc48CBlEGMeJRwT3lwcynxwUPnXMsupQ19/ZtRPVUYnH6f1nOz+4WpSbtgtVT35f
MEIpBfyrz7u7e5Of3Z4PA6fDxA7OjvlfQniSDir4L4tjvXlcRtRRtHeC4jVf1ZPeztu0R0OXfAV7
8/Lha+WHGW8xSmtMY9RGBSK/0Wv3l4X4ZWSAaUqXP18tDhs5DOs4LmgP4RdqBSFCaarFA0Q2qyh2
BEi5jszbYJL4sLGwteaP2cNlofRuTtY2z/3TgsVLfPNQnjOFN3a8TUush2pyXGFjfUgXHMQdzjI8
5h1mWJgStvA1S7VZEsZ/vbUmoxO/2EZmaZSm/AX8UJJOnX+vuthCzcbG4aRsdvfsX/i5x5vO/O/s
+HVob5IydFom0TZzw/HIAEsOtMc997O5BGaFI/3VBQRW12y7wj336khTrhclXuj7no0RUV8PlLtO
rYBW3rdufdWSU2jLCZTEvf57fc7DeAvCTtHdhXEMeC+SzMyCMDqqxuJ8HcRiutzVD7y3HnzFH134
vP2ZkXgaV4Wb+PFYuqIzR7VsrksLERK57aV8HCoqyjbD2y9KA0oVw4RsBD+4Axa+0XcEwB8rVPhK
Al7btFY1HulEg2mhzVwIi1Ap5cuX0AvXVsjtCYvgvunnwdjP7q4GejXJdIjtZL9/Ulwm9SzXJoz9
ywLs29E9h71RJhRKiwY0vNcfC6okmG4wWwh0X8yiINenCAVH9WfuUZqoTTXV/OHD9JT8zvRaza+E
TMBDThpaxi0Ww2wxMnWb6B9u9Ig7FJByiHw3FelFmQRWRn8YJlB1OQzQuqUcML69ZQ3otODIvehV
pkcwtpB6R5dpQxPafofVxean0Pkxyzai1WPfhnobLbJ2Pwzips1ci/PVMKl8GLkykTsiqVU0ras8
W+GqMoPDz3UQkC1u2r3qspJ4ZglwWm175muQkHayHRT2rIdxiNS6LwITzDJVUOyKW0v8K/fO98zG
ZIj1mFjTjEJPE2AQWWQPJs5YCvib1znziEyPFYGpX6MbRb8D7swmB9gRR/VLYhRsyX9EEvGMN4fu
3/o8PhudZbQnCiFurY0OEbkZnOXqG8DqOQCajdRUAawiu13n1bEaEr9nDFrSkrTjcTpX1BjdjKWn
mtnnC15qXQCnjlTGs+My75BDApImws6mkriAa2BTHOtGOQGWL0DaxqqnyX5bkNGptudnXXmDi5bh
XcUmOHdP6thHyqf3UOgE2mS75Ke/53E/d1hpXGIwYS9ziGN/iWSEEhAmGgl4aAVtwFbk4a3eUe/F
VgPLJiDdpsybfz0zVlXk45C/2g4ewo7OOGnV/op7Ii3FGDWSB4yEcHlxEhdrx5/7pmzcWmQjbxf4
g+iVBWBFqhkpWAaFSaUu3S0lMPKOEe5QAPAkHUoqoK9imb3ArleEXHM5tuiQhX4vidDkFghFqTX9
dJqmEekZiNs7QwnhenpE+Ojp9+OPZvanTLwrU0BUuWMgzDJ5+AHvbTOvK5Ew6yvFZtwJBQr6UtSD
R33P0ijENwIZNGe+kUCgOIziJSGtXoMlUP1wnNh6/uIZ4FlVxE8X0zuw6CSChERGnW+dtnSJulcS
uZozC5HXR49Nf73aQT9f+qB1q6ZuLa5PeSt/rurxKWn26qgIQQbWyafdEzEqUqeepY9mHe58MuMJ
jzsQB85UMdYVpUYxrT7gkiKW45V7HlwONSkBko7oqcyLKbaq2pKaQ6oR0F1l0C2OOvhexpqHXD78
zDF2hcWnii5FixxZlHetrRYKzhOtxd/6rCJMRk2drVDDjaU0aJwtTyTp+AOUgMGuSLseacFHel21
6BLCiXp3uTKyQyoC6JxkAmZRXCwrR3HTghvbKRYVIn1ReDh03JVGc5Zt6P4zhnwMZb1KsiVxCxsG
rZYS61K9/FwiCJn4rAWvMez3UPoX6FPDYtJDo8d2/WHZ6lf9yDa83TFebrtfXy3hvzK3Ay/Kd2rU
Hfwt63QGO8A+NuE0NJdaJPFLjAmEJplf9iOVJy8fDqb3+edwChqwGFAjR+w8HIzWHIT21QOOBROI
05LAG6eVMo1S89afvq4GQyFvWHJT48h/IKSUA4z7SAQt1nC7Idd9l5IDqOY60Myl83OgxlzBurwv
snMEC/7QRID4pb2s20JHBcxYjCnkVpxOVqUwfdGBnFDXSoBVXi5ZhyZbiUrIqG0r1gX6IkTCsGZT
PovhMY0+xfT95ml40SWL+yQzLc7n67UXGZbYZuKp/kvgQ9puiQbk7SNx1QWEDZQ93MxB8lR4IcBB
/saX2zehZo3+zgd+goxcWfc2AeVmnnpK5ZBmssRSdi0cl6nUJWGyqpPTWANL7RMVOEnOtcaOTF/2
bGMDTXc7SVKfCwy5atCxtBeFsgy9mNmSkQ/tbg9WIEryEQ8J3lbpfF/S5eO3BvyXgwc+lA3pApDQ
Z2uuZ9c3vZcccYw8Bj3q6tZdpyrvJ72Z2VW5IxGyAgD2R2HXBJQR1QWaZDn+OqDei1fHkOP/GkiR
9gDWnTTUXECGFaTh8CG1i+mMMnr46ZRAl+peqJ16cwaxCnNQvIZyQEp7eccAycBmFUbU6FWdPw8A
jYEFeLMVXulM8deVyc203VcpjGGUrIC25vPYOorMPtqtUI36AaKJe6EmhCFxbSzqR6shZd/9DisJ
49InZc2jF4vVDnsK2/kWsqk0KhoPqlKRnilyOWFAd3WVNIKvvV2KTggxvjKBVbOGGRn8uyMilkvb
g8tZrTrxFTBWamksy7qQ/UpmkJBaGhnldH+0PKS7/dM9IgFmBQqdTTO5E6K9yX+MMuU19x58TtS6
XFxHGuFwVLFRm0Wdz/msnzdT+wGkQC/wnu6Nstu9GHJlEyb2iI6dS7+X3XRXMuOAnj7vm8Qn+aHy
BGIij6VIi7i7fd5fVGbCvaRPYEwIFuvlQkIW2O70pxnjElw5ecNVpk40l9skVupd5HfXCscA5b57
HnMWPbtS8u1BNosPgClrUAF8bcGC8/C7lI+AlW7TB81jQC8dsm6zdbBxeqe0oR3+daR+EutoTFkP
rA68DFlDs6ikdvoYv3uWwq4GYwH4fLWalyaJhBXzFZp02auuA6X2UNABZIRQWuo2e37n4FsWwT6p
89hvAlruVT9Mi9HRKahPS1DzaSz3k0aRvlV8Jp/vjl4/q0LiQs0o7+i5l7f7u3ZiDE9/2e4gQyf0
2c+5lffEggHmhkBnECT8gQpAM9rsgGqPDOeZ2B1s3kpuCUGI56aHnMj1Y4w6cC8zAR63yKYCprs5
rI0cz+NaC0fsZ0RZQs73yeamFFBFDqbrnFoPsV59tQLr+8PtghTrybdMIYz3Ctk51ytQKQHKoUwH
SzZIXJSiasQeVXYKzGOP5eoAA4kXCY/JWc9UxkWNBOGJRs118a16Z/cH5JZzP02P+wRmm6WogMiE
wL2X64dSyF9ogP6Q7eu8bhmAJaR1X21yzGF779ril62GFG04NRbiRhBv9RPT6dNi3gVU7+D/xgYr
bZ0k/5Pxdo5nTqHGwBr2YaEt+Fw/SdEsYL9II9xUQNC06lE8Q5Li62z6Qo50K2bhcuhPu3aZ08SF
SXbi7wv03lhimHTNw8+NT1jnOcjfmpYJzwQTcyRqtAjQpOJnMjskqOqSM0ZiZCOB64JLmaqSjnDM
2CEcM7tFE5YRtF65Ka4jllzhp+ujx1sYAf+fDAb1Fc42Z2aB6NPKbgw9kREhoqBmZbe63Mwaw6lV
wvy3BnV2wHlAZr05Yx5OmlktxWSnUo09z/UzrnUjTd2uDdi3052EWDZ4y1vTzRnxZc3WlaVsI0g8
ThpePX0gd8/+2wBgXFoxC3UMdGjK2WY3lrMRMjnhtues4lHVtTTHEuvbnHEvywov6xtnrlRPbjdE
dsiAE+06qpDW2ToCPn2OhlG7u8WUI9cW6Z5FYcucaFasXMIA5/t0J7evqOpOPuGroTS8SFE0FVZ8
ATVdL+PFX5VxtslZYQvs86bu5RyvoqtcSrqT1TdCEU6n+nmtMRxvFEwIuwPWf+cer5GTsVfTeUPO
XDDbj5JXypLGG0Kc9GwpNEQ811A2yRpqwcDTqu2aiHHuFbFv/TpiOxzeVehDO5ut2njbdZjsa7iT
qBhWuiRCdmLP1AqCPbRGnuIzMWtQR0Dj4gN3BobYQh5gl6F6oYJ/qrJtsf3A3YbrHbRBKx3/EyWs
8dMLndTMfw3BpkqywGp8Uj/gQY03Uauidbexs9P9Q6HiPpyX2ZzuG5X+T+cmcQ8U1KVBnjobzNQF
izz4pi3NJKlYyGEN6WZ80lOqOnDnS9Yv6tzxab9vyijR47hDwvPi/JnSr0lVPA9bQ9tBH/ZP2Yi2
27kAGZLncRFTEhshjiFXxkAdRykrjyFM19fhlD8B4m893HqQcRTo56BADfZc1pdCnGOMJIctAsY1
E6svsakJvjuen8qyPs8eqYwp3xMTT08OjM6YImUE0eDVH5rcv+BwFINBY0eQUppYYg4D36SV9nhb
LvtCBEJrhiB+a8rLq/yGVBeTuogXFIFkPNaLfywwAjx9+ijRN8p+aiZWqgFIZldbjRIh5UTnUk1S
rqpJWtoACLV4xytG09TlYXssV3IzpucBkB6k4xZ0ewchbLOP6hnxkZiDokVtEs7ihfsHuE88brB9
T0RQCG4A8bEVzmD0g06CQA6s8GWDEd26vBfP+xTyys9r7so4rwa+zg3tHHMVRQJGFyJkanMkLP6E
914jzd9JHN76LVRh2j23MOVo95iugOVPK6DnEmhYiNNazuzj1PgfpCEsbfu5wysDpkvN1iio8ZS4
yVZxcvFxuu/6V3fH4fZddKNv0lwAK4tEfQVgwelHwOymyaHVrfEPvwdbkUmQpTCq47XXMq8XS430
rJZgZ78SEHHCj8VMjTbIfqDD1Pul9R6HEpcjZNurVV9Y6MVDW1I8bPFnrG6kVRdFnZZGtMTJiCQZ
JWUORjvd9/WbRnL/33nkreiVlDbpM3DTQWYMkOyGyBFJrVc6Fe2NbMRDrAeHC4CUQQmBTTy39KBP
xDqbh9+JG7CamGiGC0Jof9GdqM8W1JkNigzTTPux2IZ73VKnMYQ2ZZDUZzXYs9LXOjGsow0pjAA9
ph5znYdKzDTC1zYNNuPIzSyKlF2cGMTRGRRFOblh2OUcykjkksV/TKAQzpjfOF4pv8VFaS252Jm0
XTloKxP53yc/7cutVKXoDgelPS4TxaE9ScRqO2umrmaBEr13+T3dP64cC6othaPOKL7k8vrAMSnJ
QEtUbM3z/hCyvMQnV/xiJDFn+pxSd4PB9t9tblNq/PefxMX7pcaDgJmpkxsVVDfPfl1UcRnCnmM2
d/udfD5e5/mP+jKxdrr67Z6ZzfJb0HOLZYcqJV1CcEeV43V6jZs7Aq+W69uzuEj5scIM+Eb6OfFp
fn+xQc3aeGvAdnrtVuW+0irbPb9OmMocjwZPJDF4hDayWOaJTO5184jJlZ9SNoNQI7W7rQX6xiwG
1ME4Rgo6wgGILQ/GLKJW01XX7lt5uwyVZtN1NS/JtvBCPSUES44z+0QCmGCbHA76rbSZn2e1VURM
N5wP3MPgdnz/ddVn7rOBd+k1co8UpdXR49ULLlAgXDPRgcAY2u2ORaF+v/CBlgBgr8OIGZK8fqfT
4i6JsjegFxTT6g1n9i0Zv2ZZrgQ8avDdrWYRT2IavDkr/z5jAHk22CwEQ6B01RW0Fb8P75IV7PYt
z8pcplR3tdOivvr7U0Pe53+CH1JcWQZcIB3OpKEeT4YiZ9vsm1O9EZAdZI0WPZPOkIGOEruiOed0
nFaaeOcaMyMJxs2m6oSWCL8b0CcNRqEFAGbsq5eXFC5rMKQJjdJkppZYSPG58b7t92ZbNjHGouZt
4v4Z6g8uv57eyTgO1cblC8KO2+9amUeoranDQcBgWdfkK2HhWMrpFFbHwBHU1UAYwY/MsCeQvGk2
dEhruIItUgYOyfMCBhYGdUAHkQlwWCPd83OXRhndPEsmgmNt0DI0yOby3glK+F3u0+JKcYHy67Nv
Kv327qwA+/DuBIL7eva+V/iYTGpXSsN0V/N4coo3GLV5fZIPXcYFPMnNpPmXa5vW876CPRtibQRB
Eub5TzoCZIuIh9bengfztd31sSKUdIBljrBdwellQdhVkIIbD8E1DoPL7UjE9kE2x111lE+0iTBC
yrvzYtl4saEE4yYOdy1O5KBWDqP2KZjw4A/KyR4bwojsUP92QlUSFTClzJ8TZLD/+G4D4E8T5sdk
zTqwluUE5rInlH6ew1M68fDGv/MzRbw6+Rl4N0VpMHPhRVGvkHDcLCni5mp/4fpVDlo5nrOI58K7
QKwr5TVnB/JrOsTWVmFFl/kzvujL++LqP3+518sb6FAa4OuNNHK8SIYy+Vot+DUkizWd9+cdJPeh
ul/dGDY2G64AL+zGxRWMCVEl8yb+cIH1wdHkrbcppvM5ShCINZXK+jGyKhy82E7kgo27oYN89ny/
zWIPJEIcarkNrH2h5xBhOryAC+bnqYkvkO14VCfrVwBcMKF6Kw/3q9vPgSnEjC/LVQkVaLhK/8Hk
9sBEzxsUfAXNMFb79KuQsUdXVaSiXaokUItqYX7IPov/GCVjrX1VSVBlfZL+MJYzHcG/eq8Zltao
SVQU8HZKyqgyGwZK5oMNC7o7EwMLmi+VLuI9iMSxdq1vEwN8/56YqtjDCcpviaFxY7dRoChb+/Vw
gc6qk20ZGgh8rFW7e4E6MXC7IOqw8nxWavn169Jb67kiLlX663yZDxmr3j/n6PR60TDoOTcGZK/m
maowhx3zqnRM81u/hpOoI7dmCtvvU1JczJ0wHxRk6Bnl51/gnh3WOk6kwvRzLvuWKNQ3LC5AjNP2
r2vS+AuhdWUFej5QjH+aUhclufHNHDueEtkLcWGD1tekqryCGHGQ7ZmXSTpa89ZS4TNiZUq48IWe
yORa+jAb5dYeoHv1GzXA2zOYABnSD6839hu0KHIy1SZkvWs8QjmxMLOQAh7SGAG5nNcdqsgl1h4N
i02v1fSq4aW2uSDMyhpB5I/olmNoH4hY7Y9ezAkBab+BuF146H9EjFTFkekwcHl8nMIQuAgXKf1c
GOvpim2Q9n1VmakP6/SYkJMdGdnTbNmkMd6hDoYEXuMD3sDxcV5ATuoiG29MZMhWCpqcB79+Yq/l
Nt0DUtXMi1K22y5VD6lsRYnwjxqB8al+BdqZVrzSbMiuhjtjMHdMFmo/H0Xgs1RgQkabIAG2K65X
srZeYdaBWmhZpmrY0mmXGz+KNTuZUlOSmntnrCOIvMIf3gvw1TWA4BEtpivecW001NzXU7oZ2M5+
oLtX3TELA333RYAdwJ2xWphDkSYERpIz9c7Kuje0IN6CJQgsPS0dgrYwGdUef15kwQh2pG79/QML
KLetYQD7/q/IYExpf7PPat2pRpYPiC+urkJgq//NMbaEsGj2WNUK7kKbv3NkNMLmWz1z9yP3a0Tc
GC2EO5pTkQQpKC6VJT6FeBSTFrIGP3mXTPrRBc9/3/yxVA855m3BeSl9PYNi9wqy2JvQJbmZdnWL
1UCIW7H4By9qvnIm+lCmUjkZsWAYfQHMRvGQhFB7ZdAs+1BHOd4oSZ7UnqVV8WIHqJdS4Ja9gaEq
2O9vwec0NU84tD6D2dPeoU7Wy5kRWqD1wG3DHEIihQfp3qhRAxaW3ocNKANSoiyyiRF40M/7y1pB
wRDKpxhhYTkLh+UiTaeGQscf7iepnn5f2+SmLABr2Uh3+wwSH2NUIiLekqMy2WWB/v4Xttmm3ZUu
2kWoSlpRA9mqfCqI/FZ2M2DW/A9Ho9tqE1jb0F/LU8lVCrIERUvFKZYqs+NpsvW6QIG1f53iJ8FT
wGKW8V6sgwig290a7dG3NwOdube4rH8d17YHDQG9qIOA1yLF14l+lpw0bv/dEKjJN4vZXsQWHTkX
EHzVhDmZHtQbiUr/15eyA6q8Ew8MvVLilbnVPAGquXCpOHaRObPeU/fb6VSQbq3fv9S9n3B37fYB
EXU5mA3Y6fNqfnqU+yd1h87zG0a4b/IwInXTq3swDE6GnH4TxJp9Zkl+10AMalfcUdrxe4azpBjd
CuAosEyExIiQDcSBDR9qtVBbaAOVzCdPDXeGpNfw4uYax+Hf7GrMaPi6BQmXjc6J3cmrIs87Lh78
F4tY5LtN3pN1iExxTld7kAbIA36x9I3o/M2fEnPy14PPyPi+lx95JAviVqrS0CZPHAWoLkr3QQi0
Ak9Vmw33xDXL8q2vWVhsuHPy/wrgL/CD3rG051fax+7t0CSzDUtddPNE4gCRS+NxNhQ1sZrpZHLn
jPTX1UVmkfEr+LX4cbnvSPISixSzfmHRGEnZb4bT2jm2YbcEfYcVeDFAmCscV6rLwse804ENAK/e
yzNegabXcBKfBARrEQ1z7XZ1A/FciMKAa+jxzsGNBlwkSby78tsqL2q260sUykonIgao3D7XLRzV
f5bInAgx6lq/AqXHXlClOe8YafSbZLs+Oyo5V/o0cIwi4dlLWV40m2swkKeWeG8B3rN2L2ftcbPN
q0FTcHY12RCOiPQ8sCMs0AfvlYIA+MShXgAsHbx7IK+PR4uGAxe4PEeYLkl8Syo+qfv/b+Y1dgCg
23uQ7JsEBWOl1uyCmllCGlMNdkovIkM7u3fkfQXD2X5RQHcqZwaAUOrXMN6GcHSlkcJa0QwoDOpi
K2mRYHqSSuhrqhpaMc+lWNcM4LWLCSvHtg/mwqFKr6QkH2izTs1FIUiXj4SY5aLVyAbA34MqGOZx
mu6mcrnEPld2SsZ4l0SCzVJNultJj6JFrRm2bcl//8knKA6VtMkx4wYIIEgBmIejJjuFKDFn35xm
Pui+FoXYlGiatcIe7tsH3muwyy52xKzdwmjLnBSRFpNwvXH1S4/euKsJiSIcW3c5JGOM94kPkOdw
6i0xNWlgtsXnZI4/2KgpjcX+VjafALtJFHKD9RqL3Vrqd5VyPgDjX2Em/vVqas1bGAFdF/qW7GJS
WL5ZqCUI6JqUeGhqOrKql9Ml/qWpaf/w1vSm9FeapTMcuGw3RyZxr6T46BgyRkIwyqz2Fl1TU96A
4Kxg74/f+yf6nEl4K+eNCMEQitnweC/7EvwjXvQu5wQGBWwcCu2aJJ9GbyovtLioOX0QcgyZlJM2
RfNMrc0v0lNP5Ngb4WWgMyqXdvKcmhi2bDojjpjqrWLfREFcNhUjqdhlUP7B+urtiGkj6bJaAOED
Bbc4EkqlsN35rmP+6UV9dLoK7ob35nD/D42zJu8V3ACGO42uz0ckPTXE6OOMTjnNqSg3uKxZdnlt
X39EsfQ69oAkW9f+wrmTCLkMLK7oWeWRyB2yrc6fgI8NStsOKmrIkZKXbyrAczsHxYc+0HlOgdJc
yRe/2WmrNbzxyPC1XjdJ58j9OxnTTr/sSKOT/HYe9nczhCmJRfty1u1LXhpL2Zi37591BjbLgNK5
wIyR8XGeExigvvOsw/RmlrSkaBFitqi/jylkPfD/CngwXWO6H33bk747ddu71t4f067gpwEnE6gr
sQEbhafXMjMYK7q1y+O6BD43JJSDvvLmYyyuKX7jipJB/8YjjTLwDMGXFPs5z0SIZirOSjys5Cbt
EitHf96WXTkwIHGLmtEr39BKiNyUovTxg7mfKylvRo9qQxph2nnuk8T2+GrDy9SoNRJGyrRyuykp
X/5wyH1VZUfmd0Rf5aYyOxtArC5J/w7hO0Be3z0F370JgA0QA0m9RFNyd5igQs53cNZQp43rjPGT
m4XHKBMFhebdVqVhdNz6YCebw7bMJp/p7FlODJLtnVXj6ie2N9NSzg+6jEGK+j8KS+thrsvylIAu
4EpGzF14I9Qz7KLchXD8xfcuj+Bd48weVpbyItVuyABZbNB5xNl46gY23yDs+gzX7hjMuS3HalwY
nt6cdza4i26T18VzCsENAbsw+IZg70114yEMruBwEIhMxp9/2nvtZBDG4L7JkK6mS0kRAfbIQRcc
2hXvqtDldBgvopVMLw9yFm817RRdPPvCw18LWEkJ+IMytbafs/kJVaymrRRm7IVUr2JkFrkpK894
C+TQMSM8CDCm1HhVoPnuKjsOujZYeqkpLw1y98MKcr4dS/R1+0K7Qsz7VxiT6W9EO+IXuY8Egqes
ciHHXA5FGiIUzpMHZqIamJNIc/aLsPUUEpY4gVPZSSaRYabZll3+swck2CL6wAtPGGHauJvLuc0/
nwYYe9xFTlL/0ZsHE3DtqUbxuyXDAadRQu2FqC228jonZ4E5qerHs2S3F/UMeidjBlxNBnLw1V/U
2M3xWQmGOMs6Ip+5EweYmYfet8vNVU/nmnXl9TyoPHle4q09/IiDoDBOqM5n2+nqWxYiVgyIfnJf
a5kZh0m3vx3ut+zuIt3WVbK79iLArtSACbCw8dnYwfaK/Uao/cZ7DXtz1owqnzsGBMu+jDjsndF7
5ZLcT0xHwB/b1k8tkCSgTYNhaYW96lJbVE17381UcQ3SRNYJ/wrLsxXLbb0/Q46XELerdnC5hDwn
ElT2LirKdgP872tyAVoGWfBhgrx0LwapXSbKjMMf+b3wpF/+2wWVno08t3WqL/jt+BtgogXvbuxg
Zodh5wCJuy4lPs1UhrpMLRo08cViTKa68PnthK2xk7Q27vRO16evzJedT8Y72ZbTZjHqfOjdIcsK
WRVsLWLkzyz5AvBuq4BkSjRL8g+bMnxbTshhgX6BAumkYcE2cmgwYW2jtNLoWTsWxqLkGJO8BHOa
0Vsdc8xKiQ7E5aZ98uVlk3slTQmeZG5fttTizp/1WK6wRJwnHIR6atwvhDrWmWJ3SJydG8PVPssw
rmns+NzMKil/mCRAaKW4TOYnrHnMMoQszyPbi9FVA5ooOMJUp7J9mEEFSYe44/RErlQagOm7mzVf
pBxyJQTgKncAiF24vzuxRJGtkLmm/xvfB5vYLLtTZpnUqBkGgov4J6LSEvSIH2UIOTY8+YzsyaQK
4LkqHEZHVnKqzozv9Vs3pGP6ktbeq5LQwFxmMq6jamgMTDYgTO2n3d1xP1D09ooBpcoLi5lzZ8W7
QIoOnoYSicmeAq7IggufGZimIGSYoov5/McWz1oCk/DCrRUncEayp8UyMUMDlo2RGMoowi8Kxx0i
kj9tkY88KZQZCIm09W2UYBz/yJbxehaam+qr+MidWtDDNK+Feww0yvwfiH7BCKqlnbVnVir6nYxh
m367x9LB9BqHz9VbLBcFT9bVyChvw7xyscok66DHGuVKMTtIjGC+tRhUpmeupzQr3OppEUnlwqX6
trPiw0Yyo/0TpQMw58ouB9H/njVtEDfvzHEVZaVR7oiFW8QLqhQr9vyPBkrLs2dMchwiSqjeM7mz
glH9zmZztubdgsrRpgxfuVVwTJAsHCdB4dnK+/ZjRJMznVsjXUHOiHjOL0T206j1vR2IXZsMnvaE
IsQiAUIPP67nbtvRV0Fb4didX7t6rSUEZYrijke0YyAOsja1Y/6VUPIO4wxskANFKHoAocOiclKh
amlzgPYyF+rcLxwV4QPvwt6eh4GLpgGovJJ15GeZpp9brQpprKLw5tiJi4YHPRzKlqdCJNajrl1I
D7Em2PFvRlXfvEQl+HyyUPkAUsQJ8iKKcsXEeqZ4/sy0J6CqI+knrYLr6YBCYKLxEYxtQkqfwjsb
6FwsHVwzk+edJiXP/mIFzwPmykdqKH1jFED6P69x5c+00fXjpW//0dqfq/H69btuPPXQLd9MtWX1
n6ipqyrLwMrZqF+oiNGUVdqajJ3PcUHuvHWcAfwqM7DWH90yfvGn1/LJbJtJcPluSI9/ou1qR5ix
NKS3loganMVrWuVZC3l+UnBU+U6BAYiUTbkQW5y9O8OS4lztJDyOjnFOdsRzLAsoAt1W24Yi9LaH
TcBOIMMzIV5GMUJRQm1j2wz0Wavx0kPG7n104Kypbn8G537r1WZlEXXZH/2rp9mEnAu2zIaH2uVH
4vW+anW22GBDnjuM01/ix3SHCb8jxowsrohNIX+rSCTbMJSPqq4gixJJh3yTENvR7dgOukPsbeo0
q93NGDtkjY/pKhoXCY5LfSNV1tnOo1MfXopAJHahJLIR+X1JyZGHrf8YbXNfrV8UhBTm28WjCeiX
cL4IhGiZvoDzmbD/l+myybMo9aA+NKVqQ11eoHxJJWB4LMFFZCFmLuhqC3+9u7kHr4MB3eC9nVsV
nR9/ijZJQsl+u7Y0NmrJsCwt6BNYZVYvgFD9efGdjBwgUphzaNQa9oFr0lMid1C8W1m3Wsi2j/Of
mXG7gglSzAR0yXaOQ7kbAXCm3x2JtLvyJsvRWai2yCeQ9/k81X6eo4z646HkcXPMIZSs6cLZHXDF
bujgYcKkmlJL6SPGb5U4bqUVxlOUjQdPjQFqOZlWevNvFwSrz/IdFQTZL+ZIKIt1tNY+pgyFONrX
M4EtSqYmB1+HDaCwDhNa0+qD8L5BB5/ao4PB2kYq8D42M+IAvkkQz+dwNmUfxPZ6TCGmR1huMp/q
8Sh2doDuAz9bj3zIfgv5Y9wdIXYe90+bGt9QqSPB0/O4JlvJEfQs01IHWIN1a5okJmP5MnwArmOQ
aIyUfelewPX8MdjsmxkdE2Y8xdS2Q94bK79VeQFbZV/b3IP/xIGyJejQciv/oOMPra00O36RWVjb
9THCmM7UR1uZL3fPHDJV8rDDVvj64utLAYvcZW8J8S4mgxQWjJlZTJblvGd2XAMeT3w6oGSPOQ2w
L2cxbK0pOiJMUsswy6roKgLhDSML+1Ld/MSH/MDkYdONk2n1qztb1cXwKDnDQlxYeDIErAdaU2pc
CxbHpUwz
`protect end_protected
