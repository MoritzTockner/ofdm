-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ASx8Fqu+d2ErV04gP7wjZppibvGDwnjRRPnz+a7v29MRius/iykNNAkoMnDeij3fbayWVNFw49z2
tGG2s+KNBr3Z0/Si+yWza2DpfQnzd+Xi0Wu8/HFiZMPQAUreDsjr2JsbYHLve0MWUAOKQusliuFh
ITPSVGD7FObW5t6+ykCHH4DCMwM6KADfhFlL37CWek139V3RothniMBtYDAENI3RcWqo6TlHsDmu
KWruEmfuxMB5FYdhZEAvMPEivw3WszSvnISb+BU42EqG3w9fO7woBNGEb6nQnEcC5Hk1y0pAPkJW
oqzEZLfB2ZquwtdErWZ2hiNdV7vXkVCI8ayQYw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8208)
`protect data_block
NTiCIjPy1KhisRpl4vav+1VCS/hJusTPpMaeQx8SQ8T8Sxg4ZTqesSGlnejN74OO6NFkzRu8t3Kv
wuaG840SdLpKzzTqcYcaJS+N7CoWXqtny3Ruofkrmpev1WW3qkMpFdA4FuPLM7gjyS65ZNOmTh0Z
yRQ0z07K0fpG4cdBG4C3QNQGhy9CgMOIZpAoNNZXtMBQQ6sIl2ArOcKI3PIHfCAIWVhijWZsQPnX
iDgOENMbXkfMjWorib/uH46SwWwrIPiUT8uPVdROY86R+VDxo6fYErTrsESAEPSiklm0HQLNmf9y
2vrQypbAq8eTDUUMvpvTHlSitT4gVlPOrCeb/ixbjcYGTKdDvVwAASzSbJhMY/R1aShI1H0q+s2b
39+L/wphYr2AdUQYFhNrzVEUDojyaZ6Yc2Lpc+JBFOEZZpJ3u01hWeWPK/GQ0Vy3vX5MnrdK8zPN
TlrFg2KEXVepVPUh17pUZfY5WSCW9hpKI5PpY3NRqhvs4CVe24/E0b2gCmqaMCLNK5gHAk/noVzG
erYbjS0VZ61XOYu65FGxeJQNlYFSQxPGudlemYWT2T0mamw2JkFpp+srIVRAvbEDaO6ie7xqMcbm
UvplL8+sDIoYHjb1krLCictcbiq53dnHAAle7ex8gq1HxTqFbEBzorc1r8ayfWMkQVkIyAMY/0rS
oE5OcA/OQjYm9aoXK0jl2CXvL8b2iGy1xxGqP1UJuxGn/e9+L5OTh6SF7WAMwpw9tVJ2RqAXIy+U
TXtEOmSXQL3Pvx+gaQUkYCYeH6EkJOYANJv2+YDziwOUD6V2DQ87wh8xXixr0Z1tsx2IOStvctrS
W4BBKWvXLMYq5kPpoKWo8ottipYwXHAMVWBa3tzuBRTu7o5YkkK89WscGEBFuqVxtBpRgdTzS6FL
/YUhdAZL2eGow/PKQXRO8ZNcwBn6DvGhTaBsASR6n7bNvnCFy83vmRHoJrvoZ1NDMDt38Q5ZtAjC
gU6wTeuLBJo+72nhD/Z724M1moI30QqOxD2IYdQpk4ePufU7a3zM9e3tHpzb+ZQE2EyWZZ2nYZVT
gMxUfiPTuOJz68tsvWEccPEmxy4SQK9RJlsziohGNYReRWPYlpa1MI/eEMZ3w2B+AvNHWfedFGI+
RUTn3LlCkUin7F83gLqGOl//DaAkE1foqXg3kdp3R24k/GEczlb2t3jJuaArDVu/9kSCSnSqW9Vv
4M+SxkLEQpj1jlRu8ZJ6FtgXFz1QOfZZ8eetuoz1cUKfbK57zuXthgXz8d0QgOjjFtiKhKdIHlVt
kBumlw5WDJCuDkzqas6UPXZI53YjMUlmYvOUz+0V/T6UCDtdr+aUZskNwBuh+CUsFAcO77aFvSI6
k2agWGDCN6w9gO/HcRGxIIJXVFhpvf3zKlYbKLkvsJ6Zeo0uYSNwQY0ASkIGOKE/DoLL6hbmsSbO
ksnzI+bCCHDkG9eBv1e/Via8mGlot/fZx9VKRse8qQCZvqPJGIXmbuJeWFLPgHiSZeODywVcvIPE
aWNjHAOU0C2XY/w+bZcFmgcDcFjYsy68tUaohUVN0BZxZoPZb+LmXC/Ti7G9exkFZ2lrQsvcvKd/
seCM4CW20z+YMf+p2zoUq+p+m6d+1EyDkrsd67hIk7OB2dBwvLNf/OSGELHwhOQ9otlbGZpojnJX
tEzjGuPxQoZHk8GCmeYjL3Kd+n9LU8P63jWu2z0TfXyD26WB2nt7Qv4u9tq4PHMIeZRbNs/Ub7/m
Ek0IcWOAMrDLmugDKGwso7SsbhLdbLOtWaFcq5lVTjaL8DL3rHIkVAPKG763uKzRDbXakoQHtyZ/
kJOupJTkepvwNC/O+U8HYKJ3vRoi3XsRYnf/D+KptJNAfPvmtbq0ZNPWTYWf3N6IGshfdmBIm62e
rx9b6gmkIYXcnGrEEYW9VxzZ0H7UNs6einu2XkFP/VvpVbNrXp/HYXIdkwQaeS/Je+//eSitWLVh
3YYq2v0fu2eiNkym5EmlS5rpkPvl/4y9b/JztOCSO6bAokdThqqY6KSDmyM5ZJA3YxesFsSr9Kkl
W6OJaeqcYKXIh3qZLPf4olOu4yIO9UC3d7VPahMhHhKfIa1qXlmD5WloE3yLp2O5GJRh2d6j/ipr
UV/dUhS/DE3v0RMXWU7QwR7twDuIGT3/VQP5bJ99V4l7dYjVSpxgb6s+GeG8UqJnlCf0U9jaqm1D
citc3xCT6RZLhzb+n8xRaq0bY2HAX1EX42ud5kPMzxA7kr+YV6KSCCvzqeFbPGmpADcKpyG7ptT1
VNUvY8NOCU1jGSVdyu5ceZFmLeMUKq+1MzVCxuTeSrHjF9tkYrqEborpNPCrzUgjeoJfXS842O0R
g3XPRoEPiFSEHUAsvqAdHFdJLhALX99WtzJcB8C8Dc/XaM5chXeflqaefgAMXhEOZVIms/bvTEoZ
QH5O8GENZ+FczVLVEep0u5Y6wrIDDuc8qDUT7WzEA88z09qGzEryjkeUBUtKWGarre1Kc7YuICkX
Dprd7Z8o8uauts7sm/xxkpT5HzT0fkmYz0X092oT/KURvJkF1w8Sp5XGEZISHhVnU5/qvD61qz/4
Pnipt6bO7As7x88ZyizgfUSpZxlNeE9BRJ7fiwtfxr4XL268Jc40E0Et0hizsxPby1c7MHb0kMcQ
D1hZPePWuxtY7cwcfUhraJngJ35hW9wfV+xLw/xdvdg3vTjQu1oZx5re5qhAQqaMBovOTjuHznsq
7RRZaOOfiMxjU2nb3aZaBA5ZSNl0q2QmmqiXx4AE0k/tOYhc7K/HKYqeLz+kzYbKFSuXHnlCrvgf
C6P9uUfmgpaKNegm79eeqAA5h5AEy7l6hLgqIfuE3zq5zjj4381a0gZhEDy1A6kHlxa58jmdF7GY
9L/e134dpB1XAXuZPZhSRJzA+yKzaXEzjK+gAMCGQ702zEX3AyCLC1EM0pE2ZXCqMvHf4C5eBN+T
mhv53CxPXCfGDB3ol5d+gqxJo0tAIkEC4VuyWcDeGMReGUK6KBEg123NyNMJ++VqzlsQVGLSBdcV
P+iD5x5GGXcYU8UtS+V1uNu1LKk1e8e7cDCzaj4U9Dbm8hxao00dNipjJVBec6lEnZ4+GlHst+Tv
iplx9H45KnLe832T42F25Yzw4nxQhsFBsTIC8Yxtkg4pDJdgEiqyGte/8rwMbdMccyKb85mHZElB
GU7Zw+VJ9maE4XB8swVBoUuqpZjufD3lHthflrwykcxzqV1+VcbOJmS2++9so+L68CBJGifJde7Q
pXsqnVz7ovjJ1BfcgQjn+h7ZsN0DJY7Q0oG8lAO703AVUPRhBmEmuha6JUfcSgwTHtDCYvhzYhgp
eOkDFcdeylYNzBicFkB+/bntjbXEM0ycr/g5KqrNWxgUWPdk0mIDLByV7OiiCqhKeWvem5dTww3o
ro64LL3eMgV871xAyWuxxvt0fIn/SXNhqONk15sImKx9+/OR9C1tEXP/o8DL86iiz7fEo4RW5eG4
JtXeerKvoTWx/NMlNHNyrispsAoB4+Apcti3Vcf/gQOVTAjZHKVA71AD3EAF7B/D85qfebk6YzMy
ulSAyKy5BobcG1Mdjg1tfB72y5muer7o9F00Q32oDyZQCgobeC2PXTjzPLBA4+On4GdqJhOReY8t
zoWlGx2/L+GYbM4vkp2o12zNn7WIwqpPlgJnkTb9BP87GLY/LQlu8Kuu1zfay2hDH+kOGODDpfNn
HlNocMJaGAhg4FvsRyh6HOLmpqWIOtmhAyxSSxisGGK0dVXexYo5BWgBXMoiuSNtG5A3atn8TTl/
ESaoAeyftoG5wFADptNUGcO+d1ah1MPJFd9PWf/kKkGKszJxO3yC9Z1vLUL02THqj7kbXd+J9m3n
zABan/8r07tydmSMz9w4er225jz0YsV3Z0YqKiZg1FlE8NJjmbMRX9q0vYoA/DQ25moRXycTS/wD
jc1crj+78rMQsUk7k6cDQ5SHK1tOa/5n3A37GDyoTUGXxyaslqzIiGyMeMaOAGEwnZo7QahHWLik
CCQJ11T4UNBD8kDPUKthkfjwJEha7+NB4Oy83To1onZFRhKNAfu74pINdWUikVrBKw47pky3C0MT
iimh+D6L3iY2Kx66lvwqCr7iCEmbGECg6fxtivhiAdGpfei7S++8VeVWWVN8jkMtG5+3S/VPdoKH
7NNLOsdytyzysjQuWdx2JxyNZqrcuVn3gH4QZv3RM+yy5aeFQM6djFGLxzOfhPl9IuKFYCaks8HM
eXCaIVRd1erIt6sUpik1ZUcOp3yzVnCogsCNLF0zb3dGCXvmRKCtp4Jx+bNA3LAIKuYg9lQwAdHX
B7ubzuzb0FVhYyll6FCM5UcbqgaGqof40VcJ8Hwyv5bxZqqi1IgiqdJFChpJFwmxhxHhEKxIdBlN
WqcjoKF9PsSf97kT3S4exLWQApFXwmNPDgVOWJfqFlgTAyUkmJj704afp/1kNGPhO9X3vqrm10z4
NkHCv5ukb15pgtBi1xWixy78ck8iaHxJTMDIp6MsR3pOQzKqJ2GF8lN/PirnZs/isj+XqMEnbYak
6B8UqyXzrri0VX0MH4FwTJGOmD0j0TNTC3jjxl99hhGGvXWHMSud/plFua01aReSd6rZ4xPJzMTY
UsmoHu2bjqfMaTFlBO9GHAZIsaurNJB9eKPn5vuYE8sRPn0VvpYD5IUI/XPAQT1kKHovmreTlHlQ
GZ7XojeRk685wE9NJhsm4Zei1tlfdQnVEp/hNg+jhv3Jrne0VN1jLzCutF4diSWKWm1K2GS4LqyJ
P3IDJuX7jFpxBxF6TUpruNJE6h/htEVG5zhfkvLPPsiHRX0G7cEkyft9F0KLS/XE47L+q5rscEXQ
HzKgK6Oks6ceEoZkJgcrqE6WLN5yC5yNSoxGD0m4qKsnXHijoQKsyu7xKLfKJgSjSXhX2hVfjqUA
tW7MBwx4lihPlbZZUTsdDsYkmKFbO99AhGSKiC2D8bQyVaGqFoZuXlMS+2SNDzTh04KcmGslYhgw
XthITmYy1qFaWtelnNNK1Y7PoTU76Pt0CNOpM7wZlgWFTbSxk/KFMQ2IJtoWgSOSvRoBn0JVdFzE
oY9/DpwOumU3RAVjCEtANESCjKZ1lh5OEnU9n04EFy0+l0SjDnzhxa5Qu3ruNRcUbKRorlyHIqMz
8KJKYmUdBD0WcgUdpkWycmXp7zzKAA4aO3nAFKWObKnc5adJfkZ4lIHqg28IywvNAkb3dZKtoOHP
BqormO83k5LPpcr/J4S9y4Havub1vLCZZ/Tzp2GpF0aqY06N96wM/78zcRvOa3OsqrjP8ZPZ2c8J
C2G4OcgXtMrw7C7Koidj2Ca8BNyC1wPJeiCiWbACW+wEIVspMiwhbjzeN0tSC3O7xRGQDKAVgZSK
0lGV5Db7UR8xJITr8WIIE5hnYhl5VoiD9QjEjVYm9PGJSqZX23wozZpZAqCXMtFBOPPL/aNLjrnr
vdFyDrCIa+pce9WSFD0dcfZWD2SXdi3oAPw7A+aVGLvLMjCx3e/A3UyHle/FRbL64YEg5KqxjMWd
grWihxRkY3fFuvLE7rFpsBu9DF2B0FKklxVp1OCimqsLENVIAGaftHFb9SyfSWmDDoIijdhW3bWt
ce2MDwqV2roIqdM4O1yElGdLqitlCSLJY4Ti1k95UEMExWBNE1qXUc2qvAMiL1hq99pmO0lYAuRC
KI0ybqFb/b1xh4KvJir5jzKVVbD7XF7VV3cgS7jFzqBQxuR0MGT3+ZHQk6aPcslxTH8IGo4yQc7Z
CcX06W1HA5XBe8QJdOD6Xt3gxdVhofM9YX5INEfqVjiOjKh9Z+zqpDdybdxseTYB1+1t0KzVuzFq
BLOuc2q5hXsKQIvSFgoaLeoYVQDxf6xIBmQcEpa97/ubP70pzk9U6/rPpllr+pRYGYJzgUnLGM2V
7q1sq0pvREj8YTbeENOClIsFRMj0e6s86OlpzSvNm/9HfCxS2f/2p2sbiVKyROTFCkcK+v7xaa3+
wBEcNPGhNdyon/TCMyOPbHs+m9jNQnYXfa2ZRcYH/qNkd7T6C3RK0632zTl0hzK66lABAgQ+4hBk
RoTRbsnaadqThNSD+NXxKjdx0D3doIX6UFRA0JP4sOTf2srxBMRgYDnnNjuXO99u4edD6BCqR8JX
DWR/r81iPd/UCHiKDhzYpbTDjKdbdiPsBT13i41AjqTItuzCaW2mQ0rviyWYyRpnwCy/c8u4DA6y
nI1X6yi9M9nrZnOCNe84h2dGdqODBrrdQ0tQHMSM2x4cHmYlKzAjU0DVKNoUSX3oLVmnz++FXSlo
eO3WmFikN/ZzQsGvEYdmPK1J5x4ubiXogcIPTf4zIZp0zO5OYTRFYE+wCZTy506XBDPa99u7iUK3
Qf/gcaPFzyBReg51yd6+Ot4tAZcDh4HdYxjoICYwm65dOwSKfgdnvIPRG8qmAyU0Xb62PeZJ0CpM
V0MT4GES/kxY9mzUtrfz87bdDWI7uJ/gc7gOxy+vG1UA5WCGcHcfzHrU3s7uIX3XI6QcBx9VZ+UE
8o7eJr+nBvS+DYaX/OVrXweqXiEGaHG3uGWNmaGRYHMOnIE+37LV08801o/3+HLdJ23jlYVLzfcz
BRfUmg4cL33P+7mXEuTFOM0MqEUUZrdPL6PciDd9VQlEGW3PUMh5KNnQGfLnj8fEhdw+fBhc0qX+
wUNQ69jebwNbcMf0jURPZ55R57R1CRVR6Td+ycrURymPhRX86W/XPrTeasB78UTQtU3ypV4Dadom
ZRpfXOw0Gu9R5Dq01fv6Q+RZeMTfcG6CUkPlTumRBFPx6g2rF/W3WkNpVR/uR4XsRvNhhzEOXcL4
gmqFCetIAnS5xnreVfgLRaFhAhbyxr244k5hVrayWnBppw8RLiEgILXARL5mmzZRwxQAzRVjfYUi
s85PwOtnj+45hnvitPsdTjru5oUZa98laYrpxmBRZuoSBfUBLofT/TswIeqVkEj5Pkl1XeIv9b5B
1n0o7XIxajPI7HP8RPxEKie/4/B6e5p77cqtnd+3eJ0KYKTGpPNxRt1IvbNW+0uqDiILKn4gBB12
DPhN6IRYwl8tsMteVPbb8tNbkS1NYmEwGzgedc+DlP//ji8jXFcVALXcYSe6KH/SFBDODOvY50m4
qwnu1H2gMFVYiDYINGVZB99GvSgbGBEghIC/IFZ019/2x/5iEAXW6BqcNbWvUP0oURBOAk4NHGKk
BZzH7oL2u1V0y/9FxLOTSyBxnFU7cDU8FZJa3NOiHn1/+tq+EW8fXMLCMCcMmLpu0TOLzxGtI3UZ
oLz5/CYfsCZwk7f8qIJaR7T6mVbl6cFQa5/csH6MfokBbcN/6fsw9PtsxFpIL82PCNB5ur4TksTd
vc1+zQmpBQtfm48oH4CkG1SOcuK+ZmNubZjZ+8MoxjS87IUtAShWjlwIUSvZhIV+kJ6FYWERJTGK
5AuGJ2agEViRCVN6bnHCbgWNeeaktgQTrb+mJMApAam69UNCWXbhebNw8/fUsY49XBSMdYc7t5sV
jPClkTgRadnm5xy50yxjtCVXLPEEriLRZzgxsawojKPV4nGTWoYHHraxmj/XSZDqLeshr6ND2VtP
zL9iKaeXgbEg6RQMOEnH0VlZ+bFQa1baUZoeM0nPZ5ziF6AuF2sUuGZKwX1ao+bgS11dFEi5tyNb
ZjYfWp4mPjsCb8JcJGrtBxvbZclQs0/vc/T5URL80LklmBEzv4AD5jgJJWW+oUh4OienwSBbRpri
KVv10BymR3Ene93hQws3X7t3eLD2XU43OLv0C0ZC2LNdEtBhCl0bBGXBXj5FcTihleLBMMCx2ePr
w2LVUZVu5lmvW6aIkMlWrP883oaZVmVYIWS6f03RgXfu9f0HowqFW2V+/IyBgy9Cod4vFfHPNjVJ
JKCGTSzQ2HXx7nJeY7MmSMJ9CDi409Nx0s7SQPODX+6+BtAFF++C0RG8RBcP4HTideh8t7P2kf17
FAayhkbs/+3peaZ+OhRHj2m4+suOOIm2rrAb73bGm7ffKbqYR1bdpTMxATqKUoyUg/ngyD35GzVL
rvtWeTSC53N6FcvW+3G/F41bsQQdbflou6vIGyZkIeuuNqBQO6MpNtHA7UbtQ05uZy3BBPfWqTUN
NWM7MyoIJsgZCpRXFABLGKSWQSt93/UtgX55hyL4wWu/KRuLpMo8rQfiKLH7H1fmTuCO0pIb42bh
rb6VgMpYMsAFeUP7OKMEL11ei2DV+ClaXZW/GE9B4izfRC4Fi2NyzvMcBN6z4C7BeNYe15s9TEKz
+cZvitQAgPSeQ6ekiQQuWMVZiVDpWMrFeGYDpwF3xFNhM1y6ZldeWfax99lkIqpWxVMmoqTNuq6W
d8ts/vvDAhrczDrS9Wfc5T9qx/KZ3Pu8HRZ4eCVX3ezeb8EvFCz5Uqgonc7BBelU2lsYlX2+JDOj
iP6v2ETbVIHeF6IF7Fk+oFgz1dvlUpNSRbLnAjFny+6duIbYEgNJRh6yYAaKs6BW4Ec/nWLU21V/
jyMhy8Tc/rJDvC+xCFCaLNLiB709Sm6SRSxt49+KmwenOi8USY3Ikrrz6B7PJU5NdXh3TX709e+Y
4V+EAx+dYjIfJwPtS6isUmG8xqfRBhuS9pEP75m3n5/fUrah7bSLvxYSdyYibkBC8udKwSzsxk7u
fYKZcxgudYFqj1hL7djUg9bDR5tWD1Q2GGNot/zLPqpqIKuPKf5sJWp4EgzavbazCEDj6QLap/hW
f7FZRQ7BmGtxWFmltl9owp1Y5ZBL2Kty3Mo2Wuzx4V6zwKIsvxAJROyXe/eS9EYUUBpX00xDZQTz
nUU7I7xSqDZukP4IFrdzO4/ctx7MXwb8CyZwX64Yz2CD/QDtR4gU37P2X7cowz7kfZ675oHuHxK1
jMvO4zqmL3dsk9HXh+AESKGmmwasvzv2Hv4GnjzbaGTAG5aZ8cGWstnNVosjmgwqc7I7F2eERwO0
3Dzgbzb7TxmDBWcbKhDh9xs31qcj9kfJlE65WP2RnDkoAN5iDnCE8pdf278TOJ9K9oxeqdL9gStm
KbVjXak2Jd3qBRqPbV7VWPOPwnfgH0Tvx5moOEPLK6OfPwUZ3gMJyY+kNTw8RkpK6mbSRctAVNin
GDxnHvR6GftQZNRNI5/m7LQmButRaDPxmBKHPk2AVRJg+UmzfcUgYbG+VQX0dhKmcbIIjTCLXGlu
B7IWx4436+6CijONt66XtOgjikMmtyQAK7zD/ezDmqcFTEtXWu8vcpN72MC35G00E0f9MQJJ5maS
XQeOCiBpMc7NuTVzjPwB2NxFh1D8W09hZoBGoMhQjdgbwpw/tT4vKS8Ldb2TxCftIeItXqLC9NaH
yixq1cJQQdAZmcLCzvftNCmBy1KMrXCVIvPjF8bG5+KZ7O4olmx3kjuoiO1zaAZ9kI2JAQ8XK9tk
weaiiYTj9XAu87nY/xw+T8t8clFy/KZLiBqCg4V13aDflsgCMt0u/NmwHZqbELTgmeQKdd2yPQqw
NSME2Pz5sBU+k761E/s9urWmDeU5864ZbUnrsei6llu8Vm98c9FbessjJetNRcbcg/jQPLi1ri35
Gn2eWaMOtMC8vfm3y11snNla89i9HAKRCop59vzxfzor7hkgSegJ4J5s69phzs0x6wsbKtcO1NBA
vW2ffsg4C5vnsf5RpsYj7zxMJR3/TAXkQ9FTw/NOiUBNTKZZVIFMcRgUTyPnfdolu5BtocvUJV2T
4HtzLn83nR484lz8BBzANC4ojxWBSuyeWhS1U9XtMemRKyW0BQFzzprlZWXQ3IP756kocyReRN73
RMbAXZUmKj/FVbsiVDZXB8FXO7FvWJFN2a7QFsMvo092/B4wcZH4lrEg7mMnk7VK4m44qN/qlPOn
8hncPggMo0afld/tb8Gcmmt1IhbyJfq9vk4gW7wj2vILmY0tM3FtWU3ry0GrzeQpesKXqCIvaf0k
+Chv84Yyw8w+hw5BnYGtpAT/uDSqJJxAvcpzMwy6cwXaBo0MblsqS8SRnSbm6ZADm0iTJjAihVQc
5eA7mqrswfvhXg9yE0ScFoob61VBuw3SJbAa62p1Q3ndb+HZD8NyutbOCyRps/879bWt7GlLH+AI
q3YE9/Em+bisuwULtx46QeSp024XIc5YzkwbS/81htDy7ZOIKF1315K4To2uFj8nxjiq7xrSOAkp
bBfvYuNVka4DvVwVfWA3ZJ/F1akhyb8jbVOib1IqjP/M+IWZhlMF+i93EkgEVpHbQTnomYZ91zoM
rMZ347I866X2JA4G3IRIBcGGUgNZu3HD53TFpvjXWAsZLaa92x5Fnx0yMFcsFKEwfB0NSUzNnMcV
tQ/NjA1MisXvTmD7V9hz/gW7lxzch9T8phxo/dQKzlDCpkDVnvmOnbzGU0E1RLoWG47KpFqazJlk
DsQSggzlKPQYGyJLhZJoD9tTZVwj4RuCUZp0dQZlZW296mK6lm0suTsaRtmEbSbbK3paWtPH8PDn
ZJ+04bIQUX2VhG21g/Argj4/o/BqFKV/bmaGP5HkB7JuP8XbuSMj/eYlKfdJWnA4prHJLgI29mxx
M1kpktDBJtd1xwqjjF76gcwb6ZlZWGjfrGfPHk4pSVbGzUoresBiW7Iu2NNK8DKkJTW/8OT3KFGU
7b54fALhPkiE1xx4r42gjnzBZtfGwkmkiaqFJJr9SR7FD4grcOCxjJW07XG6AT1F2LCVfLd7oe7Z
UgzyA+Pt9Ftejce4oJ7K5WcCkbmiEzMrhjeeafzN8k07K8lxdVfJFWo6PKwaNjg18zBTax1/Qdp6
WjH+zan7ZPK8rybknzAZrqWS9JxRdA/PtagzPP5wP93bpTBUqClOBJUCfDVQqCIddptdam5UIcsp
rlhr1SZw1ARXtWXhw6J9Y1u3uGN+3pQE0orsx2pTaODLZopSSn4Y6CKoHqFyfhrHdGBAbkw1AVpZ
`protect end_protected
