-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
q6nPMlyDPWnH5KbtLZ5Z5Urzi4bgBDxUNHEQ/uHd0Pz2NzqxwfrPtwhGrIbWPtanzHdqjDgs3jMZ
93W05m3vFShzqv9q+ZF5XNFvFN2TEXHo8DV2QRFPcFJQNKRHPkvNC3/R0OzQOWFITY9YpdavQ7w+
yWjbInYlLW3MVzZ3K5tqJ0ebdDxAIfda+NzkuEz1SXso9pcfyWoZ+N8XjMdnWXObtWT3iDeVpIOM
7MMI1bE+st14MPAxMV6c8aTl8Jr0s0jkehvmzN9RUTQzH+VT/TUQXCFeNKmZ3lvf39QqanQF12FE
Vhx0LqXVRG9tOFynkqJ9IJ6wJn4elMsDay5AJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9600)
`protect data_block
c+gDYeHFFW91uD2c00dCuGo02lpq4dmXehWPAgBll5zGt0Gvz+SEbm39UojhA5vZVRIWwUrN+6Rq
1LSE31VWI14eNamzYJ+1nDmWRvSfD6pjrBNGDNrLanvTxMPQv1CpMWCPJVntYx6yzUcVTCJpQv6F
ipiVHyX6au60VBWgalZed9+WmIm/Jog19O3JccJ1t3yqXvnERuKwtX62+j73084PCqIjv0tB3ZBr
rq6pE5hq/Ko+9uFjqeL7kLMyHTiYN9A/4ptCPbNy2Hm4fQoYR10FBJtvMbtpl5g5YUZ0o0ez7xkO
b67Mfr3XA1XIEcHZi5ZrOambjfYDrjGufYab2W0YcEhX/zqVBMQeXosdgHTHyB4Wr/KtZeTQruaO
jAw1yLVlRz5gsqKRKXi8Yug38DqsKdD6dtpvMVO0j6TV/wul0t4C2v85s6o4AzYfi/VNyvhaEcuf
P3XK7mp5MvvwauCwLV+xthXa5Oe/KS5Vji8QVkuCjDynvD44LU4h2J5798cDYrKve7aixna8VgkJ
ZY9SoUUDvkPmO9kKRHdmrjLxOYGlMSteoCA+2Y24pY0FrX/39d0MmJ9M5rQ29pnhjdkL9xsG41Yl
4lsUGpobIVxct719tAa8GJysRaQqT7I9f9ujT+3EyrSzDcD8ai/oG97r26yrRD36LJkiouMgfbLQ
2HcE3buy2tjlcN69QLNjewyJmPUFHuG9nhAOCHuA8tQn7UX5tzXo0sR4w/g9iTz/HpaRmIKifVZ7
vW+pm344h/YdvXhpRj28hdbA6KTw8zOmYZGYEKzqvrh+ac/vCz4z5cGujS0ehcD+vQ4qNNC5fbK5
H/RZaWg4m0FuY92l45XQnON00C7WK4DaRxjLwQvTKW9bZSrFRFyMdAalkG541OOqVKJPPbaJpQLT
Ds2i9/EIk7HImXFWhlQav5Rcr6nXixxEUuLsW8bdbJ18rHdSV+O77N5XRJ96WVpNk0HXvjVVRHGt
QrpOVB6rLnlM7GKsJcUxs6i3LbXIGNuPp5Fc3Br2BMENK2ZX6jxnpO6XN8i814X6kQWfpsq3Hi8J
LHIw2P3wKadIwbbVkEvROY5Gdbn4sMgHlDUh0Rqln4s4C5985TH3h2vCGHXFgfRTCgyoI3gCk5j9
qOXraXrShndG5+9cecvQgaLEfXX5TjEKshLG8eSEGY6KJbgVuW/arD1MlvMKeofC8YqvfliOwBw9
t560sO3qI/mjprcFlFMaXpHmPBNG2UlKKmzFhcXzH4rRzAoUCKefI7BzsOzAlIiWGOJBC9ILJw7W
R2iSWA+zCABLrEMF+GogVyhoUdgzNvryeIUtr7J5uHLMPJfknidJVqH8vujQR/iYbLw/On7a85xn
g8h8/OQ/VJwJuXuxWXsEpQJvPd/igqPz565r8aWaD1WE5W0na+DqAfmZmeTVdnzz5+OSU12JO0IV
Lx1rfK5n3vLiObOdpbUjoCZb6+R4kSONm0d3EZRxQAg+Ff0B1mBpXchCkFwjrZz1hZInP4aeQ75j
xjH5DFQ5qP142ebxthyb7fi+pqgmsVMoWPT/ugtMGPu9YD/NQz2uE159w5w+F2aR9pLjLhfSZo/g
HDPPlKn7GKzwtkoc61g9vCvKxCoxDqZ1Xom3b4qzRCsKO+mq7x87U8YHMC+/Udkih11/vrDX2uX4
E6NX26WoFabO0365OkGzoIPZCWlmFRgG/iLjVCThQP7sOgcNdB4koWtQbflalRbFBMIp0avc5Gu/
bttnlQsqeiRQzH5MXDzKBXM1pTdKBmG7jYNQ3PNqSD9qjFVkzXJRlz2X4uR2Lqhkc0pj8AVkumJA
WmKZQUtIkFWErm+6++4/K9z8cQKufNSUh5u1PEngY3AqqlV5DqWHlWEZFtKBKoyn4k0dJQE1UX62
2aKe0NC24KX6KtVZaA8j/DYkR1djyqeQB+neVrCx2j4gU0DgcaG+LW3UTkXHEX1K0tCSHWAiqBdN
tRCjCW8Q0eDKQIkSvZu36VdUPdRhlYIS5FPLIZs1oL7GqG5oylk/aTY5rQsoBQMJqeKr+YveV8dK
4NhN+E9oVXXJGo+vbfvRiI/CITX7mU1zgwcp0lTxs7xNsnDRMfbEo/s5pARdWdRNzl2Zo9fhIGvL
qw2bG45apST939DAg7ljMkwxp07pIFpVKv0YekA2nMv37hHSi6gvjDSqdhRMoz2HvZ+Id5/Mwpdv
vZrWJCIKh967+4bXW2UVYpG8BiSD+vTzcmO7WiILEu34m+Z6HABXGu2T3Py6rH4/JGF/anuLDu6b
JlOd9qxCZa06gTKH5pmrhxXGGz23jlvgoKJejnRSdUuazdpcQNhCsvHVn48siQ3wbYh25AGj6q1y
GPgeGG2OhyXfnIEYdDs0SSVFzSabA2VTQQrkAl4cr5+pHeRb5wf/umMqxBmWREuzTIOjJQed/BT6
QKODOqafcNsgIJH2KjABORdbtpoYcXFOHPf6rmmDTJEjH8zeZWUkZcYC1ABf4okvMLJB0UX1edOE
l5OvN0YpyeJ86OBQOuUcH7ePj+FFtHe3haGkO9RlgoqvbwiEfFWkRKOFPmbRNbDtWLeEnCmh129H
wRks3anYOc3EZ4s1aUFgS8/9LAqBxXIDK+x6y8Du4FI2EHhPdKhpKB3PupXDH2HMTROiHP9yMPXe
HE/pw5EPg3jIKSv1HoyeG26otKNySg1eTGP5C/WrkqLFOSgARg3SHJBAr6Nj7evvY3H1qtfxcRF/
m6qt648705cAMIWGI/A5R2Mn4lIKZXlFeHTyOZqNdRaGseP/VqCzqdO+0JHczafDi+Gn1mSgIXEk
ONbj/HDPiUXWz1epPzD+4WrlOgiZQqVfodsfJYqM7nmJ3jqSFqPrbWBLc5FFpILikArQj9+Lv47D
XkIF4ck9ahbe22NTNogVNu8iLtnjPm18aOQSLF+Ik9NJDbpGbVniGpyTSy0oDsuve525PbFdMZoS
Hp9mCMGOqpi24qdgmiqAzSme3nWyTl9gwmpyQEIyeOAoV9KZhcVT7L2whq2ILQYMUmhooJYVNTLZ
ggAjUCMvAejWqA5RVgljQtsYM9G54tI9QDmcVKZfWsQPPxKi/0JJbL5K92Y5kXOpqmdeNjPJjH9J
zaOVoD0xOAPrhsmOkpfK0FWJ1s0xJGv9qH8feuw0yKMAdZxT3Br0Qu4JJUTxrn07mFMW0Ny/H89K
rQf1Gv4QY6QJLNcrof3d8pssLYOVTQx2VCJ/uyQifnoF58zfceon5L4fDV+gkTXE5pj1w9VWMQlm
d8Hq+MytCrF6Sya5phkHak9aKCtg/XF1tgSx6TkPNgYQglDgZDt3c+jk5FJnmN5gCUoSwPPDNpWL
jCFpGQpFdNzvfWzXHxOOp9stKElTd9QPkP+moUk0x6ARas1vgEuJlzf1qjK8cJvwHnWx45jwKlqd
es9WZzqtjpbi3BeJOczlluBQG1JqD5ybHNAzWZQUcHtfsMXVCk6Ybbe2WWLHV+U25EXRV75iVcIU
z/ZFiq+rqgomvNm0Rwu/FuQU60j3zCTMOquWHPVsaZZayUIJNN6PFCpp/GeDIrAbRLiI5e/ZRIlx
4IXxWrZd+fILs8qzOTIefRU0s4fWAepxYYnqZ7EOAqIVs++JQGRRcORvSd04D0rQWYjle/4Mxu8l
03fp3LFlm4XBuxcHb+zEBMoT2mDRElma4p9jYl1zVm9Rl/G98l0lq1yAvTle6NhXHPwUjRCkwTCT
fNrjw/URToA4c/DaKCKud8vm8SGnmzh8u5IXylHyvys1t9SRKTUZpvbHET6xrTRdN0ZccZssimG/
4MiQQqgzd+vdgS51NLxL0x0cZjE8tZTV97IhgrZDGneCaZRB1CFuv+qCdh82All8F+T9eyN+44rH
tg62+MfvMZxtuqyZYb0yNz0Y3+NlLGh3+adXXTRKPYimWr6vhAEuh2S1ByM6z7p3mhu3DnEMkGw8
60XTLf5ZabCOZ3TzyQIbErb5RVoXYcAHryom7+DlI0cz8UA0JDrHKhkA8N9Mo/kCd4dETU7GitAG
QHtIIeRVsKF3Q7QBMCjWNqX0fvCMjQfHYkrvpC3eqBGH8+N6J6SFrKmag7l5BtbTwV3d//CvytTR
o2zqbsnOFLlpwJUMYF4IdwBuGdJMMGS1QkYa/TyCYCqZ3J23XRJykPX+FJklSd1IjuykzlLNnZhV
lTo+6Cj1rWeFRrbxdVjFurU7Wun7cH7WQVXdQmbEMwdiIwsI0wZxPykMHzguyZkQPGfP0qH9Q6V9
Tr410pPTeya4DfKY2VChEUzlLrxrOfbe0G7743OSgsqXlE7QW24WWaDK/Y4p2fzfgBF4Uof+mS/W
94LdEKHWTXFczQEHbP2Hf3u1iLm2pdHEw6exUom7tqfHIkQR+kcTIwsFev9Gzy5IvQgX8vNAiNu3
wlgZQvtSSvPL+XTDR7GXOW4z9ENPYjkL5HCf5A5r8UqimOnvBVwdBN38NWG7msSePnC94hvKAyi1
3QokrECMbeEXJXqFyvzmOY1dRvDgxuU2XYzmOo6DNoIIiMn5W9l0hioJWTFK1FNLCdFpFHoxOSFX
bFb16Ik3oYP23zyogsC3+UQpMNIs25umF+ylk4buQ+SEvlVQPrn85MwELA0d27s+s1lgkaFLQSfa
21y9L5/x6ssx7hHZKjJ+xzBHe18gNy/XITgnCFbWD2VESC1E9NiPkcoSBhPpVudWLAkLENG0aOx3
XWjo1TNEOwLdRNsi5Q0eLAztk/8iDHlxiUjUcOdniFBXnXFmm1hsQDLcy4F1orieUQ8miUyXBjIa
sl503A6c+PQy0m7GWoTmRRXwqN4JhY0hSh9QzoiNcBtUFDP2OLTyPIj1NAyX9KcAfsU05VrJbYzH
J51oEhccTaugPeR0c7fFToaoo/5wG+1WpCHi+nX6dU3hPuKjA6H7YVIJT84Q0V1tw51kenXM2bYp
IFWIyZqitZIgWwzhRJnCfA5sCf06ydtlTd9R8TptPkECqSyuMUdo1eK6j1FoShRJmuo00ha3yqKF
8fu6RIQ2Z/NVMYcP+fgUftxKltQztddeY2O94mciVskl8vpu8OSWmP9hZovAQD5hskE9QqpfNvOm
IN0VhwbJkwNYu7nsfv7rhIdCzu2gWws40zKZ0WLWbC3eEVBSlSGxcVNeAWc4cqREYeHUQN7SFysI
cVej88UfhJV9L2tLpucT6ziw2Sr3Dr7w2DarkkGPmk82D5lAuKVja4CNbbvYI4XydPYHdMcFV7u7
wfdT5iVWIDQ+VcZHkp+U5QeEDK6o+mjypuA4fX7yTMlGUH/r3HbW7H7grdJi39/5RmMST4D96AcN
VTWXGG5lMHXQvsFsWnCfB2waHRpqsuX8xSbfjLwmE0MDkYD3yNCoWpvtWkcV5d67XS6eSZu/nt5b
XFupX0REKS5RHhoEGdSeK2qkTHCg6ZKeMpvWoppwhKTAqCPeclHI25KgWOknDaiYTLrBbRnovs/I
/p5LA7BBECJBlxrPob+QrMv0NznqNw3P37Lwd/9Og2s4dCiWNIWf5toI/+tiyC8KK8MLtms19LAI
IClOgyCSJa03GbkA93nnXF+rTNCGFuXnECIL9wqSnGNxG4X8ArJ5aHwAFIccFxK6gL5WY3cctZo6
l+bU9GfhmgaYWOvX4Kgtljzs589ovb0Atxqu3xbnKbAJgmPUoY//a5bVQiMsdjke9vEGzuzbVd0R
Qx5vyj2Vv1pg12hQQhSBhigzK4a5af8oaZKwygRkv4xO+omSMqI3Iu2Fhzv6GyajOlc8WLjJpfb1
8E84b6DRyq8JLykgdzhGKnspJ1VVR3BfVkdb4Rw9sA5ddj5yS6XsxaG0kFZgRQti6QX8nIe0y+SR
I/2XVAhEnljmRXGNi7BImFdPDdvcWj3ma5IsqQsC7eAxpwzRk8xw15ViluCRihxAD4yUcV1N5eau
6RkHMPTHznAElN+nYWRg4pKaG3zHvg8+kbPBrisD64tsWInsmJuqHlP7JNCGKe3KGMJXEGT1dkOw
Zcbsh8ou7suKObkPzdfgeNFW6E0lKsDbYyK9/lQDLgFM7k0xMQjh1/bfHjEaggBXMduaf/aM2e7q
kqo2KTOmCKJyisTaK/GSu8/N6e7b8NIulSMSKHWc3HlEwtOR1JU5BZxmzG9uuof4M02kvvNXTXsP
C37dVKGRjh3tJ275IW6m0oPVJUTy0EKGSnnHoEN1jeDGQRKmSDTETjemS8hzU8+XGtRxrpjrXVak
LqJu/F07ISx+Bi6FM35pp4GmL6dPmGOfJOV2vkcC+KqWtOywbEChYKWHa1UYeeKS6Lq3DRpmCpkY
dL9nt8KBRe/+NcJqh4BeJ+XSB9tCABg7dHp6Ugxl0ZQawFIL0nuQsTVp2N+S/v+GTSuc3s4lUOJp
+RW7zQrGi3GnDM3Gxb4jAeyB46y5z9kLSccfzJmpazSaohI9wjJCJe0DuI1biwu651aSRFd94Ry0
QURqo3fcKvU/kwlRpdo9Gha7a6lYnLfPS22UKss5rsMNbB4fqlDn+lzOBNdLTkMUVOPjZ7WtZF3t
TX1HnAUtpC2pTfR+EJ1fQzIEyjL3NOIYp0/LDDhEv8FE5HKEmHKxDbPIR2eVSvzbV2X8Z9RF7RF+
tqiGdFn/CipPsuchnGcp6rzEUbQaslmgPGaJ1+F3atSQpnN5TtSkDX9QWKQwKT8AuTY0xJ3YA4TG
cBDacBFbp1/CzNgTvjARValCApFhIHIGCXEUgATONhqzCZNu2M+QV88Us6qBExTl4jVOlZsVUVfE
XLa1t2WjQg7g2qh9MY3U69CQZr8rFnLUYnXpjMnbYrbQPYqZm1yIk3Hhrvj415g7OMFe6WqMwXji
H0b/nYomqP5sbln7MgIkPHk4c5DZ81WV+BQIPNWxB5/0cVhxxjByMJSVh8lzxzfF7ayEPCleABlO
RVuKTwqhFUNREpUFaIQA9llvEFJ38qjhLEgBjlqipLiGMR0TRVVyPaWa2sBXgtCt4WcynHmt55Em
BZeI+a6zPobGULNHyUqPHQE1yoQsgLr/agCC4l9/fpI+oe6R6YuhbXjS/jclgE/iVZljFLNj4l2q
Hkbac7slcgZ3naDv5zTqT5KpXrY73wRxcwr/vrvqhxmcKyw7TCYl+wHG6lWtObsC3I0PQoXGPA6l
k0/wO82GaqSFLW/xB4nd3P110v+QwQBT8r4KRvzca2aPUgkSONcErWv/ZrCkyvIQwhrwF/15rAE1
9hucOKY/v315f9vcloyy44DXp5TxYuRWBKfq8zf6i1SR52/mN8IVnOjP6+LCicX4CVFIkPOvhqYI
/eaPbLL+wNqRXE8C/8DzLTvokQkIw4MbsKfuLZZIAKE0REtRYnhnJMIh7UC+pskEziJLVRM3MVsg
kg0DkFMwFihgCKGvwOZz/i42jKsfpAUtCDkJCpbQq2E1vFFMLUNDAqwoYqu12gNOyZUV+G1C9Z+p
x35ALH2bfs0LhKE/bdfLkse/n+vnJVJx11WIIhM+h0UCX72JGCbc3qspNUqQUjq+3eB+Hu13Vi0I
aROwvua/OeC47oddqUiOeaKc2LAOGSVxNKdf4mZLFGa9Jlnn96oFE4JMnPS5H+g43037YPh/HI23
/6JLxA6iWlMox6O0AVHH3jTsbWzkdyTN3tNpg+esbcjUYhnOH7VDKyozGu42cyfUXcselBuOve15
HIgaN793dJNVVxyt3ZEfUcVfHvA6dl3S2sjb/teR2KDg1aG4agtbgV5uF+2AqMe9nnbBVxxcU1Qs
CIUEj6bjblfHCmaHy4vUkjMsW0GLNe6GZ0yIKUEBj5KWEUAfmeTfg1xqIsOpZWzmPzPl1hasLYVw
u143LAZiI3EKhHmAsbYBSH79gp0Dp7my51O0Mo+IY9iNYPHheOpKJ0bkCUCQiOo/5jFavk8QSVuU
pBEtK5+LIPt1N6lKcZCLp5/iriA/KWx7yHuIDJDCJYlAKTW0mZm8wuAsTXXOi7bmy5WvPWM7wmXk
IGYTW63yU+ZDwOrVyXevWxcDVmQMCLldh2P8QJ8ZQdGOuBtV2fp1vZuWogt9q2bvanIJqtYpolfx
SL6ncd36EIHUR2lCvtNx0YbF5hOnPXVMpOyCqrHf7xh6L2RI4AQx4NvT24LUMTZRVUCe6v5nM6ws
bKLaj3LFSL1lGaIyDkfYmjKnBHDiUGkwNfTVSUWaKrQsknTRXevteSVeJEE3LAfbw+9uhCg00ry/
RDYI6m2Qs4Fk7trJVoSVGF3zAchk0LGd6+4THPIme6flZGAAtHQ4LLPhGPF/UCXAwq32hipQStxv
Le3pkFHNWAoxPBNFOebqN1trCJkz9vH3+Kgy+ntkKIaytnHPLgV4gp6qbkmD1+Q/AMJ+FDZ0NHuo
g9hl4TKZBOJRSgbRBG1wxBulxfD8+KniEh/K41EubUOLpvByio68kf/XrFbb7pKHj4sH1ytVPYaU
VDTxdOTad0MqU253fsgUCYLz9umsDVilAbpYFwY4sW1oDQxpwRwN9tgyQ06ptYOAdbpcTFGp1RT3
pt87DbPi6vU7kzM2oJiP5godxmb1tWPTJ4/f+uDhw/mscFYDvvIIKzgWEESmS3vm/YbiHXvRRehn
TFrESFGPLe1eIt7sqqkhIzb4q4ywNXtnJwS5hHZrR7aTeZKDix+kmM+MV6oCJFXu4/NWw+fPVxSv
hrzOb1WZqdWzGXId0+vMMVt9qDX+VMpFAkr5HxIwSgx2F4v1uT9fZXlFezuN3Xpht2lIpohUXWt1
MNg/kcVotFUa2uc3Z6zqwlT51zsXaIHnjCAhR7bZk2wehOIQUvDWJWBKxDl63m/rh7SRksLJMOM8
kPuDH70QIiAe3dUh+jDi25kbRjnkGEvR3pvqB3NWMUgTsX9osOx9KaU/oksE0R3QUZOCRKgV8E+F
NYtUP7T4kMgv1VjdLdx5eE6c/CNAUUdN89M5ozWCbscJwevCKcqBVtBSGQr0q6wDuk96FSfm6w/3
mo0l9Wu0r30wjjmRW0pVSga/9IlRH6yLnVj4tMhcdYpPNuAUdjZXGoKrm+w8FSZvqM0znYNoWfLk
FJoSnUV+3tcfTmZEWugdqEqFCivxBI4Oo1BQmQ/hF0iO0oZqM+Xiu7LA6nQvpGKPsvgXTTWcU6gl
m0DeSqqLDCLZNefdKxOOvgV532c2u1pIuXDvmj1T8uZVMOI+2ZXus6qvUXX+Eadq2z5shA60Wbbx
dF5w6SSHMRSSWH0LOlyoKtIHNGsd2Yyj2ZfBF+Ti0OAQHce5H/Ul/bvLfMOE5cfoo4hRmCACESwN
ZWI0ABwjMVQbA9H14pXBQCnuJBsg25VHZDhB0H+L+MWADPQ9AMMkZjUopa7XAxEyhWQjffCq38b3
x6lps9ZDtYTF9j9TvMcOGeX0bcZrx7NbAQAsWz6cqdMaM6Z8Gdl7He56+RmttRtIzNgseebmRU8L
l/Zwb3w2THOgZYV7Uzo7mJ3ismNIWFRqUAY+yWr72MzvOpl7H1NN+V6aY5rR0YY0zBvk9379nmfW
021YmzczL77vWsSRJC80J9tRh6osIAZNG4kVzddi3VM7ZaPcsh4nIHOV2VDD3r4ECD41UfAQ4ysC
zppJab91B6LWQj7ji5K/z6VUogwDx582R7oKnU6j3fT6XEFNoYw8YPUuIsGbNSzkYGlR361PwxZB
g4DJ0gvb/YZ8iefaJC7pphzBBk4UI6HY/MdzUJ5729QPU+QX59tHH0zFUS0DM10LmO5+k/BHd7R3
prdoL2uP+B6JZjBm+0U3wLrnF3as8Bzesm1jXPSh3XjMFK5gAYg7JWHlVIHoPPkVUjEUCE+WKc58
I6W+mDGA9DQ1J7QkYeBhz7Bd+/CGYpVy3MwjmBSl0ko/XVx8TbHAOP6ZE8ItAxqe1bFw/Yye89Wv
E3UkUG04I9SIXMBaBSkj2fvwOVyMt52esR2oDDk5Rh2s451Vbo9aOa6R6sIUlxFhDsBPOarZ0BY4
nIuAxpVQA9fshdBNLfhewM6+kIJcNCbGeZKTcDd8A3Kv+/CXFTvqUY6bsG1cNXedXrKdkHX9slUZ
yYM7Ofqh/8PBxarpaOgX9xhuDfVJJf0cOrXEpxhsTg0hD7yD15nJM5X7xY3vBagzaEowgg8Xsjuv
xmDjMY8Q4ZX9fjx41eBbxpB2gyokl3iD4YJVD6lNIOxFVLzgCC9jdQJFpQL2bDmJNU96VUUYsHG+
nNyrgCjB5FkhmicHXW02cN4K4rlurx2DBzhSqO5EqR15cSgJvjU2glmBBthVDJZ0wLjN1FzJd35E
qHdu71rGpY0ls4T2AuR9p7yTV5QkhkyMpQYXpfiVQw7XeIgoOYjW2ewn/WdB6AlJxZhGYrJaIkkm
W3Y31DXlOZfGeGaSLhLtxs8V4UBNvTXqjLV5In9sWiNsyl6vlcllOnQBUcEMljo4h0uPeIXFe4k/
zmKTMFN9afWLr1hPVCxTPNtI4dVOOWyvea7H4Xrrpm05NDTzcDtQ9y6qTD/Zk2/Ug2t2CVOzS/U+
E8vcdi4dZg1s+VC1+qYxS3/4lUFm2t28znneyuCGllwLVQEy8ViaTQ4PFQihgHYuDqBYfTuBdkMw
O7SP6OyIueHPpYXo0nuNYQRqL03bASfixjBWrA+5C8qPBxyzRO4ouRSUDbizeEwdNWT3xbaGdEYP
2mFvxjbH834CYtqtJaksmJg5GO/Zew+ifhViVOw9iceWhrR5xuRvoIKJF6wBrTchO7ij1rWcOBnZ
WY6V7F6rhpcVjZWojEmc3vmrMUvNdcm3kjzfO2tRN5lpPji2jiV7Afo+UFPvUCHIZ0U72BdX/xZH
7PTQILXKJegIi11ffCKNtRJIWU82Z40ZCDjKjrkryp7n6F2Kz1qo9oFab3etHG/0KaStMcTqv9tf
J2JtRox2ZUYeLZr09gAtUpkyEiZ0zXVh+xa1KcwIuUePyt8eTy2SeHwkBGYRLi2GfVgZyO9CuZP0
HulnaH1t8AHQyzfoXYiZJzsQxl2edG7+K+W9MUv5g/q4A/3rEwzpfwgj7DUBXpJV5M5Y/t2w5DrV
pYxI8AYpSE207f2SkaxU84p113/Y1Lv9121em7vZYHaMNlrI+vZKu1yYou9w948NxlP1lUBnxSOY
jqpOySGFCob8cRIrmeTNcr7WF419mxKsjnWaGyld4xH3o5CrVRR4MP2zEGiahv1+GHmDsjrcmqro
tFxJTPSEZWyOYAwIUFcsQdLGAWygriT5W8VDR9OFWY3ZAByXPjpNSKNeRZWLm7DEaMeS+wcSqfXR
TmA7cNgqGhHJLAkVcOlCxqAkhxrUkjtkS3kDi+gSgqQdwL049F2nEQAjwIlmHQ09SW2Y4M10VJLx
ud1iWOQIWXwiZTAX0R0YlKoDjm5RFC73/VXguve5u8iOagSowApb/ETQOlpsAbtlx6xwwHlEXC9+
dzP3Nkc3cdPWVhLAKJ5Oeqvncq5M8Dnzgv22yI8qdvIKPDI8RRjbIB6LKIs8MuNHaPR0vFCl2Kqv
rKMi5Xq1bwuy99o18K8gfkg7I2VbVEFJzCYTK9N3imdbaHcWPEyVW38AUOVs8AXRp6sB0hDg9YXR
pWXhfpQWl8ZBFUWluFWnoCiuVrMcM2yBeRpQCnV9YRxioyOyOuRgnOfMtNs1ZPiUSKZbPmu0bHv+
loSWDY8YWD58JUPZX2kkzBWTpcSOLQOIX2luixsVXmizn7flHKqzQcyVBzgwXRroYzqpJaLHT/iz
OXmgrQUpoia45xZ5fgju7Aq/wHWOwoubrfsbIoEoCl4CTVilFgLj4BCh4HMLNNFKCk6dyRjh+lIm
93bvI5Avbo2p52q0/IVPETpwpcbGFY3c2dapMR6WjxpavkGzppcPgFzGIFgwG1hBE4qX1LcAbhJI
hntGNjEaUng9njI0MqCqwCX7Udun3AUK69X0H/2mAqSMrgQOF7sAR+/KgCgJfSN16KCD/Z2dpedq
N7tuxKa+Q2QhTpLW48Hx++fBHzTBjfuuoVirq8mARt3cklVZFb7lrVBAJHZ5DHPWAqHHlXueOkC2
KyueTwPAeS5FUzeT9Gn0mvhqqrS1KzN58xiw0HtJVVHTagzT7gdgn9DQlG2lUO767OoJNfSZ/1XF
smHK2k7HmDqDJ3MqnFaw7nYgwn7oP0VJ408PaQROSV4D2hM0dy5pvOL/kWTOEApVpXu0unqNsHP/
t7S8BtfE4DKBn2+ZTyVadRKMvmdRa9n5U7NE/C9ajZF58ey/05fKNE29TK5KJES81/KHP9ZEKKBO
n2caupiORunnllf+SHeWe/8HN0NAb8y41ub20qVUbjRa/3aJ5SxYIsP3scsc9qTQy2Zn4/G9B5jN
D3AY6UmjLxviGpoocXpRfQFmjWa2X09hxuMOuBLoFUZeSH27DgTk1xslC//XC15SEPPIWel9w5d4
MQkmhcVrtZ4DwScI+nspAuxt7hY/Pqvs6v9hJgD7tNqE8qOz7UUTLYmDuvd2gwu25sx+wNJtNr+r
7Tmj8+Q6UR42Ij9RXudEEOgwQu9sOdZkj3CdFXjN/CtDesVPTVfu2+Z/u7fEn3tLFv15AStrFgv9
X369F0jG+RLZTu+GmDAzpmPuqLQEe3nLvb/U7VrspwRkBGqKt7X+1+HcqWxNEOHyigPOatJZOs4T
d5yfErO8Fzxlk5z+tmCoktqBij8RGK64Ocqsx8YF9WaajdqlZFSjMRg+wP7NwA0sTn8ac6N4BP0V
t3EQ84hXf4Zd9UmCFBfiKztJhOrDLjLGXpE0S0tGfpkcffrluyJhjR7caid7zE/+QaMOk6TNoj87
5pXSoOQcLWo5EEL1e0aU4Pz/D9zWEHkV
`protect end_protected
