-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
UkooJwVYWmlHA5BiBN12y+T1GL5qp7+eehRHrCY1t1Uq+U7tbPhPcOKGg7Cg4yawEylqbcpbLhYc
71wt5EfVM9SRafgJ31WYXr5Ap3ojaSC8QZ+IVL/V1h56Chf++eLn/9LvDf5jcf/OpJebMYF8mk7F
9/WvfvuhSymvZDOd8LpVXRZpBTtU62XHQ+hd4rf5rZ+XbOd6JcfCbONpwhesRHr2Tp+QYrr2A7Bb
mXjFNMWpuNU8jPIwqlvn5BYVu2LcU43wzYwA1Ap7JE4UmivDZaTkMNxC5bEEM0wXDt4e9BGORaCc
ehLpMbrzFQu+JNJahwyu53/cIWlpOP8jCAb3WA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
Md41Pm77A0LYHmAD0JnQ3NfImb9zMlI4kZA0sTQXQo6Pg+UclO+/ftzFk1ixSCkl5oRGSvaqDm/O
wRIH/PrPb+E2eZLhv4TF9gefg9CAKkAFeERIpaw51MDi/eqLw9x9s0P8JPxyFi0a3k404MHrvVbB
keM053PzWyFhRQQXnvTHg3GeZ2WvjYL00y/rO4u9JH9BezLj2AQz/BR6c7aG6xPW1U1WrTPc7qUr
UVJwAQgXClJBJzLFuBXFT02bJD4K+CnUkd0T+z6BoCcYIDulNPgHk4bSf0wUOp2/531l23yuYNp6
oaV+5xxGsbxJ5HqJe+K2kBAo3fMPWheKurFwZPD0CHaZQYPufEmq5tufqPE3kEBwvIVfyB66pzxE
rj7f/2lrxLWZR3/itwQs7cKQH7Ti2gP12Kqk9iG+Uk0Z0HvpJCp1COTVEZv/IEZPwrho1FUubtQ+
CWOp0hDLHzxry62tELjXge+zVtUbYy+W4/oV9+9PjcrzJ99nQi1ieWIGZ2fQLUlxhneqJ84jjsar
24BL1G4cHXKoCuOp+8aKsuYtnl/JzcsFi4AiJCjJtGpruaxt2XPJj9Ynt9YoDJ7CRj5FICZ3KQeO
x+PVy3VNAg+6sh7XphaoVxGmHk9TlEilcDjb0NwMAp7KUR/80irox5KaFMDFET3N7f6lJN04twOM
pJIs2E7wMBd1u9MR4vtaQitu6+J1ljVkQZws5HvjA7PE1au60luIasJgPGMPgix1VCBiD515PZZo
X0k8Mie7JdnUlC3NWsc/M1WbqhAYd5dtZkWpCcV8XqrKCpfDqiDRDZVKoCc9MWtW2INECLjWZ7su
IQihRyZ6NpMAybKRLAW+ZLugA6p7lyp2/7LqLKmfeEMBqla4PfJ7Nkjt3aWxOfzjHEAB4D27Vihv
RN078lToZ2iVhyV/DVdCcI/WxAma4oscSeimaVSugQjhiu5zc8zAlaRLCWU6YdaNUZzEOs2uiT53
cf+o6kYJeaBrr8Ut3MMdKQfVEQ0FyVsyW+WkWZBJS6cQPbxPiyy3g1OoCHP++eytJIF23iDxbkD9
pEng9bu9LUvBkeyrq5BADkuvpvyWOnbI2wmw0Bgflm0b8M4Su53eHQn0fqYKWToW7SnP+1CuUe1i
MVUYVhSgf8K00UEo1btPST8bVAsO0jYHAxoQd3pcgas+fk1Jgq+fSKkT/8uBUg4wJXWx/RYJdYnF
wV6Tcmg2ZFxwhdbGXRXyYdoB6640HCqbd5maEfmsPV86QhUxYNQm9XKDDhRHvtBBiILx2eXISzjr
m5H9PbIcARbAWMKFe7p/iwEoFM1VbNqyg8cUDRP5DTGDIuTN8XI8GElSylCPzDNti0Js1qsKdkgE
O9K6GxBhZAnSMWtZDW/Ar5DG+HqUrm6mwQ5w+DfeX/3tcKtOZW15/NayptWe37f6MPnbIGxQoUDr
YXevTUomebXeH8///1GGjHL5GwZsbWuhOeQWFoPdxg7C9OoafDEVrQCDKQc4/9/AD8J9IEMsFAUK
GC+dEMiAogKH/3Hr9mkAhhMsEm6Gp36+QV7o7yEV0fJY7mVvtSdPmEePklW3OObAyPfHmC4Oq/ej
KB9QcMMuBdHosoyVh6d+Kr1HuoSR6uh+x8gb12+k9ilTuYCMRbA4dTFvRpvdqJaUM+qjD2V8eKeW
0FoRaQAgE0Lr5OcqzUaszcn8VqsS0GUrKsLbJ84fBb4YNo45o4QRLklA6jXU8C1WTptB/UqGjoLN
soVLTKE7p2C/+d9mrJTgcmUWnrRpfrhm7Qxlfs9fvABp2dGI+q759mDIAoO7weweQpGm65PAzS7v
KWB6vgXrdjIdM3r5rzlxVRrnDXLKyyi9M6BfPa3sZax7uzrUSMT7h+ZOqEkxS1+x3BB0nRZzL2MH
pkVbk8g9jmI8eWh21GGuf4Q0VGXqNx0Wy2hcLiixrLqaV0iRCmWC0joDigivOCDcy3hyW+vDIEnh
EXSC6LAi0rT+eYdpHhILcGpIg7M78f17cPkI6i5Wv9vNfcv/jEGWhdtkwvIEM7NFj4ICMVR3BI5f
yH/G+w3bQYiULdQnLV+Y1+RVZR8x5JKoPi0yUHYvmn49xCJpsNhvqEyPcyPjWUC+53xPgr1UxABW
uQennIIUo2uOhGqLBBWwobjfkba5ZIcCbjluj5EVCOwyxzHrw7zi8AC6eOZjyTSclPbZwUu1TljA
7tLeK6YPMfE/Yd8gFW3sAy09hOrUQrtG2eMb9+wefi3r+dvRLmg8dE7wMRqBdTy4yi1S5EMcCMCv
DM+qjzvJLcRURRS4SdSjd8KWghOAZkHiYKOE81A/7X6se6YcS8KcToEdkhI52f+u4XvXPrZ3Ms2K
CGR+nEGiQW2PhtOXGeFV8BT6q+y1C9GIhGfzg/i0tNQe81nmDcab0Mp2SQuhzePZZpu4uwQ7ihMm
AKpDrd49NeJfIdbRRis+cEJtgSSh6Bk0sDd5y+G1ASnr6WysAHb1OqEahj1cKCWX6tyfBEz8wato
FDeZDWUglY+Sm01ZXLD1FHZXis2EPpMAzYXsuvLKrlKAg23jSpB2HwamjYTPC437WW+9R8thkSTu
IW3nWfbJcYwvtcXPB1SyS/MXz82L1aBToVxOfZcoUIjrKp/IOQY8WHq3EJthzT5vEhKLz9TY+/U8
MC1KHuW1tkcixqO2kjIn3LLQCBc/9JUDHhu9mLVq5ZHmnNtmggHieCSi15FH2BJhUvgrqt/zokuU
uT7nWEwtAdNxCtNF65PN3zVBGS50osLiw45JiTi8uHkujiphs77AMclRLM9Im+whKDgXw7vesvKn
gQGnwvcnPalnobx6bFTS0oz6P7LnI5I+Q36h8FW4urDsSgzo2a7SmlUSO5BjS7EKRQE3G9I8csJ6
EpOJ8aGm/wi23Yfv9zF1S8mKcGf2h/+FhJqNThSaqaFmUlO4mvbdZvPRxzrQIlDeK7YPEAOAXKP7
XeU4BfiseCnnfaFAVrYzZhmZMUTZ/nbxwEN19ih5vjwDnT+VzQig9R/nGueqqrs0L1HmBcet861S
JpDdqHNZ0nZmwH/TpiDq3M3i0fG8xAaqVFnAX9reQ2NQ3Xbcqo+vmQYP8X7BLauQuIbYFBE0pLV6
1VD7j6PROOSW8nUQdvdxZbZdpCY/FsMX9NJ+29eoj6FFZpqcW5Q2A4O+gjW8tj6ckLzysaHJOXUA
46DEMYD+1OKq4ZdQKf2N+6/VsZ8OyKfwXT3z50+V57yGnlg/xkGImwf51h7a1MBcgi0GwzBnnEED
WgG4MVnsf18zu78gdCgI/wNurFh58TOllYvVL3SAagd1sK/L5wxS9DjRxM3mVza3gKNyLxq+fxIr
jO5KSjE/c/35kSY1H4zzAsMW0Ei/CeX98Gb6O1YUb3j0r5I2oRbIG1DtptMi3P8wCrh9/whpvLvh
3FjlpCPLo01SoQZcxJpwB3NzQeFbplW+P98KgiopuRCpuSg15SlQ3snVYmGtpSShVAO1TI+97v7d
BhtJc/hht7rg1BFo2if6ewyKigrfic+DFzRflou7hkTNIXkXzzOMedG5zDG/iq74K+326mOS2Kd1
4ZEiYN/VawNetBHdsfuhFwMDV9VjEuZI5tK8RTIXBG6MtxbTlEv8n/MTWtAry5G0kamdZn1Vl9P9
jpbWFXQ2tb9y6b6gOjGptKM1QDmFVpoW7S+WRP9qn/SvNBm67WhA5DyOqra6acudXc14oD4OxYeq
aWUXWuWbnB60syDeQDZU0rNK9EPasooG+5dH8DEC13IfwZWJJtbX54MLlKm020YM4ohNaJ64Q0HR
yRBLmTXcTzboHhTrMgxeUvEncKlAHgBy8VtqEBE12uYZqqHuRmD3O2EyD0dVWLKeE7HIQjQ/mGbK
HtRMP1f5MZZ2/Do45+oWhHUysA+U6E3Gm/eDYPMl54yvaeUbeV9pirllqc06SwrD1RUPPfSMPdmC
tyCBfDWoCAiE1ag/ibm6t99mo2R7YhTwBFQr3LAuuQG8H0PEmcPnUYNekjcQhWV9Bw1UcQjGJ3aX
69TIg2m6dVZgh7ZmictfiNhPYyemFiQjBSFi5EYSNVvcprQRFy6Hv7X71ARik3/Ym5JwfF02jEmm
g0bDYE5RJ7B6zf6QAUBQAi1BfJFPF6t2YMcZWwqPW5nTE4uKK3admTQ6Q4ZIuqf1nC/JvW9iB2pw
WiFX8ANLnpPp/sQn6ISMU5vazyNwylX+PQ76c50oMqcZjIsHQKqYoDIpOAbDOYs3KXxzICGfkHYN
kXw27M9/pOPZ37bSK0VDhLgbfIJ/6hsOA/HUvDTkcC5tMhrQo/PnJw60/XeNJRuxr/KiRVBGlxbV
kpM78luflxBVtjK81UkN1zZX0cDW8wZfFfZ2txoVh+c2qfzVe1F/vEH5ymF+YCE+SEuoXzpG5Rk1
buMKKWSSXxQWM/uHYyG6wAJ735kjvFWhkhiNErJ7c9InZvJOMKGVFtTUxZWBH+EjX3+GW1yJnFes
NBHswwvZYapRY3F9p9t3k5rE2wCfu1Bwm6FW9vjxbYRoPTnEgD98DZ6c8/rpmZd/jaq82SwN7g/v
yOXFrYq6ixKSiH535wLr3t7xVL8RO8c+fA/cga/gvnThTC8elrP2Vwb6KUG3Ya00RnXuiiBm3Tyk
Qe37jxMDZvTbFXDRQAY7CB5lzKrSuwk86MtdxqyxucCwvMfJsD909cx1XC7dkVWLiy5TqmC9/GGZ
gCg73A+2FoqJ7MuJoNNg095Smns2WpPS+7vimC+fXBrxj5TxpgKzL76K04Dje2Bty5UX/itPeG3u
FH0Hdj38onLNt6SE+rQq+l475K7IF+zZ9xsxKoVqdEsVU1/2nqaqeimvbGLU5iFnw+VTfC+T/uZF
GpVuR5HyGamlU0lVLZhkaQPHWzyLx1tHz7Fa6Yn4SQ1Pfln25/fE53n4PX2avCfSQ0YTk4UOWZIN
knVH1MoilX50KfdEN4yNgKlF8CCR3oxWQ9DO7bVVSbpfK94Ef0v/2jyH9Zdtqh+zIQb9yf0PoyYS
D/OmFnjm2pM1BndYzOUbTjKHq4y/n6OWzauYiHgYqVqZDiVzXkXJ0Ff9haX8kJaEVzb70t2eMx0i
w5M4kmxxoS9JJfNRm9lJn1znwFoY/W90Lbs+jDLeumWpqDgIOuLf+TPi9ES75pwGETg5qkSSjNVY
rziTTvBeiGoDKFOohjPYsF5tJWe81FCHV3HkEuGLQkOMIVbKbd22xojwyBFcMrOfifGlU1Hr/76n
mz+2TwcXO2e77qwRoCZA7FYI84WflZ5ttKPXZG0qGhicEocQyQXhgrGcO6gVLcW6shOe4KAeuL4B
A/G5GZXyVmdKRM93wwdzySN8vdR6TLDxDKFHUX8cZ55yqSWQPvPsKRmsvql3qZoOwX+hKIIw8uw3
IYSCpccEXZameuPCQ5TKJwFpKDhX++rj6ipHm0plXPPqisCjUsUAjgokhsCB7KwiCv3C9TFG2SHj
DDNw1D8HyQF/1GdQov+gGnQqSTaROOYV3cRWozKZjmTdenZIfq2DsZjCT1BuB1VMPaUwxifikDku
mEk18KqK1bykLd04k1iHSaT0Tv0PlKGajveAsio2xnchsC3MUB1nYBL8YyuqlNeUKtkS7BS7Z1cK
w5liGEC7/xNa8HU/PrQh0K2IGBXcltxdVew+KUa3cxDowSN0XNAH8j9qnZr9gGmD1YlskJmO6gw4
3E1gQD4WXasvH76ckQ0furCLOHHv4hP14gBoZJz2WHd9uq5Jf3HYGvQ+E6TXSoAJL9MKRnvM/Umf
+B/E0UB+4FbV6JFZkk5Bns8n1vLqVrpiIdjFhlWOS5gN4N5Q+pI9tdjJMkUXTFypEWyF+3jy7h6B
xjqksisRmdgLzedJA9NQE9Gdqz9gx//bN9NOubm0eimbeO3xavIU3/sD0xkC/6cDcaImDM9SHbWq
DKLC/FlyDTQGKM8wkNAKqyBL4IoxuZ5DwVlwFdh3YIoJW77niRC+F2m+wHrajXzt9N8K1oS5v/3v
JXyewKWHhbTej0yOkUJx/xKTSLMARU8YaIx5QvT0EsAFg94nT6qOHqw6RBW5ZiTY5sANsIQZW26R
eiupBpubdBC3OCZymkwxNhP2zQSKX0Zril1FJOgVMYmd3ERF3bnKnN62vrXt1fgkegZgTQURV3BP
UYXbJznnCg/To8lO21VnCUuyly+PJNX0iOiraZBlfkdVw7/iraHZetnjYIzVjj5XKqCTWqP9t7BE
RHX/F+7trBQE1knW8iv2Q1jpU8FMaAuNdateoQD4DUAAY1IS5anq4pKuSKSa5MEAAjp36o8lbRX1
JZM7ZbCDNnw0ohV2K/PzahUtPYQkgOl4Oocn8cgFFi2/PFwSrHYzi7qQcU7OSY1eFZhOk1WAPM9a
pwRBbQ1yVn9/vgJ6/ScuqlnnjMDeyPWJcXmODF/Rs6brPG6PK3KkvvW19O0Wt9GsxvU3QWSD+y6H
E8oI6gqnc7FK8MjUYH727rSAuaIA9QuAQYO2+U/cFh6Sc31FATrp8kMAlDN6q2H0cZ+nKb5jJdQK
aGaowEJyTkAFxE3KBzsP22+vSxa0uyczZNW2afaRuoy42TYah1PrE1vR7FHwTnaBKrkO6z5JNbOv
Xw4zfvchwgnpo4BslLich+JHBO3lBYzPi9XOBQLs1nnPRH7ZsFKenUyLJ7vJGH4yxkBPFqsgCUQk
8EZ326Btrg1wgRGuKgaJbaZ+i3VUDNwmoKref/3VFCTu9xtqTokE1zS30IDnZj8uNtePkHoCoggE
uhoOwZFVvzRr5UD23L2hG5BA/g4+zU7/mpfztfzaNY/HHLAJ+x9QJgtF4gsurJqXetV3/aosz4ER
lyb3Vs8jEwWH/MkvKcHtH1N5NWTHwiCqPxw+knTS3zW7hYXLLNfRhwHPqTxXaKZcRIwKuqET/r3U
TTufq+feMRdaF5D2YLAVFTSJUKLAKwg4OzQk9wcQPOzywIyYg8grbk5cNSH7aGxARQqHFrPnVaeY
Xz1kL++suPoMZ+Vdtu1NAbfCUzV12T9cWcMYpSS4zTb/mYr5euxIQhbA1bCTcCD37/d/Riho4DmT
btE9/2BOvWULJaxcV4T1jhLh9MjYiCJjqLRq7hOvzXLrhKOmyU0cdPs4XvsMAYbPew/evWx6mDI/
qpFd1eiJk7bQ8w1iRdIPIT24+kloF8A9AMu7jF8H22+mWGFGDOKQrQ5hT2uCelLFzrDOunQ/VuMN
ALcX1JAUALgwuIIziDpaycHJYskZlvZVUDhsRfaDcsNsqbUg0l8uxgDpgtffTBT3vl+2Py9ORhWv
DP1PG00f2URC7fp1s35Wc9wUv9/BJ9VuLlKprF4eW3wB8J0pEnOgdfbsHnB9WdPRBLtioou/j65o
TCszRrDr8D6oFaLjf9sj+MH4T4t9S5QkPUS20QjR0f+iA469RF4VkJj26uqDtsNfwcv2CFQPKxG4
08BAmbGZMzxCWRfZ94HRF/zExYhdCM6IEF9+FOjQCvmebv31RzjurjT8X4LDuhKYfWLscbRZOVOz
aUoqGhy+hFq1kfnQ7ib96KqElje57+zYgLcbmfHeDaV8fHm4Dmo2zMk1fjmLZa6nHbMHwiQYR/py
kVeHnOdRo36mK1x0YFsY7lLWS+kHKfm5l1KJLKTl+pewk6ydyk/f7SwKe2S3hVEj+cUcnsnD7xDv
3jAuLwYQdBivy6jF1avqsl9IZjQ2B+PkK0g5VlTwpNpktoM8nnLj87ZMgOyrkk0ZkwcOySYkUCkk
hwObuGtlzIU+6Ohdb2s9zrs7kYRmRxn3Z07bMirUA+KWbefIiLDq0WT0GIrcjgp+ee18hthFiQYO
Nsp1jkJe01f+X5rsvqYpgPZ+NHfoAaiYDIEf71V8oCaOYmg1sAzvlBQhg25y3kASxMC3va8L/u+f
B9ltkCYr3MmU6WJzHk/vvGizEeapRf3AF5ZJcEbr8UlvV+WS4JXKJPtRiqScXy8+q8Umnu6A+z+b
hE0aTBbi/Ay8rtJWS22t21eLkx0bv34/dQVW3/t5bxgtI3kC3zNlwWflKwKZqUNV7N287SOBE7VH
x/eIz1QRdhJoYFL+yBAptTHDnLLDYRtlX5/QO18FlI25FrAOt2CPLx0uW21gA3UuTt0rawsd9zVn
0g2+am4QdoK5nHqzI4Q/wiBREgHRqHVWwSW0J2yXclqtFPbEp4k3RC1BXIjyMtKX8ajYt1VPiSnH
5pbdkEt9EwrupzKjvV6bq7+fhdaCNiNMCjF2rcTWtqPTHambSiWLOhMQHx/fufZB7nUT3m6ahN9V
gD5KucusI/uP2ZuXPB51P6U18Dt+U1EvU2ZhCifRHIKGBqm7IB6k80ZjaQmBg1npKqWyvkPuxkoh
rMSnHEJXP1IqKmTmj74hdpaSJ5hbNRDJNygMu8VKvPc45bhMKqFFrhy702srWlkmBpQhTPMquMBM
JpP7Kru+1U/CPaKpHtBCaAVBvTOpxSm5v9+EtFAK1j1WvcNIpix7yu6liG0mXfWtmdYkaMvXsKJ6
iONnKaWtDNUhjwIXpsVR8MciFO+pNyFQes+L0Z8IA5Sf9534sgQ2cD/ezVyoX6mNzlNXCP+OFgNY
J/VNja8qWHrFxEabvDyHLP2AWyXutOHFCsWaX1o5lkmFVvoKI7iUlC7eQxtnWCaMeUagg5cFeCQ4
ACF5smsJp470R1CA53yPIQqb+2Xto2ik523n1+jfywrZUdA9kSsMkbAD5OOtvQz2Oi5CJ9NHuTK4
wDzNZQv7/741kx0z6Tea/+LjG/oS6Ed3XAUaZOSOvEc81LFt4nFzb4u6q80raHA9Quij892Sm/w9
wboMAg2CfWIwLBWcjebKKkRLNoNk7cEdwetYRxzShBCqPGRYAzUmhEIU7nVIY/eli4nVBi6lFCPE
eU9J91TH7bSnNG9UzBu08tDw6FhmOd8hANKm42dHRd68nurN/+zp7COMGIONX02ZWeVeaXcepmh7
D4Ri9qWYg+R6/SQ5aRVA8wfaV9war9SsG1w6+uXMxAPgG2YJbdY/T6ancSEH7sMnnCw83a8lTY74
CTPy66uQcnpvfloMG7v/FaZkVL01fRpO1GCqW9t0g6qhiwhS9al5u5l6eCyGcU14n0MU9t4ZRSzq
B2Q7RCNc2wg18TuxUPMKW1qEG/L65vBZPuB0191e9NRqgueTmIhwBLkwdGkHFrRD1aMaHe7MvCPP
rnKBdcpkodMetvA5kgNVpDzpkLVseDWg5IgfdkCVQmw3iVk4lO8z1ItCnn0Sdt/ponbmERByXI42
oYk/GNVW5Xo5hf9GdO/hmiNU8/W12W5i+M1++g6rgY446UyH6nr87mQ4AeSJ1v8VuPs9Q1FvpHy3
qHA4gEkXQrtgu45u9na3uIm5AcSZu2C+UU7c3Og3TAtC8uZsZw8ZkBUrO7AaCCZTI6IIuvupVK6v
/jT/x8dDrPHNp3m7XGUtOQ3f/gns/BfupSXERmgKcOUMQlF8bAmDHcJIwuYq+JOiWZy9ew00V8uP
I7AtwQn0oueoEL+gKAmbK0buWs/DEhv1b7ykNABmgSYn3083zqO3GmEhkTGR2y26gfbGZJ33I9TT
n0svbRzNMAWEjKVQHwl7J1LfN+/y5HfvmdYtFlbVWekeIZizti7WOCa0PQ5wRTySdRaYAOfLPqKM
6gBDBUhyeOgmDdhUyBi1L0F7fwoHGSEsIbxMLWBTbIv1axIy+WXO69Fy9nNYcuyk4n3aYrdMNXvk
EFbb+jR8yoK6bH52MewpnwMsALaP9ORbVY1ITYOPPdA0MVIlC6NVq8E4zrhJf/kDqJPwbVBhiCh/
jOOhkr7kQFoAFhwID5UuhdYUEmcBbZcO46QOliTCe2KkNeKeylN8g9D+sH+PqAp83wQSbaxpFhaQ
a8qwmNAw5rUnHON/oHy5V6IsWUBlaR0ljmw98YKbHIpkJFj8HL31Xt0dIeAEUGkYeLhtbjy9rcvx
rz2Ez8qeTA8QLVUlz/JlTMsH0FRg0vu6SLxE79EgBhxY0dFh63CI8I3vbVy+WEivEJ2FjRFv3ADx
mL3jt0yhlOfe//N/1/R0/XrBMJVGwvRxmckWgX64skmg7UoqVo1JSuyVWHuW10cbSodturLsMAQF
6uMJ0Dt+TVVkPvVCLjQe1PYff8k0RiMw4qfNmxzfTfFU4byc2ROBkXi9lW9WiOveJuHTf1sp8zjD
p9Db8s6cJw+c+U5l8HaRQidqDFfh8O58bWbIb+yb3fCM2VeFUx6pz/lz9/zY25UtmAL+3YXizaGz
KkSER/XQeiWarBzhkYys8JWDVpC6JYuYXMg1NLePJ2YydUwE4gklXo3gZB28k4YQ7lm2x24vqfHN
jydb/GjNCpTGfz1JE7LON4899tgiBiwTtCWmdX3TamcBLa3dkNlkRf8vLWADy8tjDMcGOsj8nOWZ
mjlm65yxlS6ObJT0nh54wjO5tjzTymU4N4VR1K44e//uErxGRtKsdmeevsxITIqVf/v1V05pJsxo
cC9/9O3VmabS97Lc1Xw19k8QQ8HcRK9ZlHDx8wdzdujV8c5oAwjUvqEyEJCG3pZ5s35pBkuPstT7
Z/Bj2thpGsq0wU4+SjWSAEe2hLz3zgrbsiMN9dTvhQSxbrhRBwKgCmW3bpWxnofPK2lQfJrR2rQT
0n9cTmObS2GPd39oA5DbC84QlqH07F+NU7D8opUO71Q2Fu700ZZpXF2daxmMaoDDtPxRrFTZYysl
N90uxrURCCTFRQ6eMR+2eP+/D8+9ZK7LPEJvCLt11xGAntJNk3R6g2DuseGrCUY+RQk5UvYMgCV3
3N8P93QAEO2RbyMfOwoiecPcE9zwMREgaNGgtACy9+aqRZiqAtlThucNysOwk5clukjHM3eKtmJA
TStQDhgr5ljy9UlgaUwwiIBBa+cfjy49VPcyecmJXoWx2cfti39l52/9G4PvFCcpbfkmEoFRFTHu
okM6GjTxnMCVEw4yehARetuVIfwMNsCE3e2rqE3JUJalnLx+JKFwRFHcSKGqOo0cCvVoZH199ADL
L2MEMCN1GC7lYU50gBo8RoFUhDXGoxqk8iITrVJLWFDFBx1nGiXBeuhrEtQr5oxp17U8jRpzOUvM
ro9IReH1bUNkzeKuPBnkcKrQGugHVO9+etCV95FRfYsAgcHRDpsRiduSAIG2PjmMhBSTnir+FmXy
ifiKn+FVneoeX1FhhYDGgCPyCqdT8Tw2dOylOFiFTj24B9RQliw1nDncbxMdjFxff+mFNqOrRBqq
2NQAX/nT5zNCdOfK5007/7tVjVAJxvrBr8xDq4OsfPnMU/iYsvPFWgnfneNj0OBsCgMObtXISttI
SmrJBKmPsrPHjKKx5oQMB+TD4l+3jIsigHSiIYATlPny4Ryby36/N24j+dUM/HqGcC+L4JwLJqIH
UO59csZffsMppbTko8TZxZb9cau9foaV6ljwkxj3JBECCGilDnU5U6MmAqfManEti66ZU/RHpCzD
2/67FS56bnGnfeBd3wJreYC46bOVbBhms0DIis9KkwYCC9OKtxz+HgoQmGszf+aq6QBN0uk69yF7
4KZVSgFQ+IPxnfZ+FNR6vtbrS3R48GRb6RxeRHRSkg3heFAfKvj0088dkxJjpRAL3aWzjJFv6aeH
toJeRnJRDQkJ1jB5Ncpkhy2ew+yB8ZFMHAkZGg7g9uJv4BuBE8csm+3YgGPKfy2auDlJ9exJKwCn
otDoBt12jBEM0v8kCF2oZIf0HoBldWxK7TJLU997t5CMEy56KRd/+z5mlZiMB8uyzT9mt+gr+DKA
tw2I5C9BRhyGfu0DNq6HoKal/RrGYhfm9xR/dS2lthnZtSRqNDgDH22XaBG3NiN+o9jjrbLV6FRD
I7IYVswFqBFYdat156LE0tbMuJ3R/22Y1v85S4iZ3S+A9oLMoqhBq9R9MoR+vhU8c7h+Hm+74jjQ
qb2GnLQy52VpdhEYTEzHH1I7MsPjJIW3IwWMGSxWgNmlH4euTjQ55fKjOBs5o/+uFBmRODMnC7fZ
1z1k7qhSYvC244Z5vOJtBR7wlev1WtR0KO8m7Ayb9EdTNstiT4LFD6dKB8k/qGhy/TXZRvMhAmrp
djjoEK+ZxlNzDizrcuAElNWhg7Hc505v81leLvl4QubqkfCiG8iERzlZ5rYrq9DF8JCpbGtKk8FR
uJK5QOCDWOBMZGMFhXTtmYVrO8Ah2ABcRSPX06dC3EhQ45WF40+6TSAHN7wucvgr0y2XeqA1UfSv
SV2x+ts9VtF0E1RrGu9zthoUSnibJuj8jApfEA7W6HzzRBJKEe7P3RPJO0d32mQzkB+Z3MxArpAg
DvH+rOYAtqnD+LGCJKpgmWXiSznPnn5VlRb3fdX5Vljf3aBXg3b9IcewWg0qpSKCjN7wnIKe26wl
V4U4tQ+/4zbvVLig7kEbCXuAWzJZni4SdE/RjmTHYMdAWbWSiYehoEOPpc92ciCq0iDFWAjouLR7
F2Ws36E1th6rpEHl4wqe82avxgiIsdMj45vCDQy+ZsBoxrZHx1NDmUumSLO8wp2/U2/B1wwzEDcD
j4/Eh6z6e7JSP5E7n7kXRR+0U356BIt2itCBPK30x8/Jx7XbPLpe3G2Yv/LS+eQvvpg4uNNkC7Rb
5OyFRLiVMAwuCU9Yg5jTJhF63lzIcHS9uRwJWTQ4eBm74FNytXJgdi3YpfdHgGjJPwZA8lCI7Jbb
z+97jtHREqN6DSxRVUGEwnFiWWENbHEq1AoZb1xn8jEnh3W8ciLpc7gmvRVNvAETd2P548CNrhIS
oa1ViMeSit49BF9v5SLjG1xlw30gAvRsCz6TnmHLEzrAHJzN1bSMGBEZfhn8e1vO5BZEGdOO0UV8
MDrOyDyfn2Oa9tCgsc3nmMx4n0kY7tvKC5F0Pzt839WCv7HrFuGcLWVAM0Y0eJz5z/2hzv7yhYit
yD8SdnJmi6kIDqC9TC7VRQkxZ8FN88sVoxIdLAbuFsOVvCsF1TUCXDGqMtb/ghV47YzzgE1iwPwx
nNFkDqDKE8YIOE/c2tUFPLB1OEAWfO7tqemUR6GjuYYNjeAJUxED7tGmxVkReamPXVu5I8wHVJ18
6ESnm+U5amqZyGZpf/4r+gVBuSkDWPOTi8eQCA2Wz1zUGR7VOJR1ez7i2x7Zyl2MAsRJ9OIcJltL
KJlyujvaExYA/5P1L1FSTMs/abADP6HuWh5o1nWoivBKEkzaZ3pyarSqF1nH0RfsXgrctG6QP0sl
82dXxGntDKCo7+aP+GGx8IAVeF6HX7cklmHmQuxE4E/91xO+UHuJgI1jwC+G9kJkca4tKQwv2D6Y
dgsWeUqUa9d23aT0thThvMhzg0m8GgW1L5ceJAOmdEyYzkQYLbQUbanXW1xGpzzB62owpop42h+x
+G2V4jYU+JafwwvUq/FW3EQG/bGe3i10A6afzhoJg4uTlE4YjLOPzR03zOkf9IrVprH2yBM9+I82
veDnIJP/SyHtB3vQbE+Y+mRxsq11oTvIFEknHWgl0P+YemhOz6oSzG2uyCyAP9JvwaJyChrPuJl6
9xFrA9ILC28rWOCud9ji1GRLKt1vdP/kO7bnKqI5dnOXbQNUhTByM/00DydqRnut7XDr49kECQTr
83r2FCeMpehxnob597J8qL1T7otan7ydYglFqCVuVgTeBffSfEei9027E4SEpdey38Zb0u3vqPvz
Gk5+weJsGsdipmBk2U0nhDySyInops8Z0WHMTP82sNgPCDuSjtwCpZdUbFHaujmz1wErnxPZgQ+u
V7xvut6FKLIY4cI6m4A7PZ7P9U3O41WiGKEBplYssd3MgySCqrfnvc29Aks4Xm2DWGSxgWDUnVPV
2WkBBqZmSkMf9qieunXkBvfFuODaOalx673nvMGbys+Yse8pJNRsTAB5wdhkAy2vPpmuWHrSi2Is
ZF8nDqfNWxH3KzhCkIihlvYJZ3SJwjUqGgBEnDisSExdf71Rwjd28JdJI/umk4p7UnbL3L/CZSHa
13rriW7xik66YIgITOsgdB24Bx0rf9oRUKPoVBLzcq3YFTsF82dRh53/eyPU/frPhPb+8eHky6Bc
Hs6vIgwxYY49G0OryYw2/zADyBCCVpxYs1AEJnd15JCjjHjwERqbxbvBaAcwlNjbWww0LlicdR8k
w1VNIMYtMJ3mwl7pD6JD3hiFS/1voQ80mom5i0p5+mZM8bn4nT6Vw64LQ5JEzWlmcmafMDRziAf0
z3msWG0PME+MA8IywP/lL24jemIG0WOhr1guqPjpppEMu7tCg3DqJRFQztpDsDuAT8YwfWWdVxaK
5nPZQI7/RSC3j31KhKlU7qTzZmIXanCSoTGz74+J/+5K6Urpnzf9IY9sT70TO0q4z/onvtoui4Tb
zg7iDzS8EMTDSv4b2nx8MdCQtnn0bUui2wTIaepXdGuXdFm+COcgnUt3NMJFO/cWWTA6LYfIu7Sz
NBvyc1evTgavCP+PTjzkdXuEQNDloQZNVburOHqPqyn2LGkLCS5D0fAhR94HRJcqIAmunv4IYipa
2O4iJxBH+6d91N2unoj57wYxQQXogQcJmvvcqfboPmJr7WZQ+CxfyZlL7m/4jxhy8NO37kWZHsaG
dhSSdfvSTDL7XGx2/x0M7b8Jd1LpJfaK5IQDRH7bSqbIa1LqOSWtpCZC9WMNuGGPt47mJu8Q+nJe
Mp5Bb5IpStFapopHYsJPc1Bqh667GMzrqQV3DvNkcbfwEA5/GcZUILlIWP32gewiGvMGwBEQVUUs
IGSrhbAavUj7edpWzXBYBBVj+GP/zBPyIGiX2rmu5ocfVJKzD67efEYA/x55aue+P3nrSFNiuWu+
NCoJA0ZkN8GKUEdHo6lS7MVXl4iDGlj4ojXQZxqysCMuwnENSckKTNgu+7zBzOamBa9ZXl7UI0Vp
rlFCp3TqlQzuFYcKpOLoyxgdMmt7qY6bXIDDQTkZUgadPQuzEfcM38GIZY4uQCztETwoW9YoERDP
wZ3i99jP6W5wsgfX6rfdAzzSPeeIHiD3fh6TEYkfUJsdfK+OG9AcJqzrStqD1Uz/OmaKfXz8PH6F
q6shInR4a1hMqHEao0WabQ+2M2/HkMzo1RocNNSTzlZcjLzCEaruAK2yb7aYFVyuSTbe7FbsCzx5
Ev6UBaz4x53bdxE+b+vcUZiKTqifJf9TKxXvFPh5h+5d+TMMC/4EbC99S1bZOC6k4wIpcqFgUvjE
8rqNaum0USlRZ9LwEBCGLu7kRK0/GultbWk/60EpYxzwB2ce9vSseDIbdKD5mK9FDVLdLcA1Vfmp
8cerhUTX8Mouq+cgFoQkgP5O3zhj3T6e2ChDhZS05D8EsNnqSPMYtZWFIa6vZlyGBZBZyanRZGbB
QIpc5dGvvwc9UdlkLCMMV6YwZMq5wMnw7oip5q9PLnrCt8e/cw2WTOlxTEyD2n+rruP87kIwaBcg
JlXqd9Vc765eGqFBCN450pVPZswUh477UaQwuzdoU9BZSRZ4UyvRjmvlVNokEtdvMlWikdPc9mDU
nL6CB5fz1r+B+otxdBx+Fkw8Un3Pghq+DRb2cDBZhbe8DShcnSYJzYXOUhN6a+/FkDPnJtY4Xwdj
vzL/uuzJUHmG6hLjxEwgsQAToxc7NFBc7BJA2XVgEh6Pi9zR056eG9qFtS6/ISTU76+gboFgfCp5
NcKFuwfYE2uWWdShK0JIh2rRM6iZ+T3eC+J1vLtxA/XQuN0qOq9g4q8CPoa1WJZKEr6DkGfOj+/P
CZvo88RNH4805Jvpd68nCndTDNM2ceCEDEDTzrQY8s7lZ9rwsHhBL5mtzzk6UT2b90Jqg7dRNQCi
PwAvYmwau6zwXtjWacd+8BCTiB/6lOC4aTXLvCrUvjRJII5+Q+AUEtDTwKipIjuewi/EubR/3LsF
yw1hQIm9IQdN2wxdp1+xmonfoFbEb0XdiL54MzANDdtrKCGXtGbq2X2b6MyAAKmAWtjovgdms9c+
kuo5EGtgFcoNHotEkxrKOQam2y6uqaLOo6Nmh2txsrg5GD8Fk1Urv5Fxe+/Ka7y+6tFLPtZVRgQF
nhRs3D8lAzcIp1k5lEWDT7XWCa8fI3CCxfvLgJupycotkTzPF743eJJ0r6Go0ZkXk48+K+Ijrwuh
ka59PC2Jpk5JSCBufYc3nD4AxHMDEmNoTv3wzvU/AcRJSlgPE9lx9rejLE2+o8lcHDTpHJ5G0QSZ
VO7s2a783IzU3wQ6YZfJWLasa6LoWqVvsBIKrIRhQZIHKcMJsm69pVG8QIhJRThdXHm8j8ZG+F1K
I/lQBhcOyn4J9mfqxknzQxELa9usWUrG6/sk7S1zkIR3cuHsko1aWJcvM3uDgCNESwKqAWrr1n33
gPsZTy/vyoJiGA4R11Fa+pZVtGyAV0SoT5RAtcp39a6z4VuuBSaJszbymqF0DQaUFQk8HVfUD3sG
T8IzjMg3/lA81W37pUnrDYuD6SkZa1iU4IIxN9oYkGUUjOI9RXbKncNdNoqZpD68AS126OE2+s7S
bdqvgN98UjQTGiJk3rKGnXLSr/5hnGsL1sS9DJtnEbV5GCJ+EidrMdcGIFpA1GKi2uBGNR+75MwM
rorMXDCFc834W2vYEUi7yiZW0mrQO/NhGGJb1iWmEFTAXl8tnhdpCFkDl1TS41a/eiEJlbSggm/n
MgvTODG457QWV3UyfYZmFp7KKblojmGiIzxfUT5mhyKkwQe3QKb0ztcsjEObMmWusmqg/+yOkIkN
oSw6VfNOJrKtNdXH0PSgQLzQHqUiZaZ+k29wZsjNDJ+iAjpkB5tyswYjtzmCFiar6RYoLq3KWzqc
KJ256MWPewGSnq0wx5JNfGPacS3hqHDYQZIx+4HF6wIIX1DMXDZcK/cYPBGyblaKjrEwmFYWRm62
4Zs4u+qL3Tau+vwU+GdJADPab3U0OrIBmjmRaVsQLIFpUTfkXb6yxm9Ej4XlfgvSzDhPtVmWCpEq
Jjd7xdk01V92kMOy5L9RXQea9sSILw47Lkm6y0f/yjMOD9VitQHKTBi55SSCSWWocOyKDmkhSO6J
CVE3mKFTdA1lNn3VJX7jQRwh89+i0mFtx0cwSbNg/9/YugnUrIVzzuUNtgItWv7WXSNPvzn7I0jj
EB9ZFg95/HrewgcC3Jl5cavPmEtzpLW3cynmbKtfU/PcHGvdoW5IlcwqDkWm6NgEXnht1QokIFS5
yOOi/FnlEGnM1ibjD5hcJ9RmzzU8h70YDWMU5RAlCB5hOSevClKR5mk8izg6hwR4WskujZk3do7F
Ef0mdhJKFhOmqEit1YsCNg0mwHy9tQq03nX0DmOLsp735zT2IW3PkgdyZWgYcPvZ5n0p/jaVKrTC
GszvGr2xNYcyIWTl5paKvE0g+u1Mc9EKnG8Ds+8FwTEOgM8YrQSQnvMQws4tYH05WTymX07hiFns
9Tv98Khs6HDV0AafaVSoWTb0NCtKJBE2wUkxL36MgTdTSsfazsIAfiLLrEMxI/0XI3uzbOV24NrA
LyHa8Pbi9kxkuQnJB1bG2OIjMCBamEJbbSFnFLDoDj0oTABWGoNjDZvJjNxOoGuKYixr6m5pY/PD
IrzUljNFQDDtTZ+L0ybpLRu4lmLmSTyML2F2BcQE4RrKQnR88aP/zPXJPPD0euAyZTNzMTv83jEi
BjVJ58ZEqwM8lHjNIwJTDKg5fLqyFTBVAn5cKyXju2HbucvLlj1ZbMOL3qs/HYE2trrrtRkk2nJG
FIzbwdWMhc3Viil/ZhRAVTXL2Wwkv+UKSmYqi2DceF9L6NralQMc/qkEuBCSoEqrYFXpL5LwhFt1
85aIMATZsnTZGiCLSATh1OcqNO+M2zjYiVXRP8f815XW3u855UD2mj29R8CzPIZaY8sD1kEIPCuT
1hxSvBDjUy+3EaokshaLwKnFreDcgkhSsWYwFIxOlTexKFVIHbqwWXLsakmuU6Ske3NOUrYfodsq
MzGBboTIRqxwmDmXGWCDa9QHEUKzNuMvjP/0Aq1fkjAWt2LwltOKaqKEwFS28a91uJLKovQZaAbc
40Ld7h3H/e3CfXzsMYFx5i9Qu9oWxLpfvA5xNZqqY+iV8n/s0eM0DK5ybs8v3LOVaZy/CtzN5bg5
pwUySnMW1Hsw3kbv9AImfdbHIxHAmW4/Sb9TVF5hyN39PPoh8KjfjcMdaI5Mnip0cfHV8d5f2sD+
pjrryxANxoKDIDjoITXXNI9EnUysMorSWuxdC1aKOXo19MDUiZTFTuteVrAFXo5DqwuGceai00jj
UxP+bEVIh3V34rvqr5/XJ6/BSNod1mqwNvoodS/r3wWwLeyWLSaDdta1cGpfIpbSEpFQPXSp4Jow
VUxgUtZQL9WcBulUZy7rmz6L6lpMUNAfP81uGKE1ydjWnH07HncR2D/Tb5psJ4r/yB+jX9nGn+QG
07PAnIbhdmfSzCh01BGJaxQR1prc3lP4LtUIrv1pqzitjfZD4h7wM5q+fse8Bwu1TpRm5SVEsueI
slg9Bs48B3eb8+0GIn1T9xmTBeL91e7XleFLolH4g/A4OzwYwlaDRXKkzvzFjfA1WJHSgApWG1mU
yBgamEMbrh4uGmyQefOj9iW6YKLuNnVARhJaJM1WO0+DNHn4j1GbihIVsaB3uJsPS9ywE3lVftPI
Z5pyLzN7A0cUf2m6otDyqNN/amRjt0jHwNu9GUfQY4KvanHGZ2Aj0ekED2Cxx2KKErE1RXIDEho+
23Ep6F6McXuOspG03inaCjVBVmNAmw/S837Liwmtod8jlYbbOCW7abipOmGoSbCQo61VV4LTy/KC
NOgaHzmeAGAPjunCJsNEkeCREuNi9DfVEQs+bfEqocyYFEdzXtWSDgHkRk1xJbNSIn5T20uV2ILL
hBXBkZu915F9NCU798j2Jkn5G+fVg1iOEV9R7D2ahlWkatvNWgHFPgLp49JqB+VLh1NEQngrt04Z
a+X+g3Mau+YdxccWYV+lt/gc0j2i84UVnVGjCQveBcWULnGPtPACzud92WXuqp9U8eNul8q9GAiA
Uw2ni7o4SZdgywUxhTp9cz58QlBXZYQfkv5tHfxuJ1J9ThlwhbpKTBCIPiX5Enge/erIff98NwLE
omDEcha593SjxVHsr6tnB9UT4QVli3TpkFtwggX0gwvmJx5x+qn2E1ZJQeD9fzYyEveLnu8Zips3
vf/me38i3Ev25/3NKEEDeSa26LrWR6MRkayqr4E6di4CzOF/LdSMzP4tiSSZHaBLslb0QIbQkyOe
0kIbXupUxT2jyBQap2szjD/Vz9tLe/CmH3QVsqPnQs7GW6krbGmgBMLxXKFzmhUGamADb6fqI2Ka
4H1g9RjATN0vzbbZYdkUsCoPAdVlUCedIbk0tzqsYWABpITZOX1Y6PFk8c/rY/56wNvwLONj947G
I8GYZSNyYEGsf1X6jeZyh1B+Kfjte3Sn8AhsCgpFm27iQIdDY/8sleqee8d+kFw+osrSmP4qhm5o
cLTSDiM/mQenL2M/0gamDxZDWzEQrqWiZUNMlDxkpsYaRBZGjqUjh5TarOwZxd1QWQx/nMWJjEGx
34lt3t69TySY6AgecXaOZ4Ef8Wyus0xhTkqCIqegBzCsUh0+Rk9F8h/tm5FlMXv9+11/nUw5aYAg
q+meSmtExtAFpxYeMrrP4/52XwMbZ9RqE1vujTXwTUP9YuruFQby3G8P82LcMGmBgLeSvIQQDwdk
oLknPjwwyD7WB2FYFClTT4E7cHxH5sllwms2zQ4R4rHv+ilpWoMG+44QltZvj1BwYQYTxLIuR4AY
o6jHeAbRO3R0I0Emsl7so9OZ1CpF3fzjToiTEtrra+fVM7WmS14zpFFaa70ExZB26w26UVPfMHCh
taZDvH7ARLcEddtqXEmiXqFVgQFVThRee1/v7uWdlL1GRIRMM8cW/wyOaC2NxaQdzke1BYwCysQP
p+VUaAvRgeNdLjpeh23Y3LcoGVuN5ZXsldU/x39JW78yM3/ol1AyLjXnxK907sL4Dsj2bpUcnD/C
h7gxqw6yKShIFsR6Ei2mcugln5DS9GewoWoyIHfIRkKghy38Ed/wgOflPqRSm2dfstfwnSd4EG42
Ca6X+Yd6RHOf219dgQdyH6Sn9dM0aWGroCWiedgEMlC6+upNIa7pt/KbxKolCWohJubEIVBU2q9n
f1utrf1pBjzeRep+kDg/QNYLm1uaCTTQRrKWUZhqpV2t3z9VZmiQWGDLZJfhZyRtItpIooHpWxo4
nb0mBwQwA4dfg1FJhDBL4xygxeMqEGZB1eHeG5anqo04VT2X6xyLu1b+KbgIcHvWITC6nnG7n4PY
3WMoq8KHA2ACfJGbNzz0j8BRNSZvOZ34ls6SgObK4kchnOsLp5weZWEeGvcz6l7Pl5Clu8Pb6ASQ
kaVJUP+JtfgKO9m+7Ey3vQHTdyJvgJlPoTlXH6QLG8qb4FO/f0ODkZIDwfB6BxTkd+3pzM2sfCgi
/GraGnq/cxqLIXcfemUVRvk1KREadhWsW58XnBTsYiL5Ae8NB8YRTqYqoNEnmuC6q70UD4QQkfxJ
PMDw23oYjKPHMzQtjfw0wKeZpRagceuuKX266gAC59ifuaXqo3khftgydbyMWCIyv3ADyrPZV/JQ
2AE8u6+GmAy11LbNPlFEmXDIoFI8e1MIwfkq7lYqN7quhzFAAwPe+nmdrItwm3Jpxf3KzmWnbMXE
cD5dEMVbyoQkna39tYnS1zT3O8O0vuO0VLtojM0ViDmPbQor2lwu9+9sNVTH3Teps0n20zKJ1nPY
exhlyBae+Y4aD++2vQfFNwCasDgn43GsvzSXnB8wYPA81TwWWelLYTlX/FA9U0KLQ4TVFfdSGskz
kjpLa9cHSHFUX30A2+JYWLicFPGLQBy0h/L/G93VjANY1i7teuKNrOtdIepaaegw1y4jCU1DhCVh
J9qm7GHyBZk/52z7VWRznvCumebtI7O27+a/2o73Xj/P9+kE5m7iVyrs6h5nZqaKS0yFCBAglxTM
evzuDSysY4XH28UhECoeYaCpwTkkPKV+Qw6lkEmhRhOF1USbaQLPK8pzbW12sxHs2XGO2OZ/7KTA
4bJsF52j1Z4oo8YUVxt1yfQKsqEaDSDFO0XsdsGn+Hkz/Njgdu+0fs6KBX/uB+0rHe1dmzLCDDKr
mjqM+JSmxsZpcfVBLG7Eb6RatZ25IAutCqlQMlVkJsxGYnEUZ1kVjVDYuzLCE2iYjiY0vAgrBkCs
rK8CmtD6L9DVGaIznks+WSRzCUN600JtW9eyQMSbUbU/yxMXLBuDceJJYzBk9QKgFjkN1ORIK7Mt
DmZmEhOvCaXm/Y8BxI/6e4HV1ngWAFp++9y7g/MmYrl/Q2kuK/5dfD9QHgGlxfGpG6r5QOa+WqRw
SXbXkzgE/L1efHdJzQ1OH/n5lrNcHT+mtd8TQbEq6H645bm/9doKBL+llxmnBPIRRRjWJrDoHZem
DSqMn6Pq7JD+QStqAQuwxb5opJhrz9ElkZ7PMyTKIftlirLUhZ3E2w6n8KRtQ2IkC7JHoSUD+E5A
/tU7BZiY6TARdd63yryT77piRcVCFkVbL9qVQgVKAsarJEtgLWwiUnRl6QzVBxbCDpZSMbbzqKN9
7S0biEcHNM5rD2xHyyK+2jpbHYbvOM4YJJucg5YPq+vHeHDZHHUupDvEwIEh78yrTcDxSQfojzeD
c1R8lazYkLNY1RFn9h7Dy50YP6ApDnHsg680OAWStWvFvwIQb2z6x6cQIXrtTJL4PTBJKUcEDNmO
kZ38ZceLGf6+KpO9ofbaUiUGoQMWdPhEkCI/lxpI27FbeK52V3RI8rJZj4MD09rYw2eH1DxNG9oB
MV48UZUAkbBDDUiTW0PRn4CR1jkQGkPWkqzWXCrEGqPo0wbGpDsYZan6m63aztjrU5MAb26QKXVI
2qZv0OqSN75CDjPojztgZmvv/Kvi69lqQqkC4SMqjGZZwacFzblBh7GC68OWPzmARDSWdg8W00Zd
LPorEzwjuqiquPwiFNlML7zCeQhat6joRP/in6MdBt1XILRmPG1MjMsUTlGJIfw1zfCUPgnS0tu1
NVR6/WaSCvycxEhL9hosfUN+Ze/2ou0oFEo5vfNpEnP+oe3RmldB4r47I+NwW5NYl3rG2Hqfv2Bs
9ahLep8C9VSgBwGEF0GA4kW7D2vWGKaIixOj0YMIY5pzSIq7ji34W6htkCLh+yyZ+j9G9FleFx54
50wo68MF7QZi3tcdjY9vsjJefe8Oc00W4uw6NjhUCZPee//WMyHddBz4uDvT87IhdgUddAKiHSoE
0vz2Mf91IfnvT7XnnHiB9m0AINp3SdgEm8/Lg+pb4kdpKV79vyWEnqLwR7F/A4pN95wM1X49fh+x
8Qh3OA0icO6sHBkVET6nqqc6ePb3mqCJq23MjzFqaJ+Y236aFzY91uevdjLf1d6KHyRvS5anktls
ZkTYlaWlOKV79a2IHl65BM0L3YPiJj4cYCtrcf2HN2Xy5dpAxDrYLwdqs9LF4MV2Z5zh3uQw8+7B
IRI1Ptb2gsyIjQCTapYGYOKe+H4xlH0UNYPQipv4m+nli+/yV5cWkpUGCvEmLVoq98mQK64+uoTk
/MQyutCktiPNiwHm7YrCa4PYFUpoJIdsGT4m4MaiHERIyXl35MCt2Vq0a7uKt3mppeS9uZxey+j/
p63gtZ3p2mf52H1YsfAObMjMJb87rKL9EsGJPvHR7yXQ9PDaxsH/YJ4seGeA1HL3gnezevgYUQAB
qjR4sgD0pLjdIccQVavlJ8TIi342MFYOCMKGPKfX5Dw4WpOdaSfstQ41a1R0lNsT2iwRH6lWBN3R
Dcfhr2oHUSPeUqYgCSmx+Lxt8fo7o5ndXh5+QLgoYQ2IiZ0j/skplDVgNl51Jo8V2RfnElyyY9Gd
Wi60U76qICYlcwx0fpmFGpsUxOqepF7mMBHYtmP4VeSr2OCXkgj4p42qQCdzE5b3T9gqmfRr3saz
ZkTWStD/c8WvxsxyFNQdHx2cYZkSpyAU7qOTPP1f86Xrdw97vb/3J763dgcrSzTsRE2yXbBo7VAk
dNvWI8KSwqXWjVWfPhWVYSt9Fa1dD2FnR13DLM1Sd4IqCHXbguQQh4gxj9u60T+wNewmjWb8MjBz
KvjlBea8mTa5wsnOgW5ryyFw00GfagTq0k6RtDG+CAHBy0BkCIO2te1Xwl7WOfCWvA4jZY1F5B+y
XHgaK9ZCsQD5dJ3Xq2+oToVOIgK7fn5UIctSd8JWkuOtSbux+aOIBSn4ONkho5nBmD0GrpFhWg5E
LXmOvnzvjZJlHBz38wf4vGfvKXA5sFZRljjwfJhkg9c0pK5sacEHpKPdfAS0iyWWMRTdFBVAazOv
Dk7PsHqrQInpmFBotbG6rkRR7JJR1bRVPng1bny04DISG21/69xAXtWjx/6fDeRyW8M7vvamt8El
voiw3A8piyi+BSdirt9Yz3sYnI2BLAht3YPO9IvcsMggkzufKmw51idtfHuTHW5kobZy8ridB+lx
qGriMq7T7z9p8Wesnu4vNHBoUOwJAHhV4B+tBc9LoPYr5552WJFYaE183oTAPBthwxy65XqR4ycR
cFefq892TYoBAQ2qZ8KtAQjRsg8GrKuD/QtPgQHx3uKq7bckTIxiATc37qoed9LhC0of88cr/5ow
8Mr1bqUGUpo4hFXBezw5NPFDfTP59AVJ0bhg/8dttwI/5V6fAunW1o5cjGTCRXviBWayzPbayolE
ZfTPKScMhYzh5dOTXOd62UmHM7PPjUi6eG1kEBu6qV/WoBiuwuhx41mSRMb7xrZ0ntbi12lUMvNp
xmnxgax1V00q20HjCBM/4erUWSIuapGCAlEX/S1tt2tLJ0ePkFdNXPIDlUtEg2IMar27mCo0fAkI
zbm4To/LZ2ybm7ce6ov1uJXPw011S1ZxH2ka6ER8TFWpYPNUV+/X0KekraPqT15nyTc9SPb6jZDz
WYib1OcdmUnKWyN19ofcRKvSXtGE8kpA76nvqAPep37eoSriDijyfhSD4sDGKMTWRfIVazkU2yx1
OY/NX40IlbxRk5NFh838uTC8T+hoWuKLsIFdDaM3Pc+BSJWIBqO1A6z+TOu0/HTU38+E+H6SaeZ8
JP8YiYdkdvcg8bkt5HhwkyFYeKHf9GbDr0CZEtVk2bOxb0CC6ROK7oLbl15sw+OqqzMq4PbXOEc+
gZq27O1YQEnti8v1+rptcz/6cqqBy1h1HUhLA63jIg4Fp7LY/Y9sNq6Mvf2bsMJFM3Hsmyxt/2av
zCBilHQwymXnPeA6f8Um3pfYVxSJaRe2v+mSCGO/POVEXOKp61jJ/iTFyT7xNGdDPCR6QVOmE5Ly
bcBNxj75wZSAkxJ55cNWWTsvzu1NP5VvV/ldxMYeg5OvGLIwq6DrDmOoBEQgyqehecp8Rc/z2IOz
u6pyhuScX2e66YRcVswC0NOX28Qt4JJxmnMIh6VvXx+IIDvmM0p4tlacttVsEl9CNRDBNoqAc6PV
9dVhw+CCaWIjBThjwSmB8sMbMAxK8vJXaQu/0lzEDr/0aXb4Rr/K2C0pROYOc01p/PH4lVWtBvf1
W6m0N80MwDBxeoleoU6S77U8JSLjT+tbSJj5NluZQKNjZ+bx/RAJk8wCCu1rhHe9/RE7bwtLfOOp
5F9izpI0Ae/ElOwiun8x+ImYz2qvkYjJHEtXYFuMiyObE45+Fg2IngDPnyk74eWYCQC5gbo2yhDj
AaSRHTJnPkh3Si1dqbfCGNQ1QepOszNMeRq4tCXbmEJmTKrmDnGk7/MFmiTO5vMz1o283BKtzJXL
r10A4ySJtcA+B1agS9d+RTR0uQ1aFKCeqLQreG+gyZipEa8xIclURmYh+7Ujaberl0ivaDsb/JtH
VEjE8jhm5Y1Sw7JAQUnObF2rd5MvuupSzpYVvYURKNzTwNAahtq3RQ1RXObKB3pfhq5wGfb6hucV
QzRrhJJ4meLciwwIiIiytKA72sERk2seUbzjScOfsDrRvHcXzbIw26nSpkDKXgC67EgN+3tY9iSu
Lq0Sos5iiFiJ3nWq5ypY43MHvytvyK+t7tVHzCFLuggXVWvbmGAwBOGodp6vXup3PgdBo3T5r4Ke
Hd1KmiaBdYt+lSfnqwA6DaWtLDq4CDSQFAw+2tEliTGYIguML5tlgGIiHNCH8RjQp+GLnLjiTxfn
W6rNhQGQ7ORDQWaJOp3hUQmU6Fc6dKT74/3SK5CivSGDRbFyNIXVEdlmLf1KV0yRXMy0C0EoSsDb
COwHiff1GByaDEFfpnBq4WzR3nVBajrOCeUgGdMDn6qPSYnYE9aJr6qM/N72Sj052iy8XL1t11a3
L8IB+1qPR7NnpSwkxLldDDf+OR7KboBE9+0tSJTRhuQtsKWjazPCMmk4toaU8z2mQ3vEajkM0dNN
qNRKssP1IXYLssfYZIWO0GVw8dvf0uvsN/0XEbB0Yk1VRh36/M+7r3uJ5rgHOtfuIIKPA8PrYw4n
u8jpT833t5ogdttqdmc2/ol/HMU5fJr2HxgiKGpsiGroGZqbuZtV86+8r7cY3FCKWbdcqtaGqGj6
sj0gzKniOFc92A+EKJVyWu5wl7rruWhEVw0zzXjiUUYCQnN6ig/cTydW164Khi98JCYjgF8CVm/I
4/NPvr/sqpndxHvzp5MUwFUiKxelrCkRbeFY9wbbIkKvPZaMwNGOkCyDtE8ps8xLOH8lodO3ZEUH
S3sFZMmVM7lReTarpSujQNvnCk4qZ59b3naI138hHmWfsgxIU4uvcmKR/7Kp05VaofPkd8bJ7VWN
0mSmrtrINzFNyaOwvzHhlDlQRkc+mU/vIBrZ5UkdCu/GD5IbxasA8UGrgcXwIkTkRIXEajclvGxX
bt6EdzY5XYCp2Nnz5adUS7ojZ1eYqH+vP8CQ7CR7+siq9lQ75lPEwgwE/kcpfRFUrd+IRwyGK1ig
Bhx7pzeUzN51lDz6sq1gOhbw27tazMcKQT2EM0gF+8uqEyLCpoo2opODjumLQeh0fIBn1lLgnwoJ
c6LpyrnIF4LTBJ2qk1vbLvv4k2mBAKiBJgEL7GgJpNk5mrKgH4HCUPjhh4TVO12ja1pJBIPdo1RU
6exv60sYMTmHqH7O8TlF9ZaePRN8jDUuK9XJa7bs1iZ/13ZeezsR5bao/edRZ+YArpWb6OYUNcnF
c+qfmolE1DMb9BLwxN9nEJ/X3q7y30l7LfjRR/T9DzMp/qBK8+kKMsOS7hTHzetLxC8crbNUlAHN
Wb1bH5jEpdaHFAx5CTC0gGLCjRfeF9PoeI4yF9gs99HUd+jf74FNoq/lwFG7G8ydVlMkViJaEsKe
GcDIZ1GBRN0f+y6Db2OhThB/KF/3T7U9sItcxgDeun3pxKGQG7QNMrEO8BUaoCGcvjzYZ3LzsK/A
3noOjHyJzR5Ts0eF+z2S+pE3bi7dDOrssstJLB+HH5Ugx5WXMci2TciMoj5Iq2iEZVa7YlEwglCU
gLLI1J5HXVQD3SW//utcvt4VwLUyupfrxzJGGohadyXuGXxlNN0gMN1aYlC9QyRyt3q/2kfpPNIc
CoOwO6FN4McubwGsGjqc/0aYjnpEVY8v2YZ691FJHGPLdKvoSbtf+Y39ecKU4qGyMY60bCgdcivj
d9/JD0Whf6LJJ8I5n9sFTxWVkSx0JwdwzLwNXo72HoVRwcVjWKwnB11AEJIsET2m+9XuVYh2bkV4
E4M4YrXMPc1CSk8dn0HmJNQwR/tbjXfF3g4SWuhZfgcpDR6nPE4ea3+2hiFDeUkRElKsJgBzWVRv
GDjN6XHzOTL+QAU7UuZyzQ1SBRNEJ/7W2HAd+1Z5uOeDfqjn7U/HaUIS+ZCEZIxrmxT2SzGXgSjx
vz6hzDctgiLZtJOlFFsSfR3rm4XuGeNXFnoMb9ds3QHi3GmUTVGhKnJ/1HXme0IFJHduaX+qaTIR
rqov4dJA3pfmGdvTeNZCsX1op2baTE527jVROnxnLDaGLYna9hGiVFCAXHpibSFrTAnashO25SmT
E+0GQf1xlzYMOhAJZ8WvVNLepZflWSC5N+Wuz4OHW0gwAkUc5YLozgyMdtvcJaMhyx36K989pV6D
PH6XXZhq9InYfY5IkC5FZhoYlT0QGHmISHu8FFErD3uLAYpfnikhdh2OKzvHgFABYDt2VfPTHzXV
ZpRQlUYU0bNrE+9ZTWmyPbdUqS3vNPFMf/xy15FwmKrc0K8LmtQm1zrgr53LebfGSZg75FmjLpwR
5hG6X0b0hn8DC7JBIjL1hSw3AcFVxAY+V1PAEqkg2DSIY7xqaWaf18Cq8yj5HcKnyhWr4e7vrHCJ
lOLVfgOb9Zx9AXt7ScsHmjwyZBlLWxNQsf6OE1zEg8pps11Xc3MMDIq7WazOtVRnogaALlfXqPHe
nFsw+49LVPurAVmfw3685cq3jZgyHZE6bY8KUhHljXD2fjOc6vSWFJrMZn7tlrNHR59rq25XcPma
LJ+HmOQq13RBshcY28ZZINz2CorlKBJZL5BRsDCM87gwKtDvrAxaSvXRWDKCSGcMVvDjcJeU96s4
iK3hWV9lJT5ncLNHLl7CYo/YFBALUUa/jP99OB/VFh64UrA2jLKjAaBreTEb+xm+NTrX1fv/2+IT
jmU08CaCXuk6uEZbxMuBiHTJETsc/g1ODAlJ2VBWyHHbY5tD8u7WG8A6tYMxCfDrC9Zq2TPY/N1r
XVBQ1zG2yVK9x1UGQK0sDFuTvfPOcTgGryXK6CG1KtQfahGkz+oXR19soEHrSjhyTfkBMnoJF174
DuAwODRLidWk45Cpk4CRZy9leieNKj2vxYNUGTX364mnknZNRZySbXkWzhT9aTQYGnjkhwyEBq/K
k2aDwkR88Ul0ZklXa6KkZsyGCz4PjkyVoXV0k8OQNs8L3Img/uWDol+fn8BAzKqiFnqtxaG/tpun
Rxz3ba6JWOsgFpA96EG0UxCUKA4Wejgo0u5tQ2axZvexZrnXnh1Rr92wjZ27CJSMt+KhCqJkb6pZ
CIXTdODXDV4l5L8eUBIABJctd1hTK2b3dgS6sCjYB7DxiDO8vtKEZXa2i9Z29d12ZhShKDukpf4N
xJ6uzkfTWa+S/gnpB6nMWW7RuwXkZx8YzLAUFaut0vv4kwbouoZ+xRk5l/uQ3hySt9EFQMd/Ii1D
zxc05j17KA+7fvVL7Pcw4jwBsnxBkR2i13jdh5IfUGfgR8uGo5/qz+NtNzMSUHU0+O1fBnf3HjAD
4WOH3z5m9XSKtwNdhAWFAAev8iAuhFv8psSiTujmJT3YzApzjjGz3H4HInoAq6NHiDrNojdmqCau
11nYpjJ1nxRVtED3aZsVWcaC5tFQjeO1BRE9aR8jrXu855S6Tn9A2GuVlL+igdJZ0aS9oVwktYuT
5i/kdYN6xqFTd82+7EOQKfOOy/SgMDf1iyj+tEFH9gFjjfuZPiCas/OPOoMgRPlEsGkaFseBBMI9
mMnBOI3nDb2illkrb8ns9m/Bel4axYyIMH2/Fiw0d/bhXYCXB9JQUtZxE2jyzP8FnMyTq8fSweM7
DbbB+8dZ7gejcOFRj+VfyWgp4xMFk1mxx3C56Nd4ebKpgVsJ5IVQjY9SXPAs4TaFPR5yczSjEMwU
/VmlJ34dLCHb+qhxr8zwxwHXyl3DQllVZBaHbSKgrkFYLeKQxnslLeIqPdl+XFVjrw6wTvjOz+Ol
qU9iHVp9ksk7OVCq/qblFg4T6VhU3mAwLirBmA+8YxnaesqOJXCLSfFON6r3RbNQkFDkatlF2H0a
G6SEQcTR4P3HZz/Y0VvrYYBMXWC0oCWyOpeGL9ANuDClUiKR07VvEQxsra9ae90aSZ93BwsExhN4
BMR6NKi5AxPVZY9nBPdDV+V7k5xUgMzIvu/2UKfLA3FSNAIsW9n4MBPhyg+xfmXYLAAx7p5uJXJz
VN/pMEGUZ1UKf1RAPKM96odCS/KsWpKVO+aU1zX/GeE17al6QEpJY2dwoBfB6tQS5RUadqnDJFss
ls8pldIn8pA8twKH/i+W/rY1LSa3yHu0+PluEFPppiKx+gtSD03pvVQVEcNTvBU/mU5rlfIzfxpN
ha45ZqJ6omufWz0yQWOjPPmqKQkFFhj26BV2qLf9ljbxvgOpCxcEIltz/oyaleyXDU0hYhyc8zgj
niRwWQsjztree0cGOE2vxyM29YzskDluLdb8BXUHMq3ekYM6hAVibABJJ0uK8+/5OrNI38anobLI
k9AE+dgSplflREsjBluvEvQuye0y2kKiwrRiMRfgGVbUtHAIXhvZNaz21HOsvOo3KsODoWb4DZrm
VYcvszcH0Prtv3l/JXq6WWxbcKpgA7sZ+wRw+OZiVf0jdwbiGjJefjaGb/IZ14CmA3YFLwGfZs1Q
M39uNRssrxhWCa3ajUYUnNqaMh33U7Usg3xgimpZd6wdw+r/cR0UQZJVM38L8v0dEJ0yjsgorboN
ptYCKqHIYSVtwFZITl0w3X8fOTwk6SZMFadT2WJDo5e9hpp1VXsYQRcwA7BISSRggX/sSBpDRKsq
3C6JWVMDxH9OJ3K4FfKbPbnRMzwXkfmS64IEk1prbzn7wNLSDKz8zD49geKarWN7e62gjvT+Yavq
Gi8GngHHnQ3TBKF6STASpr7flSli3wfND4YWERe8lupgWJr61Yg9rwi20LHhhJGUt9fWjbCB3gcj
6ckIhLlnnr81jAaJuB3KmNQoOZ45dSr5iNDxJJvmVi1/g8m6Jblk3fDrOZoGUOc/4h50Z/1vvcNA
tPEEVRVlzayFqR3/Epjcd9T5MhuqB0A5Lsa0VQlID5dy3GdxA1iwQneLSDg6ytPnmRN7g5lgN48W
CGc0SB8hHp5sRCqE2BFX5sL4ui1ihpm0TyyfW2F6Dz1j8CrMdc+vzZwHOWQOobOCZIqV3+g7OQOr
Y7AjpGIH+4/0a26hMse0Rai2J8lsm/dbY5a+WFDN3xdL2YZ13IcZZ94cZDSDSdkAsSphWF5I6M/k
ohpCG9W13Kw/xejQq4cCc7Hh1XAmF60aK6GWUSsfZIc4EEEjG0rqJS5p5rfFLGTM7Zc5al2N3Ko2
VBhN0B64m759/sebwZwgImPV1kUHmdQLNfvTt8JiuqTw2nhUGLVUd/1AjQLFGfNN+JU7fxHWq2Wl
ja257qgb+x1zqfCStNhd90bhUCwEVakwjiXeGx5mzCCU8HZ14xcVReem7xd1MzvgG0BFVqloB/to
4QuOlyhjKNEMIfgN3COMop+8N1j8Ui30Ll9NnUodHOh92lSknkXULBrWCRpCnvGmInHspKNBgH6U
YGgKohjyvcXfxJVtuXCxXoh+3HGlOwz3vNx4bKmRtYJ4T3LDLR6MJ4BVNfobiYcC/HRGT6xHhFak
sd3BtcosG0SJU83bRqXrDs2Cn4mq0v8ubDiZc0lxjXsI1efGvr0uKUd+8g5Ip01k/OnJTkw7m9qA
ekdc8NEspTQavzlAHUCZPJh38hLjE2HBsU77RfPa9GxIahaXZAQUxCJlER2jRX+1u4FLfHTbgk7m
HWff88o+dIMUg6Eghmu/hnpgbe1snEx/XiQtN45IPlfNYt8mFXS4Z7PzIayjiJliDxUk/knAx0fG
xmFkwKFlSSqZnuyKeTtCW0uv0Ze+UtJmmjy0DjYKYzz0qJT2r9pbnTQbL9n1n1SOonuIhayRTZg4
PbkjwyqLmuQYqTGnz91Fx0Hy/FYeBnUko1I6z+BQQDfkxKHHQ2sCDIvxne+2H2blG4cqed1UNc8M
Mf/NR9oqgVacQB7KSQRgdPW3lZLfe+HKPIDpdXkKp7Uj6JgkD/rkwlw479tdq91q7ckFlyX6VmA7
j2pQKPt31YYArhvVTkChP6/s29WQdU6K6KZ14aHM7qDCfGld/wZi5AQjzzR1Z/p3KumP8wIZJi+Z
pcYNFOokqOtuy9Fo/3xZbKhZnw+s3CF2r6loVwSEXNDXmorz9sPvZi3BMCtwXYK+2ByKGf71SuSS
rwrGnUFuoKHOF9Jilf20qtmE99HLh2l2adKa/WDqUbD5ub6vfDVMtKstxIFPhcotu271kaBSIFKD
4nG6TFQSaey3CKJRQOu29fak/vuU6N4sYZhBm/mTaKtdvX4x1atiBGqN/QJxaumhXf7p/nDRHd7F
b/uW0YCKsqdjJsZ/NSSkTU+PVoQepP/1Ts5Z72ONhekkdf3Stoq2qiLFUde1OgkUCSC0G42uYBuj
KhIKvtG9CKua/YXicn67RQMcvViZV0ilRYAniZ7t7qwAU8kZLDYVV2J66M1mbZH/j0NVUgrfNEcs
z2SXPsMq2Av6svqCy4NjpArEKgG86WSMiu1/rsoNtCUEXXiM238GjH/aPhx3ig6jlii7lAAleq3/
NVFej2x8sTh2t0HMNSwnB6mXpFmbMpRfLxswDQJqt9BUh1b+mLxXSBuXVf2rmVEBi/+GndvFtPto
9uo0px5FU3fbxXCg1R8IdCdJbtP8iGa/YidRTDrsQc4FjcaR9NK5zOteX4Y3gMfsu3tM38Z69FNR
2W4LJ70u+TRZAOfOcbwJSnayE40xX4F0aLaa72EJihg3sFq5dhgEjNgVa17c4zQ6CZK2HipgaMB/
lcBTii552PkkanwkgrPyxNOWdFEVCHbnDZbpeCsriEbk0rRIpC38en38r9INw+m0LZzJV9T4FT76
h6apJbowo3TAaRnxhQyQVPfMs1wFNfek9PPgd9dX1e8TWrwdjXAzwPIH3iuSgEemBK5O7+m7861E
/Co4OUNs2wDgXxSZC6m3U3E1BnAocizlPbMJepSzE0UdXdBz8z7CAjinIOHmtuj9G/P+0gc8fjti
psbLBQYNqCot7C1uVHdbyKsxq9AYoEGWQ7rbwGOzKM+CTnfY7fKHBszJzHnp4DYax5yc8LaSqxVb
LuZVJXGTHB2dAmOptbkmaRCkZA+CpRotjygS2mjMiq0CFGX2oZyQL8XFCEi+CUs/BtnY0QNpFGE6
y8WX6rsDHnWiXHeJnOYOXIlXoe/spZYCfsshO6NRQ53soEair1nmNqF3kSr+/L7YyC3lMizCIFMx
h4HvhunTqyXNS8wXKRtPTco+JwJutOemSQJaTZ0hOCHbyQ74Od8rdN624YRnw+RPjlCf9U6Wedqq
sUvJvXStqfc5oNI7H1IANPf20REQ5+bnACnsigwpLtXc5Ksn1ilH6715PBsW/n8nspLJlhgs/58P
uLlW8La4e+jp9pxMykWqGB40JHsICS+zde21sf68j0q4GlmAkcJey7WQy22G8hDqXizLocZTvhGN
SB4KRGQhT3mfHEwauMIykZ2aI24y9QanSv3Qwy2hNIPK1bcHvoKB0LVbJCtd3GHq19CbEWJrj44u
QmIhblepvEwUwp6BBeDiGdF8SXCtlbKbA5dWPRf6UfhNsvdCR6vzGdq5eIt7H3Ed+FNyMroSlThv
EbahZYyR5UEadwOigQFmfmij3lX6etqiyP/WG8NJMxu9oywVzqOIQtCgIqdO+vRwMsW7jX8HF6pW
9CmQ6OehDhPrRnzJQY7Ge72mbavIzWGPSqU5I4iKt7+TISBdJnSDicFnLwNQjOqMPnkHaZagNbA7
tkPew9HqmZeZXD+0x5QihnVq+gIUnYrLE+wK7My9g0zWhcnJz//5zwgmi/Qpa2ug9wjPh6YDsvoL
KxokOxix2Ix/7Sh3N98Ii6mZKOYLb5YQEv+B2r0fVLa5PKRtg2//jno81SjkNJencxY1MYTadFfD
NOPIArZPgD3lFMMhqRKGPRLn31fijhpGZ3ZfWhv750scXISwQeXb9XjF4Cl6DC22ww9//Beh2kCl
81qvzRlXDtzFG05fy4WcdzsmhDBAYV3c71ONeQFsSWsuLZ+1tpr3zoP4lqKgIg5fNC2AP7m+dKjQ
oYNva4B3vS9aJNuK9APtqnOuUpMEaNg8KDVXn1Sd7u97BGmMnaWp4K2xQuB+UIpRaBXgX88VuBMP
1Rgfam4aFt8NIpbl2VUi3Du+14R1UuAva6/stYwyeGgQNtzx6ZT/HhBFt+ICOUSSLhdw8FZmX7gf
LyUBNGMc5/6U7fgNUkd9leOLGAgHkl0dhaeCfZUtimdU7vuEyDEiPc/b5k3rawQRdPph7/GG+Wao
JYz+umPJD66L/ezLpudnDPNzgey3YWEu1vO/KCGgiUoYjSLhBiWIaD1FNNIZmoYelLunZXDGoiTM
WpbGtUw8iO0miLb/LWCqE2iXkreY3fJiYElGxLFO/ReRur0iUUs/Y63vYOGB1U6OtPcJWq9j6G4Z
0vXO7fhlbTw7WmePorc4EowPSW26hvcvcKmM9M3GjeJx2Wvou8F/wqFYWx9gXGngh2XBFdQQI3vp
YLX3/6YlcwawfmJaaaMGK5hXMagaZld53ymdOmbiQ/lEhrm11o0mz3eFzSvcFlk+V1JYoACsz2rq
lCDHmM2LW0KYOdUn2AGnfr5+BwGhYQY4cJMYhql90ONzTpgAy4Lj7f7byEP6lDQR+vq5+0JM6Ic3
8vHvSqZfA+6kuqOiciS7zQbNZCJFOfhI49iRv8be6P9l0R5r47npGYNaPsOCGsN4yWd+r6fjUZle
3ESVsR0r1DXH16LmizwwVPBCtwJ91ROnkGWmq9fV35+KVjK5UmabNzuxFqZW4XbKTkNm2wwY3FU8
sZjW4x8X58nz9a2abldOnFYzstBIePoLQkGO0iSwlO2/MbZqRaHm+sevXE917CNaN00GufRXeqAj
xRpzwbBB5ciRRSs8x1kMhRZBQ325uQCsP61LsDyhy+ubevAfQ3yRU41Csv3+Zz1b9V45Tm3B+3rn
F4R2Gbxp/ky/4wY+W1He0Q/YrH/u6rjTFRwvn/kw9EewtstEmifz34mfKUzCm1HziqANThFEdScl
NgQg8q9frjgeo/0XTiM03kdahy5MtfLUK7dK+GQlfrgX7SyviM8SkA5yBxTN4Mzn6OQWMPF3PvKH
AOYsutDUlUOhirXn2lUOG/+3vd/ILF6pxVT4C866aboUkM+us8kS9gF3ZR19mYEsEG+oJBQ8unML
ELMNjV/RCX08EtWrX9Wt/6Q+MBYAQH9IxWcD/AqI02DfShP6jZrqFw6e5xgInXldZV9HJExvjQMa
/WS+UtQHht1NU+O4UlT10U8tYthmXA4E+QO+nIqyUOdKQvNTEkIvaTuRtn6VqDMq0zv6rEfprW5q
+nPuhJyCjMY44mK9MS3kbFo58mzNCjVeirH0QCzx1kEsaRZXHwITtE1JkuDDp1R+/Hu/tR6DYgt1
JJayIAsZ60cD+1PSxRzMB2j4htmgKME5RelmcZOeblGaR8kNb8OP9QDLkZ1T6czRINPpawuQACDu
5QZajA/nm9zQWukz8426tkLTZA0wxhRTz5YfAJgdUNUHp2CXrV/aLo0uzATuEKdCmNoIK0isFRMC
TAAsZgqpTZDc7DM8fkZYiS4hjzLCXof+MI7K2gj8HUmz8ro7SVwEuDEbtYd5eeQNBA2eobWGNK2w
YuKkg9+d+anTXqCULQuFfMnLUD3PwX9FnGog67iHaxj/xKEqyZqieRUz54qtfwg0BgO9fhQNONYl
UUfKJebjqB0FZvJ3KJbVeH7Qgde3OlV+Y2U/d6JmokxnnlJLY2S6Q1YWhAB/gLj9cdtCAjrpdoL+
0jP3Ai6C34vnX0v6yu0Uy8JGayIdLD+WedXADDsMNlQsIJTut/wxWZMbr7BCXdzLwWPy+dXsGR1x
ulbHMVNdKKNrQ3XrAyWg7QfMG0zIfna7tgCAauvZbpSYz/qmfeXASuRzNs+JDLO14SmLUoIwJ6HK
IDKMVlBzy7aKZiB66h0i4fhVcROiYVUA0KknUcK+YKsjVUYza3vJFp9Ydx46P8ZkeZi7n9+/OJTX
dmmE4PNVjV/QqR40riYBgmVa/YlFnCSfdBpuzMSwN/jWzrKb05Q9uIOb1SVIn1E1tYJ64H/kV7df
DJaGgPIlLe2wsnx9JIGcoAT3dJi+0BJhWZcOmQkTe8fuJsaW+qq6FobjPvtPe4wZxw3ivqMJEKtx
LgxtetSFfOBtPHpizZtnm32doPIQE+6foOyjXW9zCvgd79m8CpO5hBrZRWUPc+PJlU1+pZrjAFX6
XNnOth3cIlO9+e5dyBEQG1p06CcGemtd6cnj+W7yfKp1JiCcW6jFxZ5OObH+xFL6nL/WweoA5LI5
D9/+k1AYhh/rIRXJrkxJR3M1jOvcVVags2uBt43G22HfirSnBs9nt1C9fGA1ufKnHSrJVpMLrt5w
UWf9DUuuHNsyc/RhlSF/qqvM9iANt2xLsPyg4S1r77QWIa1bHx+xHlwHMCDVfle8wNwFkb9lXulI
fPlcRydcKs3lCOC0NXViKS/8kYTW/5MRCQLkjAAHcvDOfmchHHCCNY9kcxQdIIdvjf1tVTPXgqHe
Z4gbdrwPJNvZxWSOJoXtjqRzpKT5T+wpbOzguyvx6qOlN52euOEOIaInKEvbBXCbUsBmut7zEMe0
NuZAKrztsH/a0wBCUB8z2nmGwv5nTmyFT15hYD9xqXQbZF8L6i+qnJTxBRyHL+ksWPCUBqDpO9j7
Wmy7dSXAv/zFKuuP5Bf7iRcWFio2SQ98eRwmUY8kkQ4iFL3dOHdfue5KHdw3X0GkOvEzOBh2riN6
bbS6zr3/IyqLOQoUimOjbNmh7JNHF8fqquFLDjJxT5Ud5Bk8F9D4PYocZZSKD193LkfbYJJwqN+X
5upFoH/taAtOAlsG416VXXGII7rHfQgRmGqP+J2twoka25AbSgg6HX343FNbPr2spS4VtKs1Ua+I
kFHrpho9CNxhXaEKIzCS2uDgTAEm9z+V4hQnISqAQ/fxkwzwbQiiGayzZfPVI2sCMF8RHfE06euY
NmyBNzHdnFwI14AEaZPK5CMvGVHqX5EaSSH47QgSsZA7Ntv0FE4i7fsvcZRlwr+XNXi0GWCRGQPC
9jKAtrOCelMt+/MPSrUxidXKTD/CVs4VIuoUx9YlBGxC8r0TDFagej6e16DESDyT6MY7TQdnbYfx
zpWNswIDliV+39hM62lX/+dXFju5UfZ+AensjasGML6+3KgN8FsNjlKZI1uTdrc9p1l2IE7yPoFn
IODSYPM0COLUzpYJsoDQratRZ1MfGqEB9UpgFdMEUGj/R8RsZre04KhapGS9H3rElHiN6YSGawzy
cA7N/+vl2+BtLDtdcBm/9bBa4bdUKxb30sMC8y7MUm7eB0Qx2QxF9EvqUUbqohaNR0aAJuCz+Lqb
778QdNzgoKDhwnEx1LQvl7XTfnLceTXNhAX/TfNg/3R0S94oxQzoyvI4iNnUwvfnMNeyyWA78K+P
fs5DO6I30+FpmpTk3/vT5ATXKw6eostD6UhhuoAjdyGtxIL2avVRo1HSxkt67OcsD+VsfaHl2Yr+
gpx1UbayEmvbHy/DI6pXeOTBuGbGiarScQnr0o/vvp59N4TLHDuJ4xw6ZayJkL4WLzg2dMWuhT4b
DESRbjl+HfIdRXTUmlbk/OAReMK38lknYmCbKAXwZxeGJLjw42vHXHDwQ/8U4hISN0+C7V/UTigw
tK7XbxIQAFI5hYcp0ogV5lFI/pn/YcgyHIKBDmYU6M65LfkGbkyGy0WaQqxBZRI4od86KC2T1fDh
+SurOpia6+cuH0FGhIXgHV0PvG6zdZl0GZ6dMdoBvFjEVwfeLl8hkDiBbQ03r7NAGBhi8IJB9j4o
6LBQIZ19/4kMdgXcAkg8OfYvB31ZNt+N7sZl0sah0uHoPO2UCpUSPYNd3iW8/KIS/FPpbjsfcH05
O4hvpTG5ttPs/EKpiIZxLfLyMMm55pZeHSLQ4hgLQnIVyYXNagA022M8wRF4d0YoRJq9CQ4Dn9Mf
+xR+FMfSFnU38ARZdlEMOm9Brmp4pfrO8Lcc334pA+FNBRMOApbtggS5uJ346I9BgDx1fAWLhc1z
2NE0Cl0gh0QEpBqP3mlB7z7DUqAbJB6oieRxPg7uz2BY1ZUZz1AoPbtxHAAdDSJFr7bAdJ8SwAsp
tAEvZsfTOzO5/+9J6XL+sVNb3udmRNNqbrTh3n2igysXYaIxNpr2z9Gp70DF212/WUQ6oJvNBRCn
4gK997pKaM1lau3JEQgKKhPD7zwY0eTMavJRCYtWfZnQQhQfmDNuhs3zPqWOV+E6gZ1lMwRUcUiQ
5QdsUvgdvml8pGRb7lIuMA8zcMRGKks4adk1Cr2t/Sa2DLuOgPz/KZOCUNTXcNYYvqvVHiz0LO4b
pnEESN4OfpLKPWwUYIKHCJhD5I2wU/Mg1Z61WgxTvlQV1NJYiKvcxWzEdSD7YCEu9bmjRmzSafuI
fgNzP4VfMgO3DY/n0ibJJ4iq8iOS9TeFrUCSKVw6mcn8vR45l44fUhRv/LapOz5l4PlZvV1jEiwy
zBrFpMU5eyJiKGOSdgdjiAS7BHoWBxCTW/AThgEkMXFWfuV1+U2ungDXOnJJv3mdub5py6ZyOGq6
dsLwNwtUckX3vehCc3VI9OzSE50opBV4F5HFyjO9cBQBTNUwBJflD2qc3GRpvrlTqFdmpAEIZv5k
x5jDtph5XRTiXdWNjnoaYR6BycNxkDgbz3xGLLekPZXOt/HR2eFm+4OM9OWaT908pBMWrbPiELr1
VdWQ/c/3kf4zO/Ki39Mni8lxOSdQc75ajM7PPlKYYCOx3Rndul/mjm2yXxs8bYi8yrQtW+N+u5VF
2bRtg2qEnR1GwGMa8CxAX2Pfkd7yFRgFKnHsLpeA9q9XPOxFB1hNI+B1DCXbGITZx/QBxtpY5UnM
cd/IMa0tmXxb1hVRvPN+P5MRxhpibHKlZJ772X3Ed7udMLdjUb4+xDXAEba8UNgH1QM6nmZCJQZV
sgxHYx/JXk3rh/Fm+iC1xCiLibp1n/mk+7pWYNd7lwN9BAsA9/9a2tFjUlSydvijtA6zepNnBHDQ
/z5ky9jf1iXYEhvNOYUjsY5xTZbOacNAOmlozyrhjRDjjLPCD1pqL6jESkvpe47O3ZD/omKVJO37
qAqJNDlqwnWoVKbVd9F787RCuNWo8kUPLWIwkTukYQuV7LuUE4KDtJDFAPgXEUYbVfzeV0UpcdsH
de/uSzDuFA2kkvKwHE1u0Bn0HbU1iinl5AINA+3dBkGj9WQSL3IANu2UsPsGiWCN2UNuF/NCB8ZS
Z/vQWZFwg71K+LVTeQH+Oy8PkL4ro3WJ4/kKzBIX5iyKzMqwHMvUDU6eiPbxceC0SvJHimSZuwRh
JClktE3eTGs4HKROPGVsOH6z1RIlygZdWfjlaLNHsIh79/KzoH/BfQXn2JWxDJvZ7cNoK2WuYkhm
9DFNKxTD4rz3fBs8eKYmxevqH/i3jFO7Kgz119eF1rmrptBSzheVMjo8KFNmumwTVA+QiXNtV+hp
YJlO0Mv9Mgc4YJQFVhkOL/DVHEEhtULNytH2R3eKi5EbNJUmgX2T2Ii8B2kvYNpXCvRDl32rL0hU
jOOuv89X7OpfSfqbDoYGPTE+hQRNgKXsFQGg43yVPgHRnhN0aFUr74sYocnj2sugU2OTzL2y13OL
3PdErDDWsCqEspfI28dOZ/8FWKZwGPg8vmBPSjUiya1WaBBHZOsW0cuLZ3vwakWq5AhzbFmfio0Q
LNAJi9fJI9oKL/UIeIbWKE7rrXUsbDe1ZGhUdHZrHzYsAN7yAYtvkuj1o82uOlYBTq4bsfmI7DaP
XRiCgSr+3nHPNZPZRJj0pr6Ln/xabzgsx34rKqqSb8KF6XWNszEqcVWqYrV3gcIH/q2ACafxwvJ+
EGFGo4I/iWKdDONiMkS7Eu3ne0fs2xIAzq/JspGxPewaMig35bqH14qEo3hcrEODLdFK5JTEcwhJ
gFLUd+lyIggI811sBCQQsuCtNLzvLJHDnDq780dCDXk9w8zGTwBmk9yLfp6NeYQhGu+GWKhZxO+G
RSdg036G5Yz4Fb6Hw2+UGXA/OwdsN5J4v6J2r5O405td23w4sWLdyml10x4HUYomkQhATQpxCy0R
SnTx3WXtOm2pm1Qhwrax7DSblx1r4GMoUBR+BloFBkmE9hZAxko3yQC52CC4ZcjIwzq5v0KEItky
MhE8c71No8EO2o6xxzu9WT7wspaM1k24CMGzQ5QIzfxkXC1Qsm9JlaUzU21DEb1yox2xCoTjiNU2
lN1KgGKjrHOn7M3ivrBS5ufU75Nxf6ZS6C66QnYT4+jZgtYnQV8FS3W+aXxvWrfCA/+APY3omu9B
YYVaO54cDBTL3VJFx3IfkFtcufSpN9Hij6pug8586SbsT5R3SXth2Vf9CUt1TXtzvH3kXSQKoiny
rlALheGcgsVsBDSKf5epgH0/dWBvGVLXX3KkiHcFHH/utq4Y9HrDRX4QmX3XypUptaup3yMjdvgA
pqcvLMmgi33x0k/1Ct3yy/5Az+339e62fY7G4KbAsTR6qxI9sr14baltVb7VIzDHR4Jr7KNW30WL
E1TSBHyW0Osakg9CT3ti4XY7VeJi49ftD9YOIQ7evJk33b3YiRDlJwdqJo1PhbMXJw797/Gpywm5
V9nTSWBvFMcdb+e3yy11oRNk7Gr8wci4b3Bw7EOvDiN+6/9Ywi8AU0qBKDduEXW7r3ZfkSmch7bx
fzR9w0bsm5RcNRBzn4uVBAHEohxBv2lhaZbVREz+ox3ZKHCFmCp9SYmckeN71pZ/sXHQM+x5GXRi
k2v67DXBpnLj5GJcybFNZ8Y8t9xh0VZPUBZAEVYJ80StFXC5ZUBe3We3yISV+kUByVZ6+EUVb60S
U48pP/qnldxVVrhBStdbzQjCV3l0wNIi4A/CVj2fu2am6KmiOtf9RYI6QnMc4AbrBjGzKVKm+v0E
YTf5ZYfHr8g9igWx3e/1r5vmu+G3ssBbkfnD4J99dEuKgrQCxUFTB+5JaQeEqsALlggQ7nJ/vQBz
q5Ebwk9HRwvaLsZ1Hq7R9l04k7W1uvY9Cwf4kyY2ilAFTKgvCuvK4uVu5LcXnWu4wyb7/kaoHOU/
g0DuMs/xeFmukCH0v1i+OxHgBZAZ8hkgrz6jm+NXKmU9m44oVFT6XoibUefevOkYMuGFWXx/Nlh2
b4LLm0j+wmo8VJX8qOv5yFfj0SFfhAZUaWJHI1T8uNUKaq5BZI/g8Idpuq3BshdQ1iu4AF/oqkjk
bagcbLDcVwgpzaMRMhmo90k8XuR8ZRuJB/RiJW65siHQ9cnOGE5IzOZDWU4lynu64vxuR8QihbT0
uT/nzEl3+StbdXc8doUDOhowWohhdw+zUnd6cpAmTl68+YP6HXqsn+kRYzzrhZzoeBz7STIIcOQF
41F96YQ9ocA0LrRd5aK6MfYe4uHdaRz+/PSSfwCb6aHxEzqtWUzYfOlxrHc+V/fN41FJuuErNK/1
SCIgtyBnPsy58zVTrdy4W8vWvgc3MsoasaLykuX5iPidHl6eL72Pj+rPAPP+2ZRzoDLWr4o+M0ut
pC9afInJNc8JMrvgWGb7BfRcF12R2Q+Pr7u6TMGZYdcngIOCAZNO8eGSWQNo3ziLvVNu7e7HEbCW
+sQ9aYFm25W+oVY5Xals0bHH2mvA8o+F3kmq5uf4H1JaPURbrjOoWYV02sJgL/vBzNlc3NjgSVjm
CqkuZEkZeGOt+r4dhP51Q/5sfNfCxdb/r/GZjMaxqUO2Op+8V40+DCBt7szMPrBC9SCcj5u5/OA4
aNoUWKJZnEHl9qM2SiNJ0V4J43n2DxokePd581JMDWtTfP3KTXwKgDIk5lHoXgGa+3YCrZRdBmVp
ZWQPWo17CaSG2Br1Kp0hRBX5i34cY/yXJOjSeytkEKyFIlxF0d3LsIyhfAGl3NsAvb0fje9ZhbR5
65acZ9M/Z3tEtusw1atkuqOphB/EY8U4/K7xxIn1E2HX+H5xQ3ZO+7FAwxEt96bsdDu1FpsjgD/K
NMnX22NXXLT6XohecJzwHiKznk+sH6bcl8LAfKBMRONHLJg5JllkDHOlOrr8E8cdRv2JQzEYmFBj
nm+Hj7k6pYtWFsAFUmCnjnigwfp3mr87Jt7mzFuMAbURL8ykXPdVYVHsyF0vZ29J2Zsa9A91gj44
SMbhG0YxbUx3w1IhZZb3jhgTKgm2SJXROEslRrLAP12FQdZBzY9ghVXykgW7qH2W0s/0DJ3zjMi3
OuLdN8uz1zv/hM0N7orbv4pJJ89+swSfiNyoppi2UxTzL5boJsDHZUXvO0X4Mt58LtEv2YgFfsyw
lO//JK3R9kyA+4jwcfZPVpq0//lR5u38DGNrQzmYUYEm3DVtPXNYyc/g4EogKqutAKgUrw4r9kur
B7Ag/NzJUcnixGFFVlDPzyVPK19TLZdOL/C8I27VUJImZdwb2SDXUgG8ArbQ0C1B9a3JM2UIF6Px
EloE5Eveob2eUzWQa6KQxTud/z2Hn7ZKVf0fnNHqCo8P678d9+4VPXMcERPsEeSc6q9HBK2S/Bpu
G2BaWIorGVWQIGEurFcmZWiqwHqOwIcEe4YrFJrv2Soi5vF0RToIQdqqUHaithI9Dez/RrCCTsjh
YA24H/X95urnt3PIFmAsMiHtb0nSgRPRTU5xO5BcQzSkMkriMY/WIcD3r6FYWZ4gIaYKj1Rs3lV1
sXLxA6W1UaXxV/tAJAH+zcZHswHffOKLttNeDdrcPIyrs3IOD7m0zAhRtIQjaX6OjnFNStYrPW/z
xXWWc+V1g2Wn67iRntbaqF0QBGt8ZEw/+Cc1d2JeUKWTQOu2iodETS2sw8qHsonta2z65cnma0ZZ
8xWOhkrLpP5VTgBZ07lDmsAOoos38YK7RyFiLZim+ZhRD+FiOyE7kuCVHc+eMYzruCspHqZenKAW
VSoXY4/0nD9Js0fQzZ4+C6NLcNW1BYTng509c0wm+PqU3fs5Syw/iBIOcwFfG/niaxxa2/fU1VBW
1hGWIma4avQtiid4mzLXLWrBZw82Eq8A7nux2REJTErgDVrvud7Rx84wLGZEIdiegWgRhQG82NCJ
j2wKbYDp/BgniKzKZLWFn0OJ5lJbQp9BHGLnbhaRC4BnBFxBP3yf6EzM+SSOQEjEWL2f1juPuKC3
Q4sTc4NsGo8lyc3iIfo2T9w4j+e0xKXO+20WU/+yi4ZrhD3AHdlGT1KW5hcLBT9uw6XTN3Htvsv8
fApSCyjiXiN7442A0hk2YPdmpqldIU0mGwKwdFpHeEtHcnY7rGoZh9xoOty5Kiu/9vsRJh1sTKNT
fA59VaKn9G1qLlK9iLlCzdcEp2VzErTF8g3kKwtyiCf/nrqaF97efpYK5sEYhsf4WXCypWoez+dh
OOx/5NpNr9upKsxymp/3K3vAFQudLGOfha94b80a0vABbAcqwi6qw6p96Ozf69Cr6apjPfsIE7x0
8P+EIZekEXHHDhTQ2MFvifP7MJnhFVqzjtjbWCAyb0XNFp+vMC3asLLN4h3uq5J1PrtUCaiOXQX5
a2mUDTgXMjgRCajT3HhJiXAbLCtLS4Gdtdm0yOqSMJp02iL2dWIQajMCHRL+a2Kgd2rfXqpUU/lD
FujuGQHJFv/v1kigLxdm6yrqFInbvr0hBl0qV10damlEXKN5G4eh4n8M9bxESEQzxznlH1UxaBaE
3cMbWJMLOQppEa16keIpCvtvsWR2yPObjf1Mgc9rPO2TjLH7eF1Bk28Ex5dPNryTbCvp9qiHoZ5D
GG0pY7WIxReyAH/xFp2g8A+vszP8QmzSr86KClpAGatolrpElBKAGcRI7lt7fbZV+0TJd8Nx/wzL
89sWYEj7ulC4RepBJJaNJoKP2QDS/VocalL+Ev7PjSKi0F4I9EdZgEfKn5jLTvp0CGRCEQmSSXJi
Wr69h8EfIMRy7PiPhX5HmEFE87CEuz2XOolZuM+gj01NJi0ob1VW4KTGhRgxEXecw1s2nvOnUI7c
QYxVdIh5WC+/qtx3Szej/2doR+L7toaFtGJv+EyNc+MPBwFkbf7up8bshQMoYpPhex51xV3Lb2qo
owb4uGYE6zCM+Ce5dl+7SONnRBWfVosQujSZAbiLPvzoWai1WNfuH5ez8F0GzmKT6y3MPUZjIWxw
atdULukvXQGABIrek/WdbwHPN0HNlJfn1Ms3V+GEs7DqVQ3K5lrjU4uC/Q+PnW2LUFatItYHgPXz
5qBxccP8ivkUC7aVy9EqS1KQIBgKmsE9HTIWVHBWNVbFDrMTJ6bS770GvvdUM9yFvgzcOEilC6Rx
X/OUoCGARxU31g8M6r16fSA5iqNDidlYcGPE96RRJESAE1OyCZG0QeXQ3MBb9oIfOaWIlDgbUA3b
ZceT/OpDdVB+QxeEfa1vpDT0/IIQIlFL3ETSwUV9SJPpRhj7aRNnmWdnDsKltdQ9oppJdub406XU
+sBjGIOS8Emtw65cu1qiTVuPhyY9yntb867f4wndS1jWi2PH59EZ/Qw+ujofj33Mi9ruf2wMW/fE
KL0fjxcvVEmTquJBKMJ+KAY4vtYEidFtHJTKgPOzim2QKmTZ7Fe+YPnIDDNx5C9r9xg7btr6IzG+
+bdjdIjm71aVmbimbJ/OsNyLqajCtGI7djnHx5gXjRiApt0Af1PSxPoHij6XWZejOGe/KyE0U/80
j5IHV842tLanm4/cPFOGCHGBMzOHWwNqroP+UsVuqBnKxsw/xdN98JE5VnvnLHIkIkKfFWq8HgoJ
SFnQbidS0MzXlUDK9TmcZYR/GV6RLntV1k5TOqT0VzOHw0HdIpBkCMnwBME3JVEX57NN785dHoG3
KgvDkLehacyxK/qD0TEGyQeCOQOCiUaJm799QbJo9BQtJmGJwgb+YhjU6ANZNiusSS13Ht71ylHB
Ii1DRnAVq8J14EDBnUOIo3mkChpdNrn24sJuKiv0iwXX5dF+kvCuaBGDWIrcr8laLMkO3lqw2Bz6
+1PmKH9EDru5CXSdMnTo2+YCc7aesejH0qgl8D8ghl2jJ3WTwCxmjFq//lpjE6kcnbHOvbtWHdIE
BAiuOS+g/B0enH+xac6kza3X0qMpWhsuJT17iNWIaEe1EKR6Y3zoxKoKBajp1T24Jh2SONBfP5Oo
9Hb96VaqKqXfyX2Gw7HbTJKetyOkI9nIMEmHSpoMEbq4XFOfEOg5+FfrljW6l7ur3YU92O8Xy0SB
z8dSHKUXgwOPuFxY8kptrBKlRetHq/0jp7+8eUO17dJnyL06tofCA8LepqR1ru3ZdiUDj7vZZHsD
tL/i+alEUtEG2r8TbYo1hLw0NWtHgH2AnkOj1OHJYRfXE8/VE0vbgPcyatD+T8jjOjFurC1MPisg
NMOjxy6WMDnsSf3OuqKpz87TK++1SCRK1zoYdXi2G/JdDmDSY+a77kV0JeDtzdWfsazYZQg8bbBh
654yvKloVXXjKvpTzJX1eXFkBPhAXHEBGC4IF4+wgdQeTAWRB8cyYzvQYFTaAQGRsyjPK8T7LF1Z
WUQwBWTvmcBbjXNNIVMCKssqGDectn/NZSn/tL0n84uEakQbCSYP1cZ6yw26zeNT7A4+8gWbNf6A
LDLSMCncUbuLEDYTEod4KDMWa/iqD8nic7/evi092g/lzdWKE9WWG7WxkJs+Era9jdpOv4m+ykkx
xKXO5xw3wJo11ykTn2oC37EvxUbtWitin6RYLI0F5O6WBSTgBaHgfmuuLTg9k5EQCkf+YYd0A01b
hwc6R+oAtK4+TuLOR6nfzbdgE/HnnAuusBWj9eL+ulKS/VOn8dsu1RLqClwxK83JEQrwwD/XDK5Q
bqtiFlKImFztOK98UCuM9H7eSfSaoI9PxYsRUPEoiVINGAp4Y9gef2I3fRWSQIrAPY2NgNfpafKN
QP9VCyhUw9kOuoeJhu69VcwhkseN8el5sxgeanKkiwbNRUkL9yH8pkwBuzIv/kOQQMLID8Xmb1wf
iMnP/8XXLsH04CxvhNb/OZzWZnW2Av8cDDQ2OYFqvTEx4bOPA7X6GVAPSoez/ucWJhnlnm/e47Oz
gLisnEGKu0qKFxJmR061mNn/8zRtRwEpveGPuFQUNUN7D08B7mne3l39SXhwD/HQFqGmG7MwSbKq
RY3mkqMyzHr34lNLPpnh1U9LaSWRjPMTXouDWWpQ+xHaGU2sUY7UHCVIIxh7hcGpyKBs9W+V165y
k32OPJLBJacxhQnHIuUp3nq367uCKNXJHWGl2L3uUyCCCOxbre6nvf34saHhclmWtdxpsTTnDu29
Mhr22v1HcO+SS0VmIepH6CCIsyfx5LyPPXfoGgqgWxMTmw/l0dnK9S1gzficQGV7TWBnaere7gZl
j/qhyVS9SFyPymL58sOq3aGiDwVmQmso0V0U/KIsLxkNXUvsraN1YbFwKT95zOaQgd4/Syl7NW87
ygD8ufAxydGNIeS+LWu/sqbaTP4Je+Rd6oE4IxjSW6lAIAD0fgyzWWtuKj9Wf8Nkx3VtHy2IHGIr
QeIvdhLDe7tyTSV+1qZbxqX+eVU9ec+Vy2Ec5fV2sAssH1KDBYphDtBm56/Ey9BGSYFsQcBrGEw3
RuECRdVvgIP2MKW0TZHOQxata6jv6Um71QJYvWNAcM2Ybh8G5uSiYO+pAv2GXIEr9J568EB5oCzC
g7D25HBzMvk4RKngCngddCLj7pGi6f77OpY3KR5s5QwaRD8AD7lWc9PsrstxMM1/JeBYGGkB7Gg4
fELou7GjtrvL1NxcTku2g8ddvH4OorNeAmzZNegi0vTlXBXe19+NN5VtBIU83mXK9uwstkPDTz7z
T6YPYftFWlxsZ8M4BOdNorJ0FigapRyzz9Kz8TIPWdJuemeMbBJZibLYy/kzVf/cTFJmsbLm8aaK
EQ3ASszawkW8STh+UilGhE71bK1HVoEH+wliWN/wt5OUsTEFFEtlc0yAjh9ZUky/k14tW2WX23MJ
xfs26ny2HbTjRkDOBQh2W5G2Hd+ArPV3w5u0IFKyDxzDKpIuG+57wdx7vIS4trMQox9grcqv6LP2
GXxfAsDr0UeISV3wGzWeH2BuGpk8BMuFxanLeFstJaYw1yPBwvoJJPNtlJJqBAtw0H7DQzoHsv5Q
2G36kj8BvTe2W8pGYgQ66W27JaVDc5kh45ohUMgz6Mp6sgVszXP970BZflsuFeoykGTOUdysqqd7
fHrx36xwlK9jozBI3adQcXQpFGA76WSIzq1Sl09N1EDaqzuFJfC17hAYqZmixat4XHPH+SH4Uf2w
lLfECanDJnlvKKcVJGmcmKtE8pMA4kJTVpQXFb1VrsX4WmSl3t+DpCy5uFTEuQP4fnp9DCuYN8Vr
FYesebaXy1T0bII/MqTA+IZBq4+9T3Pf/4A3BeAWSo5OVqX8AI2tNYTnOd06rR8Qkf0GXsAfCXsj
TiQL95OSYC3q6TUmyxIYzWuZXvZuxBRyTOsruBBA3i737wFZyaC6aGTMevwHa/AJgWDev+G/NGbb
R53ATq4oRhQITRjBnKzjHWzKCTJEFA7xSTeY1Rn3QQhCalgnuu+bR3PlMu9+clFIFdhODELHlztV
1Y5zBe7eUhkrL7CI+jwAC+6BdlRMiFhJDA2FkEaG8PJzBDKT0apXyBJRUHGbpWk8qTPQOgQoXgqF
l+E9x/kcoPML8f/9wyRNvW5q3aWVAoyD2K5OHIzzMZ07CM9Efw+VJ55jBd1f5IOk6LbMGNSEx3em
D/PLnxKUYDHGMIewhqw68HY8+gBATnIXAryuLrli84sn9lLgkH2wbAuxu142n0yMkunuTWw22y33
D01bkANKM4VsVcSAYYtzaxJ3zjVizNAFqSAesz+Ko+U8AKKRjd5g8xP7PExRbYAm+M4IYBHU281K
Li6Qp8o1aeX2px8G6x8KVkwvV2cIuJ/O4OmTyR2DyeV4BYnqkPQS8iXc0eXXDUOLSjWt5vuEkpVf
2lIvaSvEIY5TAhbMPu1/8aYzPBNr6qxkR2VXQBrX9ljCxMIf+NFNq6q6QxeSTnbx0++AEv0C8xgx
tSIhh+eMFi890B/8oyr/Wj1uL772l1/PkVEuOufUPB3bsSdKsvnz1CQcj3JlSLV/McZzx5Dcfnhn
O5e4qy/+5UwbRwHC/VKWk1zqnWu0xU12d6L14DknDZYncmwKy/E5r2jG4jEvGNZqb5F5EOig1VaQ
JKOYAFcreJYAMqQWRDI67812DiyOL6oMqP4XWn+ZK9Jw+4rUxI0JwmYuWKPq2gMJFiFdk3qSVfrv
8yqWH16ArEV2KH8GVsNPjlbF9otUVITJG8HPGe3h5yuW64QAxPwFq5rn8nNCxqI9sZWabfWrr0GP
3/zEMr1ynXXj3BdrJpK3OY24gaB83b4iybwc9QU+OarqK3LqQ2gspRSVo8ft5sjMoGrElTzfR13U
SWSCLqhP/+VDGALdTDjqe4pjlJDcdem6VGdvsTlPJXDxHJty+1XrL22sxUW8bVp9X9nKL1ed7Qzj
hxH10x7F/PJ5z89QEDGmNslxDoIrG1OEX4s9yyp2WCcJS3TKCxfUcs3aAOmh/426zJOZTP9R9Tbt
vgKgfr4j0LAoAHA1TVvLglouY+NdwehAUdroaKq+62IplKu5oTIZAHsMC0+373gWx9w2ezt4P3YK
dGvCvF+W49g4lqg9t0NwbnKj8ozpXo4Ymq8IJcaEGBx1Zye0p6wTZG05jHKuMrlz0UiDWYc8Domh
qcOj3Rn/CLzxSdgQnaOASyzV67GU1Xr/t3dqCgmcGN3yhRbsBbYROD2Nz3vlUtQYS/StEh6bzdvC
r4U1LmXeMJVLtcddhJRghMwKK5dtYGZhGzZ+I+oamgYoZbk70lrfgZDE+s8digqgJk7d8+7mY700
+BAlgEX17gaNrlswmMdBtzjOc76AYJEQua0NOucITDfa+FRyCoO/LfMzHcOO/tdEIsZlwPedwTbh
yp9AZOoU22ucGdOa0QMtehs/9i8RcuyItW9pvLdFNFowSu4n+oL7bzGA0pxDz8h8Ir9d8u4PL/V4
j+FdINTNR7wY3dZ/8dsQK8AI0AJvLrH2KvTJ5iWu+4jZm0fDhl5Qmc30cwQlPMvEd8SqnTsC5CCY
gIUu5cRbHbMriIolXIu76aMKw3eVnHVJO4NTxF216FcGpwK5AclZqzCGWoHIrgbc9dEXVzL7Q9pB
BD8pUuNPY0U6R8CKBL6f1EcEpwkum4oFCb6uNfAvhhKGtJEjRe/TTfoU6x4lewMtkZ1IBwnGyGf9
pVcnT0eRc9j8vNZ8y5IUA4uy6iI+5Xw5llfG/jeZgjRYIwJISLXhXZe93uEG4zmOj+pbNnjie0s9
u/EtMs6Kzc6c7hNnwUq6ks/EWjDvshTudQNd4jN1Dd/FHGLZxfvQQ5tbijCoZTSzObejt15CygUx
WNOOsVpf6/G81PMQLl8uf5WcJWy73C9lfiXYuPxyD3m0she+3PcC7j5d5NPFcH38KOm2wSg4P3jV
3WSVfvTYAyJfNfBcdXSJL+m3h4FK8irNl2Iv+Yd8JVj0fHzI0Zr9slfT9ZIN8pqET7hBcTU+VHwb
mSabnpc6ozhpoIk+Q/lDIg9gdW0RQ3yAKJk5qcB7bdjilsXCOX6c9vwrjzn+9Z9j3x8CqHYTfCQZ
3JWwURsl/zdeeMa6AAIBUIbRRt+VR9bgjPIA/4lO5jiRDcdMZOiVn3euJEttqt+wjfoW6Dht+8z2
wMfCCeaNj482Iy1nXFpzfmn5/8hhoZrzzfjAI3sHGHTrM+cLkPnFqJUZLkk2eQqPPF3vlpEVsmi0
rVnvoj1sphplHVz0XiNjHlWhYeptLVVYFODoAKpIPeLE1/dnHfGKvy/a+oaDRyj6uc8kwECYcNnA
CAXic3l1yvx/2wo7FUEEQFhh7DLVxhOM18IkHOF3rlr1JtMhHDQfFx7u8nH/Lp5gTVRjV6TX9rxm
XOquc3qa2xDYNZKFQbXutt2qN17TTXhAR6grzgaiX3EW/5pA0n9JpCv/Sfd2MGFDZcAv6v0TDcOA
P/guRXYUwRye19wl1Xox9w1PLpcTvDo1G9XAAYQOnjoaQlp1Wt2thdbQIJwG7JilMhzz3MiD1vqn
Lmh95r766CXn1lTDdTPbBSczwUjJDOyXk78QPkc7tKh2GqKRG01SnSNcaBBgpnKvnCWNE4f7+JxV
k+fJxvwVkW1hnB/zUi/pPq7uFeCNKZOIe6UIbPl0fDoJ/Ux/6Z2//W+g6MndYNwMraTdDisEpzBZ
wf3ITBzJrmRMZylGn+fcUfl+6UHDDzQw7Y93yDGpJjYMry30zNCWZpGHVcYsZJrUblO0Ix36RIXK
cKTOH1XzveKik+lAUhsd0iDG9pinlZRpGxKPM35vKxmCiwVFMVHgXsHCQpm1Wn7bu+bfL3PQ8Nmh
SywTvgQWsy1EqP90jhYr9amo4TgUI8y1qcogY0QfVeBnuCfzCTb4XpSrXv0cNN+sBi6raL3QTxQH
Aq0nh+sccLYg1vTVhvHjOZG0/Ep+XFBsB6FI1EXrnuMquEhkhlVUVn7vBQFsmD80OoxOOkZR9wuU
O0SbDv86NtgS6tdcJF26FNr507ePwqpEiZOmHT3RBmu+MfGGqCaFAxzgzfzDD7/KiPP9d3maiJ7Z
Z7VY/JmpIPN0YiZJOo7P5gqOvIrasB03pdNIofZ3W33CAgyF035Xzkd54gTmqfJfTAUBHXf8sDSs
jKNijLJ5PA3da6WP/EomzsowW1PF09qN1Orax61OPF0QxM4bE/YPZ9/aI7wW74BfYzMdki86wsBZ
e2BpGdF/o1GfjYzXReDi6V6NtRJM6Pd078sM6x1WM/79sor80/InoPM0gDRigetFnowIie9roHrj
IGfwxYp7wCbG2B0QZFOrkc1Kum8gb3Htf5YfdjEBlBKa+LHbECVd494moRMyBebNAQr4gU7GpODp
ibJiG7DMwPLpQnBTUG71JTn86tE32aU+oZI3WDnyWjfITjZuCIUGgnBmZzmIuBLTeClelP2eWcFo
PN81PoYMJYN3RGgEfM6ij9ODCo+/IVjYXKBPhnnbF6EurIl83F3VWO24ggz+5YmYJlk+NFJ/UzmA
lF3mkWNwuSH1HPilkO/z1TlLrfKGvo139RB3aymbKu+wMiebe7VG5eelF33itfCGigWLfvOS2Sk6
o8XKAEutIPPIVw7NzJ033bc618yQgwpA5U6tGFk5ODVR/V1SOoaRcHGWtcy4qaoITfOx1Oq3m4VP
kMdtm33afWMDRixEuinW+h0IPajvbb4y2mXQY0ADmTM2WwnWsZ0lT1SWKV0nxomwxMbossESDGJG
giIbNIfIMOzAgRSoVteWMhzc136tB5vm3FQq7uq2z9x7bGKv7SB3CEgtSsMb4dZEc8APvdHDb60P
1ORhJrLAMLgQcDVSHuybtief6Cw68AgpRwQcvEGqEVaTqUygnal237/NjHsSvgBjPhR5P14JuehC
IZka+qAZAkAyK49zG/OltTc4vhtV/lGcsSYW8jf/EDN2xYVz5uYGnV2spvR7pI7q3PCL2AknXWws
AZDiacN7Hql5H5ScR+EzDi9NfWoYHfS5oVw6BBJ5G3BjY/9XpK4tW/H8fJE32dA+NrqSxKGT69dc
a2TlxYx6JpzuvR2Ah5Wd30qxQMzVOgwK1nWA7WV7CRa7kRl8QLIAoto6NMFvwDBAGWktT5AQ46b4
jp1HxA4b8K9cOw5gosjuBo+yx+gmaaFMcezfg0oznXwEijQFZhuy7g4NhCg9HNIedfFh8Wt//EXA
abeO7cuMMOYHcbzBB0HeZRCZRK7gKK9jbGivut/6Gix1jfB3/FXOK4G2bkBBihCkf1Oezahrmr7y
mddGR76lq/LpdgCqZZTBjV3ohKSw721nWjjYNCZnyD754E2/VdyyIogQEZMOQ0tSSlaEEbH0G9pj
Hs+uueQFcbD0rluxrGyYZTmJfVlWnVqEmaWmDgQ5h8dDFod0dsv3pJfDcW8SCcf0RtOFNg5On17A
6INWK3igT4wXwNzApbpB+RD0Yhob8O4eVu9hkhXkh4c0BiUdEKza7FMkH27il7Jye43pu1198tIr
oDN9jXtHXpO+e798sa9yQA03FKF503rWRKs3w5bOGA9M5r0y1N4BaR356RClff/Bu6lRsuFzi2ci
ML6gw7AyF77zYxzzQDg1zd0XscxmptEWy8dYK5ZZYEnR8VWIvwjNSEm6jQgVmIc5bD+jLDDvRMV5
m1hwFLBNJY4vr+qsD2TWVp/VZkuZT/XMGYlx0JrAV+bPuDLKgDvhKjr3T3goS3eUd+Zbbl7uPquZ
/pRzWNnZXOfWcJQ/UYaoUQV9AHRHYnqdmNru/Wl4xHRF6UXDTur2gke0mvTMU0IY5Ap4DFP63A5B
X5Bs/wVuqW0E+sIOQu0ilWpL/kCarmeF0wrkmsPAd6IiM2cC9J5TY3OnvcZne3S04C3nCH1CH9FV
2XjPcIIvqtiF2lsLtKyEjKE96LS4Bu0lE3Bxm5DzmPtljdtmcE5fkZV+jt7EhrwXsmMbEbmmQlK4
OX/IzCpTjxFkNmnGJ/ofR5qpzpi5ZOacLQSa+50M0Q1dSTwrJI9fxAomuLWXISLrDWeH2x9xecbd
CJ+6pHGn9LJMI95eGoax4BeJscOuiIXHM4Xaf640G0+VjbaFitk66bAv5cTLdhDYfQxumszU/lWM
elsrwx/M6T00hz+SI2yuU2Ycr6uY4dGje1OgksiD9tauHjVvW1jO4u7NK8Go0x2SCInLYEEyWgnX
Gp2kH8HyssxLMXWeUFKlfOI72J3UiAQyX7fjicmgxy3QmS+mfqE57niU6aySv6Z+cu5fTnJkLx2c
6R0WP/YMEoPgf+tLNiCf4pZEBDbCAmc5czrAxO+NVGkMFDf1PDZGgn7UErQQKWoMlqhw3MH6motl
UBeXxZ3IEGU8PoKxMpYjpU8dHvQlN/f6AewRX50LY1CuE0g4F9Tua0R3gT8HybEAJTWJMNn/AlHD
YC2I/Fj1dbjObcNiifHd7phA367PPlMWMUZv+lzH6ta/ZwniLVfVb3hepqq9LNlx0XtW41pnenTM
TMTtXu8XDIaPfc0gtsOIr0xqMNkTpKvDoB/COxCPJAZNQGEC4ml26+BaLF4Ddun+ETXik7rCZ/qL
4haWfslr1TxPRT3Wfb1NP770u7/EL/JvfdgZKeTBVaTpyYfrxqWz+eUvUJx5n/Co2ako9gSmSQMA
WmHBCFofNeT9CPU6+rh+XwZ4OIpu0XraMC/ZWP5St9btb6xpVcEAcl5dCesbRSFQp5FmKre40O0G
OJQMSp9F8/OEDz8ooZPWrCjQiMKhrigDhNw/esBpfZrzuskiNhruRRcwpuh/s6SfDFfPcoIG16fF
V/Fx2sFmEUzBITzHc+4riy7rrLLTEer7n/Egjnrf7wCct0vnJZWcZpU7xUAv3KzG5CqyJRmntDGD
I0dGegMmoO0lWbt00/nUIbwqtjfKACCpfAPU9uwAU7Sp9FGF/brMynK0OzFOUv49oyHJi8ZOoF15
qW3LYApgYSaiNoJjPBTyYt41PRR0OB0VFLYYVDo1A/bvhYq2Un8hpJtnUP9XHIPelaTtCX8OBkVD
xSDDQr88WAwGfLWAa1E4UZHI+0Zj+Zu2sF4xouycWKTla10IoZwfBQBJ021edH3eUwum/IfzeyRx
y1co0q4C8l4/Lvn8Y4OTEyng6JOdCI728SBVFx6hBwfI3dkAKSY8qGrNgRULCH0NKFnlZgjimnP6
QLqUtmZiyD46HtR47nnSev1Y1I8rh6rLJjoLQa7R2rTiaqKsi+39BEsZgtSg/yRC0b14HyE17NTM
cjyHJSsB+h/9avT45HndJhXGkU5pKtq4rAY/v3sM/TuRM6mZkQtkTzQ14GdUem4X6rcIfZBQuMHT
ypTU1D47mWRX2tzcyt+W42nrhLEshhPtB6hV4yNz2KwBGOOcwIUTPzEM2am/lUFI2FDs40y+aJb/
UDQgttOJ02bKuwu8qPgIBhaWXDXCG1oRViP6F4mmM8/Cmht2NangO0v/TLxCFAr7h/9ONMIm3crR
cCxYyMIT0pvZkSs+JpEzzuvObUx4tf+OGiw8cnH9f5CH3vAMwi3l/+2mju+V0cCoRFeGGzQA/WqF
QCQAFpzH/6mm1izzLGayiqXMrPFxNg6CzVb//mUHw7kmS0/yEjjNT8ADEaNTrimcbxHCoF8gOPJG
1upAs9k9FWfAn8FRQZzdtMU54QV/qVaFVxGFIzutbwI8q9bzstpNKoHoOgByTBa6asTIQ/iugLrA
BXN6bfDnd6k/zPtADVdiUuW9DPByAIpQHMMwEQ3zUqGV+sir3dkBdTRPjjeH4XfQiVGKFvreViB6
o5T8G6uDScGvSjUaU8tspdx8Fmm4EAFxK/xt2E1+TVfLffC0uVy2vBwV5TrRlEdzfJy5s0AtlE4y
VtcQF8xIFG30zCEaV+DGcDRABMzr7LZE1+dpgBDk5SUCIKzsv+7izy1DAza/OVyeUudt9oBP0Kj3
VW65M7BVqyDCm9rRuOikyaak9IQi4P8stsO9E+8mxHNt8HEI872XCM73oSC3fSETGoHkIgCAuCae
Ia9Qsx4XvkOXt8JGaj9BEQZSxUSIsKUGV73BZr1rWODrMtSEOAY29ohtefbV/8lhKdK2xYxzRu+m
slLBlhDWto1VmBWRgV9k2854I/1Mo/tCofoR8yNM3YzT11dqxx72OxjNtP/spQ3Rth75EP1nTGrR
EYcRUcoSJBg2hzewQSeQPGFUqEl0fmzJCwz+5D5kzVPrklr/sGaGgs/857FFt0L0qBm7+Pm56rrB
DCHEGItbslAGLZSaYhy8ufiAHHqfOPRKon42WlVxixNIJms8qbdLKR5QO5H5tdBmDRIBybfJU+Zb
7sVtb5wYi9bnk4cdcGpGgcxkMRkeN4Yaz5lf3bIKk9fPnZIUkNRBQdCYdKsyjGNaB95a79UTuFO4
hrxwVPfOgVboLcvzJF/pHwcYkim3o7mkEavJZe3Olp8kHMuLbAO4No0+Ql0ET1gN0psNiZjr2vM1
qmSIzR6pUSx7erEhL1NO7I93Qy8i70+SpnfsSVpE3cJiOg/E3S+3dglzBw+h9hYoShotsy3gVemX
0XwKOsjeTnhpGcRlt0puco2cyx/N3lE18ql9f43Jo2Xm6jyYjWSx47epx/pZ3uciRsOlqUiu+31W
2ani837aSjbJaOAx+SFRS0Jcl+V81LRyAofpLDsEHUEImVtqhViSztwPuPAxVDQw6tpdOA+s5GhV
xoMZYbA9ca8p58NnfTCWTEdfLF2s94ur/0W2ynwj2xCF5msg4KT956zyOqqrgRtiENeada2YOudQ
mrd+O+4dkY/6LvVb5g9IN09XFSAOlM6Jc1nS0CIhwWRwZlyFngp0D+Xx2oNWbzvhJ5Mc2IOPbMbu
dnzYy4bKgqx1HTqcpkNhuV1NTSC+LEOts0oKPmlagYc5i/TDHp/Uijn1NxHyw7hkpLpKgE/UNTqc
XMkIzV42e4wKFLXWT7+7miLlDgl0KuE6Z4+vTZteEahwOIOG3kcjP5y7+2ABsc9C7x2y7AoJB8SZ
7PmlS8Yc7NIkL+yXXXTL3VOxkaoDjqBVf4TCYgioNcOmnmNdm+G6DOQO1pTIqkmGNZyRgcoFBm4L
VVi2zHq1pjHomer9ALu72xY70yYbbZ8aGiqRMQjrlu759TUmcy59FwlFF+7+shUW2GVBDiXHk5f/
rQkxben7X7RBb4wYmaIHEzfrFwCh01ro0botJZOgiXClx23bduXWzH6A2TiWNayYBYtHaHtRo0Od
yzkxWh3L7bgqx8nV6BmGpIV9dmLG/tpyo87coehE1slkUdTABAMHKVci3VytFf3dUKTV63lFmSDo
HUJBeGDmAb43ra9/pLUbFPQOX93L/OhtqR6gRM6J1iwxjy6BoHNlWx3Fzgog4QfkQ68Mictvacfd
V4vcDm69wk9jntM12hkfmGYN4MbSqUelEsj+VNa/wT9drn4Dz2hh4HvBzOCl1Vdy6jM023l5QjGa
apAFt+B6zDzlN7T5klRGstQh+pej7QcG0lazSRtkcVjpxuSt2ES422DqDCwPY4VhqfyQ6gQ2LrJT
Qx9eSO1ePFQeFUbxjUkpWPR+nXiyBfbEnk4ra92AdM4zqR8am+dh8aDhBmVS+INFAgb9YJlEIZLf
/Q6hbLs8p6UYpNQPw8v0PGjhSxiEVDncBmrKN+suLwcCwTclaJJ0mFJTBL+cuMEQIL4TQ1b7jB1f
1Pg6/egzyTccYR/2kyK2xLRRAc7O3O7GX3mS3zfIoJAUoIPdwt7hdpNbj70c6PnSdKKnNp0lyXrC
lNMcsNbLZP3ZwW4vDCSkiM9H8ZZ2szZpJ2sGkROKUuQ5eNgmSTHaW9MNeoOLQnI+pZtetYHQz819
ehcScJCEIxM260WHu6N0WsRuVpoPpWj1gYs8PLgbJrYLhwTz167QrZgGzv9WmpZez7ydeNU8RryQ
WnKZj7uLjLxSxo8vR3Z5CXECymKdv1CEoktvYqZqo6rA7tbxj9oN+KEPrS6WPte0vDZNBdV9K+cO
UfbNFZIKU3fULsJP+LrskpxNlktHhH4NOObnNbf03X4tpCOdCqfaxPi3VA9ZRdV7yND4WYsx1hs6
2rXk9/5oGRgmHMyrpcBAm8KMLVlaR6GEMsbNJzMfky2+QJNcTmOZahOGhLI3SZtkZVQ+IGSRtIR4
mTC3bU7pgyxL6uqnXGn1aVSoUc+s+d37sVpen8JiW5xcDVEJbYGyJhzQgwh+Gkb7ny342S6sq925
11OzGhn7GwWFQTVRNPHCRlcxzNvPc6RZ9onX0xDSu5tfqimz9+hql+/vw+SlzRM7kxGyJ4mZSd02
0MguwzyZOtcOAALMoQsGLicF1VZuU7UpcQ2Ad6SebYe30S3gnHT1H/Hbr/1Rmgu8LoHxYTNlFJvu
dQOuTLp6id/jHkRqtukwcxDyLnqy3cRsLluqcN6OdoiTnJsJS1PfGzaMnTTTOCjMNRHeHK3LZ71F
j3yW2cwXuXTFZHWYAAV0Ji633EF2Sd8ZcUUEZJcKmrO7sxLLrJ+yqEWfftuZn7Fx5D18asqYHP88
6XeICLNCr1Y8ekltStRTofWcxksgR/4tc0B8DK45uVxRYL0wl0i3SrYFWljP32br0/6GP+GRNi6Q
lXBMy1uCOnqiqdrjGG8rxSUB4zIE9uReCBPTnBsOrRiAl+bzLrloHo+Z01EChDKXTU8SNgoAwVXP
QIV/bpx6nLc/0hms5t76Pn0UQgXc1d/d99+b93q08DsOk2hd9173pmorFea9uf2jSfHaVoKDZYNn
Bcm6m5bXkU97Szg0dtgoFMw/g5joZFFewHm0edDNEdDxzfcLXZIAt6srh7UpAtgV2B/K9NI5ewjW
Ne3Yhb/7Kecy8pAEg7fH/QsmxEzq4cNGt88tgbooyDvgXEmatYNhFbLNWoVlzIirPRoGd1B0Meju
T//DXGxUmQBAj8JfK8R8iwWQPdTD4HoL7o3SEmW4qkK6PqW4D0KhtIcspvx33V4JBSwD3xytp3k7
+Bcjx/TvsTTttosixpoqLxBf3tDV3UhxGQyIAGzxFmVi/lugXFtCLODtNHCD7mctaOvxuf05b8dE
ykwYb1gtrhuiGdPZFoRuztSMx0eOdU30okMoLlTR4VQJzWwB+qzoFJVR/AJuvaqnsz7YaN4S70jC
idX3upE3CdYmevt8I5G/1mIIrdSCjWX7PKwlmG2pGuy0K82Ku7JAiKlExV7GxZCVEUgOvuZoKXRT
iie0t7RVVSoftlI5R70H4D5aEkQFbUqeyXvo8jte+d1/hRGTJ0imhwcA+fZG8M3LVUn869eWWkPp
I0Xwwqv01Lh6WndGHXYD4d4c00wczW9V5GsRqCwlcoZMgtzE+2RFhEwdOlG3LF6qOdrYisN4VSq0
y4pB/vgN/riCkohEKJu1vng6vxgKzC296hXl8QyBodfxWC72Tw4GrXtbaSVLCovMIMZSbY3QtGA2
laAb0ZxYt/54h+cahhOdG5gba+j2W/VlLDUn2E427RAIwXLZy+FDfPr/p+JTmU1mx+CqOUyMxfY9
4MevhqlaF7sYZXcF6t1eI/5LTcLWQKqqoeJTFW7RiF5qq9G5dONZti2mcNqgegxgSVn5hmBz3sHp
tt62bKz786G8IdASsjpdnsBMcwHUydi5gEouOe4YLUPdTIEeHDMuzdfYAu5P4xAIHP2j4kzY5tWU
+Utgeeimk5VL6galJYEvgCwltMTVit1rAD/nfBrPAb9K4p1gGTld3OSWLSmVBDnAKFd4Tfv1Tse3
W1BCm7XXV+5CGLjtrWzZA86AicNAlAnNEXP27UxHzOvSGf7zjveSlGzxGvQWN3I0KNh+aI9H0WdJ
FfibZTttfn+FK+1quXmoZ4dDg2KfzUXedz/Y8jBHqyqt7ehRkChw/gfD4T9/Lf9CutiVNXsYqSK5
ynDsWoPzlD0MX4Rn0bGjyTMaLh5Ua6oHntrRdWJPT5S9KUp9QKt68c+ljODH21iRR8mLjXkWXKRj
8pVzQ4TJSAyP6GFiDyoQ23IExfYsY9eupeXv4jOsX/a77oauxFnDKT+JLG0mVdtUXDu3IoRTRce8
qO5XS8XnvDTwtFavRcdAskvdpqUyx/jHktZGY5XZurFOuPa9BUoULZ8+7P6qAyEq6eywewfxutp1
N1uebgN5J7w3Zf0NkOtUbs8zQXQiyJtT0hioeiALp3gRhXIOjbRMgrx5lCYH7CvPHyYzkpCrL5Tp
OXek3P6NUB3eAkVa7Rd8fpoHxLqwoB3YvYt3C6tlajTgQjAKmpOzXE0odY7m5XJp4OEP85QBzFf+
7Z4tz8QA6FGMspP6GgffdM0NW3GicdqbXoeOu31AuYHZbD5Amt/MCcznx6mzjeMEg0Y5NsSSPcpl
GC3S/CFF39fVF7a+OHAJ3Q5/Jy5DTZs2b+g8ctydU/Ufqb+i4S8sJLEs6OcvHMdPbzCjmUimjJxZ
bx4D/O+weSVR5hinjkTsrEbKIVOtiLd8b/JZRGGzLYxAd2RRAr/p5rComHYdilKsksWQl9FbITF+
TA4Z36MbTzF40DsclzsIvGej0E6lmVZo4TbUqWIfeWIDuMKnWOCtluLu1H7r2E6c9AyFzSUQF0Li
GBMICRNv2AAeUOIiu3zOzTz2CrQWFejRZBsX3ONEIun5GEk6vA9VorXzahm5xBps0Fbf8VLPpyu8
T07Epr5Lk+gRJAEOu6pnIqevibTc4SGux9DOoS8p3XoyBxSJKcNA5zlqcSZbf1dMC6ZSZxpy2tiW
mdUSUZA1vnfcYv8FTop6KibcVpAgQL1Ik8i7YeCICuYpxge6J7tGmkGHSeQFW6qTl8n7fGVoC0KO
yjcYqrPtMZTRrTyQ4T4Pzj+J2W43U+rikApRW3/iT/WX0eFqKotNECo95nZ2D60JimtfX1w2Tbqs
zpIAYVcd9AQCFvqRit+TDAvAPMtWbPbLM6x1dj9RbHv5crU54oSPXT9N/we+i3g8AcSkDU5asl7E
inJcZJX51Ep3hc7JF+SILGF61IRkhf3p59P5x5UQfuhNoWr5dc7aBI/dyzTeyrucZFGaMKVhNuJH
/mgwLzI7CJd3/JfjJHN5Kq8OzFvE3hSRcGP7maPIebz1LlYMTQddsbRgupNtCw5Jkw9jYdHZo8TI
10uhAN0z7mFQoVDxvHm6Wcr396PLRQkp9/FXvrqYRCsoh0pIzFtMjfLbb3+xSth2TQG5gL5a6K9I
kGvlRzV1+g3d1jjqlAx0K8fFL51ETfz5PHZbnrA/gLIlfPeFAWUIgMsnbfi5I9sKlstNZeDh5Jo4
5nJfnqcK8ChqwuI2uy+faiLpnD6bPO5/KVOrPUJdJrcUi3QGCw9PxWvBD0SzjF94DYlsV51QrycZ
3q1oU2c7OePpsXxGvvhm/6PpZkfRy9sgB9q8SDbl/6rlxEy5GBYfmklGThnlHqU2YFWJdlOExmkq
VN8027z92fG5pX7n3qWj0TlGd4RmA1L9Cy7A0X6jlilxGyOTZ8cjk1dpa3fNsdrWcZtu/FxzBzZz
coJAr+Ib6JIoG7ivwVjlRbE/C0gO6QxSg75vDq0wikOzFSoPvazDbM8fgObGNxgAlJc4F53lMhwS
LvWWrMZ0UxdQWEEi2xwTFw6ZHOmqGQfmAsmI9WvKb92Uenn2Bz8kDqQ+szYuWBFtFOMEjpUsIWbD
g0nmKCjuiTDaAAlO9ilOGedEXhHZluKqmpxIJpWyWOzlJEMc+8oc70avnACxN3eebxICdGEKtuxd
7GWq5G1fPVlbzYwHFBq/ELCbOVvYw5SXb636hfCgpZA2kTpdgicEVNymuyeJlMBeD6DGciy73wBO
IE2c69ob7yhUjDtklzvn1qKV1MJcZzAgcXMPmq1m7do436FsIP+ChSLZeqV+uQJLAZg/Xa1UV0rZ
zXFMgW6mJPN/OirSyww7FkJV1ajrnx25DIa7nT7NZwa0aSXOwSpnzcvB/onQM8/fcZ5KkHzpDQQj
OpmXPEsIMyTHERuldd0QJTCWMDU3AYUuGkNqbOBg8uAbrjVtgLfK7b4wFc8/ySux5mMn2/i/7kG+
3b+lU2wO0f8c4FZp0VhcL2hyyoMxPL/H5habCOiPeRI5d8EnRPTWBmH97vEDq+jzH2FcrnHYgsxO
f5KzsIE3fNAA3bDsoaVUgQrmq3tH+aiN0bl3hedwiN4vOcyf+mPztuVlzaL0K7cphyjXvSKr6FK3
HV0wisO9sNBTBJDRhLq7tY7RvvHv8yU4Jo2nX3rPLlL9tNX/nZ2m7Af5Txy818KO/q1caKXtbHHj
HbgfJ3aM4tzP//QGAYMCCagA+6jvt9Tk6Y+tIcF0pPjDHYIoTghpP3psiY1rTHRu6eIrke5CQlNP
mskqA+lybewYmi7proWTyymHEiI22OOMNhRIv5Ejwp10rNlyuyNgiJkqlqmA3RTepV64+ZsLpz9i
JKSTB2+vd12KKKTqF0LPThPxxOFKQHy/r2feFWu6Dc+EUxsz07W1lFYyFIzL8LThAfcx8n6yV3j5
1R+u01E1i6Gbw36nw/pwLetXBl+bBtS5kQ1LtGZW/CwSOgs9Ck05jq4KEfeBl3zlBbahjGzNlMrY
h/iGMIR0ipKBxFFYqqiFN0Ck0pF/3lSDpyJNc3rvgE0dJHgPbeM4tLFze4TyF6lxEBfIBZ7125Yb
PhfnYeiZdteF1L+XJBS6oTXqCUqit+5Kzy0eJbAOkbfTJAlG0sfaxMP+lGaSnMHep/44szHL03ah
XW6jhypvgft1KMW8zTYrfSvRgOgecsSVARQTg+yn7ZqPB+g8FU/ga0eiwD2IikcFUaZKEI2d2lJl
NfrySyddHIqD6r5ERpD5GqIRxi4uTTJtUxWQnj0BMMLMZxvNFTsaKNQP+yHCC2cEJFqZ88IHvBVo
4nnQ839eXNcclM5pPHNtiZ8riiffMHJgnpV0zCgnEIiPPjj5X+9iCmulGCknJSOVoFeUu8QwRteC
e9FtilUD1iS8/Eycrm8krDRpesgKsGo+RAJFZRukZMDPnTe5HxebOd0LmC/EgJ82HTrLdJjAZnHR
vn4uBkDXskn/vodzNy2aGJrxE0v929qH2VOmVRmOwAfPLrWgFbzJw8V6LC3jXCNNhAKSdW0GlaEG
h2DkwHfa0KFlykYs7KFnr7x296rKGc4b0VeM/zjS3BKDseKRDsuvroY3wnFFK2qa9lmWRzcLtEsT
Q/NNWe9+sZudbxEf39SRFB9g0LWw+Br3n0fPGiHHJA7I55oDu5Z20mEGoNYBYKanCldNntzw9Lay
U13lzA/XDVwmKGuKrBmXPyKTX4/kCczZaTahNu3DjcoCtviHmwi5OLgmBdIxq08sEfHRowYMXA/E
2rW35C5oSVWDVQdYHQESN/z1Q1VI9isiqtRHwlQtnP59wkKPIjLcQ0V0eEo3lUxuKNXZi87wod6L
irBbprp8YtHVfFf4AWZw/AyXK0F1MzsEjevd8PCUHfrXlWQiBtcshYi12staUr8GHRWUulUvmMDR
oMPn/huXwyCSHZBD4duD1vKoqivEGic3f911hYrgLajf6rxUgU2UFHj4aVwOpt8Fo6aG54rcT9m/
p9vu6NvbMudb4PvNGfrTCiG1DEKdqKIBqJ4ypwukk/x7zSc84nSGSPr+jqN9wu9y77Qd1gK4dDOn
8u3ZUoQiX4GLPD+IfZ90F3mQLOouqDAffDFsnWti1NsX0L57O1EkMKyrKYqRomF4aEs8fMRFDyiC
8/N8/vneuoE9bmUfvwoDh+vfmzzPPO3Jrg169rexMB4mKq/CBbqB5ENeccS1VeUYHmedtixhCMJW
o6apuyDakh37Llr0LQRKq0kDy6zoH+kYAQ+wcJOEIHMgYf8s54SzbmobA7MeV7UKuq3sW9SiJILo
iBQiX19wS3Lmqy7opfKdVFMSaoB4v84Fbz1Jt4TAqaK3itJCX9wvzUBH6Th93SrvKt72adZPUw3c
/7j3JZWztEHKK5XeDgzgvTmyieI8E5TViWNTNhV14Js/1iNItcmhRiVo44SKKUUeDWQ4XTOfThCJ
FkKJ3Kw3u0K365FtJ0zWTZC6pSpfXbwbIoVjDtZFLlCEVjwqNY/U/3qAoLwd7mfOUSzUGlsoZIGo
ic/RLzjCjM2nI1hDqJ2ogzhrVtaNloKluIm5JdmIrsQ6eKB6n1wJVt/G/i8jV0Zl/VpqSFgPGQ6L
mFTZw4jNetge4YZoF/kTZSwTQV0dOTGzQFsF1EFwuIxwuUEJF9yDb30uUalxSZSHWXJj/OzcpMqn
fzWY6VsPcw/S9rLwPGc/cHju+r73aMWMbFBRqcdHAu/Bkg1vXBA0+ttjAUYXZMICN83RW5GwQ0f/
yn8m1w3AW0/xQcQmQl0da+xTd/StC+rPrIlXz0m0LaLenHgXm0MwT7O5+pOhJbUmUE+5jbPkjI7W
fif+hQ/A0cNavqSPPxTTmED+cAiMm4ALEPWZaMiqhwrCodapUJPBNVzOZ7O0jw79uyGfB6kZrAhX
Wbw09nl/uTGwXlj30fmwRRZynN6w7Zm0AvdI6H9z1uUsVjIaprkW/JYQCWWyXuzEWJTY6iYiN7Uo
fqdg86gTR9uPORuO4o06oenaz2zHNhMwOboojLAmX6Pam+Gxr/xFqBER0isKJQmoyXk26/wYYTFI
kFtk1hMW2y8whazB2LO118x/DL/WXMi4sakknXC6m2vBrD/TV50ZWtwN0RrLYuqo9pAGdyHXo0vu
wQo+XW3M9FiURXZndEhG21x/ONgIJjkwFgrbc8Q72sH0VEdKda4RJC27jYrHBwUqkSTD6H3iqAmt
lRzBEEyxOMqURvH9XQdWm1Hvb0r8ABISXcg6ZNh7Gpw7YFof21AwPcsx4NP2TH9KYbsTQCzVU5MB
pGqYxXl/1MdzaD8UDafZX1jW7NFWluUvLjGb8ZFMjNIK6Fcv/xAg2ERon12u3eyU+5mvmxxfgU/Y
Z6tTBzC9snu/d9GxeA/k3DZKOZorqiThEA1kcvS9irAUzEAIefaYvp3op6AnCRmEplef8JI3+ypx
2h/tbkU+VRb+hStWXCcSNK0K7J6szf0NASuZPZN7PrtnZvEdX+1jPlW6zqYseQ8pAYLebJOxVX21
UPL3kTPcHiZEoARYg2+ysTuwT+29TRzVzCYytWA+2iiPYNE2zVuWpYsBe+Bhkf2z2IyGrqvarmZc
YBq7Wj+R+taNPOTI4WAq53ESg9fH4tW4/GMhIYuoTlwJcu32hjE49Ew+Et2F5ksWmLyf0g2eyseN
FsdPlGDsKYFtfuJ7Lm2FvTtiH4qyd0vCG3JTAvGmE6+35zQFdok3VGHw6650eG3yPgdRsN+P+cjB
x8TIYNgK8Lg99DuTFGSHwJtpqheHZTqXJ4dri6sxT+z4tfYZ6/0ndKSJRIrvyniQbHop6Hv88RnV
ulrrjvW9qzP+kR0BbaDDmbN2wz/pOOUV8OFbK2R3Xuv5cLfTNi4ORsvJ2rVmjqyEowc0hB4CNhm1
e62P5VMx9WtH/TSl08N9TjOh5hvau3YTbcK2sPauWNhDuU3Nc1IRSXhnfHj9mpRk6CGT7yCrYWN/
dncEXtgpLOgKjfX9iGaZa4CKeWjY5JWQNzrwZGbZhbeudt5+5fSmltAG65fuLJnPKJ3BYN2Gh8MZ
XciSm5H3jsp1dWhMBfirTI3zAxlryoIFfKCj5enst/igTAzrCQkDs9TZNCMZd3oONiPiLm1galHb
cJMnYSVn8N5CAOUVZDqKZPVWOxF78BZMGPfvWVURgRzFAPDjXIkMqbAjFOj2K0/rVOU21cNVUjem
npQY7chTZVW0b+1gA4njYBU8ibAa2RYEny1na1bCsKB4HbYOZdSbI2RkN5ft5YMHf8GGFBLVKLf1
gCC7HWA0Qe0zLw6UZi1BpiaL7m+3hRcrQ8Zo7i9a+DeY2eWMNi5XWEyYA1e0o5Z7j/4iBtl2cuK9
IFPAvzI1jrbrWI906ei/FSz0H37LwqDDbeUt7oolSWlZcnNLOzFH0DTEYDreQJsHZusRbRdWnORu
z5f8tJVJA+BZB/IEv2+a9EAFJ1ssRLokJ/8kVJzP0Vf/tLO3WQIxqjqUfMPIupcRBmHU4Hh0koEv
vKfoQr38CJcWT8wakGDdByaxFoM0qq/0+7zt6oQZ3+DkjekAy+wQoQAwyIrEDusfn2+h6yZBZgvs
ZK7z5LxqYMOEkDLRhr66XkPWM7xEZDiYCaHmXjlJtXG/dQ2t/nX+N+7XpW79WxXdXOIXYFP2fqpV
Ki8d42Xr+u2fgfVaa8IHuSplnG1GT1k1Gz3Z5Uh9MKkK5UCBCJXmcyJHFuPHJ3sxAvoDuo7GcDvG
5RyJSzFIxUy3ZGGOvVAPcBGIqtfjOWd2323LNtDuuvqmubZdfKAFGZlTbxSn9sajkuELeIRf684a
ET4sSESbpZXhr1pjzk0Gfo9X8/cy554mPS+4fqaN85hdrOt8pZqWRkx6MymjJSs4kE5+L3aFnC2s
2xIkzXB/BRPQenGBPqEHyEt4zhiNBVNUGGCDHNpEBzSPEt6okQKmvLI1d1zrVrguCA5TFO7CTRM6
hsjyQvXjZUzEk88JTwy+F9PbpzkuLRfdsRkZPGdNy5TagQ7dsxDjYMgXES7aqTI+ahjRnbnUjcG4
Joi9t9SNY0dDLYjX4dNQCg43W3SGaZ4RsxmKZ0nbVK+wwztJrG2RJ/InNO8jqxDgsqc4zuIm9e+e
j+ldjU8SLJO/79XjrYyxcQJ9NuHlZl90WnzP0xHS5OUslf95VySTxMD/xzcxaOCCJzsgduWdeWN2
ZxEbLp+9viK1Zk93+baMSqx1DTFeq2yZbdBbKM7JaQCJqkmJ09u2zYi5SfKbD6QdM8Yo4kVq3yU5
4y2jm9xk+XivRxopzdz7maandn8W3YN7eYnzl+CKarkY+SXiLiEEzyYiWS9kSlkwT/3r3JX+v6F0
ac2ZWPP7z70huJBGOHs9yZZFdYKtKUKq4f8eCf0HlZQXVYRyQ/Ccz4brZRSNwXoWpughdC/Vl3hw
4utpr4ZHywuFr1j5BdH5DmgSlTWhUyHlQBrcY1nqjnyo+ih3rNHVt99tv/tx/wZAIdxve7mNZk8O
xbbTdi9DmXScMqiMLT9u1S5cyYpnxACDu6Jyf+/0yImJ7ZGG4vUxKAJw4hCQ2+hR5Plot+GBT5WY
lPhsi5KOa58knSu192mm4CWvZcPd2J4DO+x0mD86Hx/MQ/RuzAOg4vHTIvnJ+/0Kdyc+hrow2YTu
7OpW9q0eFdao5RjHuFaVgM2XZn/fbh0RWrR2i62CBzmyV++qUd6sOGeqanyTxK0dYmIPCPA5gD1M
HQDOSJHO23uKmwogQT+mbhEXTm+obZp1t9E+c5OQufkLRhynumua6A5vl7fz7XJclhfKTapNNomg
qGIb4tjOMKuYiuu3N6vc3KuZnmZrpg3jTiUCQ8sSzcEdY1ELUW25wJRKfyDeYfSTLDqsa0l7TwKt
XrF9upfbvH8e1kopgmmqoQPJ4Un1NqyF4kbgqZ0k7HSTbobqatsGh+aC4HFxl1GHWU36StSzPL4D
9UIXAYgvkm60uF1DbhbIDSUmhGjvL/CC099qmtM0OP1AECTcao+1ESctChR6wqRV8ZYqdh0WQ0s7
1zpxH7zUGBBKpPS4pwDhRo0zXW9bMDLABDJSdIB4EMh3XPwzQkmthC16g5dsXVMwYlOzAr3gzuH7
gspcmpRY/P86YPyQhVxSSJHyGx0ZyNL3HofEP105R5skmmVEjVQM9RTeE/mXJ138VDgXFHp57w81
5qHFLIwuO/+F/ume2iB3wPUu1jCcvM8aVcXKpZuypmkScgDH41cjpYaNKAuCRAJ3UxBffpwtpBUe
GHKtjjTeqZQt+dl06c/sJIMvvBupGbQVTlemv0WIru/gyBVT55N7DMr6qnbwaeOBaG6PsqvaH8zJ
jSf2+BkcWiTpEkbOCiDm2LxyqgXwOtW5jyu6dNYRBqcsIkBizDlMy1FHYqd1zPKSKG7XbC4lc4q0
kT9lLbhm1hAake01OUCfJOz5x5UsVI+d3z/LVTzOtNm0eeOKhpquPUpmbT9xThiZTpOouxpPw5MS
485Gpgx1ttgAG4TDDgKzBO/vRCrFddbk0kPFy9v9BMWoxQyfDurHADdemcu5H4xabjvWow94r0bg
UGCx5ORwpLrf40LoBdICE96vZs/a150WC7jziBnWd1onINFvRzNh6Xv9Bzndy8NsrbJwctUWt81M
H1+byXkJlzrAysF/BTTgb8+cpryCOOG+vW7NJ3XXOJYrJi6czBOWQCWiNc505FDphPgAD9lhNnx2
JWg8MSlqPkUaH9d1JCCwbaS8084mi/ovHzcVti2/wtGhxiRfugFSiW1vkAIThWOfpu4FPJqhwlbX
H1/gU3V6uxKxg2J0esdAfV5qi5L1BB/J5t9iy1MJ7psSjILes26THwvQxgKy9AUpMMVJO1VrQ78W
0Ao21dG5y/gsRpPioK47sjU2E9sLvieQCgv1DEs21YSRe1ZrH0OqdrpbFUZngdFzodqRLPr1vkgn
lSwTdxerh6P8OGEPQ+y1e4p1+zKd0R6AhvqN7Lcm3Kq3cp3YEp9AW8mvRgk9u629r65S7Ipra+Ad
NjDAG9qye7xO79/ycUVcgWBSgvO7zOh2wRtjWcQdmfK/pb/k3SXVyihzaWIolk1/JVPoeMjNF7IG
3jBhOYxzO+0No+AVgPavf7LxzoLi6g0sLw9rCMpNwx/UTGEohj2OFVQjytoHnvUf7meXhjwqNI7A
m/fvnTDf3W6Xat1A++Ngew7xPiL0P4Q/Fdpufseey0f5RwcSJ/ioKrYHOv2soQGRdnASgG0qvagU
p4oLlkZFEteaCfZ+Oyc0eeEHbX/m1+l6Eo7xlVxwAYfDs1H4domj8FcfT5cjzMho+qdwZ9gzbhwu
Bc+zAyofpGvT8JEWKk+TuNQMCzXEk5arJvMnKIUPyeyDtUE2o7GdUf9ZrZk+zH6eBrpwTT/GCefe
g6cNwTUvPjW3qN6484gv48G+pyikaBzOmcezx/pH3pwHCoQqAOgEuKib8UE+BYoHzU8oR8Zn44zq
Y33FzA9fslsWVxsOu3bj+gv5Vq8MUiwjOPfmmhljs6aoEEd+tfqUh+U2apSzKgPv/TcA3srefJ3w
e/TmSrnGhW3Wi3ULtwxHzC/5fxJ3xKSu+81lhc+4smZoB2iP4gRYhgcU5NxElDI7jTEa/dE7fp44
+1/tZC9RM4ZoOFYDHGGbEVQZ4SC1LfvN8+Dy+cj6U1NKLK/BvLB2cAgFCycq8/aPCy1SKmKYVFWO
1BrPR9PNd5In1dXNeRuVryo5UAJ4V2YLzndMdUX6E88Tgid6c3lWl8HRIjQWKZoMvZra/RHBXYhm
K8gWhNQb5CDprmJIxN5PdNEgzbytZsAC/XGHV2wbb96nB5JGFxosmIyqN+SVF+OmPdD46eqD4OOv
8wLN1iebBylEZgKBfNEJP20N9dOjCy6Tumll1bUySWXdLhpdGbqaDv4oqXJBlhwTvOHN//1lbIqY
XPujzW24uQKmnsTvPKM9+vene75P+V1EOvB7wiccxXUP2pqA2FYwCV/cN+5I2QyZvcucIDb7j/xv
4jFUxJh0iRVHZW0/xn+tAgLjQgP4RLcvLrRpYE2lEDs9qArF1KdjGx3I8MoJzm0ZP8Y4Wx2JaydK
6Fkr592X+Oa0PZA3Nn6eir4wlN250VekXDqMqxfGNsAa3JFDpP5itrd8G4m6Yw1nto3UuYklQIKT
pJKwjNbD5kXERZEz9fCUd7KpaJsZweTzJWP8huSlGESb6x9jIhWhnVcXh5LJh93xQcq4jAxWi0oL
UE5C8I1mK1EafvHA8eF9g8yj7zYg574swYHFrvoxljjlhwPdvE1nNhZRKs1K3/jcfFYIUCXyZngR
MV18fh70aYajft2yyOEAXbrq3QCl4GuYJRPV0WqtEeKfNHi1Ogqc71sVlJcjOy8W1g/MsAEv2oMm
h36bapSaKzFsKTAs0gVQr+q76VMsN00BCfBN8iM8NKo4ecinRooTaBuaUa+HuTzfB7BQ5U0XQlRn
v4IrUp+/Jmw0Z0ymISCinoySONg6OmdS4jdL8KNaWlvKDgWAXgz807I2L6HMV5lgs7672hik9WWK
Cb9RL7k21BHfQQdXFjWmjAGSR02ENVwmh54lJMMdFLmCC8zP0yRofJGLVDvGsIATFKbckdzXOiD/
p8b/xJmB/qP41Dkjpm4uq1a/6GCyt/eGhPoc0tftsRSSmEhg3wPyJWZqIRImCkSXSrlQAQQYjyCZ
Eo6kFc9Ci0SGu2jMdorwjs/TO2TrVbyFNjaTT0JxHI/av6WGqTdQJXx1qy03jCFe3WFPBzwKjtK8
hN0VS1tzX6Jhiyuz0Mb6/EDk62/DyQx0kl2p9F43zk3BmvNHY7tIsZ1+r+8hdH10WlkLHy6xtpUV
M8Aj4WtgK9o5kSEXZKmI856XYrZcrMCRBHINP/DXJOOEJnKq74Z+18LGZlEVhais6RTKCE8lsaQ7
x2YN7zQrHN/oDBeVHftrwl98b8eRV+G9QVEQDUh4vuJj850XJDWW1nD+gTCfVwUhwuPm02oqM33J
y24RQoTrhcbDQA+9AibbeMuE1A6H0Ow+76wlp6MLz2RfefFnf35Yc7YaeaY2rHBBJf6ex3hsrqWx
LN6pik9Pg0DWb/bMKujrs+iDDtEapMGacQRKjDGoZs+C0pihtwlZN1fYuOeX+ey1OTJbvW0vDVNf
YE/AWRFmIS7EqieF8J/qrjnRp+y+s13Jalkc421/Xf7lOYQqi17QVITQeQLs3L03D0SWm9PF6z80
G3gu0BXemkCH8yGarqmAfs7dlYMcq8RjYDs11kjjyVWJqqReZkIi+m071VoZb5EqZOJ4sddtaqdF
+J+6mKBOdu8sxZV10gBE8nUU+bmVP/I+QqHQ2h8qQXTXdJwn7lzYR14Gr7RNrf6EesxKjriL31gg
dpOYGOnqgVKAlwaFNYwYamjV37zIE7ZlUfCvEnif3mRolXqCgiqp6qpR/LqpmUxB/vCMV4FGXV0n
sAru6UeVgIacJT7XhpfJ5AYN6KtuQbECaxCWKoZstUqYDBe5SqFF8x6k3VEb19Gm+3fpVhEca3ps
Nrv52EeNXvUjKLY3vDzCIDEglxup8vw+dMivpONrXhwPdm2nLFnDjD9gqZ4wNNJKqqEa6bh2xtwB
xce+xzJ6MKtUH7MXaaqpwrXoa0OpVDb1xbANwDfMz2WvE80O0xt8W4ajURW36bA8dx3a6Q2M6SNG
lFcMD+cMKuffuOZw8ofnQBwmb5OTMXjqq6tCXiejwzzOE2FUPP8X3a0jcARCem0OzZML0uApBiB/
b73A3At0wRRDtoAKik5qvSJjiE8QgXWSZqPVNeGORodjdGPzq1oX/NbGwN0cbQmsgzQZDuRGx0YS
jRX1Mqbzy2C27HlTMEdxLvr5xgV1EFBOiK1CKZ3q7aA68PO7D+TSR7wWmq8Y1rlqXi9OwUP+sBNZ
67kiWqnxr/ZpczsTUgi+iyhe+LSFuO5ZdNAs9prIblk3/OvfrmRkF/0FUsvuALEmoIIpKrpTJ68K
HIrd3DUnyrHgWUf7vejGiwK6mLduAS7CrOIHz1xgTTbhWXzw9mjiQUelW/pTvT/aLX2G3ozFyu3o
iEBSa7Xzfp3fYF6Ebj57MLUlmza0rAtzynrD9sjaNn0FWW5QbV4eHchIpNPW0woj/DtmGSpFhSMG
C8vwVaNE1Eii6Iz17ictDhHmByZ2ROjnMD5gmmzhltxyoo5W80JbnZQng1M/HR8O2fAUQDbqFYxG
bhYLhOgQNFMM8zt1I7S3gof7ugK+71KWOTpyGrVS35GgCtoafnwIsh+4fzlUsXcdhLZY9iA54KDm
34VIyLEd9XGLhPzzpdWQg26IrpTbs4S6/nD7hvEUBfPHcDS837uOnjHW0IHCsJtfhNQFpgmRzE7E
H01bF9vZZ8tnsvo8ZCQR3WhkUx0/1u5EGBRWVRAi/pu3hjjOiWEYp+lXDG+gr3hUqZ90SlxYTCnS
iXVe2XJcP6NedN3oGmL8AHG5Xf9IIpq3unh26WWxttKnvPwF2aP3UUVvMLnE7o6zB6b9vU0Kes2r
Lwl+PVKHjYRAHnBDUh3xFze7sIWtZy6iB9xkHKrsBogNLujqd9C7ZW1D4tZgces5bmwPhr6PLCjM
fPAa4/97N2y/H5ioI2pK7bNKxtRC6lerummYIQFSWi9f3WZtKeUrpET+wgft6jW8lpmrANU9pSRM
2sK/X2ZFYsh0Rp5bjpLM7+VSVDbfzWo9LvU1mwJzLIEPYzvZjD75Lxkc3JQeBLxXp0xFmkQjoIJm
szFFuxGPkqZUz86JjCKCl3SJTPKlS4H41aywmy6zQ2S3kMgM8H8Hoi4IqhoYZJdiQHKZAiIt1aYx
2ZsKSNwfm+Bn5fqfSrNGYwZV9wGAaalpgn+uomefCP58MRaFrtB5ODMjLIid3SWKKY216gPxzy1l
BvbMZeeT8mEwPejcDvWildT2fu07SMVIQApRVqpy2v0Lo6mTndFoMM+nLg19mU+EMaRhYREjR2JK
fbSn5cQDY6MVSLtYkQKrabO32gUH2fdWVvAfVsFewXmKnXFrsesJ0QInGsNPydNBrYt/L7ygay0h
IQ0jIsSwnKnHPUn/DphzpiMyUROo61i5lTSmRdUeF50pGzCwBS/exE4IWawseVDP8m7p7jJWKVQL
/xmgag1EHDFp0ayN8/0628QGKVom1ZxRxJu8z0Wv38Bk9OSWCjX4tvWhAkll5e89KvOcE8hiDQnX
Vk++PN5tGDZ9BtSzd6ZtJzFLrT20Inif20xqbVQlKaBdd+UboMcZQcfeqXwtMWgoTRuf8Zq5iszg
uS9u271N7nSTI3+Dy/0VdEa0JxJS6aL2hYupl/x8Rw/uEQHy8GY9MC6GpoBsDxr0g2U2AJxBWEGb
ikxcVpLYHjUuqVwmWlQ0ZFyxrSTFwDs6umM/hvJ7asuyJYyOeFx7ipzqGeyu5udzno5R5xYvrFdN
GxrwCX0t6uBEHS89ks4q2fdREses1tczEksWBWHOnY3KOi72y0CZmqngX1S81MDBBVhXKC0UloDf
akrGFgrb1eot2HfM3GxENNLgJCB86AoitPMm4Ok3pE1Ok0Rdd7a7u6PsakSXkldP6idB5I1w01zp
VvyYVIGzFlDbYanNMC3fMbLCyGT9v4NPoYXtrSL/MgbVHgtYqhlNmdSL5WEGIzLu0LSN8n0ngaK7
nVT41yALzG91w1oqh6dM6bxBJvyghzFOGH/UMrbzZZdbpQlnseVSyshYRO5f8FqaR/AhUF0FekAc
DXVUEWy80w2CeE0F46zqtWQYglWeXyOhG7ghpZNyWGSHs0ZqlaD7bQ8sKd8gvOdMn3cY4/xhOffL
jw0Dq8nBi1IBnb52uIq+lw4WuQx9Fvb5f2SaCy67Q+TUQbXqrIU8JZls4s7tRCze6uT2CkR/W0Qq
cjrZxE0P7LuXKrxYQ81UhLODWKj2QUU6e0Ajt3zzP3bLtIEq21ohr3ckzXcy0eBidvXQ6t3BMTlg
qkFJQ5vLqh3vHN7KrTAWf4JP7EbmppQzgwYraO+87GLEvmo52PYArEMbTK/G9e9aVSjQAgQrVevt
RbRlIBHIViPtKnz89B1jpF4dg2gY9L1b33GoWjC1SUT2AUl7hphrtVoONxeSW9gh8RJ9pKmtyrcW
zpgUXOQVtEb2giGWU5r2vfdal35SdLqpuxABx/Xi7IUz/sX6p6N5zweoAoJnFdIjUHhRqm2DED2i
46uMQg2DOePhG2wISOeTzNeCk7+RxnLKAKIs1y7rHfXsPRhhOAQJOTyeV7XGWM+RPmZ0iw1B5vP1
Flj2qE3neA7pwP2sPh2KPTu9FNnwjsGgSqSXb+e45Jzknz5QCGk3ujL8RuhKaCtIyB/yR67ElFTI
d8H8Gc14GzLvceIAkyWplLl2jE3f2Y4BewY5/+uOxrmpzH5fODkHv0T8R/vFUhCIfCvOQ3Ne/2iT
esWhPNubuVRx6NZWHAtctPmHqS4o2fygzdJgiYV3iC4Uv9WIBfGe3ktfGp1YBc1tWGQPvAZD/wg7
tqdb+l47hxz0opi/oLgM++ciF10FGNpMZnk4UMIGtzax60XF/w/YSTQQ95sLuwg5Iwyer4nWi2uZ
S8i6FkvQizWcfBDQ0owBRUEljMpayNrY5oqIp2kfjsmO+O+7fgyUde0b2ytyDuML0ll0S5iC5d+z
iTTS7hxYhKk3ZkXrgONFcH7NyGZa4ZEIEcCi1FTDmJpiUfdH1afQViVrZFnHKu7HRCYzwutjOQ3h
bLFG9CsYpPCac7j0rRlQlqOoBnZfmyDWkMRZcWbjgWXE7TMG9f9Aa1It7VtvhfeFmyWSgAJ7lPm7
Ljdr/yboq68BBHNcCdqfPc7xcNY3bVsvJWYEzpffx+p5ciad/NNxXQ8DDMkvpEUrwKFedJn4WdRY
YpmfBGJIoWSOqsQHGVUa1lEP34NgMCWMcCnSTWqUJONe+eTHLED42PlKXoFeu1ZO6HWaeI75E3x5
lLdnYpk0DEL25ny2e1Czy4eth2BAO9XEUSDOuVbsSsXCzspH9tzwRXel8HAJh7ubWHDHXAXRGfzK
XBly5oemLzv6oByf+UqrdXSp8XokHnIKls67IQeJHdZ9ZkdhLQCL0W53pmJ9VMElccQPokJNvnBh
XYaZLOj4l76lbqhYlexdZYcd7cLX1UmB0Bm89jkGR6przOgerHrL7y54HcBFeP4uRQHV5nrbLNcB
YpnXBlRGMqq35iTWjclSn1CV6uPD0baOJqXArrawojZpQ+yUCKbARSSHaZRyPsfw9lHe0kUkJQiP
OJGS4s5g+QM3zL5hJYcQNyS2/KHCCdsYUdp+2gHDY/6URi0hT5yl1olA8IOqwNNcp8zsCHgqEgh3
agSPFszJn+rP8lHwzVGVqJ4iyZHQgHOBAd4hzLB/gcV3+kdeSRgRKasygvsTGxz9pco/4RpSRuZl
6pxXSLRRCA7GtD7yVX/OSuSPkWIfa4eUuVJ0Isj1RC0WsuwCqAwtHsFxhHZcxYngWFn0Dqv0zQKa
RbQQAXRLghJp+YIhqZ4LfzNL92kkaDnNwEeWcMmXMbHWWIT2/vNEbb4qI3QyvvyZ8Hf78ZkE5taU
jr+D3DlcST05QpOmeMBT8bQ499iOXrsyTNmZ0xdS4q59fyy3g+Kw+jN3+7ihYpIUOXbeWu0fPoco
cSMLvbrX7aTr4GRgf37LonttbH6sFnDCosXAQ2CHo8WDsTgxrmwTI31Gt71MhixlXx8OLFyTUGO4
xhSp6dF0/s/NCViQvuPmTxWetim7Xa3S3JJQu3bCAQKE+uadEQxs3jRlKSrWfQIm8af8tl60hCH0
+xgDjfZqXW0KL/R81E5ElqL1aAQTuhREZPXBwKJV7taiLp8A3cpySW7h/VZ3Lh0ektW3G34M4nUy
zNbKLZvgOnjBlhjI6+h63UtCltxfETYlzYXSsWJfZQjK/AXX01T5mObCZAmfmjz40nhwslB2UKdF
GN4M8jy3omwz21srhhEav8M4T7iNctFzWb3OI5zYL4h98A8Purm34hRrWcAkdvAFt1ogB+l8ZnzW
j6+5ry9zAkVXjTRvp9QJfO/9ojEpbmDqn//kLjubXDQFxL1+c+aNmkShu/vkaTARkK8c1XYKzX4C
c5NTW98v9xZvXc6ed801oz80nDIajtUIlRERLIsBbDc/FX7Htuhg22OD0mYEfbwb7LRVZG9qHfuX
NaRQoaJy4BpgBMJ8DMhm3Cez1acNMuLQUFjd7kbGDwFGW8vMNy4faecVG6xjjlP889th7+k/rGus
MAYdzId7da47+hbC8sMhyCH3TzUdElsETYsdNPo+boEL5YaZZrGmRzF1QMW+/X4jN6SkSq1OTB8n
gFKtFnv+1oRZt3NNZo9MEBqMlLlNETZIjbBsm0FcGHLIxl6DB9zlKyvjQOKDQ7y/Mvh9VYuUOD3Y
+OGVmGglcCzIDvRL9AbcBqMj+1MEbzZUuyL7fAVu2GZ3bXan45jpeWe6eMhDhsBIQTTrAds2Gnny
cqfUkftV6UpoxuTVCqzzutGlv07dgRdH9SAuTOFEUfSP34FWGNt3wPtvQfct8hVbJkfSU0L2hbIS
QQ4sxjZ+qX4AUn2TEoMC5nBp8eaTClzLXuxguLmKciHMXqTeC+YnQ9tUEejDGG6IDg9UF3JbJxkS
T11XI7FiSRTzyp+Ns6M3eLyfgg49ZQErrWofoIhlL3rp8ZYvNf/BZv9oqYRR8O7km3dWml92ykJp
nRojrI5ioqgkLIk+RjKWQTOWaGiVhyQ3IyUYML8vDOjmBmRQrvmLT0X3I5kM8pGvs9KehBRI5lQh
J62JcWGZAuhiDtyYoBZjzZs0P1K9nKIhKIggCH27W/GAAARN0Upbz1mPgw9xozZEpi9ZZCvCMhF9
Gf29nmaxtJazz+dUgpO8A14s3tvtzwKRpeO0oNhr7VRCgrc38DYa9aTAcMbrXghxEL9BRNwDVjiS
OGaGd46ZXjmfZv2c+5QI8JDIdJY7sHxg+jkT/y9GuvFI7eZ1s4OcAZ03PCVty7CeGOQXce63L1AF
LPZa5LEBki1pMZmSMRHDje6ZPwy9tjDDMwD5AmCQpPG//nBKPR3+0h1IV4pBGvxiQSQJWNQxaA3u
ZujNgnqv7eE8GIujh+NVmFtT9xsNr2crtUOEWnBMsVAbXeF1ofWqURUMtgUuW/dclRaL1UVKszqr
G1gG3Ev+M1Hin9WAZC1wjv8lsap7+QexMmEPRiy81zk64PftlY//ZOiICg1xF/Rv/DNTbdQC2k+E
1qqPW44x+S4Isl8d5SGUMhZxW558PUEpLsNUEH18as8+yJ0Aatn8fp4iZnfGU5CReYsTmdRm6Jdf
ivBbGT7KdnwCVDwgCQ5utyMgjmdjTiyE8PMxj1G+v/rJPdrkvQ4tswm9SYwWQpWyhmtxuKrMgs5O
fku/FD87CWHPR3SOIcfVw9FDCT84i7kWL/69kRgkjVuOQW73qgun0bXDMi5z7guU7yrGN51W/ojH
vAsODNDWWOzXAnVt93QpNkWsh35QbdTzyt/RxguDqBp7t4La3jWQB9UpPZPjJIv362/CHeBooQiA
p771jTfqw0keOoag82x0W2y1DT5I116YvywINwYrB6cJbiFqK1yX2yBB1/TESq/xS4j9olxzspAz
PpkqtKCTaH1sjsWaF3HsAFFE5IEm8s0x/hJMfIWGT4rvTRowdxCknrwvOKwr70oVnI1HGkYYySEg
r3wG1+lCZ0svHuxFivMHh7ecXU5vnP3X0WiR1TrPomO021N5Lm+XAozztH5tZxC5RzPQ1e2MiXZa
0C8n6P1vbpxnA4Y5YmqE7L0rQLSO7iNWCvwgp542AZYzWha5yH4kd85huA3GEhpPDSrYjhb53DAS
ykwmDwaUnPFoORey57V7wn8A/DdyjNvUk5X7Q/bAY+g6EziiTZPUN5bZw2Eikrr1ho91G+wAR+2V
HafA++NcFBCX+Dx0/E4iFPydPJOyWqxCaO6J/xVeGJHTilRsIKgWtuzSsH87kZyzWa82tPjDqINr
ALW5UsOYI39/JrXpq7O+gGuHXvYof8UVjVSFEUwsZwmK2zFvwbU5ikKRJ1PRgUt1CZba3hA8020F
qtkgOy7RY/qb/ffKItoz4QMFBVz4RJVHPi7m69HgGjTaT2L/bCHaUyshaIOi/yZPJ2ZGC6hpATgs
u3rbthKiJVhNqSlfpDaBkbLy66gEL1i1Ylcf4UTmNommulmJXqhg1Rt3KhfB0eVh+r++sWYSJvCl
I6P//2jhaf3xwtXHCx3AAH3b/eQz8xjxJjAPp/ifxPo3MlroctG9lnExzSGdBNNdz4X50eEKQSbU
UVMGz7ccJH9Ks6AHUNZt17FdatWsg9c/VkzTIMnnqH65KgO9zWQ1MKwQ/6QJm48P/4fSo9901T4g
IsknbjelkMOk/8usSOkg8hIeKlmmeBm/p2DdYZRaiVByZzC1NVCz+fJOszjEr40lvwAZQqMyuROn
OoDTUNsdHGZLtBNJAvleh6th27pUu/Z1eIrVC5fB3dwzk5ylddisIGHur6PSkBVHomfkcXgyMwF7
cQSlcbYVJzgpDzfA3WVkac3wopX+6czVKiY8GgIZpWvK4+EnxEqMU8rs+RvInOXpiR2NL/SbdGDP
1Q1iGc99fghVwGcSC+LTBMB5a6K8OC/LVJVjEkKU4Sl0cxUnjZqorKzfoBRRM308gWofKqVduBsf
uiJWyIuv/u2mwy5S/ZAk9zFX841dqZs1xY5NXPwmM1yObXhSEBbse7AhGfqJyQJNcxyo5b+23aey
oHVXQH0348AfeygYCSL/Z9Ob8ZIxsDDmFVyLBBrd2bV5XHgpa/5OQOBblBowhDGu6FOUlDov80Gx
/j9smBMuQwzSF0FsIDh9U1DSC5NUks62ae3Eoi/Nr6BDAaCb5z1pKHS/JdHmGKyDJkbWJtFkUBnu
cxNuzOzsYlk3ogQcA+HWQ8U3YAB6IWwdZWunlyT52qrAFzoqQMYYahkCWOhDKAFu4vPXTU2ctzZI
xg4MgfxgIiXXnHtEOtzrGK2ipMfTtillqMFgK87jDtaq9P9Putz7dmxHP8MiBU4DeMFvEMwiDTAD
M4QRFSdrpFSN9TAHTc66sG4IFIrvT6YdyzC/TdtV2FrzuiZD9t8I8sLrl+ieKiZ+1qjVafJFwkdt
O14rp+ZSPHr9CFPXQnbbqU7HyjFtAmkub4HM5GQaOrg6DXV5Z0MhpQ/HAK72C6l9LSLKx98e2vFb
7xCHMrtrX53u56Y06Zjw30ulUHMm0I1P1pJ4odATq0XF0JHxpi03wbBrJvvPfIfkdabuS3R8MgzP
stES16WkTeXREFXh+9zw/pzIOyUQkr9ZiCnzw3GywpZBOelxLSPfIrB3wNrmImfP44ZkJKoedCsX
h4JWr4GRqQLYZg1K9zgbfgwbbo9GbuEL0fG0PAswNL5D1W5Uy2DbQUj84dxvO5qUaVt/UOha0ZcW
wdkMuE8Ufw8e/7WxgK/rUSKSFS9pmrth0IU37NPQunU7iRzXzqcXmf6OQtUq6MDmii0+y1gDOUMV
vidXiaCQ8rX1oHn72NfAU/MG9asP2eFK+JOywrxKsHIkCGF6jYcvDdDyfyt3qDGO2yRZHs5VNiIT
k3M9jSjbTymKqE9b7dw/5es0g065cwLURwltJLuyvHV6Sfsshf+trktXgWvmJBfrq3r3KF3J0RK5
6b4yzbOOUgvzprthi79XPz9RQyverhQsBluWWW6esl1Vfj1UNOaPCBMGL00W6zDtlyrmweVxlZWQ
e0ogAlyiudNMdXVrQrN1rasmtkqmXhBjXofONaDt6OKAUErJ6vNxke+XLHVBQv1Doj5DUZf0BHcz
XIvuBnQrf4NKxLMLpUS2x97KGXsMIAEEnt62eNQq5oDiMeDMTIRalgDSP83POYpyhGbbqj9Q2n5F
61bJafVd4kaww5l6PJVAXYm4QQK0ISrnQBlC5J1bWaBc/Ft3RnjEuE+AvUVu5BssuTmWkcyzVe7r
BYYNy5mOqPFLNzuf9I2C3TnULEWneNFZAJjAv9QmyxcRM+QNAKPrJX4B+Y64NYCjM4y9EgcQcV47
C51ZJ89kmceTYeEdQTxzEb8w7rz9AjhhXMtXJ3db/MrgNqyNBVyq2h4L97steEFjGoRf+aOcEMgp
VNeUr2MZ7/Xbvixl72t+Wqdow/+LM9hlwSk2OBV5peke6+nCJ9GfyyD60FrejnQ6Kdin/n2QlajG
Qy3HcZlyrtGHDy0S4WkLnkRWcV+5uosNeC6Ljn54zVbrhtVbZPP6M+Z8bYMAhDOvmp5qdb0DRrrY
mEOVRR/7e4dBZcMl5FFypqjkKBbY5ZIcdkMC99E8POipmlw1QL0OiLx50PD62D/rfMm5UktonfnO
YG92qPEPAJGJudhENCffMp4vHz2cTvRPEYIQZHb9U40Bo3B3Gh+O6CmIORe5ryqK1d6drEjAfmPs
nB/ha7wyZus9DuY5+CR0ITuEdOhvXIq6rNJtQABpR2o9W0REMbSIl4basA5MdtXI9uuGvKjOE5xs
BU6+PulYv32LkcuFK4Zv6eT7bFPOkOM+Znc4bddPSieGMhd8w4y+vIj+vnDxDLlzXcDOO97BMBzS
LyBzeMZX6J63q0vyxI8Nx/2RsXpY1gyXEDgwhu79kLLV8ZKHAPgJd+VFtZheJ40KsyeFzTEzmAV/
nh+AuuBT1MhgMrsayommbzGaqNzArw1h2a7yWFUSChkK8XxAkwFxMIgXn5zQ5ga/KF4tCHaP0QZu
viEk93/b0Va4uMFeh2tyl7DkRg3I+hnWHNaIWkJADBBJeOzuEAftbUO9FGcFLcx0dY/0nmDq7tEJ
ldXeUB6QtoDV4v50ov3ky2HYkCVzfPhc/Y76G//ygYw8o+OUHl89RfrAunxWHYyGxAygFpybZIf5
CaLT5NlnmFk7Yz5PYyIbcPgRPSnDpogthbUB9Zx2zIuCBCp/4ljfK105YzPl3PD2xjaCf/lleXR8
hHhPjtihXc/jpP+W7t2fVqJoTI4GkGmIlWoyRemfKxwjO8y54cE/Gr0eV4vYF4J9DpKVbCagTlLt
4+mpqO3QOA33LOv5UGoUSJ8WYOa+yzOd8+vjqco0PVTPdgSirmBWsIHAGbP9JnSkMmhaKBAsQNqt
PdKf0s1xyft/BjzLo0HEqd2b/ZuaWpovuzd1EG/aGAeE7opN7GVuhE92nnbdiIsex+5Jfx78UIdK
V/2S5ErV0lyLY19QGJFweWCYC9TG2XfRPMW3gGURXa6B/ah21/UI1KbPVzZ8x5dLm3xRZk6eozyh
TIjIPd7OXxJJQ9DRg9pdfB7TMmltmrLMZnawz3Nx9lkpejuNae3hKxtD33Q8mJm8Mqx49l2DDacN
tibH+bmVFaEMLWIF5jo9DqBlKKkTLgFJEpdQKgUajO29/55odsWRHMsv1Tb0BFveakg9P8flbwFQ
V5y7CakL5wrRK0WwV9aCVmOmAM27jU9okXTVX1MMcMbwto2aynezhhn9jimMsny1Sy88v2tw8UzA
V0W7Eo0i5efkQM56BGvK2vCB71ZUbZYFGfQbPY1K6T+8f+npg6BhwnWm2NFabLHeXUmtT8oojgda
xQQ6BVPTc3ecmPh3cLr53MLXjoIycaKuBbxvFq/p/k9RWgDzLhqucByB1cs4+F/PbiSN/9livbzW
lVdYna4oIbhD2B7gRfOcRImABSXsOZ/NXG8Waiozt0KfpMTN9WpCiodArxOeGdZdChwi3BuxgcUh
o1lxLbi9/s3o8glNma+UZyDtNSL4IkQoh/1n44+G5umagfUiLv5wWmc2fA/bnPWaRW9/ZNoap9wl
i60E/VBXXXymYXsULFg3B/Rx1dGnZ0fsIvn+zI7c426uCMOXPpAuwpsWB4AH5VNCs8VaTwrd2X7g
KAZRZAcHVG5sykqximTrW4GQqPKpouqjbN1eudj5w00EFfiCXGULPlqlKUM3DIxPIMM9CrIiNxva
cLjnvbZtoRA4hf3kjB21KkccsxJzSiZ7kOPAlhJQc9neV9tWRPRNqHkNGSJKIKb+lNhP5SXQi7NO
fkEuCOHGnQi0Hj83vo4hmFsSY9eV0nInijCEgSAN2+PqeGp3j8kk0TnR937H0ivhClZhIYXZwdPr
PlwA0i0nwjKS6gVTUx/iMF3mP8kk/jah+nzCO97JxzZQn9ueYnKdygsGXTvXDjeY50s27cR4EoxR
Kbh9FbjRHWtKOJOsTAWDkRsKaNOM6oL9oKYNqPQRrXvaJYYQTCDg0OfKn+0CxWjhLVtB34Dhpf0Q
mA1OmNePNwXjeOwvYUnapG1DRBgwMFbqNnIdY/myst7EahP7GZZj1Rq19E7dAMjo3fypt5W7OGa0
ASo9iKEmeb3d4+df6BnDHWmpDoY2PbC/ad1Gp6OcwXuVwRQt2wwjLryuxO+vNxatJUpZExUmaxRz
k9d2OuGEdsBoO18+cwgw5GhAJcHlf/RcLuOHKAJplpx4j8iw9saROZlAnmotkvCKW9ulDGhyjVqu
8z+HWGIdhKWk1lh9Nj8zgS6l/VZjrM9INFKvFQCaVphterfWMbDoOArxikZKQCiTqAhgzPk0UPKz
QZSiK+MenPcymklTYVLYSqPEXF53kk8w+vyfQvpyCuFo3XVi2rn5bmzC/xcMg5+jTN1mEhp547i+
loratm3+Gj8FPDoar1Nv2vC3XZC78/V+GBJ+tHRhGcqVIS6VhuUtnM7e2/HA7Hxd5/04Ua4oK0QK
Ho4/FhhAid/r5s7lHxsdvyGjoyCzkoKLat5b95XUGKABayUf6AiAGwEPnb/7ztXL1FhpDSvBYLop
UPuUnhfpRJj3SG6inilEc/rRo/FSeIXK4Mr6oJS58DkEg+vxcFHY0BmOlmisDhOlw6SebRhcpqeY
/j/3XB0BamjYgMdtmfNuAPILSsvMsH+z/g0Z8t7TV6EqfV0hPRMgB71yheEf52ovfmk4IP+724AF
dhT6U1L6ZR/OOC8dmur/t6muvQSjP/45r6+uuMBF0PvLCyfrPZHFaukOA+a587UhNoqQJ085XiRw
X+gH4MWHy2TqLxr/4UBUQuEDRfL41W+vmWb8yQ8w9d+ngqKtS8UPWTx07XF4P76ZPWbw0ejVopLE
YLu+mGAI1aL3RLoQ04JWoS58TL4hlWqTSOL/+Cnez3Uqexi5yFvsLWB1bWhG2HI0MV+NpyW/4//E
uxF80zbZtWVx+nW2fx16fR+R1R1BiWi82LHHyrKr+857kQTWtQ+WGs2VOuwTXl1nqtkEGbeTXBFb
HmjHgUr3Ngi/GSKWdoWQEIgVB13rOv9dfN1bWq5EFrpJIwgrzmTXiD/x6VeNQ6oN/heIoU+hH87r
hoLvOECUlvwcxBKLcmV7Jl7fiNVPKstCi3rTF6jF3AA0rZEZ8ExPs8I3NFvQ3Lz43b9/AvFTA+55
5gXFGJOZjrlKB6kxM8Wr8cNvnWJwoOiSfq54wowfO5oELH6fQ4QXSnsI7le1AoNJY3vdrbLbdS5S
M1zL4UBymKUvN8pArLyo5opsxLLmIxTb1utouIpYN4qIAP1StGqujWNuC2l5ytRL8bApOpt6SzCZ
DbsUZfvPs3cgtJvmBJfg813+I5yvHvBj4JtSXZy4HCabJnDixiKx0d5ihH9PDEWMMExaKd7lq95F
HjGxcgurDi0+thgoAmcHw4bKOGpL91wlgOXSi6VSetZmPUn8lrgQsYtFsju3xzg2ME3sy1Pvm76S
9TZdwJNjr7Uxmi46RtmhsJODf/BPX1ZQbSE2AoYn/RzxvG1FOCFU19CSa3ccsuVr8jTD59FWqV4b
Z9C7yD0I35ppLex2mkLcOLdopFux+r16ap+SwhCfeT77EUT5lZIhrJ/mgXcupM7eBwdsXyP0NKsM
4A5t0D94sy7DAS5OCMwCSiC3sHAOF6gyQpIUaqvkZnJFpAgZTPKs7duJS2cFEgpekYZWOYOrOgSN
Cfugu/Sfp6WG1+OmGXgJA7UxX9GrYfkePUkB+G6EpY7kMzgRtwk4yWpIjCVfWTN+uBG0XoSPl14p
hNQRw9uejHCSvgqjvV5Q+6nxX1V1atge1z1LXj00JyI0wedsR3tOrmRJuQe5K7CFzKG3NcaO6kGH
l5PQuRuNa6EuAlvhKbCU0Tsq6IUEvyExLJPwKeB75n5qkR7p30dXbR0xZK/PmFd5iGXx5f9D542f
pMRhIZ++HpCvZMEfH1JkMv0Deqm084YLGUUKurBB9BrrFo+kqgHAXqIvJLzEOsclJkKkB0hg/UAF
F8YqLEmwv8z8U4s6yl5ZaL/lxuNXRZCDD/7iDjgs3RE6vU0z2rkjp1F5ows/9hXlWpcTN9kXhhm8
qBjUO/em9IxC2KdtMFWUs0Gk6XO3vVycYUzzN3ncmU5eQ66Aqi/4zyL/JW6RAsypFGmLRnqmshkD
mN244at8hUynS7891D+l4yKPBX+ROGv2nhfox23GzId7bMTXF1ZH3prpOUY6e6DPuHm2vnQnhr29
YkvCNFPVG7+9z/AmPq8TVUgUO5q30jigukMqJM8gX9cxbz9C78wVNDGduMsZtotrtH0VgHAUgKUv
RhGhO9LBQJ03VPBQnGzSgkPKpX/RS/RfEabJLE2h7ddgzEt81Evs4QFA3KBCq32MmSv6+0I1mmCM
l0oU6e2v7U3nRlU+UymjdDFvNNK88/NiGqu8l6qF2ysWzwDGS9Bh+MXH4jZ48paZvdRA0q+uD/ff
XcIJeyw8Jza6cDRo4BSx1oI7M3UVDxMMn9BT9d3k6Zi192sKknUoTCKoCr0RnszyzvtI6U5PvEpo
Da9LProZqj4dWgf2pg5Z0de8YR8agMq2W+8kwh/SY9t2OprSZMmvO4xEzTNQL4FoVStgcGeEp7jQ
svDnVyw4tTO97CMIQ3euGF4Wc+MbR6ZBDZxU/r8OgO41CrQ7MYVWBSwQfsqJ+a8U8shHnDT6Lb4a
/rrfr6GL9fvTnJSBw4ROT/yFjIqTWbXxCYZfCa1CdRuBayu0g8C8UTMt1CFb3t0ZTeYQfiD8LPCT
Cvw1TZ7+JgbfNP7C9BYEWO7w4ngXvu7JGO7+aY5pTHJzdDWcNe4LMj6FB+tUwoUM4JQsPapS1yQF
wxUZsPgOdYt3ff2TQcs6DWW1Ys6GNtD39JjWu4lORFtsBvX5PTr21R2tGL4wBtRwWMAIYiM6smvg
4xMYEM1dtz4yhjyfG7ivuxDAVnEqXc9S82aN77T2iMJ3KhZKc08teuU78Cn0VXeqPYeEMWoVeF1R
2jsW3KXVFqlKs6tlPWfJoZP2mwK509UpsGGDEQxcqcC5R6EGHGDdQPGtjywJwRAeicUqqELvt2jt
+3zbGEo8F1+DFsz/41+oxiLpp0cgOUGksUj87dolwkNR67uPd3TNicZEatngNvcRPKdtKYmO7cSp
gK+lrXQWvzrw3FW339AxNcs/z+c66zWprrEAKfjvQiMK2Y1Yfw6xALAExB0wTYc1IODM+EkK7hu2
0UEQedbtcf/lpDkSzzyIJqmCFFxa/CtkC248ns5x4gMsrmttRqqRoXDCIctvI4elVvCVrqAnLCI9
Hr8EgV4SWQxS7uKWjvIqWHXbCaK4f9DNJnU0QnmoHIBM6jxy1PevC6BD0cqApAgkR8AKEvGn0/EK
3f0O/etHDXo8OE7nPCgrxHO9mPmk/ee5HlsjfivW0f10w+m77QMzaNaCREycHJhN/cJKQFsJiFy0
SMDVBJn4ASlxnyLprf0Mj2iF2GHxroL2GfUV/eOvdus6JUkdJUPL5+NGhNw/JbLY6owYGbNYLbK4
f3dQ0/HdKofBfD7RKHphpErCuld9S8DiYhmars07rDO10zuPQ8JCmqLpgGkJ6LEgSQAmAlG1pZfm
8WMP16+7+YQbgVOS1WtNNTw/j2RwWQO1HLnReuQ60BaATXX3J5v6hXeQycuuKv2qWeYWJjJsd0RA
3GulTpXLsNcbCd6DI/U1dXNJmmgv3Bve5WcEtxbXx7XXjjcDAupde5odeCG/Z07Sphmb7lGrR0I+
EUOVXi1iuAL8S2G9DOK1AlZR2TecuEZ5XY/clNnmOxajabWdut2DAiGXPWNJgNnxbe/2Bvr3rWhR
H+X8VpRGUFYJNjL9GzPY4MIAdeYHtqRxmasmzqbygAaY2CJlIZllPPBz36oY7VmufW2Hb/Uj4r/f
QKvOwdNRfTFHjZF5Kx8s5xDa3rl84M/RXnLew4vbfKpCqxd5EAIR89gGrWRAJzsI0F3iYTXjvDkZ
4MFnR/37nGLnA5IJXxckWSYZEa4g/ZIHZSoLatgHElc5cZCWE5UlEayd7VT6cKuPm5kosn11Fsjp
89w+Q/pEu4fMiLGqtWAAGxo0J2ZhtD4oXz3XgPSM0pME5uvWJVGtRJuzFFNRYi96gaF1uEeCZNU+
G8llWZ8ucD4SVVIo+kMlKxj4h0US2biE5Pja9zN3QPtIJzkmgdRb9rQ0S2JM2rFW5gRd0dAu1PMm
3lwRfkmw5ghTcQLhx3ihaEV+HeFUmhmGW2+RATMVKpHsVCFSQEajm+FmPUlvE0Wi+wPf91JdVq/y
H5Zx52VRiOnyWC5+3SmzVrgsveX81jneSZm6tMZX//KHk1Ugk7Q6KFYJMpZe3mMgPgRcxBYhuIse
/G9gpvTb+5iNpBdwKVuI3z+PZYk2GiKw05KGsiIRMdZazFWW3BBqwwGk0+5aCiZ8dxXlQmPx/kbj
inDyLuQn+hA7wACne6eaEg4cwqVcciXcgWbve89BCFbKiJidnLEIrjocDEjZxq505Nof8FNo9i3x
nDK1Dq/mbQhoC7oyhvmDikBDRvshZAp0qXiutqwU4j7d49w0pTV9raMsyQXfywKXNsb8M/OUx8jc
F/lz0CycWM1TeBfiKoXxPX8YbJVlYGbd6XZ5J67EeiBAAtQG8xIlCADAFYlyEYXqbVEXa4WL3cVA
578FziMBLM6Koh8GALB7TFX9NYUyFx5LYT671Qb9/+uPLQ5LoFoSDBivMENfNCwwlv5huShO7Ris
mujIx1fNKvDv+e/Y/vo+D4vck5w2V9r3MvEMfcNEiMolyka/V2PgK1ajIhD/FRRuwRRnGe69dr14
OhL3ShI71SSGvPV0Vf3UBlJStdfttTUFbFPaNg/adpOImWMrlnMLedhNY+aZkbMf1BeFgYuQpSVr
pckY01puFlGZsx/SSk27nTakpwYD0jZlO0wmsTq3MgMbvf1pVltfIlZFvhABs6FX35U1LyBEYm7a
RIlbRlkXZug49AFW9v1YjUKlLDkPdHfTLpaiBysJMs0iF66ESeifIJOoiHQWRujZkgfpgkd4AdoB
Gc73tC832MDGX2B79eCcQB2cdgHROfhIzLFY6d6x0PeTDwdmYsLKGE0o+7mYMJcQGNfv4GU9IMJq
MRTxSmUeNcT5ZsG9vrAHn7ItTU955hmy4Na+JZYmt10vYMxPiSH/sx/0iLFOOCsPIz765IEJSbsE
7CVUQGvmE1QZWiKBGtfBxYPJY4dwDnXNP5y4KjX0pakxFqbOQkL6vsed6E+/zjKf9iosnRmfO7xz
+dx8G7Kb1aOTyDnRso7PY0q2yL8Wq0KiQpme8DdVTZBOQAVnbHdXklcoaXl9IFx4RIqXduZ6xdKT
RmFaFN16RMmtC50KtO8dW4n4P4ngCd6pQkSpnPirRUBEpwmn/ofmdh+Mk1Rm1fFg+UqXQ2xhae0O
UId4nBFU4y8Xtrk8bnB+gCZiwBnlGlCmy8DCGRVCxejoDzP/95P9eu7KYVpB3yzLf3PZpaiBkytb
59QuYJYUTfDwYUjWd6n5Xu8+WoVTQjzZNyFp54mPQDcF/lFjxJA8RRR6ltXAs98LntdIDRm1u8ZR
7mR9kr+bxgqmlgFmWFPpHAUrBukr3dgodUgWn2IFxf5qDCcvkfTXC39qAtHmNGAqmG+7bEyPAQ8u
D2pKSbpn9jLFe0yNEO67gEnsYdDvt9ijBib3wTJZhddfeQEf8f+yWkFCvH+M6ciEwAoKJbMqrHCU
fRkJYOK9yqnjlt9kjR/AgkidPcFvk4OQZPlWnGuccZHZ2UhgclEzSRO4DT99CvDu0dsv+S+8jces
mkrdSyxm5IBgsM8mIe+Y8YmYHTbiXjA2cZWcAY6pZoxgn3pGWE5Ts6sTmBtnIsG6HgKf+R4OpQxM
ChL3FV0R4Y8QYZpQXby685grnCtvUiMrc9ml+sizAV+nCwjutO4H73kppWPxUNaTSAvwPSc3l+hu
arHzI0L5dCEwIqo0FPCsFIi3s84L67t0XFAHBd4Gn+IXoRL9dlJWH6xl349udG/b5NutnCaahlG9
axkugCGLniX1k+vRrXQt9unB3Cutq7Z1N0I9dHAdLhbIHSxFRxgtPg8Kwaa5odvO8CeoJ2Lp7cCS
STLLI6i3o1IfHwAtOLGFNeD6/s9PrE0eTj3ABcgPH2QrPVIXMma7I36fSpu4/swRWlgs6qHymYEn
T2WV8pJvuKQR8oZYMWhZAK5EfsMWdeVjq0j+F0I9L+dGWJZ6tP+icecx6CZ33EWfOsZzZ/1Xn94G
ofpLXLobYdSabqfWTZ4hwglg22iZlRlmiw9/v5Ct0HLOO3zQed2DYSF2CjwzmFzBcoSvV7kt0Nol
b2WPaqDLZFj7MOY6rAhX/KYxowbcYfhW5bsQrgpSvMkUWDIntxYhxxVtMsHGEgg/sBepRm814KYL
Tnz8UHxMhcWpBe4XrIuys7o30g9h0rDHkcBIrQbsFe2CihFt2nsv+pH/7VHtH5W/jK5w48n/fLis
o3IecOfP6j0UAMu1V1DkkJnaQ773zeBZ30NCVlHpeVN1WStguWcuN2+VBBgrlwB00wfmT0IIpIsn
lPvZD9oHDbN8JnzxHHgHGe8TzcstZAqzH0PI0BJcSgRRn/Mt2+3CLo7cc6vcudPpL4UiRgTsBqCu
ZMaD7WTDIe6bhFaHfQDdYikkC9Q2/Rln/fDwl+FwOC8GssMZ0uaAbmwS6iX85lHh7MaIVeFb4PH1
XSCwsB7SD5FKgfYKeihwRMM+qzkeT2Ju2HroglXIB96MyTuDeYlHMTy+V//7CV8+Wh2hoVy98iCg
RoNO/I3PI1KgAxI9HXywjtWq7+srlmZM3L5i4oGv6nXwCk0Elp3RugSF6nIZXqG5wnPlrhn8KF7A
T2cb1sWEobyii+A3oqXHjBswXN5xcCZBXZVIShkNMpR+NYiFRDQIKnPCRD1RBp4WbBLyrpQzjwZp
sjvHzHQcgY2YfVVKARP/RKEW0OUChjuf9QNuvy6B/J5m8v7FMLQuhcJVl2cjD6Wu3QgGnV4RwVBE
9+sMyJKtUwaIP7aOfRHM/KeIhhfUTgs8fOoKTjm6/FFcTO5/+iYV9vFUBB1VMo+S+AYaCD02woiL
JKuwlybK2uvRds4qQNbc0VjiK0krzOJvUGrqiZ/8/0shuCwdyZn2TTZ0hjjJg6YSTpsO5GYKt+2X
E/7BothBF3YIhgAqIueFqFANU+THT4Regi7BLhDRJcA7bX1GKw0NLENIlN7VlQjtm9SpYNsw+eqC
gmqLQ8qsyUfMPGS6rHtiKNMseNUE9bVgxjBa9OVrHU41LoxZpf3yfqxj6lyQ149nrF6JCo2F2iST
CRXkCJqyNLh74bc0FCmZr9aIMecWaOsocw4L123M2jQcMnfYJ6CcTDGBPU01xlvlxv0mXEwKFAxe
Z2asHE3YX5BtFdZPpAhFY4iVywb7hx1Z2hS5CjBSPkEheX0usqsaxQGvr1tYL4+M3hE6wQewdrGd
YQbWzbMaf6ysYFpUsDzm4GUD0zN11E8P3LRYISXkGEG3ljntq+WkPnkU2p/as+6dTdgcUmJPUW3C
HZL9MuwGbtjL18LMxAdhsYVbhS5tPpi7CXfMMfDw4AanpIdmYlPB7EQ4zuyeGTEBVTziIs/P97vD
emhP1/LLm22AvzXsGEpIk7IsqfcI58zBov4sl0rsHn1Yx8TS5cGoO3SEZWnrXW1Nu6pQ7+eHBj6W
fKLI92ss2UOqfyujdTJmN6QmIN1n1WxBXpJRc6Ow6HNnM3aSAbTu7Wb02W9on2+sGdAxEbhUvSww
1H+mBDo1lTu6W42kJnbEglMiVC4M+vYl8g7fYw0SfOBww74bwfeqhKWDHzln1kyUKEASK33iio63
k3bMe0Xi2iq30e0p3OUaPNbrYI44liVVXbtArs1SR7llEmV088BxWddfkDhYpd39XnV3BEdDsqye
ZTHRL7lc7NLkdmfCw2TyUBrsRlGPnSDjruxyaBCnOBH1RE2iW7V5dZd0VThmKn+KaOa5GWu+ESvf
AkOy1c9hm/OpKIR5VgGnpowehkMz0eQH+B+MskRe+2D/5pP5k9yTTNI7FO3T5BGpmylwc0R0NeCc
QZ/lbkWMe7AX3G9TKlP7kcFxAp6HOR1bsi6ViYYKO9ljF/B1vt5x2c5RIiFjFsf5rwPH8Ct6PaNt
TVNFgpSxoCzXYlegdiVf7CmJ4aQBQI97cLWSVam50wCj8uAv2FhjQQGODj5OnUsRawZMVbMCU+b6
ly6/a0yNbnv3217F+AybUIZfm62rDGP8pStoPAGwIi4+7pePuNRWalXBPLnWl2l/hOJJXe3Vfm1S
pZSARzVuXreGSnbqraY91PH0D9ievKC/XXa9AWHI08En612jzov6QzAaVYDmRP0gMe/SAjTk5ypu
Mt55Q7za3BvAzvmeX7aCa/a3DtU9T38JOtszuIkS21QnXfGmWiYCgufA5ay8PPC5JWmjMMfrNOVu
DgOl29g30c2j1idD2GNhzsukOebpV5OwoGUHDQQAncQmuhB0gyR30x9K5Tw+w75aFFxINx7a+bH5
C/IzAwvJusmnUylFpDbINZOWSNyj8MZTUlwwdzIMi5V5g8dZLrC1ajIdvWjQYJQp97HQHEuc9htK
WT+2pKATB2XJw+uNTDnA33cTuo1ryPcyYFAzvv5rJImOx+BF3++M2N9CMP66kHj4o7OU/3NTi24n
DL9FRx7teXLZ72JZesVEppbtJNqlHTlrWOO3VJ9SnDw6ccJJegDQjZvb+59YulmxFSVQSiTuOGOk
5JyO39CnI6L/1vs7LcmBuSf3Ixx8b/MYwPwuGHwj+AgbCpB2IRnHTPibVIzWXDK5hbx0yIFPxkAf
kR2SMPn7Om1yUmdBnfmEYtYVQLxlTG7x/SJblgV9nnl6MR4L4U0aIDqJNP49QOSFTr+itK0atstA
ULqdvV2T5ZgPnNALQmgY1T8PImEc86MMZ/4g2PEbjxNnplTDdn/7UIcSQpJIus9kAiW0y3bnkhpV
T575ZHzmVDDZ7uU7Kt+78vAc2awtG9mVA9xslkCj9h0BFKp5xvsvkfhrdu8SY7uWR3lcec4uuCVC
FpejFqEN8QZtiSkEvXFZ0D++JBimCn5LdKjcr2rCFnBvg0zUc1BOpR6BH3LWv8xgPfomdKipErka
EhcDTnMV54CHlC4GmABHquz4osoBTvwTFQpvXofdDqkTo3+rqxjlfquBYp1k1yaia1u9F0COF9rx
J2mvr2atbNKY+sjn0hb7rz1SUc5Sri/WDCGu1r8LP83/VSBiBmh+vWYlc49lXrFINPoBVuy4Fs8M
MbH+vhCFsTnfIeBClPokvmDSvRbsa3UJuP6trWsr8J7hHIT68UAnvoXlcxGfp9AHRflMSecmG5zm
8rfTTT1rRzawaSPF0Pir27FQltCN8iRIl28r/1Ujy4hUYmImGydZ9yUhf+dPPol2AU/lzLox/yKd
P4tUecZ3OwrJwqVl7kNxYmk68uAQJyezAvqsAKwZHbN2dG6W42I/9cRHWV9UQ5AToeJYc8rZsCSP
ozSxRtEWyr6qKOZXoF7/IfBPEIUZIahrzF7mRMM8IeQJEoCpfE30nWgghslh4bjx5//50SA6A/4j
7eD2OPH5UCjyiplKOF7eqiTk0NpxUmQjS4UNVfLgmm90boqj+ZIpmpDfPJ9S3HazFKSaJTC5/Sop
wAh6bmTIyPU1vXowE1kIawKgkFqHfzElDSJqOIZGW2JNjCvfzO/urd6T1EdB/KW+7X/N1YpPSwFd
o55wl+ZPq/C2cI72ljS7Cd1MI4+RTKn4s1v8qGmFk1UiMDSHIC/1UZSdA3QN/XjO5LPqtGztt1FH
NIOGFho0GlXHG1kb2IF8XZVsFe00LChn8cWWIh6Whiq2lE4gd0eChXEoIcUEaSq4ygqJ47jElo7k
KLca1ZmiHWP4OS5tMkYIImOdHmOdnKNdVLXLHB/8JarQBzDrao8WILH43WxsIscQVufGTX3/BwCV
w6RCVofZgXn+FXDJT0yIpBftvop8JtHklS+X8hbpr65rQ6Rtpvsl3QiwIRjPY7CfkBUCPHJ+2A1k
TCObslT5SGOwG9UoUIiETijWfV/SR6AmyRulrVvcg/sgeAfNtiQZrvFoqkFWWA5DYyO6YAVe3DIS
J6MihN48cZ1RDQDMZrwYJpwHvRCh8cELCoEPsWRiYBKJ2/N2p2KIST4U1TrNTytigWRkmgnk8Zr8
ynQo937QnCeiLzEnPQDnZyEc+jQUq2V/PxALDTKKBJ+k6iz5MOgsWabrYvpXCMsT3feH9jHEVYEy
qsXvYHxFEogCoB7jUmHr8CkixBQS3m1cwX8063Xr3Hze8VuSVu3gy7BWdulkGBFA3/KppvtiuY7a
1dlp3GIDly9dZ20u289k5e5t+Ohve9Kpw2Ioe3OP01HCbage95HQiHBbTce6SAXL606CRW8Zl2rP
lRrDopbVWRJ2TGCFESwSKVPswLb4N1EinCQsLy7sd6lo8WOIaU+v+3/uH8eTwZuoNSBvqtr0jRjm
bvB2KKrORv/iUfLNmBCQPcqC63wKZhUVuusVepAkCH06dvtPaZLomL37aPP1mZOxTQHQqnkk+IXe
NIOOPTjUo1mIwRXSpPku8Z6RJIrcGJ4oQ5KIcr4cBlEK7T3ffGcbnCqEwhibwpu0lIfy2MdqmwBH
cq3ypD40NVBk4Y6z6wvZH6ETJEGDUKxccYCN9NnCvnQPbR1vesNnUBMWbnLr81askqAEOaBQsbsK
FaZ/g6U0wifvjPyv0VV9cwdIECAQrVOxo9t90fRe9lWqCAPIdBwYfc2NcMCkVSSW1QvlS5PvF4GF
dKE7zya91wa8W7CBbIERvmS0IObruykAVsbdNu+ikMtejn4pypp0MABsAJlMZqrjFcAFzS32lcTm
5MObGZwyl55Zyf3wVWkpkgOt/DbnrcnJa03k7j8NYGt6nWE34Fkhi6QaE95vgVr4HaWSRKWgFNZj
KTQaPPq+OXR+TTTDBDGJxY5NW4rsvj96DYvGU389sfC53HldKIHfEVwamRa75WZwgfo1TbGyW5f1
mvlLAKdzCkRfEwn1x2Z1k0cVqbrtrYMa3ucPnO0irM+7H3hwWCUGTYwI9OY15oKesjmstUNW3RYV
+aCjTnXaZdyvvCLu44z/zIa82VYEfDihOVhjnczVQWAUSH28oBtOD3fyablrhTAOYmTZ5YmbaKHa
uITk5tVvsCQ6zhL3YvA5UbYIsCTY7YYOsNkGR1rFYFaEKZghDlXc2uA9exiLEuXmxbcR3TQ2Ku4M
aqDJP5CPFwmn7OSdjQr/NLwz/UUKAouy2CfIdtoev2vJHhd+mq5AcrHxNzf/BAJM5l9G0OUQzWOt
aIAxi/HZFyTJOA/T07z4bUbsv68SSFXSnCbqSl5DmmevYBOvqincydgQwZoJK/Oe7q5hMpR2KCk1
l8Q+5k8NCDDvx5phqA9BjZ/PJ310fF5nUSRUYGtn0nWeDRkyoN3XB4si5sx7yxvtSCbSGN6IWLUs
AGSmzoHr2y8G6I7eU5roGlMVh9CA7OLb4UBrFzl7pcn/FjDg/WUxqm/8/n8vp3PdfQn/zR7scptR
LgkEH3GSzyoPCLqpXJ4ApW1VxmnYv/DPzUANWw8xuR6TWeCnzmPsRXy0bZxWFoTrRHpmr1TV22xf
rCKvGvUcFN9Z0ulSmTmvEImKrmFZj1nkSV1982yx8nmj56MImuC2MhxyK+iIqwiYVFvR8PlLeSlz
VmGCu5nQjDO9hVRt49fpleUlc6Ag36Tm8Vz2KBh1ogBRL4OurCdmS//jo6hQ8aHy+ByunRfDa1SC
I9P2LyyG7q1tZoVMGHP8FuSYb0ETp6euKFD7RmwTyBPo4H/JZUYJWG/q/Ygf6Bm3WVGffB+5nxT9
XIZ87CEoUuwfhzfreFla7AoSiT3DQVX+JjWwjeO/XYYlRWsLIanF3Aj7u+4yByL/rvyk3s49LPpi
C4kEf/PVuD4ZuNaFP7g538/+XJGqB6gvuW/siST26ddD7kxUAuNthx7zGhsV3IjS3wegJMnnvtb4
48ZloIn+/TfCvQLEHd0PtxNeXww1jEKB+OgtMKCSnjwy9LaCwBy+LT5iSs87r5ox1PC3oaNGlKgF
Qe5wehToCWNxnLYwE6vftKCZq9Gud0RiYH3bQEnHUf8eh2AfrdyJZJ2UG3nbfObRSeGk9aGu2V0S
N9AFSbEi7oFceAHEQUMc7I2UgLuXMr8nPmoAHvxnP9KLLSJY39kuESu3iAe+lpidmFd8ztrdIrCM
XrzZM7Qav8TTU6Rd2LuNAH9BOAkwuHwLGAO2PF7WAv258IqL5eYSfgPE1dJdHgFAdrEaECkV1xsp
JE+6E/4nsjpHMsu8r0yeEhDWap5oJcNpvZGZ4jLUDOJDydw11QFArlqfZ3rse68AngzTlWZMN7CU
Zi8l/VyZiBzHpfGXUg9sppokAcGHyrf93OXi6xNDmhXq8/XjOxy8SIhPNVA9oVEBBMdRY0SuAdZs
ADCXCcI5RUUa+ZTi5dYMzQ0IFsQxD/2EFxro0wxJtSBmg3XHQGKyvsL/PIKbJkkuqKIyv3ykSCv0
pICecEEJusECvzcktf1VEt1HeS0HMgMsL/GXktEXdHGmsYg3jBoG09mF3oB4C8eACRdaoeMbUE4k
4Lgqg9ST18bvYj8Dii2Z16OhY8oftEpDcYBQjljntOoq/vsnGIv/KCzu5r8z0FwhQUt+3bmLAkQT
MYdemYWGRg78Cbx1GJquEG4LIklg2gWWO5len6RqXJuVoscMFd4vR3ev1d2YUITvkiRjqaoHx4ZG
yvvu/X4vkuQwF84MK047CigtfIgtGvszU00l5yvWYX/dWXAFhkAKQlQyqvpsjoC3e4EM/7hiCM+B
wlkP64yGdnB1o6qY1ju15dgFfWPY9GIzQ/Vh03Zi9s59oycSwv7/I/pqlgiXJDHhiKr+6JMlf+ZV
0CJtzBehdIsYRIWMrruCCW7/x4kXop7KvKZxNutHcvcT0cTYFftJyG9w9qsCPFNxREkS1QtutBqy
s04BR8ns+pL85dwQ0TMiPGz4V+eMURKUDzNnFdrMXKLW+J2PSDA2QosROHJk9aOsIfmdWP8NDFDa
ztDUDK+beq6kxJKstB9LZiovN3rYKajCf8xon8aOOSoifW6HvSQKVlpEYK0jso123UV37AEgmv3k
1KQZAcKgixiMT5p4bub6aOnjoN7z5WEIsP7PHi/YjIBXX+7AW8L97l6YCvi638LvuIBADbThD0At
lvS/Yt/d/geZ0Kk6kB8qeM2SebstDdu6w9yOXOXl8ex016XlyOeaMf6wsJiNlkMzghGIXjLqZprU
SN1UAta1GZjgqkcUx+X2hStcxgSl4dSZljDI6EK/2clGKs1Jotw0fkVLKp1DiGROLDLLVJvotazf
V1QSuzDYtRId/UViZ5q2mqhWR9eODPN37jWjIsmcbGOkirNWIfOfoCLeFOqPRRlo8GkPymBBOoiR
tQD2EWJhDQmlngOG72Gg39099hG9LHBjtVQbf85afa20RPV001Pdo+bzOkhxbGRI4f9/D6auZdZY
KnWLs8U/3+KeNhgLsQdGHUB6Fum55Zci+F5Q8DrCkRD5Uvro69LDloz6HelND4L2vt2GWW6rL/wH
6jDt/+lZSlBVXoliLu0QNh7dGxhPtm6zOophCAKPg3GLWDaHnyAVP94zLrDIojYx8MNn6xXDRjg9
43xKQ/Oi81TUT0wPV9smyYN89HKQ0ZEKglJsroh8WrU3FBj2I+PwkLpURqdcmZ3SnJXW5t+7GfuB
piwXd1F+sktOvonFLgFwfizI/HXKJKOXm+ceuGMY14EEw0k/XTby8ynd9zoBf+FmNbKmtqw4SaGR
jRiUL0zooK1eXWCxwz36hjxlgNTh32KOOYDDdxF7F3TrFO7RDLV0FVlL0PzN0LNajyicAucRMT1z
ew9HvLej57i/ccwBAcPGJNWd1+QVnnlm6ONjPpKDrAesuzzw8Q4CDrG0sUxU9Awifzt9w8zgolRc
CwL6VFOQ352lfdKTrVMPQ9BqPs6cPNS59XRbsy28fFCVCDmSZV6fMeTkPzn6oj6uU3qc8g7Di3Sf
ZAMy+qGvUKXX2wfgnzvyExOJJvcmbqmDPqy5FvIQ1RwIN36Q7+H+5RwK/EMXxFcPYVkdLSjPf6Db
N0ZwY9hwHqIN7MaYoj4i/Y1XoCH3FSkRTsM7vpoIUAdSNw21TebqM1OrswPr3Hu7enzsprxb51GT
G88ibfK2mhubkkZQTUgMJXjrPhrYKOmHLEAxwHkJCUXbsxRoA6GQgGfEX1xq1EXPt4nftO4SKZ2Z
L/SLXptSAACGVP5GQSOeNtxUNBspyhnweSBpY1tCs4mcUzjtc9A2qCI/w/vb/ofc2Q4m7PuexbWd
Vz1IVKdaFJ8h1afe31VacQe/Uz7igVbubGlLvs2N0npm1MEsvvFL8qzfmVVyxmYTycDuiHbs0P8b
HPFVcdFFMV+1E5IXWUO+YbDXItOZWXVqs/1KRaX0kJcFr59LyrDVN1MYD0Ww5s1m9J2w5Lko/SuR
HlK5Jg8oAL8lzdKn0aN8hvmdznAMJiD0oWzFkeWFDfXLOTgUIEwrH5ZkkRxpsWEkK8QF3zNq9lAK
YNfZtTL/iVEV/nH0Ks3e94sFfyNKdXKaBcETxU3U6q0pG6kMC+b++T2gMdh65GQ0rwWA0gEKXkFA
siimwkxGGhdCKnwvjS1PdV4wKkPveRQT9d2ks2AQLPYeig8ZkmrFseXlUFcT97HGiTKpqDidxOCt
lft4W+8ILldtlL84jFbBNEmgCvXDbkP1mpvIhOLuBXPAmgLRrP7AjQZJeRUmKDvqz+kGrEsjDIRt
THLYbbWHIA97qiidf/gf52Aqs1tW1EeyUDD0mJu8fwXPEHpf5Ap0LzkkJbs/DvYt9gfwDu8+2nSb
ZXvGadG0rWySRBkxtu0ICdds4lvOZIZ0FowIwQSriiMh530+x7XdVxa0NHmVTRXogsziry6h0avN
mvJAZBXRvQlB8JDrTB1axyb4hESVADeLQ5JYk2oX5/yhDcejNTUZoTlc/sc9zaZrbdPUKwbTiEYL
+GoNmNXjZNg6bqFWdA4NN//m9eFX4mSK2uzFiuHR4BFNgzGf+0cVRE20svqURpfkr8FKGr/MZUIT
ytVzeIllJhtEh0fLYvvcjNVmeuNLk07TkgckGZH9WRjNgru6IHFxsqyfqUcnLa9qcBa6Tf31X9mS
ehS4rk0fJkPednzBR0rkzrtyvdrQE6QLXdDLz7sIPfAJIk07quXdfAqu2TkmnG5SFTAjRrC3QeU5
99U5MmbH0HpSqq8vxWx2Ra8WH3kB+zhCW0C8suh3xgslatxq8+oa8xt2c2Zh7uhvSyONq+dbF8ia
jglDYRAb6F6SNgzESCuLqvu4qk6OLnO4xvFVkEFKaz4HO565FzZFiMdvg98Pt9zCz1ZoKNkUyKBL
M7uMk68p5juB2rwc0VQtMLK1Xkwe9B5Hp4nrYpQT/JUkeObSWatLG9FiQl/TVUFVVxAOiE0J5NXd
cjxOco4MtwQcvwLsAE55UWR1QiBZ8R3AVowX/MIhRuNPLDPSPYq5MK1TGfDiDg5G38y3BTrVblmZ
i/ZNyEvhFbzVz0h84QzDoD6hsxTEG5GIzB48HrlDLNfNZ6n7VQ0tgpuyR++Lton0FOpEMgs3Wngu
BqYv9sExHo0RBt4i0HFZMMUTqKkiP2SjNhOt8PJ5x9cFRjUTlinCid5Jxq6FVpcW9sQGTpWB0Doj
jQpkVjcNOwyE+f6TkT0zdnrqNo5N129RqYi1EK83EQJEQMKKe6ONVbpLePNiILP9VHd1aLNyPBZU
nJHP6etOXcC6ZijO0E/flwsbJGHnIh6Lf/LOmTi7jv7M5VVncH8YJoe4AFGaCTnCSoXwwwlXp+qq
W3xXtPjS/dfvk8SlpqeqWkMbGQvRiBrRwPkpDyBfljLtyyNmuniJIg27SfAib9jcYRJoAblHdUld
lzLA7X1Og9wRa9B0lZqbolRVVKBwjH2YkMV/nygLyVKNC/QQUO6h21DBwHpBMtw2S27zb7xJcCJN
9azdj5SUv6X3/3wB6IVjY3B5Mjl7cCbIxwdMmjB3AJeLX/xbttW3TwhMwi0so01BAQQaWE+Go9Rn
MOzitIyJJTPNBjTHOhwqxf/FCydPpGsyxcDuBtMeCIXaBPWXOHFuc9EDfCFvOSKRwfbGr3QB0C/x
2WHC1ONGA5VR2TH1JkXXYmgSK2/iRCoDc29lkeC0DHidycrHsxEKnxRXDYa5ROruSM7jeysUdWcu
Jx7IlLV3k7Kjt3vsUyTqspt0BQxjBZbsnPqKdTlu4YhEfeV3w92dTBZKrsjPfEOqBLXcmvg89+qz
oUo5KtEtwvXHLDNl8Oyz5jmJ8tjxm33Dvusrxth0gyekjIzRNulDN6rNV+fipfIfLXeScxsWkjRX
GOAZekTejRCYzlwiJBlr46plpyEkaNza70Ajlt26d5M4wniDkxBpxVRfDE2MNfDOL9rLUyubHzop
oTGDE4rHGWdoyYbocQO+cVV5gaBe/KKMFNxXn/ESk1VdFnPnyGJy+dkgTw2WS5zFZ36wA5P8hCjK
GpGn2CDCGSlonWHOp4yHwo9864px7dMcuhdaIpXnTcx6EYul9wEw00fu0MO1CyWuNM50j47ipZmm
ZM5RZWXtRDAHBG61s5sm2v2E8u5EM4oYvKsI9SKZiQO3yCQXr90RwGbFES/HvjR3JZDkjNXx0UU5
5xXHOiXnKtJa5pQQwaHvSgxosu5rTALm2R2B/snuLCxDM7iayxL4tE+rli92h8R65m9DWRrv7raL
kNnQCtvq552xkkeRMBrGxgdtjZLqkvSRMkghXkCtcTulgBNi/qsCjFao0N/0hDTFa4xhZfYZdgIE
cit9fYeG2LDRh5NGyg9Ad5boAGUoGba4nqRmI6K5GS8nVepB0MffUS9tFzMtPMhXGyHr4OgTF7or
2O0lHT6LMy8kYfA0HubiNSfGBhW5RBexofUiXkDsuMfAouxU3M6QUzXQOm/E8OAn9i0B0deKM18u
XyrjEvt40hqOPgXjsHhbEATmMKSy0BuUYL189SWnAMnn7wOzQ06H3TyV2WwyUBQ5iL4fhl2m4tPm
XCwTvTDOL0zeCxDDPR7JJguTeVmV3JEF7okfSsvsHQE/Xv1zxB5TEPaSbbVry8W9sHftnWapLY+b
dx1O94m6POBCaykalj46L/rV0OBWRD5E0xVS9O8rkox4WZlGVO6aLz+twXzG0Tyf4yLWGXlEb5fP
Jyf1tpCU5JWi2Qb0PSNlonaZcTIyCei7lxbVsYFU6Fra+QMflsTxpj6J83C5VWLRg6r6PLnYJ3/g
8lJSP1BqQjLWFqTh+rw0OW/qqAWybxtFxin/4MTm02El/JF+5pw0Kcl12lsSnAr8V3L4MVG8+POJ
XbJ7vbqOsKUj3u0A/tACpNYvZv8Wie90lQuHegXiwWiWuBEa68CiY9wZ3XMmxmMZ/7KcSoj03A6m
gt1CcWx4jJQMgsuS6sxBVEfdl2yR8xsnnD5dmvWhnS9Nf20W4e0RbpXL7QeRYSo9M1LE2Ukyv9JY
QjYo0z+QlOmpmSsV2rULFQlyfWqc6msO3aa77g53p6WGUbDB+MMAi105zu/Erc00D3If1GwLj0/d
7QjzT/uSgstzXdkEirk5wFxanHm8jVKs6d2iUsdHeAaYZ2ZB7+a7OF6K0gtMI49O2+DTMSTTVHhf
wUZI6U6ZwZ5PsnoPII7N15/b/4Nz/ZymmIWlIDh1VRSQN3OLtdsWZdKLBbmfGo9DwqE/bSeuSUW/
+qEIxspBuYdGcAdxPqLIxUqvCty1Q24b1234S5DY1dsGMLgycUROm9c9y05DjtlMA+RRYD5/1/fi
vaaS5jszzK+kmGahkdJedfAJmdYgYX10O7rv5Q8NTdcK2wOSQI3Rc4nJAah89jbIf4SS+Pl4adFY
JRJvs2K91kUDz2FOtR1EiXXfUa1z2jFtJbjWmgXHjoivV6KhqNj6cBV6Wg==
`protect end_protected
