-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xO6M3CmWLQ4ASaiVcOSYmZiQz1egTfeF0N2Fc8uOkwUkbnyvIXJzsdaPDWTlOqb92FUas+n/U9Sk
jTjZvYL+BR3wjESpwX5pNySHiGGzSvXsKPcPZj4qx1/ABeK6xIoEa32bD7DIMx9A7yw5gCEOKpTM
A14iCAInI7bk/6eFBKSDqllNjH3kzOneX4ZxeABfvid+4ZJ9P53NsZUncw93Jh4O4OhceQO4iI7d
/JQ8AloxD3L5F9mMI0pR+iFnPQq7uFYpdwvBN/AQ/Byt789H2P6gzOvIUwbiu4ETsSOzhN/sxQpZ
SCJ2810zdaCq5u14+ZTOXehgI/vOfLGj5LntGg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
B7s9GOiEzbjUXtRcHtCm49w61vo7pzbodwrGsQwDN1qIP4vOHLOFFGz1IX0mJgGxeOeZ3AHwObiy
94iBAfJ2h17Rki6wwD3vc9Hh4AOMs9VDSnhxtGAeAWeSzFK7Tww9bmL6E/ZDdRZav8VFX75uZa0I
7TnoPdfrc2HkgtDtLVFrr9lI/KkKWwNO8o1P50PuIDcXAomINCwKcBYXjWzybAKiO87WiXKdNo0c
Hbhst7eyH4/0plZunVc+H1+VoKHm2VohgecO0/ZyUcJAFgj6lIv1FXBvUP5AF/oxMFNs65Bl2UGX
UpK9GSOKjUQl1qAIUY3uJcB7/rqhhHIniQw5gJaS2jGXSCds3z6ukKoeKiVo07tQ5ex77oz3KkAA
jGTnu28w37vQzYDgeLtSSBG1gar9GB8AwdOtMI6w8eVga4iW5k0SgvZAH6E+Knqua0kwn9TGHDLq
O1sxx3MaQT5XGwkUxNQYm+8rKQAiV0WWuR4/1SRl09KLM2uYv3sxb/f+UR/av1fTi9yGE6p+2VaA
SHQ3oIQPWhcgr/rJf8OvHcM0e+NSgakRGoj7LG4/5caCi6AHL0eIQH4Sz+MUVgpArkxRiG97JD3J
j9wHoz3l8iApPMUUVrZnewxWSurJt6noHVXB6+BgWP7YpNyOkJuB57Pmia+Cbgz96OvkakcUgWJ5
Rndj3H4NdHUvMdQCOP/Y/GYxyJoCx9HcZvLwuL6q10i37jFAz8+n/GicMgkpFWoJXmXtBZi8K5+V
wB5yvZDVw4ZiR8/UpAoENPFSlp05uosEZ7jv35hoxD8X/KiIwgfX7RLKeZO5a6qWDUA6a48+jww/
ziFeq5eMCx82qUVImoILdSEvwYbtZr5a5Dremv2z2J+ibtJoEpCmfdXYUQ/ge9g2og331QkDLNCW
LzGOyr8EzEkjeepB/Zca2U6P9qz8/Tll8GlfSd0YxFrSQaZnlOw6GMumD2874tg7hmeS8Xg6J77e
Rqe54WwmviOvok+Kuaw8k4D2OMlSwXh7u2123Tj9Hv+l6JEugPAXSud5I1q221exu/CX2i7Cu4rL
098GNzBwrSonxhlKa8khfQ8ijD0x/x55qX7E7na3ulSq3r9gyOuXmik1O/ctSFHeFgN5lDB106ZH
+zKXD5Bd+jl6nHsbgc6RelTCoO1WJtMtIAzj40G8cd3rjT6qYsTQZCnNHZKObrHDqhPAg7yehdOr
bHaJGJFR7+iFxD4VQULs5hyd8MSOG+lB7QwHHNCsq+ZZ+FA6mVw2KMLx3eiW8MCxyWXptrGG6V7m
gTxkEpVcO/v6KgEyNHUpXw3scPe8AOQXxNqkHWbfqC9OXnijJcJV5wq2BenJCan5hL1LG28IQaBQ
APXUUQxonAK1qmaj84lETEa/Le6DKPaT5rdqmX/giZ93W7/sdUXN8Qot8alj1lDF1420iGeLdZ+N
g7E9J7JiHBsl2/4hq4dNVYcocODZ7TLSxV+VJH0Cqu3DAtHgHu7m2RflzPWnTouBiFId1cb+swY5
sD8RLyJP7HvmUSXKS9ESpl++729sSki0h12TGVmpwK8sSRxgIZHSWD/1gc3VGV5L+d+4LppK/UyT
jmAZ856SqC0I7mPjvpMKHo4wQ0PCgx1nAnPkzwtnPGLc3P9Su/yecf/yIQM9zfcca7YFtM8BfOho
nCspQbCiZzjesvNbML4m8eSaDgziv6RKlJZzfzh74km14tlyx2zKJID/oMZOnjCWwkecXQPrNZBG
g8hH6ltWuENe4qvKHtoG8/BDoe8w9E5JlyMZr+9Az3t7nfia9ZaNc1e2xZ10ydDeFdxjm933uo1e
Qc/3c9cOsb6XOg7EIakCJuvXvZXqOez+WT383k//3fB2U0IzBE1WomG+ivkP7TqTSqseCTM9fbEw
J6NVMSsGAxpRXFR3uyzXQS+X9xBsj5yK0PZgh4OqJSN7s+ECfvDhGAa2HCbogco3MiQmK4cl+ihU
2debGeOOuQxBwElFeWT13D5vPnEJuiXDikVqZPXBi7phs5dMpBJG3VV5HkC+0l0DIP/eTm5f1i2o
VOOyS/vBtYgCczSBnJxUCB7ZANn1tTUWnKq7Z/p0nCrBxCkPF2r9Q1HKD2xrLv3Ef/CwJByR2tH7
5LmTFzxHC4+cmqTG19A9k8j0B988pCwe6pdYpLSGA8Vq360bnSZ6Nr2ZPldcEb6vBXDH5sHEVUuT
vqcHdVENJB6cP+au7qWETU4IV6kfrJLccn+hBziJ2dUseyrvbN7o8UusKcLIcVxDDlolblsXyPTo
qdATwJU3RNJcPBsqO3uVPwOcTggWFQuc5CpriyGnVfUAHY0I5r37HyjKIjD9QnWG2EjsZcPCS6De
PtTRZtBFCeMmb6uDI21xrfyFht4fzD7UJEikjOK+Ib8e7ukZ5lEwyQEA+ex53pCc4eUXcb1+11Sf
mRT/Sh4JkTdgsZMbr86r+UZUOtGCQUk5E6+j0l+D5ApptBM/wlcgkwrOkPckeUfHoh2CL3hqEZe3
E1F9peubMuRdeIX5mIBndBjI468ApeETHx2mI9voO+ZVQ6FNF4RgpdVmQAwnjCWFbpizXRM6wiig
cxjrPvI3uZTfc7XKPpuq/2uLG7DzV/e1bkzzwzyO1PCdyp/nHhBkyxZIqIP6pUplhkSEjXnuhn9K
9k6zReVg5MafhIOHbFUNGPQcigmKY82qlIVrhBtT77NPgpN0mEhr8Wo+MXbRm4gPrYI8g02PXwYF
chRNb8UBXtIK9Fgw6Xi/EuFAY5ctWs8MqlTA+WkHw+6lNuWn5+WF4v1RxYT7YM9MDoOKeutSL2kI
FzxePa6WnwbeT7grtEfd2UeNQ7dig7NVTEL8/hW4qojfKram2wqe6k62jEehRI6YSiNfaV7cBpV3
yBN1y/I3ZpX+pQzuMhIr0fPM+2H2WGb5dqAKBnsPT4pJ2iMTMLix5fNGo8x4iT0A7uFPKk3sr/n6
V4Eh+BtExQ79CvlZZAd96DGz9PqjFA4yNXo1C2VowIMGS88rCQiTuPwTPQeSl+P8aIeP0q2PDBJj
46OKV3NYz6qiWscCo82zscKiH3rwg/BcEY5Wpi7qbi8mZW8ujvL3n3Ti1cu5tew+0WrKrmciZoDA
Hrj/EkWFNNrGfb7Sj/SSYdEeGQe2aLLUcdkwqqsRvsAMreOzbSHTAfbeiaBCUCOv9EKdP0fbp60S
H9I5ql0ng4/ggYvWEQQ+w5u4Dok2qrvwAmMrZMMFulXVyhWSbF5DIWDL782WiehlmTmiiwTyr/6T
MGaEtvkGuj3pV8dTPo7nj8ickB7Y1yB4DSAd3Da3Yo/kknIHHpkBICSuHHCz9NtypUbUzkBBNX5w
2/d6251TzLaUeWQ4NdQMRi6X8Qr8M6QyvAo+WH6jCw0pJSE0sirsXt03N+K+GhNg3kLnuj9ddYEi
d7DJxgjYLTQBKmsRL37MwRAEVnvd9FuHwUNr8ee+6Poot/jJ9xgJ753SAPvDMM9jXaonJNIAtg5a
3isCOMOthRxI+6fuSjIbhbgTwvGsJdVy9LcXrg1Y0N4Qtuk3VMwnZPLw35efJgjwEozbcBsnSxBh
4ZN7aGmYDVYTrUfDLiXaiZ89ngF98ZU1sP4k9CAI8xv01/98TmLq6OXap1MnPH2+FOcZZeYv8GcG
XigKgJ9DQ0vIfQeqzNQ6nS8/pMNGNJLbONzVyIgycXXqvMp8vWxDFgK3HeWA/ugPFoe5HIdKFZy0
w2wKMOv9dEzD5L3afQ37Z+VzQ/f2kClaF7nS5fjzb1udD2LoP55twgGvei/Xg3Z1RcvHZGp120mz
cZIgTMkodxIxJJcgyukkp9HHDNX0lmo9+nqdO15QMwqcNWO/KqbSOR+gt/j590l/yEmBsBLfkw8+
Ba+3srKacFw2GJcycmKsm1OcEBYOHmfswcK0tV7XaowgnkB+NFYJIZcZ/a9kOcfq0F0EUzNXuWoO
3PPxEjHZs+qygN14S5VndZlkqZFd5Ka6dj3B058C3hKkcEdu69e8VgKwv58sICcO5M0SD/cYDCPV
Ek0J7LD/qQgw9Fk8TpE54it96sq7XgF5O/vXxTL7wCmM1dA3n4WiYYG8CRV8MIlnp0HpAW/LpBBt
JJZKocAbK0C8aqxHd8w0+Hs8IakCmJ6wGITToCN3YCOaLHY5EzlGuEShaAPGTOi1MqoVzxw2OyAa
AJ9D/54SVjPzRrHnpJUvOis4ShPoGiD/gAOzL/15ZMOvg/khkUUN+HvsWPFo4f5BBIVjXKuEsKWX
O/3LkR7hIDPcniJVHOfqTf0wwHEG3RazVSI/JrMWRvW1daWwi6i3Gnm7ZCpDsERzBmeQCC/KK/cp
d3MP2gejc5TS20/DpKaNWwPry0WUQsNa777QcQX7KA3uPD7kGcWSIsD1AnOD7ZV8L4iBNsnremP8
s0lK3dFJPs3RZctxKbkY4IIJsQZs7025xp5M+5HeYVAyAbDxHzLjCZ2i8ke+0m1Rg1C3dNjGj+IA
OJjXlOkWzdLr18PwKIAbFS0v/zhKxuK6Iki2rhTdaahRTU/gPBs2sGk3nxYwATEjxIv2FbR+4pe0
worVfT0UIdsorY0Izw7WYnGEOup6cF2dkM7S+u/dZCkCDpfGLlF9G468w63s/ZFtHl+QbDm6Cl5C
ozgfXcOygmr/yZi8zrb9WxbElrxiXCQD0aXtIXgXz+b8srHKAdoVKNqggkUY/mVyavDRGSNWU4tW
OcT9sR6b4NzOLGwY8fjTKniRyu7Lq7ok3tYhSL/ofaVsGCZSRK/tOBXDGK/+x/5UVIoGKXp/gbfZ
xtSRXMpRLZ28JKcvGwtOmYauJvpZPXDw452oHhqsGjmviGBsHHEMqxNLDa8JbRrGIiJQT4QEcQ7r
aS9jK2r3AmxokULZPHlgKafoqUbfq/AF2BrXuWxxhDAbxRNkoJrxd4/WCE3fZC0T2CSEP4q4w7kt
IOVPKB7or1bxkCl2281eQoMfJTXSQSjVVjrL4yn50wYIueK+sJa9vuq2FtGPHmmATVa/Yp8NK5FK
84IaMnH6zc6jUFRmMFVXDVYlgRz2I+w9ALupTD7iLmN3EmTfTLoOne0Rr9N7N+q4NAEm6+OxkMT2
GIhR0Iuscp5/PJuwzrF0HAPjuRM46ZZ0n7/aVD9/P06dMcD0qbKfOIBvbIbZHhc3EbF5qvqBSoHn
Xv7HcNMz9ua9S80TG6ihKbibKe+XQUPpUeDPvgO1quTCPcGNqHbT1zmtpPkRSmsVp/YJpOwq0xFc
c4j28QP94pyM2b+qFKdE0JzkVjTbTxIU2vlYd1blPPujWUfzzRahASSglBBMM816c18dLP+PxvIj
YVeKGmkSIXif1aILemFiWmouJQINt4udf6LL8zV/mLtrYxvlEpRcvZWEPzA61ZqPUOyCO4TsmJFo
Smdky32QisUo2WzQCVJa4RrV9SBoJlUA7UnBPMQO9kCZSTz8/cN5hiZgaPLorQTS/4PTIGkR7HMr
Rcn20ttrLKSbrbe86+20nYzERCIQfiM1K9XIs1H0SyU8veJegQz6tRQJVpxGObFTg+uJDRGwknST
oph6jFxqMZtHO7jtfU+c9GzgbVXWqaJT6BIEA0WJk9QRFEy2Soj8eJlLJQ9Kb+DZ/yPBZmbujFQF
ZYNg05Gju5Xv2S9OAdi9TvLZVqw2TnwPBhlSpe5wEw5HZGZiN2SWtCSdJziaMYL+4IMAM3XfdA6/
jgCra6lhSZkEy9adtAswP1uGC/jTjk3gokS3T+JUvQrF40evdlfv4FWpdGXuKNjxe25hMzJy+9Y1
2H82ALb7fQ6WPknSwF/E85iVi1KKC9yxgVDzZolopKBamuWMxkaUEonOd29EuWcryMOK+DD2pVSC
14VpmUgtu4fF51bMK53WjnHBNy9I3z09F+txNZZRfB/QvWI/1Xgfi/myOOeKaFj54w7kbqXx2wKz
Rkylo82zszKoKXTjlVbdID0tJdbVTVdIFMA6DjMFwQlI0KwHVpphoVyqpumDvaABDxbhhZHO2MyM
fI6qEMXkDRgcFB30Wr1Z2F150iJ9Qrfaz/HxPfpDcKyRjO0z6TSJaIno5xw2ETMSlD9vyVy8Jl6K
GhBr5kJAX2aFW3d/3FmZEt3zFboBZmxSZ2V1Sm2pH/QiBDa9jw8jaWYFGfA4l613NqtLOYcqGHMH
xJyNaJZGZxPYvKynVf30EoMRqCCNbTFYcJwMoKeYsP6hfyBHwS6YwdwYuCvNV9lU3Ka0A6dDVLJW
j15IL0axXwEnuJVdyUng9wz66KxWzvKB1sWAbiGBpsJ9BJ45g4LimO1ZfUN6CzoHoO4GJLPraHxK
L4hG5W24U25T3xNjh4962xKODnmoHcJw4e8yUrE8gRo93nNcuGEbdAYP85Wu+uqrk2kUYclAdKMH
ZM8ynDCD0QNBoUZtxV47+DBH9r/M4eqZ+oUpu2yfjpPYuTO9KgniqfZyB5j5sHfSA13CidbluhfI
H5X4QFm8QSLd9fQfXfHFQ/CVQ2b08nmo8zpYwWRXO1pBbf5WMat4ecPk1yVUUbmanBZ5uZdKV6dp
QDdFLL/Ac0i/m6OAT3LlJ1NMcmdPkWVjFuC181d3ysKX0PHgoIevmVTNAB0nwUyhRd/iS0UDF9BQ
ZJNF/ZubyGgicq9K+kFPag6UaMmF9cFiUh+AxOaaAW/mjAeM7Qsphz1o0msgK3SSaPg97iGpwNlp
UNLTot5ICQ9ciqX8QvPmfnZ/3Fj14gCQk9fgT69HsOnuOVV8KSvkHSX3tdKnMlgxdpdO5Snq9slo
PM7RYFZTP3qkNiBDh5hTc2tutkYpVqco9FbXPjVqmIELek0rb98Q+JjkBLzVb/s6YduA+bY8lfXR
tbZNX1fmh0UnU+qVzLUqznUDgDjlxp48Cfm4ZVMlQ4OqHE5xsapeHHeMOi1C3gJTucWCB+ZN88Dq
kEGk9uCo8sMLpXwbQgxGmnmpB+5O404BVzLBeMSpV3eO98PRZbPGSIhHjyuXUXekN2sgdIpj5t0L
2RyrTka/6ABlzA2en9Rw+e4o9i7G2wKRS6n/CPFIKL5PEY9YkxMMbNy5nAwhmCyTiPpSmSKsg/dg
mFVbc27XSKDqU6Pt2CwfIBscD5uCoxg1+I0nO3m3MegFOezb7WDJkA33C4N5DXUGmUwQ7xcfswq0
NXmIqDt18TCf1loNDWprhkNcHT+fS/yXMVnMSSSuQunFC8uKvx4ukEXAK3hCDF8xB04eQytztm37
oG7x+90ysFzZuy39dX8KB+JSLWZWIJHkNUZC2bF0AKHTKUKExYwL72dLDusNjJitAmRSJ8WVWawz
u+1sC0gZ0au0idUvu7zYDL03RqiALecnVRkepxW8y+aS85vEynmJcMxicDFMpR2mGcRUGG20cPqH
o5Io2hl3Sdv1xUVNeUshJ5x2Q/yJqqWmA2O/AL3BWdEJnKrbz5BfLGreDHwmPlrkm5J2H65FfDRl
OKVNFGfEH9t6N4dSIm/QGjE9NeftYqE/06W1PCtAVbfMrhZrNHo+NMq49w8ByG54UooNV/WaNJAF
meIg79VzfP7jqOfTp36SpKgckG9lDoIsu1s+7t23VU/3kszBdQw/WEB9Ld5dktW93Rk6WaUBukww
Ejvuk3udufMVsRLPBRio3syKdmZ7DN631fScOz10DfyfEF3wgMcOLTG9hYtzmtrPHwyXR9Rq+JR/
SnPDwys9pWxwJeAUZZmPkiTgMDTLoM7SGbf4Ewry7wc/3MmeehpbDDDeXYmx4pl/A+diBBGJWidG
mG1wLELGf3nwa47JjA6wXxVTarJwGB1eDKfqUfb2KKcZaJxHOHvrpSsDlUckpzaA272No5fvcNE1
kmwDjFBUe5XlDWUrdl9YhxlBEReB+9a/7iGRjnX+8Un1wfLyFX81+IxMKO3rV55jmqAeAX68Czs6
c0RtE0+lJVUjRG3AXg1v5vlxjztr6TGB9Fpb0G0N3vQy0Ye+NXDD/y1dOcn1ytTZk0jx1C2aDW1y
1/3GZyAo9/4b9ibAj6/kWrvgGPLkzj2Wtb0YBnaz8eqadj7ItUVN6tt3VQdMSXERd8gzr2vJ/qoY
w8ATqm3fUiDas07B3X6tEfsIjKW13KHW1unbglFH3TTXtafAQAVSV2kWADBG0RawSrH3plciZ0ux
UtlgLP+MzIViQYWCqkIkcJ6x60pdxqnLFFId+Dk3ITlmrN6J0jlfeav6eXwtQrHkJXur68Brzc0o
X8XarfPrOPVzZrAGdCsy+lD8A+rvr7WXGOQPBFdmIVsnnzPyWCpQpZRYpDE+epQYO5kMEXLo4+dP
+HfpX1QIyRYFo00wd4O+ogULrKYk37gZBmw+ydF919q37Mkqo2ctTygV/pPRaBiu2YIkCq2B3++1
LvczB0XVP+lWpcpQqfdkieCPoh3lUX57jVqZWglEOa7BXk2tTVmUm3RCNQz417VIZP01lsyp1B5l
Erbl1RiXIgjWdwri5l65dic6pzlgeCnhtPpBwvsfi9sA9SgFifWtVkznAMfuhrl6zhur5egbA5IM
YAJvEo//jk/FFUG2IJcBtWu2I5F0oXU65/LD7U93t87BOiaxGd+PlGuvg4CDzIWooVpGby+SEJJf
muwGVlXN3v9dh08CwtTxjCXLK/cLG9n5+4uiECNqXg2QvhCTiPFCr3967yUz4hSw/pysQ9giKEyF
CW+V7uUL0q1Jr7TGLxc4FlgkiQolibJK9XxDzw//18bOx6SVXvMWVqaETsR942wgwK3bRUWSXwro
+tuufA8LOZjt9QRuwWuLUMX+22KYfuETQ71aLcUxz5c5THKFeNv5wb6AmQbcP+XqNksK6lraYu2C
X/qqsFqJs27Jny6GWhGw5KLkJ1DBwfkUNY+hK4fbo27nGaB5xg2O8bhBVkJvT3A8umbDvwMDR5bs
U1E4hdFAIqUVxpKL8D5C3xX4xNnQOM1Snl7K4PaRt9pk8Uc7ujKYO8CNfcm5eJI3S0bqxKeChMW4
VuMKd7kyhfptunDzf0tJk3J+XD60eAoS9++XROkZ71hzwMN8jofwgZE3avCf4xpmbXA7zxB0NGHB
iuvDqFdr/4p7FzI0Z/0tmc1B0n9nfN+nei8onu4FR9X4ge7BdROPegjOcDGJD09ND8HVHfSUvm9P
DUD1H/Ko32ihv5tWJ2Wy7Io+9iaWyT1ivoBgQ2oWV2B+YUQKYOUOo8mbMmvYcu6dl45/ZdQjYtpN
X++pLm/UxLjn2xZN2+w7VvXq2eV53KgXuoM2arudQdpwx3Y/+zVGS2tq4L/4WLeX1bmUoUrGy0Eq
PdKVYneH+KWCd4KXToKbqJMK5py5GC2dlErOoG7MDZ73gnG58ZF08xVn7SCbokSWpaoRln3N+W1T
ECEgjXsiptxjNg7cCqeKYM6A98I3t8hWjOCAz8Hu8b1+ARHFMquiipjsSqtgKywmI36QaaF1d9YW
NgP9E/JNCPaYwkI2p1K4JGIxwZ1Eus5LerAN7H3mI8Cf5N8FizedvCQQ8OTPauap89pOqhcLrXnb
kXASPKWE2xp9Ua7ij4rsRwX/++3j5V++ycfQ5fvaEIQEchIyrFpYTIIA9V3DsNd1hZXEAoDsnq2h
4x8fedCr6vvpGsIvA3CbFa+9jPNWPFmX+UZtK9NMMNqeZSWU8/wQUOWRpNrSCRtLx4obkuZUA/+h
mj1B9+GALnJtP+W4QPtQAVGj/M8v+TtiEdYjrTFKch8kcEpWnAb8/0ClXJGgIaewEyotDJHsL9US
ztOde/iTy+CusWr43VRpln57+xdwifN994KqC6P7bjkPf74rDuEDiuDuqy7MakgIbEBaIv2LC8kN
GVqDOLCzSzUrCOOc6aA1T4oQI72V+VlblUoghCiqZ44gYy/Jcalym3DfUxWrFUpnfiQATxqs0HQL
7vEvTJShMrnR2sRaAJhShHCq8EC4ibr1Nlt/FT0fEcZFeXmYeNKkJ7lfuPUkbPduX4CrJxxWxKFF
NX8XT1ycgWPLulkCNaABFFiFolpdv0wfyA/Rj4eLl4GYuPCE0x2h7Dh3ukYp4OLvNTKHWqwdOIpF
T8yDUKNjRfII1zdEAKXORNUwVIw45dvPNTINIrbCFtmCXBaihYlJvRamDjz1LCChGK9m9vaI6k2Y
biKWUZg2/ufBN7uqgk+LuvOwWgCO/kUihj2AOazz2Lt1h1LdV1tGABTH9ps2WolB61wsonrDgB/q
oJl0eC2SZekLAXmqSEusgd04kljz/V3SPCqWqWWjcd5Pqv1yqH1C9RTNNbHRPxQHSZpL9yFMT96J
BcAEfZLbPNLg3V/opIOd6pGTJTqNQ/SxSUaH1L3eVM5iX+zze83TR6dV0rXtPWylJVXP8/UP/umq
csG1q6hkucFVKRSgYwnQyCLfkX66Xcdj3Hl1iOs6mwwvDnSDDzqv4Dvm3GUrI3nxnez7UsTexzNO
CpfTBMdMhirBV2tpAvwqFbMAKwyasj2fllsUav1OSXjQhSuM9hPnRY8Fq8CjYtLGi7EUGNnc+KUe
wQ1+ME2PYAeqYXPfbss3HmIcliAv8G+kBlcQj1WzaB7y7891ltItJq95u8J+amZKTK71cDehhuWo
fbXN9prkXvH6LV7PBTmQUY/RE62xe68VZcm1/pA9j7gGp8MPf4RYrEomEHQ1fsCEfdVaClSLT+sQ
/o8+hsShzEBrFx6Mo7amFfItvHvdW90MOLBQv7JLJ5ZqLkiJYhpVcoiIaHaBkG8L8gTeJPtNlZuZ
06ZTK0XDqlE1T9/uKWnwBjIUkVcoe4CjXzxLmYid6HXWJhJCEIkB6H9+L6VxU+j0ZFRcK4wCMS6b
sUEJshbzIyQpSNShVOxfjjNNRzUFhYimLmdMUHmRRXyS2l7v3IphMyXplJtBFSC8xNy5c5nuVAey
uLhvvZgINAj08xGjn38QojoquBX8xFk/GkMLYjWod31iz2kbVNAmmI7TJne0Z0EFW1ka1ty3XlhA
6eBpNsnrznudzGJ+YmZr5D7ch5XSzOE3XEkrv5O47f9jIcucwiz6IQwEGPkPk+AZ+JIxImz9JPmF
LA6qe9dnNF+Go0lni455pFbeCOPG0ETz0t1O44o2/j9+LD5vvOKmhdKXsfIrpVh0dg9zB6S1r4SR
Lq0Wn1doTqvFiG8a/D04Q7VXpCuXw1nBWKtnWtAwr+Qvcyt9OHUEXgCMFRwjHfs46YJo+5ZTaNaJ
H46Lh6n33vtmSBUGSFawMc6iV5upJAkuMHKfqI3XQJgiYjjakSn13nA/dvtorunZYyPB80ACSA3/
2axKTsE8loZqp38Cx67LRQXe0i9ztFrr4um8rgYER61Gg7RX0/eAH4HH3Sd93e1b9646gu8jDIzd
RyuKpbR/aKIDYAmCPlyzgWCKhVJ1DHoBnS7v8KsjRzWJBxJMyYqmwyLww/fit+keAaScrCqec1ru
1ZzKhUvu9Sx18jSo4vd9N0SawtRZVr14tkakp7VX7mMiNHdb7WaQucpsWYX1IoJK3LSVUVqwFSFb
SOjW1eRUtcNCSZWMISaBe2ZHkY91OvfkfMBmfw0WtlGYEbKq+7KIagI5oHTpQIyL/GYuz88U1lAX
7CSa/Twf6vakuoIB/8ift2DaaZ9/ONOUhM8XB0DX2IxwTs1nKLXN6WK/bZl3kKKGPYxBbhhlb+6r
V/ZuyJXWX56pu66Dhi5kBoqf/iRRSmhzuFA1S3NZ0oZDMWDazZPP1ikF8QqsHWGjYPCwErc2lfsb
S9fcN0NOMzFay6GnnuDvG8kH/luHMjfyKnboai9QTDI47vImEtWTPlT98CnM27AChCRhAn1xLBsY
W00PgW3s8sqkMK/SuVXkVUJ1Ii1ty6bVNoQU/rGhpIhIfAtksrN63eOXtPFFVmZFmPEQ/LSaQNIR
1SCf77gTyohUkxB7EhMWl+0FDkt0W4m82+rq37yobV/NW8XyYzlxL+niRNmqSAj3gaj38JDWEJOz
ZbJOUt28JPXOxpGN4LDxnLiC2H2u33S70WDs4YUcE6yQAf6MySIFz2eN0mEOXdhi0yfJsVdGjvyH
WMDhHRiF3duDRrH42vq4dLMB9yXiY/W/Im7XH3QUNKMFrj6PopCCFeSDOG+D2TevZdXnr9MChdOT
hyWAkSWVITDdcisLllqoEA7mkHwH2yx+M3O8tsy6DS1yg9O/5QXf3nAtqki9K23/lMSd8MaV1EKj
njEe9zAS/LGxELdJJWwgEmA7+lBUpMV/klX/Vt3N0yWwuFLlUeSKTIaieAOasC0aYh/TGXL9zmen
KVL/mUW+kcu2gKE3APYIrXJxHqzqTJ0w6wi+tli8iheR4ZAyLwXf6vrl5iNxQHRjimLEXW92AZcq
fzynhY2CAeXO9tocnXYy9MDZtv2b+/Lpunbv/DFryoJGiUGhYzicjZtnVx0YLGU+nrx66whw1pW3
vhvZT+Hjsg8Fd2GwOieso9XJY/pYW/I8IwoJgHIaPcJj6Z93BdGV0ZQ/CwURa5pCw+nywzErNr6/
9ZtUKZ0GZ+e+TXUVHZL+Sbz3HuVlMJKoMAUB9Co/6+El5ejDtk6H40Tp2xcivm8hEZkylpVX8Hmy
IvMLk0bctNKPxqrA0/SrjbHZDx37h0CjYRRIoO4+qzsmflSSO9XBEcMqgW9ZCqdZnF6+7XcwX1Vm
2r9F19jTCEF3OokQsOa9xZvltNw0f0w3NGtXPiFb3i7DTc+J51fxEeEa3cLBkiDMmS6Dsdm7DPOf
gbtRllc7pZGp5yVzlFFVrVmA2iqi7mIBTVWaH9FavuLaaTlgoDF/WZJe7QQduv6VtpSzgFhDt8GR
3zSvCHiRvhrQgALoqjFstY0WiLRFz7o8ZAvKlPV90eZ8MrLNACdRC/CdGRMI/EtBFUw+xw4AKph9
JfnaIqSCC9gJk3rBVlLX5FPeQHQspUAzp32JTvxMNo+dAHe5vFxAebYoUhogLih5DXxuvT/VGOWd
6SFLrn3igZjPsA2qNpnamov4DLFV4grFA4VyJZxXm1QKU53lXFE=
`protect end_protected
