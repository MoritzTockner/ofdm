-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CfSekdm8mgfPPvRMKjy2UdeA5tDOO8RskHhVzNPW4bsC0iIpqQonTj2dN3STaSW0hL69lpAbgwsF
riVO7XVF/VOEX8cLZ+WztNqKw0YYlRewtBsn7qix4Nlf/6prFSeqsIjZf+FDp77f7irQ6SM1hQ2n
4HiwcCTopUffy97yIxxnmlsY0Ec3ONL4+Oqq+lkV69Uc+hF5b543LICsm7zB4b5Hi3HLDr9QLbL9
nI8iZfOREMILl4esnpmIUgxm1T5jmzXtKQywMeuALV39GJ59cqqJ+7EjiJZ7F0KJ52ugXzmUaQpk
Fyyln94Ivc9cB5YnNOXrfSweWXWA/qT2vLDgNg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
S/kH5YTQFZ17ECb25wq75wzYUKd5Zf4rXsjSa5WZ/JpNh06hVjtl7yYCFkoa78pctLBsc5OB2+wE
hurcL9OpnD63nLISsbINITaS5QPCv8qdiS1lylMhW6UcPzCvf/kfA5sP/yQggsDLwJHJKBdvkd0Y
qieCNJCMOQcHgOEk1sO886/l4gtMq6f0ATC1f3fdXxbKS23gQP/qYg9Q1wIY2FbLftMypYoXTsF0
gX7k8NvcOKiAkqYnODYVZKekAa2TxOC+EWgP1aL5w/Cgf6pqnpZiWui/aQJ2JMjTzcS7liCzReMa
2pJXXJ094c9vjOuhMkI0d7VyT3GQ/gpNprvv8YoUsZds4DOpymx+gto3wyKD1/M6phgyJ9IuIqx3
J3NXKHg8lP+EqMfBUdpPlTR9zV1jLMuvMaknFVRSRImRs0XvZaiA0CNJPcCEn9SA8J1BHa7My+Ma
wKXrrgA0KJojKaTa9Mhrj5yA0czcLqv/eSqkgdfkSgGiLqxRNZxdhqvF30GifwS/4qEa4FQMkeK1
/K01gGefNmUJXGawnLkp5K+shMbZMjXqjIN51mg4QhhvEjs0WtPreFlAxO7kou0DN9GrLiBeFZ22
Q/1M+HJ2OB2M2QXRcGxoKN9FK/LPvYyJ7VdB6CLGtIYjKBUBFyX8kmbDO0WlEXpi7aIWlCavagqG
Q/ARw/o4Xt19T4qOQ8PpADIrp/fO72/aH+E77VLCqn2Ge6VG8OymrLfOmaocUx4+5xfJP7Em41C2
8Ej27U6hT17qYLJu3uNwwBtW0v1KWcw/TiZ1IXq7JFKpEJZR19aD190LSvf8GG8lPo/73baOwx4g
OgeSUB6ReDAFqDOScl834et9Sg6c6egsAvANewFzGw8QoZSZGobPfiUYeBDsvcvBRCAxkyC+uCrZ
1b7R63AwYamDqgaj5KzjsZelMh4ZmB7REzTlOjHUz4L5I0oTNqy5b05dNbrmLnQ7ShJJPdLn+EmU
0EMEG1iXRWGuvx48Ov+knbbfxcOS0+Pd6pCPu80oaQo3N4nokzPDm3fWfbhnIsX4yvs+G3UjLgT0
BhY8jAK0KkoFXpWhzChLjR4aQAKYLNdQzhAn18UBBFJrFfK6jDDUJW5LM0/oz1/HxAwvcL+1pSSZ
Tc1zK+TyP4RDuKc3uFnYHhnJv1sjY1ibCcOmv7LGAPCr472vOAOPDe49Jlao16//8qX//1ORTebW
xsHvZBlLZWZuKBcjooydALyiZmgIAz1dVSadkgiw5qQeJM8cdwWy+6Si4dTwzozxnUbj4pfghKPT
ZiAYQQTt+WF6eZouOxg0Pihf/+6k+bfV+T8WNvmV8ts1zt5Ntt7nP1BWzyoRjUyQsuK4T/of0aRh
L3o/zXSj36+oEo1fSiqj5YTWNFbWpuWHLW95R976YW/JSdvEbYpkVE7ZgqExgvf6uiTWV3Sb8aJW
AyCHzUBrWxQeuoaLzH03gzQgmPFr/Yil36DFXHcWQAwWhq0z+GlLQZ24nt+D4YUoTVaBhxcNKFG1
HN0Zr9eDgQKEFQH1y1+dM70N1n6lFU85mYspYZXc6imzn+LzrXFFCNHX577p7ftbbHyHjyFAmGML
lrpXqPB1GNnnnH7ily3uoFKwOykZY625INki/VuawNDbgRh82S9NoytRKT1tlKGe3HuY33x8OqNQ
RQlHpnH82OCZg5J4c+XMUdciAqdt1jXLFBpldeW8UCrqWTKybcBZreltuajhceR/ucp33HKmqdGO
WHfD10PYO7GS9GlDj3UehW8o4op8j89+ur0YWkMRAr6CotkE65Z8nLqZIbQXXw7C0ATG36eZOYU1
4Ggr8Fo+2Ubf6Fr2P7n5DcQ5Jek6PyN8zZOfHp3/A/KZWJ2CgZRmN5q47YA+ARBPp0vx2TE0VeSz
O5+5g3w6np/G8Rj5D7TYwWWMUEyMXMsnRjKOE3gM6LCkzs1FGcSCuVsYb0Vy3hMmxiOEXLW4uRGd
eZjAtqAIOhkxNcHR5OHOmGM4r+gFrFPcPvnRdj/QpYpGTgSutLbIRYUUcCdxtL4FTG88+ImTIRHK
N1Dg39i3e9UwI3eSScxUA6aKi0Ql6bSIKszRmTt5W3uPpipOUs8zwrBLTQGPr+P7E95Jr0lmtpJi
ZZ+XIfSWOSRoXn3Se8ivn3e2zKeT51P0Kn065OQNb+k0m69zC6R0lgB6XK8FIH07Lq/hsfJM7+rs
mxLhaVr5PsNLyxGWiY4oG0jqpxkMCVoMFTVKya8DyLKQBy/LcRmB59MUJSYYuhVJFN63r79Za0oc
OzChaQUsQEzIKwgZ91XPg5ODwBeoat6qH3Q1ibT75mpO1IzCtfGr6Fs2VX8foxyJbzhVsW+mgq8O
9QCNK3QxQ9R8RnXDEeVoDpWTv+EO4NvVTQLLDujtM8yaehSuzntXkzM8lZhSxKF5H7qqC1gR0MP3
8PUE0oRi0nQa6+R7YraEE/f9r+AJlFanzWCVRC8TZChxOTQnzwEd41vPVlLF5NdhFvKP+C06dlk2
G9jD1jAs0NQ9x3N7AuhbnMpH4978Gd7Yvm/J1DHvGECcEvctHVC67CjlHkDWCaNWcth2iblKHzGa
Z2u8S3aI0QTD2QtK2weMq2VBoCyPr96RhTphfVTxnJXE7y9zgxQX6SDmf0QKw1yWYmmX8wUclrtr
3ZzgiROmv4T71VcnEX7T6xxybofio3pdupJzNC2O8sfsxmc1g4pu8wNywio/HRzovN+9lLKF5t3u
s0YImN3kg1EayqruYMDDvKcpZEoRsfES0+hKpgZNZ+SuZ9YRgLeiG7XhbmyR59KaoNZTSEQBARV0
fbSXjpMSH3kEv1sXpKpiwBsmZ1eIXQiUOfqgZol3vBi8ns4sBuTwFxcJAix+5fiKRoiF8Tnr3uGp
T/5QEsxS98cSt1RMt1ehi3n/+lxKNplgvAy28Lb9YMOg9cxZVGHiwaRc0wO4ffY255DNcO+p3cE7
L/QsHhKi7a4B1+o/IiEAb0hYLWWs/6eeiJVbZzQeqjFtyCf/qaB5W0xFmEK0AVfPSk1Ai4xy9Cl5
aZbtTskPWuGm4sLE3wMFhoLhHqdiRvUe15R5n85uNJxgYpvUGBCEz2vCDGMcgawUsit4lQo+voVj
WPv6Yuva2vE+htUHv/Ttsd1JgqNt+LZUKb+ymwtwkvIg9K11ThIFvWCUTqoU1ESmJBHqbNFQ9BfB
cfzxrBJE3xoDayD9IpOvmy8GCbh9KU9eS8ls7eMtkweRrF+5YquNQQ07r+z+xbpFNf/LniVsU3Tp
aFhXZ9OrvHGs4Oemv2fWq4S78TzEODg0MGJAbrOyWA/mYIkoO3IVwb9AemFdmyZnMWeDzzcTEHpK
r9f1TR8Uubw8dbrnVbNbl/m2VrSFTUfKiA78WwExOXHcxElhcIoST4tAFHW3L7o4pNzHIdM3OMLj
xXbTQd4hzoL4XyS6ECLbYtJp1dfwpNCyX5JLkK/mEJXyHInBcgv8Xo2ZeRthp7AUGX/fo4fOwVyx
IA4PVhCeQN5WztGTUfn+k9LsUQXaUfHLv5coqoczB3DxouHADVyi4MT2bEybMxnKm7zLoAE3Ct75
4bSexl041yqZThEK9OOpEe73kpEeTveAzvgpRinV3Gp9usa6QZhdKZ30OfMCVUId7B8rFjy1K0Ii
J2eCQ3/hPLjFUZ42Fvv5bIPIjv6CrybvkVx5xYquMChWOZ879Tdc84prTZqR3LLp/rqOTLIO2f4w
DeLjeeHUWc9vCJClhNsuQnEiVumakuUfkxpuqp/llNnO4lW5A/ENkDD+8niiRrCZLQe+53qD6wvR
UhoZMhVLZbGIMSbiPmRsVahVjXQRMVwPND89WjmOkdbBKeunikg3xTHb4mwq3Mb/GGBwOigJrDRD
ixKH2b9z54IMySy76myUoDOyBHtTtrdBndgFbrm0mJtkGxKGaQhSvRqwONknogDwqmwP2zquYgg0
1IzdtVZcGyBK25V81AHTzWNJyrfW34Q3I/7os4fBmINARn3SjFMuGfEbXYROlEkl+0LE+k335EGv
+/IQD3qUW6ByzKnYprQ1FFuakpiW0og9dvdEMecaj29YK6B3nCxbHb4fc4KbUmdv3pT4XJnkGDkD
ZqX+bgha2WuCnYod+4dN+PHQ1LOvcZuWVqkP3IiMW5NoMTwh/jktQWVtbcuR20BRq0BLO59s5rTN
crf33lo2vQzsXISeQzpu5JbnmeW9SgI9dafBIQi9I421hAtVBN5F0TCTE0i37lF+UGQjq5l6rNJu
ywMwft13s9QqTthmeR4sioa7L+FQtK72ON0bAGk9veGAuWLGrpZ0kKQeZSHIM4sUcwHGqpWLgg/s
c8VCrQFy2xQk00Hso6B7MiStPAZm4RUM2BphAexJSCq5UXufVsWo2sTM4yTg5UIAnL4RXaEeZgQY
CcX5fqAoTgL1B646bQAcmAv8SP+uRMPJ/7R/F3eRf1/YINxYMNIdjGsrLErfNu+o9u6mqF+nyXmI
Alf8dsKYMuhEL9iXwm3lD2Y+UDNfFSXXMSpJ/kIC7sXRR5iL1WIxsODf1NXCZWyrRYpkLUkNv/YG
QaJ8aVbSdItQCl1naKYcy0FzWgkR1NRyiw4DrHb7cIixZSBuTLjQWK7vBNdYYn/LkWX9zOmYgFq8
iOgz9rRXT7lF9Q0Rz0nDmFcFoan1sqCUjcvCQFPlk8ZUeQRPTGLQfJkOkwyZ3fKeYintv3GRtlyN
ao5i7toc0W983zw1KS1pBUZsGq7kNHX+IRZzbq7uhjSjmNWVvXz1zZyWYP7XWBq4o7ngJxncIA9U
PWlXw3Bvjzr13p3067KJ5uee5V2y9jrnSmqR168DGmrOSlxsRy+bRWczQkbr3tUT3OU4eavf3jip
XIwJS7MzJ0m4sTaIuZ/8PB1IS9yorRYxCdnQc/gNwcVKaliJTx1rzESNs9cCxNcGVTHC3lYAASFJ
aE9aTVsZ57qZ8+4Z69GF+LfqUypd20vB9DzH4JPpaxJlbyGeN6fnJbK9s0fWK7rcd2kAgx7LIOYo
8GDzf43AHtZrb+738z8mroEWr1YkrwmPdGt8TSkoSxhnYTO/p04FKqE5Lz8HNfWnH3C90LLbC2pO
J+1deBElgEfL0uoj4Rt4aCcRKllO3GNlm/HeFXeKikthzz8UkLWBy4Y82mpQRrAfJHHhnE3ZY606
OFw6+Qy75Q+OLkL5e+ySUHP9xpjHkFetnXfUgMjmKHFjtXhYabMgt5EJcQ51i7oOKUkZBd1C6Q8S
JDxhDm9n7vmtGW5cBhZzhjdkKRpwoSsV0eXTiqth6ifAPP8+dqFsHJ9VAGiBcyPiPJhdGvO3lig1
z0ZKVRmpsxPIxjFOlZyWvLGI/VAzV82GiDGlLugfOUyKWfTK5XbnqAgfMGkp209Vc/YK7CwF6QG6
MIIquF7Jo0sMalM2lueJKPyCey0EwPb9Pa3gpi8kF2uEMI4rPuLdkN+weiABYt/QE/rhNEFjN4v0
T/lmGO0RTjN1w3VuB7xZMn2IbJOEjChb71vpCEgJKWNr5e/MgHzXIaz+gZQ/w58C4TdQpPsk5RgI
v1N/wzLdmLenuql1mAdyWWpUwsE9mUbMRFzvsRiVPFqHq3JVNiR4t8Jz2tQ3DmUiHHldjkr91G4q
Y4WfwKvL8dw8ymB7Mtk5KmTT9Cpqyn2jsRdv7ou/28fg2J54K8mJJ+lJ0KvUydYBWOiU2Kht4fIG
wXz+Wj62ZENljYamqjy5l3Zxyt49gMb3i9ujC+ctQfG9jiFS1PbcssmtYZPAZ90mxfLmiZNFNRnT
lEBJIihwAJ282NYrD2tgQIQ0FZcXk+6/mKOC5bg+HRG6GPsVipaW91WmVQ0kL2d6Son7Al8IQ8lT
rnGEVcGgf7za3XSTHNjChJH+XhJA7/WUVGWl9Gn0G+JbKmKW4iXX1ci7NYvNflJ5E3P8RERsyPKn
Jc8qpi9aWwfoQPpqsJtRvFdXUALG4NZeTXl++rOlwnq1FjKRmK8PHIOXH6sChv4jMzaD+TjMguq4
OOjaCdBpnmxoDNFpFSgy3b8ClqQAJdGjuXSebWYTMQNhnY8dpydwvaRyVp4hF2wceqL6sRX1hHSM
KKKUAyPqElytbXSfX1Gfseah1jORDj8/d+pJxmsDFpCkOYasqyMIYmUfZGg3pV8bpGhBgCRYS/Go
XQkxythAWgBr2pI126eIuuLS7BnPcAkY4LD+vZ1df5EcEzAWJQAFFZAmQLZkxqoqm2BFbUqAHoo4
mDuG6f5HcPEPH08i43/sEgiRb1B9NXHqLt7QG6lXdTZxpOap9se5bxKNv4ZJZmq7005KYb27JFs5
JeR0gZUAtSexOynW11OCv1PpyZIcwB1ltGj0QJVzQZQTHT7teYA293nY2Uf0KqYpTGGedttzSK/b
3WzDs/XOqfkN9eRXXPcMvMUIaQwIOnrL9itkuI/qMhGAgb5fRh98wEG57JXXaD9KWT6QRBER/1S+
CBOwrpXay9Enta3PVRa/gzsEs2fJ2QZw8FNq4q7LrYoGMPgB7Oxti2X6EddEbhZ1N9Z3soav5vSA
58d//x2ZRbZTQgM3tdwh9MWG2QZEZIDKtLFJs0J9Vboq3Abxwmkf9MVpIOb44wxnw2zVBh0HniMl
knNHUVqwRPfS2fwIjHG47BomxrzuyR0aAamN9WcUWVP/zmG2grffeQ8L+8HD86sJszOSXoVJIlqQ
eXCLI61zRin/QJq7D+UeVr49TmnND+jD6WJDBja21geSwf/iaMSkjyQXdKBwvQdcxy42NxBx1ORy
Gh7OKou9RPrq5k20Sd+HRkwtuBAmvHTaIpG1waI6E9j3n7hPmjV78kfEq8urkjpDe932RLCHdh/f
OZKXJ9ZxqMOe5khFIdQ9mL2TNb/X22ILSquPzC0/jS1KCIPzNxgFs1cI1MmpSikvY5cprc4I+1+F
KbxpOnwNZylhnGDzxUfVxB8aG3ddyG83eK7Ad4kOt6HO7byvLvgW5c2ruadRkBgsPXmI1ypsQ1Ko
zExvaZ7yoKWN3cqSDRsTKfk8Rr0jatnfTFd3b9GJzWARRYdMtGt8CYNn/L9e4JZj6anv3JncY9SD
PcakphM5xGV0XgwzczhpmgKDmpSChg1PYPTHrkriOYg8DWxmdhz9Ut9k1N20kMuWRe0uIbDreczR
knxD+UWolSLnXu3bRFRVmxeaTluDdNAA9qp/DGT9cHX8L/UuobTTYeDVPnyN2sgfWBhJGN8JvCMX
fjU7otiq8cWnM6L9qCKo4/L8J4nOw9nOMDJDnKhafhE+7syvaN9FRikD7Rz1bbn4lJgnUirhDcT+
ZXAsuHBKIJ6GIuc5vnjW3bedmXdvaqLh4m7I57SOQesD51EW5ypBUZYUGWUd13mycXkPIZ3kpBOM
+M7BHk8euQuvMYx9IivZXlzZLOtnb/QgwuCRcgCSyJyO6Zi4Fam/V/7kXyKNeov6kGNjzq/hheZC
UsEaj5tii8ueAW9DBrT6hiyP1RBdBEuMZhbpP3gK7CuTNInudCFrSmBYPLMrdPJEIui7cO81vuVN
U+0G62vqbDqAqLcHTTL6oAYyYQHsqiC9oPWuO7QOQYHyV1DrUXqRZcD/siQXWwYV6xOuk6VT3VQX
H22N4OQjkV2liLCwkek3Rtg+RwKHw6AicN+KTlxxTVxZnCRt9N4uXqU/3UWd/IL2LJyyzBsxTdSP
ZkxifXWZeQxquYabYopJNlXL+Fv5eAbDCFn3wHIffhlXbzzswDJz7Qsi/JReq4rhXEOn7KqDO1tn
9eZYfkpr41Yg2TrMfwYL2Y1COhZmeZ2olai03QXndt6sJWMEQfNTTwFkI4+ijJDiOlaI+JDk/N8R
wqxVYvbh8TxHFRiN4c6A62IUJous+NcXOQyOj/qt8xgeQg5CPq5InM5Nmo0epEHO0A89LsWm3hkQ
lTbBVM7kkpUmWEQnRmOte4tLP07SD5Bz0q+J6Ljs5mm/m9RtPTX4caOHVO8oGmoUa+YmnO2Bl8u9
nhMOIMxn3jIpRtT9sDeKDsi2tX4os95qERLCpM3U9QiZF6Q6+P5lXNMDuQnq9O6g8M0sQY4wJezt
bAeQ+YXWYFBfnaolDZ9iaXn5BDfTqDoNBqyWS5iJpwekvNG9JyqoGAIhpPIVLlQuHkG7Wf7q3yTI
BWpBI/brG3QD1eExFFACQMerPtpspr5MF3U1/KEn2SwtbU2nVcOqbbohOduyfNYQWo2x6bFkzRyQ
r/BnaWtK4PZ+QpjgaOjQXRjDuGOzTsgCpflhjzbSVazEcvDCNUaIpRRmQc0V88uVPEPSlZtN/u4M
E5VIm3FqB6p33WmXMwtKFGs6GlEMQu4SsmxNUgdTQElifUahtCnCTjt68cTTIoZJRMmjCsyUPNgx
9f3y8L4ToS2v4hrA8sG19o8i6t1jnjlGEfLtJk0uzoJDCUjdwNl/Urt0PAhIxZTOtmaIrM2ckjg7
Oe3noTQ2EZjxFWp2YvKSyPJXTKVcqbq49Fj9je6jqoluun5XOe09slWayoo2tEvF/f2a05oIlrU6
NOEU9wW3v378ex+kx7K703hLML+5yPt9n3o9F4aTXriqDZ0LA+9C2tfgsJ/qeCL3RjrSAyKB3LvG
ojnSIRRjssMcC7D6YzHOIh3l4oy4SQECnFJhPLpdmw506hio13gFVz5tWiTAAfOGrPYPdOF8ltxL
0cPOpR/rQ3MFqbcPp1deWxkwu0wZZH2kYqG6A1naBzA8aYbbOY0+TkdcNFTo2jN3a0ZPq/n2U2gf
0o4vtSoCKcj2qh0IJwpIjkHalQbsuIpb+FZ80dht8rgudTvOcnSSaCS4nox++BULFG1eJSTDPJIC
uK/rBIyCvIrD7zuZBvPMMOZswtIJlEe9r0sK4TPG9uSE4Cw00IqTF5jyxddHvK8+OuibYxV24Ykr
mCqJ7IuDMQQ99RSWh6YY/UdewJAmZy3yVK8d5RlUynMWTljy4lOPAoC6G5CwBZXMqo4JaLZ94cdZ
BW9k3muZt+2X2+iQVqrzg6jGbFbz0ELIvTfycIpymf0qNwAr3TpYsQxIM0G8GYNohSWtY1n4oQAJ
RELDCrmCZowC55TfptCYhjP2rRJEHkMBIh7+jQp19/owIXPqTAxfBePmi/4G3Ebi/X6oeOEbK/zN
QEwk/z76k2uooV9pMC6zCjeMTMZs88L7mpoYHLXykw/EkS7ilO7f1aHJjgsuaoOKLeKOqpDdp6E5
ZPeEtUt+nYQtSSnROBbB0bQh1d1tn2wk7Yqf0kDByhktCKJ6pkXsndohGhiMSnqTf+YTczeg0nHn
kT57Stg+ZUZUzzxQIanHQYydPz+sEnN+KT63jeom3VEofbFtAVVupNuu3HvjmD2P3qqsaD+e1hnO
5nqim0cNwmC0BF5v/guUBUbckynvR+3GPLJvGikAKDuLjw9ItkGSQaAza4WZPjr+AgnAAJrwkaHN
ue31Iu56tD11HfIoIIdI1VK1XgPCTRaZ3Lmpe4CeWppnRCPasjdcKbsakHdBD31nUvJYM9tLY6/L
36fVHExg3vvjLyHwOsLOyo4oZT0DeVLtkNyCujUxRT7j+hpQVRqYC6vodh2vLOwWCk/VaALI3Va3
R8zOQMb2Ns+uFVi/5cCSpQuRt2teNzON2f6sliTrx4pHkAYlSguihkK4S2dbfI/sR/75EWLuT60z
zDzX+cjG0osD44qPjVHObWBqoFZGV7bg+rdGXs086r4sg2x0EGamAYddc3k0LE0ZMd6e/adWfULw
w3Jkf+TpBaJ+J86vgEztbmZAxppkjTY1v00TAwWBbGfXj2yzjvct4Egt7tk3ArmlkVBB5xNzlJCM
EeyF81gzTLuAx5yf7Idk7VhHqy4t5W8lPv75lvbliwq4DqIKXp0ZN8r5UB/anEorp8cZeCeWeEf0
El6nwfvotQJeVX0YNAY4vi+MqEyXO6hyfs1T06CdoUe3vVpdtHZbAwfn/X5uldwpf3Wk0WOXC7Yj
RzDir0+yBTTIrzOYiQXk4P29svbeFZl5lHqSteWva7ZraCY0EUhLHAll7HDu7j4FtrB6E+ofAllG
CjZz/4v6piT16zFmwFBbtkNORDlUbcSSinqfGrsCXsDmZK40fjE9eMCuBNA41RSuqVlcClDQqtB2
Pp38kT4V5pl3HtYnieo804UM8Ls8lX5HvzYqZ0wzP/D/lJBx4UShCK+7hDGHUqB3tVr4nrLopEJS
xxlHpYWYBrdWwXja4wA234YNKe6r+cK4I31glE5mzHtbs1DoT9JIOaAhsBEFizJjE4jWKb98+ELn
972+oMbuKm6xLTZ6x0zF7lCU1mEKrF+caizPYQrxlnFZCvv+Fv3I9KCuBhmNMCG2kX4UA03Y3R0M
PpwxHc4I6D206THgM5tVp//+enrL4wep0s86zWFyIxXJ2n/R2KcDrwuv6RFcIJlVlSFibQeYVyfs
JlwLM6T5dxd70Mp2sF/pIMH7O2vWoh6da/xy5DKCcNQQ4u9yPKufIvwCJErIIDsTW04NhvyqVccS
xF0Q49IHeSMY+Or7UL2U56nZvvaHJH250nEuW0Q11Z7TOSXodhiJKARXyCH5TQiuwLauclcQPgLY
jhxjYZZax5tDilfbNRRuqqJ9iGoAiB+TK6Ecgs2t5BNll9wKAhdgiik8VRVjCdaVistV9fm9N9qf
bShvAu9vBbJ5vQlNS0Npa9U3jxkuyn1OXPvQogrcD+FOIDTlnwdNQgOZmPzkhKbKWr27TyJtVaPt
7rSMS1eT2t0ThIXFa53IU19H5Qr0hdeXBvnj36nUIGPAKnSdK390RQ6FZvIA+BwKDkDd08sBO5dO
BNEanUNtHgKT7N8asyQbqZnJWV7oDfFPZk+zq9Ofsu6DXKQ3Yp9gSj+hT0qLeV3cwj+Saw1cM09P
9gA7ejLdZpbt4p5LKiG+8GR0W0g4AS516qScgJQI9KWVnGE1rrn4OV+CtiBYYawtJx6CvLDjZ5jL
90qpURXZMLKUZ0sIaBdGfhKtiR+I+mEYbCm6UfjjmWKD2JORd/8r/15cGtZkUvu+y9p8hhj2Bprj
xrAIdRieE0D5Oa0+21B8p813qGMwfpaEAFtTamLy2zWq4c/KCT0WJpUIRha6p8D/68kfDKJjreDn
8zwSRPWO6Mmpqle55XqOpAXyac0Et9pEs5rmTSk9z+WD1kTsgVqaB+tIznWMsug6xwJifBinmEnl
YDYsYEyh7+yXX6L8L9r0vjJlYF1LjxGDdyyQbWPz6Zh2OS6pWldkSD43/RPg7NWNGJvGH4RMc8mZ
Bhus8a5FAUPYTRA7a0FBzBSDcfVEXDnTKT8wVkBI110+81FjJ0fSCndftet2G1qJOv3l6x8YQhk9
BmAty+AiHtLJuXEbQOVWMCLj47DK3n/rKZwIJu+hf1AIhuJ3+X19n7xQatYEG+P1L2RXkxRleQfd
rZRSKJOEGSVaGDD/Agh4hwKHFZIzWOxqcleFtnEtW2kQCM2zaIfWu5m59LEdkoJgNxTQz+ZF8z2S
EJKCEbDQFyA/WzIeQTv2zGEQBw3j0dir57FjOieCaF0pkS2OO7XUncSaUjmrh2TQ6XJldkIc8ahn
ksbSdGg1PIUxE1JYet7fcnjAaNAVu3YB6AwV0EMynQPrO5IPhjZYk+WoP1zH9+FnMchcY5Eridm6
FsCgZi6s4GB1NateTrTmbNCTVzvsfQh0TKittTVZJaLDYbKk1kEeYO/KqdVksNY1rT38UXMQBRf+
+3Y6zrZpVL97dAwv0wXWODsMdG8KP3fejOOKcR9j2tr7Lf8UdbXypo7vJCVP4jb3Bc+k+OG+sFB8
qfLwz331BGrPjwL+aU5CK1l8uHz3BFGGsGAo+2yh+ptFyWyBcslVgjiT3TBDWMi9236TJPjmuezm
u67Kf22t18VHGzhZ/vQxxLavndyXwEMOOPgNCeQ8C6LF6sCch2CyyD0/M7Eh3YWtdMYisKY920AX
uoYYdX9X/9b9URa37es9NUzM8jHQtx6+GWPEzZm0wUYAIgwwSuMzKQ+rUHLMumAFdXPYtnUGwMRs
iF0JrFN/Q5Iye3kBCWKoCpp73fO2ZszlfU+0bh54puD0aUHWLrcCb8BOfoO6jeNJIHLylpy34R9m
9LaygQ2gpDmUdu+MIqGfU/eTb4HmK8u7K+ZhfJq6h5Ap7duFQ+u0abjCkIyYbiYbha1/PyYp3woU
eZIPJh9N61OhRcTMghNUjTOE44RT1JAOHOJRc98zo+V3PYWz8O0dvxOalkJpdlQ6ejaw/CbQCcxy
PpMT5Tvnfe/MUDEqrKPkdUji0DuFw2Hu0dkxwiLlol4f5XpkMfXTr56Wu3IrWm2zvl6nIcuz2ArH
bkOMYjnVp880RXiheCFEhB6VH2SVNS7uVzcfrtbvP7bmsHkkmaE5/njBZnr66XgXfhaL3V+UIi+9
A+brerXq8zjIVt1zQRpGdFGOpY4oTXyraTaH4Vb6OpToiVsoXhHGFR+3jasf0JAXxffTDGhT6a4W
13GfWhnMHUeBTZSl++3MxHSMY6hboEw9NSe9UrIXtG+VU+HLlgcgr9MKpjK2trXc8VmzIvlSESr+
PZ6nX6/1B7QCAIkOshwaVm9sOXQq0UDWr9dkN6QHcsqu20gbJ+9fus9eOTvhiILMl3j9oGQLAwGS
xjKGx241w1gdlCHKxaBs8WILezJV7xZjDWfLyr3Jp4reGusKIKv4SAgYWxgPoO0kHTNE98S7kotU
76qaTvLaMU1dPK52r+3E+ESSBBQ0jrtN43zluhEjidRBOQVZYW6XazxXdiG0fh2P4kbbApt5GUMn
Ldwk8zsqVL1n0CuJ4Gy4gWgZwllq7Oe8hG8fMlO5z2J/qTHkrrK+GnNp2bpN0hwcCCxQCA/DSmG/
eRM1dNfVYmOyDOan4XeUAOR7TLKhFJTjxB9MvstoABqOZNLTVipeJhFWRNJePjV3y8IITZKv73pR
shyP3y3MNJdbdFCFUabzdXRC7A79rPoNrb1JoyUYg2LOQ3lgh+oez/F6U1PciCY8TONJyFzIl0Oe
xRkN/mDamvoLddOjJUB5V0Kv1mdsFB2A3wWpckkm0Be0gi/Og/YgZ8wfL10xR9U+8p7rqFWpo+Df
arJ5zy3lv5tJjyXGXRZoxLtPjmS9IFP10iM0NrQtLu9vYzyE3heSDy2thBIVSOWgDebPpg3IpL17
QP+g9xZKSmSavi3FB0jDO4dYGjJguFwMvjWmZNtx86RXuyFd6St1+QfuBy+gTE8atW8eTn+UTE+t
0KipNDHyVBZQ5/11yUI2i851ZCIFm2dcBAHP28MlyBStUSFKWrKPDz2ugPIoMUIywYofkos5BdDG
k8vyPEukqHh5cuEh+sNwbyyaYn1B7I8aQAlNw1pfgHe0NI1UANTWXJA89b20Ho+4guKhKIjniUSw
uUManz2WS4Py5loucqDmNjwW5bcD1nZ2C7++CXAVJhERYRSohNZbO5qFrJMLrjSyZZwZO5ILMwJZ
s10oJiCQaqsyn1fPDJ4wiEzBQ8AzUGONM7PEIDNMpBtARdv03Wbgm7wnvHOTih5WHX+8W7bsYYnp
ls0x6YszH5wOYAj9nNZHn1q1vRntQUr0fWcqAKIV05eXrYaqJv9u0ZxldO0IaHfd93sLQI0zL5v1
088zvAq2lCFaS+4Vn61+xAPm3SfRf0J/56FJ/vRSpswOUBtO5aBN/jmBfBkDAt8+xFkZge03vo5Z
7nwUruG0K6KqxozgPtL73r3C/fBpS8ecJ/5yDm+citd0sQFQ87lbHep8bMlE8nPE/zVCyr7Gvglk
60P9l6BreyhKQ12GpdtcMs6RViYT2wTmJ0qwWSp3kmH9psTrNrDJNIrrdvWilUu9X8yGvpUzLtm4
3jrbNYl7Yew+Bu4ymAk4rXQoAsvw+dm7IpcjA2GcgW1elxMJDhbtVXn5GudWg3e5WfOVindev1dh
zAynFq5sP4W7TVnPSPJ34nVOdi+a3C3bcueMc5GYYZucKBQwCofaG3EZFVP5aXW+xBo85+3qN5/C
AW+zbW4jyzOchVGvEi9zf/5tzXmpFK5KCCDw2PkeRLFAhm5zitJdWOSreI4Tj88cGB8rvA7t++VZ
Ij24Wng6OwRLK0kM1cnZBHIbeiVzGcWGXx7G9Q3MFRHjOnh0x0vphojZK4Littb8utUGl2M+nO8q
baHldF7F7FTfuarTil2WFScyvTcex3Ntj4425bYHKwDU3vcOP4YCTtxnsGCenNzpCntHi5JoOLFO
MCv+pHdB0SW3oET2othiiw0IOgUG+XsQK1AIEku/0IumOxWhg9pNNlNYnurjr7FeOo8+/3olUYOz
kGaBP5A1QSklwwv3mqOTgEUGjswQEN7k8QQD1+G3PAQg+Pk29/BnHpiMWNoqLmjIOnxhqzhADQOx
y7z8ZpdaA3p8uzog257wTzZ9CmPKRXEdaFNUvVEC3h2YoDROsZ3MR/+fcRa30BhNJoYoIhME610z
lsdaBGqKhttT7moUdCYJRrMo/fNZ2MEAJADugeD1i+zTrd+UuE7JlPB14sipUI+sxStiaeayk2VJ
M8wTzEGsf3hTC3lohARlA7M3O9DTNVsOK/QDR1fUsgGsEr7kTuywSNlStf/ovPHvpVvS0uuowjOr
oMEP57oG/CDpgKedfjwQytPPJpMO6/B9n5VsE3Hzmh0yIhJAfuvBkfDOGX3ImgwnRh7Jp+Ttq4ev
iSSfOW69E0LFa7JQMiLBoUh+gQqMCfc4nPNbVx21lH1RPYnTwLEr3QSOq9Rtv9W2gTt/xiZ85Euu
AqV/anNllx7g9IibQZokuLk+ncQZb4o2RG2Qn+uaGieb9af3yNL/MdVisukRt59/9rJHnnZfn60J
M36GDX3K8T/MnUlyLoE0viRTmsvn4LkXgosTbHARqMoFALANgoPIuekOxQ6mbJXLoRA/dwh0puhI
MWODuY1eTitMDYwFNzPGrBOjCMnGS7WAtj+E2UyJPqVLR8Tc2jR7CXKMTRquVfKyoESLqXLFS4Ye
keOERf4nMNqIvDyPj3cQnSOc2RNFt39oM56XF7e2V5ciIk1OrkNy3xNySUB+uh4A1WemlvWAxiEz
+54yHqnnrGE8TN0C/FSgOd5qj+PACuyH1tn7BSrEio6fZpyIr+um2gI4qrJqfRt3IzLFYNAv0yC0
zdPoaOKxmPoEUMqe26gDuNVsTLEv4lghblK6av/GzfGIBVd+CVKcPixM1OYQgp7rtuaCEAmW9FAU
5gQmbXy4KECdDVMcaHDgOmJpn1Cjz6RrkiyV7ddFMVjU2EwKDxSP444tTBrSMxmqRCv0LRV/a71b
ZJg2Dg4ghfxcmdaXGObw5pmN2lZU2MyIUPiU9Ka81lzq6IIYOEIdjBE1Ek6l0Msx9BFJnTbnm59z
bn/EihAke90/wTiKS4ye4+fZmGQFqzpNNX+SFC5u8Mrg+NfkAgrcr78nCJDixgWwmN3UmCEacMay
VwN78lGMBokNnA3OjRDMihLaRnnydLDWlNQCRrvdH5OBLLyydPMtDdrWpt/uuKtuapszlj1t7Y09
FbjHOkKqCHnlye3roi5YDBnb80ZoNkChS2W0bqQlk+jopjLGl5bHvitqKq0WUmmSzrStFUi8OBOD
a1WqiVXLpWOp9OI7oecQoRRs3zQkB0Orj79xrOmn2GCgqO8JIWsj4wb1zopsJByzFul+z3Vj0Zqn
KDa/oEJHTkO8AHuqMeeMtpiNn95TmqJKQ2saNH8427C8mJ1R6aEoiErDTjMHuuAaBg/8qOBW+4AV
SMXK+PeDJYVuPLMByDWAOmDgh1rbH0RhBjRlFMRKr4vSgYASUmUFbSvntNLLcwSdfPntRVP9nswB
Wqp4b6mBOO5zdtiG+d180HnC/Vk1BEM0f/JNDzKB2WMZsgKkFYITWjBuWuf7znMC61hniI5uiIZj
BPJtQ/EcnGJbqc+UNiuSqYyYaWjw56mPao74Iu/eAXD+Z4yRlS5Kr0Wdy5g4FPSDSsYYPtMto6eu
n2hS5kXcxaNY3yetyzb+yc4OGPvJ6n3bb+6RqOd2n7Zh5Oa6eieQom6QJV+jldSqXrcJ5DPiBhfx
hPVq4/G89weKmoEyKdWW/fZEgtTd9zx24pmB1P7xEjvY48TwWbrnuC+jncKXFhcOuLyoFvKdYtVz
iR8cJk19X5UbRUmTSayARxHvOY6c/ky0Jd4JwV9IPVeD8OYL3fMr/6sa8ggPb3ZnZo0Vu6hFtc91
K3arD4nFXMd79BEiIbdPeO71XTZkRRJQdam/J7Inh1WM3sRF2thgLK/cfR1dQ2r3rQJ+hKe4xEaj
c21BDrn92KnbmIOij9g9lf/djXBI392BYT1P1Z9s0xCG+aF4r9ltrlN/Rldnp9cSBcGEWoHOPMog
XAgWDwY2lyjYKt7RLvZNXjLp9WspIqRdIpcAX3j2tgK24iQcR9c96iDA4BJFxnpegIbVlrIkdZpg
8+yuBvM30AtoTmu1+PlII6IgIEVVNXK0Zur9KEHC/+5i2SfyfCP0ZCWgUfLcYvLyBko9Ys6PdqTg
k+eNncSuUeEnb1IzSUOLPXDLMCYVB8mVyQBDVuYAJTsRegg+JuHW7YBI++rbMCp8epRdfcg3JuBh
+Yia+UbF2OZpdPIYRzuk5xD00eok2l/wXOse5KABdX7S9oYioKxxoJ8at7y6QjLbFOTMCp2GTTg1
+5VMDlbt+z/VG0QLsYn8DNXewqba7SRn8KoIhvd8HcOTv5fUwBgyG5tRuIUQzkMZnLlEhq7o83ad
T4AamWHsOpqd9tNrqBcpJDvU0KP/+1Xpx7X3XUjX5j073ueMS7SKucfgJ476RAGUFjPlso0y0Fhw
2cQd/S49Fm6P2TSsGdCcAv+hqaTe+PrQAjdeBKYR89zVo9PQe8nF5Mb7DHecrsiO4PCr3OeSg1q7
Y0/4hOvT6cz4Y3EbDNKpDD4wcO76qOj5F+WiCFfs/wfz0uiqqYL+aLEUCB5Ye1VdY6OUErDFR1BG
byRnOP2zIrXUpM1paFnpn/+PtUHVzNQVz7SqjPllpQlBk8/coh70RxMXuzN3E1DaVwXN/Y3uKZgO
DwdPAjc40F+1ej5b9ENwYOP9Ws8xk8L8ghcwM5C0olFgCXnnVfcy11BFfZURqMMdZx80Qwt2EgJ1
Q5sOZiookj97hmv165m9mW51++tbNcSUYx2p3AKDvpbdCuT7F6I8F4G0QGQJnm3HZPzoZ50MArLN
99u2XlzDXmvGvJKcz/LSg8g0qzpZROryRXRmD0WGSlLx03rZ00kiZ4A0z6BezPpgKJ57pWVcNIdX
r9QAKrFU60+FqYNS5qcdmsAjUQT0MB2SLxyfbJ59+QvjBkbgKZqPcHtc/EnAR7aki0aokhHpGaDo
SfUj3sMSeaA7XLGzTdsTVgEww2Ori53mIwKA3Yf31dZlgc+gTCZhOSXpevpzGWGKW3ii0Banx+qJ
XEPssnxzdIYnvVRnB9QsU9TS370s6AkKGKSvHzxR5pncsY6Y6oF4n/ihCqL7wQofOHYUO/ZxTVWR
ZHSeP1Bqn9tJW25f5HYD53zjoLZdK1rY/gCqWvRyWdjKAD6Mj72GkTNIxQj7QLDIUBxH0d2pvriR
dYWfNUbIF8Q8dE0q4CMENxTFgWMuxyQjr+juhIqrh9yCCI6ORjhTUlMqudVnoHp6U3XwtJLsGzF8
zD+Ry1wr/if8iXmvxUw5uiZmoJwlmLgmETMMsc06I8O2qIycBCGK3E7H87vaBLu+GaYioO9FfJcO
SpIh19W7hCEIzkDSoGSIOhTOss71bfkrpveBjyZuHLv4H81gJTNxWnCbz6U6B0o5X5i2cBoLgzh9
bthS8Teao9gpgQhR8xL+S5e0hJ79x0WkONLb9urcnnIFw+y/NjAv14M1jhueU9s9WInK+aCzyigr
fP8FKAFoqg8tFv5Pv7vu/b36d7qeowylV1A8trZ3kBI4KIURRdCZWFEErrlb+A1psgrSjRRvElj6
LZHMlCTl4DeRGvEWLX01ERGy9j0uf7Ugjl3yr8ypFBp6wbK5AgB7h3z9qKfpWzSMCLcJiqmVPHva
ZV1xTypr1431jzJH5FctKCzrXhVgqzwruGEp3I6VizcHPGVtCn0W+dIj7ErE8iE4XX1+fWzPXSVK
GVILX8V8eQGQFIz5mEduzK0GAPKAzjOYAeybomWnsXmFgZgB7xsMBJLoe0V8lvRpXR8Cw4SsGGt3
LuRhb35pQRwUlwHJCnD72MkkxDlXL6jaO0ZhptsEhgl4KceKgLe6FHM93dmI/5UtnsVwb8VgZ0aO
6EYDCr0zXSE9/xWYiv6RoREUvAvfPFiqeAWH/W3MgIm83zBDwIO3YFvgRZdLWqytYx6tbnkeReAj
Hc0aKgckT1k+Yt0r+j53GRJLD0FgW6gBRV+La3f253AgasCY6Pn5Q9zIGkGTTdhJv+jY6a60IFLR
pFK6IQLfmI2JjJtgwaYE/yECVfLhTmmrEEnKjSTaLOUvCN4VZZ7jWn+QNrW96OkXyfLZZ5JrFeoI
gF5l75Iv028XpBMhBHnWZm7sk4mL/tUAQCPUK6ACjXdune8DrpMJTwXvPJs87hJoICQ+J67M8i3v
pZU+Pz5uxYHtExAx2lyBt57Hgz5Kw4BNBmmUxoC4dP3KrNsujGJa9d+dCf33FEU7BMkJyLeo240O
Uza3vP9ZMTFOrawWjg1t/5vzLKex0CKgOjJexCeL5AUhrlRUVJT2iF98DqAfbryXK9YsTIEBtcuZ
SxTRd3C3eWOhoVFNsWrXoM3CJGvicA89dezDhvI1tdldjyzCixB3xedH9kO76OQUPs17gaWVfEfo
u+W8dGh/E154YqqcUDjZ8pBB0nwB0Ic3BcGsmKdg9JZ14zTTrxwNE6qtDN/YbUXFm6bHMDndvt69
qTZeKQyhAEs1y7u19LQsFShQ+5Mf+5N5MloR2SBJiC/MCnBD66lfafWuJ+HeiwBggj3R/sFdEpMx
+DhwJOhMEVSihg5VIoEFVvghGc3CXENHYkk7s1e8Go50/K8pfnTwsygPVNC3/s4e6HHrzFyyAEas
ARe+7TI2NGL+LdhNSKn7um9LO/MLKRN+8uYL6LIi7RN4kzkjwWZQgR/ep2tiFneFYC+dXmNVY9zJ
pPYpqtSpgDcxtf696YA4fT5Uj66tlj5jnUDtI+JDVnk3OtqUt88avbypp078eztHmsReptz3PN73
0i8fdv8RB3TipX4iKWMvu2k7sB/WLE9KbmvR6kxa1TmGrywVPy03GgSkMwKsYIPn32p6G9Bb+DDa
Qf57Lxv+binWiWZlfbQXFsMLjXq0JnTe1KOWBgC9x53IHce8+avCTEatuGCoJCJIhiVQqM6kKwwB
L6N9/djjZ4amACX3xy4KDPj1TBx//hjTydsEch64XyHdTydmfAOB9xw/eEpR0tRq4ANkJgNAW7Nn
QBYaVHGyLJL4uPLjl4hXt9GGXPANVxKi4TRM6m4EYLC2EKWPPTynCG6j4346no1EW4bvOjpoBbp6
bTIdeAhtI81ho+N4Rw9zQMXRZUSb94LR2u0pBZmsYE2JbPFbEWWtoX6caeVSNvcaTEVKrYQdi9Lh
Pm9gB+Rz6eylz1DxM6dKsRqEKmOQ89Znh7Aa0QhRzVUKbTBvOJgf/suZ0geDrOM8zmdfktw5pRoO
ZE0mFmvmniKO5g9ZkCYsNTgbD4O65zBJZhErqu24xn3l3CaUknxL6xCHIGhRiuTHve+rcX070Ka8
ZN61IAVXP/acISrkFQ7QUgb11bmOHN/uO6Q+FSxN4WvB+sKF6tX4cg5wa0LQd4un19mjspwdZTag
VPxj02I/HxxBHd8/V9WgXNKzFyT5sFQGbux2NnKgKA4IChODqhuXdLr7PJmOJyQUvNh2UK3mTDoq
urwDVD4A1wbKlhCEdrRqvf/8tfnx3sc4Jv5yGKPWXNpl7PhEwve8AYpkno/N1jfB/IGqThyxSoy5
pGhPWxfxJ4APmPaVwS+HJdVALXEaKmSX35N6iY948moqES83mcfUumjlZPD8uVnRklm+m4MqwwCM
MpvX7E/Sxk39wHaOi/ocQtu+FEMZd4aw5xwgDZ5/ZB4EyPq2EMFgIN35YVmlq/1lYI4jdkKTExU1
KsYZfiPUB4T19GqB33wbq1CvwhSqLhQpL/6ew1sW6vr2iG2ZDqq/yS7nzO9fjXEsbBfKcYfRu14W
n07o+qtYd2+BPH25d7+sy4GGwhyBhsUFgZuCa0NKKUFYIJ2biqhMNvbu5eHobau14/d0XA4AMcIq
JtxsNwYfCpZ5zbJLNyuzB9zhsPTIZ/l3RGhW4kxMxI2wv1JtXiU6WoAcSAzPCDZmN5/a/b46MlLL
96TuhhNDJKA2FcGfLEIOV5XeuiqhIRPhBtQFfWgV++p2atKe1iTly/uzhQajMVeUSxKDI9C/znfv
7CmlQQnk+VkQZQNIhHeOz0Q79SPu5dWF1jCNQVCpGuVqSd3RRyZgKuFH0N+DLAUiXl28Sx/BxewO
IiC73t/+IUEGr4nqHqN3ZczG8sGG7BHIj6y02j852IcYkKsdz0Nzq8Z4oXSRArBDaiKY+1x6sbhm
mCUzXRtLRTA5h5ehd5+nPANPFYzBJOqAcw686fq6SY1bKX+Lgw7vbhK+ax5olqdlLEUu7Zvum/pO
KBJOw8A0gBthXXaf66b61Jj3Lkma5BcZucYVwDSb6x8cRti1DbAm+BjoYPACWhx85INmJiDLH4F6
5V9G8qjEONsO0K2OujSPPJL7mCQv/F9OeynDgZypeRB1j3p9XBNqHK/4gVIXr/foHa5IWLQJLPmA
kUvXMVnFsaJkVrKotZI6JoCvBsIP9MqxWGfebzpxhOgl3V4ObokIY9DMhCfnZ4N8xECnC17tEUrm
AeepTf5crbXKg/yVDw5PTXKiLtkqjGYSYAaC3cX44bE1cVqPFBb55ghET6S0s8XtP9dpH4A1ZK8b
OdLRzckms7dDpvJ3keqow7TbwGRRU25Dts1+3s4iUb4SToVT+4IE2h8CuKR0Y+I7yZuRJFCdoTSO
+urwvxpvRMBFVxfbmh8Da190Ncs28f7Vu/XUdcp2W34VZbHPOQfJLfIkfGz1joY5RUtwnKRO8HDM
zA69TJycy20XaKz3iJy4PBIt+V1gVZ1ZX+JwFwlEa0hif3Q1rHVg/QXIlSHvovGoNyPZErC/C9kO
JlyZ1RnW9FNJfQfJJqxCqAujvZkJU84mlCtMBr6cUMJfH0oVV8F+YNK3sWHpit59ohH+8GwESf5d
Kz+eblyShirF1ISe+x1tcf/C/bEar82wVx9nxP3ggmM4nZhrk2Z1MFO3NvOcb2+iJk0GUJmcI3HD
u6vSgKq1LwdqbPDjCJ5xvxz+BAnV6y6YSBlshAlPbOrCh0hhmY4kLeBmuOosYRwR9D6PNiq5OzRe
g+hoK1b59cJsCaKPSyC6pz2DD2A4LF5HycjNkfIztkdWbEaH/eVyb4a4oftMhlPXXaH4EL4rGkTo
MWD2PckvSvSAjZNdGF6MQcssckbJhAEa2Jts5oPEuMGxR7PPQoMmrG4W+za63q9GUegw2lLTrR9/
tU46ASUND70wo18X+ZVJCP6ETzUkk00PKOF21BnfGb/ItEnZcIwSTQ6MTQLY/XbdCOeGsmvhHzR2
cnexq1vM42EQ3dKZi2Z/qlnAyBj/ola1IZ/Ye1kN5HjWxRr0R4BeN0TIHsNleH+Ih2IXIemhckcY
NRQUNEZjiD/HA6fUVgjcZbpBK9ETlQh/JN5VUqRo+k8udyW5gIjttxWP4YIZtPKbxEPZl1DLxDaB
GwqD1ktUCi/PwR/7ei8cuFwM4rjoVTellTzCOEf0/2oWA3g08Ez/3ACGiIyz+ZNgCNfnafOI1RX/
3JVq069MByzm9D7i99ONjzLIvCMpVuc6LOnNEGstd2wFNUbdTFSwSAc5UK8q7gRQcnYtQ+FwYYTj
mqQkLQ5uKllBHfPPRo3Smn966WfJo/tML2Mlws7WsOH1hpzrHC7PaY9hmHzFbIs+IDWVOd4yuitp
jOjr14sRiUSmVuZZA6dnCkE2o7VFvEdp2tG5hJzAJQpZB+RF8gqqN+2Ls3Tsy9e2x5cp2gQujqMP
gen6Au/Uu11SjcrtoJGP2HTJZ/l65djf3rWGK8EudgrNoNgWhsDpjttBTuWWo5uki2YODE5eAD8s
4lGVH5ZPUwtPf+Vc6/MKkMXgcXOA0gS79eO+MLFSHhbvmNT4NoS9B6LDYs0qlnIp4mXn5iQOkfSs
/eww6JOBFhBScOBnJXtrHVAnGqLGFOONH0u0GnPInohAWTiiZfOzW75UJfzy07KkQ8S1pHjztLjS
K8g8aqbNn7srvSS6rnO9wV4/y/2Sg3uS7C0mh7fP0WzEfE1vOtMqkUwC/3JrFogOYnd4OfRmLsfj
vtw9n7Lyq4wzP8YfYhblzeHe8HWobum0knBgpVSeXHxvVbc6ZlX0D2sg5TA4JMaVhRZPglv4/2dX
AU9zTUn2995ZwC7LAjE3YII4F56tqkN4kwdmg0zFapcvNb+tK92HTmcI9t99clcWoOjAlPwGPYOp
5ehZVt7beS3Bl5PdIdxtG2dtx15NUnEv4EWsqLMB/03Nl9UOdXMIAqfKjXKCek6bpk3C3EqT0cDQ
5njqfKmEFQ+vNblL89tKpqTEg0P6SIfehJXFC4b54eXm2wUbtzRU/qfZl+qSJXwsDSs2dlYOvTn6
Cgj2CrRC6Oat+Wmz/fjIT5ilj6/D4mwo71Z128mMTNrFUQi879gLcM52nKwuQQUPH7u/3NZsotp0
6TtlUVvPPcqZoyT8W+yYqaolVdeEFjwTjFa06lpvSS1k9V8Uat8Gx/wHxOPH2bdZHrnTHIXcHGNW
0gqKC27tuD9klZjU8pumaEa5hFCRfN3Lm2ZK0Xr2lpXb6BukytNMn7KHyCaUfbm5tL19DJryVYn4
sx/wmb3rsW1CCOAu/YoZ+5pdVQnE9pPKUra49qSLC5NlqYN82dxPNpWyXiXeK0uIKZIohBicbH1c
OMij2PobeGp+Z1YcmUw1Ml6poeujlpp9vq4jp/F4LDX132vfQ0MT0KZyFUr2dnpp5QetouFoeqsn
X7f8zq7JAnSLGy2Vr4wSorAGxVFFV9SkXHcFermwTchS6F9D6NDlI1v32Pvwfs251shQyK62grOy
FWnwExH3umJiEKgCf40A6ojeL/Ry3vPTtkBjchjcuVL041XvCz17eQu+CpRHxVNivAbLAPFxHiDZ
i8CMszNIM+CMhFXFUg3afb/jcPKUzU19x9ttmqT4AgAY0716OVJUlEkmPvB3/7ZjZu5D9RpZFXgQ
W2UAKsxS19gee1OPOtGx3Tc6rdvVvh/PzTA2YWHcgCIx3mmOzcrun1Z0Lr/WyA7U/98/TW/swvCO
CfQNIF6da1XjYeQuj2aCvx+dLFembGNojP6I1wGGQjtN3zQJhUvFswKshNl6Z1/tVPsMXCL++oJJ
QFf06Pf5gyAUjvb8OaStiL6SuOfcQEyIG7hAD4KodTDINQrVf3X7zVE61jc+2WAtBRXEf3RC8uAO
G6g39AFbpXGrJQh71WdqzUYEz5MvLYluO2kk6cBZTz0ZTOBoyITWujTUK0/bz9cL9N6EUwMEw5s5
tzKzjgv4WsKdUjNR8XmZ6p67O2nndwl5W7NeugtM7fgY/KWEopIdOlFkK9HCd1aspHIYJmbOXU0a
sQxBmJAJOffiGsdI1m9xHSCuLHR60lLvhhNP1LeR0ALApaIcZ7Q5yZXy3WxmoQtqbRd4GFLg8XCS
WjzT7CyXzjmbQxpWKgLPedt0tUZf4ahIknRKjKWLqoYoNtn6nVK/V+hJJnQWyUZUyEQCguSghU47
ej6XdDlYVkOtijjy6xq76W19sIkLp4fNBChTIBeem7SI0RuFQWdEMgyfJDX9NF1Qde7tNzkLxkNt
zj3amIoV4UQXhVHOzF6Hk33fkw0gBqSBWgZVRdQoq0D8pL+yT+m0DAXzYDVmA6RMdVaYn261xWMF
RN8yU4mg1opdUyJlev3pVG0hJSS2ptwCBs4l2oPRiVhk8SeCI+c5T2fsUlSfmMYXhYvfKfaR3xur
eQ8At/ikmzE76Ain6AT+62Sb1hZnwcdo9rShTbDh/n5qpzR8O/gbwcsvv0Xx/dicspCvmJS/P/pb
4XElnhf6O4fsKtPSOxb/KnZfr4gSPCZukdnxGi0ZSBa1Dhh7jm6u8AmDej4Z1hL5lWFf2f57qR+9
R5hM6wmAR/xAH+NuBk53U8ZovRUZYei22Dyr35nr8Mb2S2mKfANaTBhmMzg4mALuipnMgpEA6BbI
cfr8euQ5CnkSny0i/z1SP95qh2qHtFzduyk0d9iMi0/6ObYtwkAhelsCKIVgEN3wTIPCPC3bbuMZ
GPob+M/aDMuB5wTulykVu895DCjAjASu4yjxoHNLRPN6cPh3NUq2znKCitkSfxBdyUvWgb057Bd5
lNVKtjSdr1erL0svPWm2w4TCcV514tQ/y3hQA3BGGutnQpSbKkH7MO2kVYAe+sqJsIaBXwVL0J85
L02kyA8Saz1urpuIyLrer3uuC2UA6461BNGE8dgRGL2Kj8WPhKtxAGV/2WjpQ3dyIzOSmLAZSedw
2a5YSkSUHeqCvsCEpJ+oyrxN6nxpMna11so8r/gWvGGp9oq59Ow3GPuglbR9UpWxmaAyFsVGuHzK
+1oDPOV2QiRQWTEbpv8Qsh6MY1Vp5oJS6vjA2fvEPM5oXrU81sntCw64VtHZR1urTIhO2icEFjvo
nnZdl5n83Q355hVm9gi0LGEi9/Wr3zErhRoWFVDJy2kG8VPOrifBJSRNmIUL/802UNvfC2bw+l26
YINxZ/4swKGUNwPrj5RQMKKcl7R7UGgYgHYr/POLef7oRBnO+dLGDxAxmm4B4XlDaOkTZXzjihYl
mrIKD7nJZrXEnnUDc6aCVmGmSXo9/GQCyFlDq0GcjP+QlInVHgErnZ/OZkULCsIvTO2MuDcBWjam
31IX+NGvsxWNpvFToERNs+Eqi5qCVuIVIbbWnvbJSXO1YBlZczD7EQvJjewHsOfPs0Xr7ebH5VxA
FoBcnatrZdQ3ddJhy5pnCtfKHGlQFp2/3GxoPju2Ar1+cQIBYFAHBAjuc7Ura/1nFwGygIJFz8d7
UYiubI/2iydqvoiG7Hir5IbMVLvw+Vmt+IGSlulG7zXMPpZUKjTD+AuMZvgQSMG9Pb2yMHqnqFgJ
vrpHumb5bJfWOl5NuSWzt4BfJTsZPbt98nn4/8N1lytxIsVE+7SCL6r/xNDcM4K/aypXlMQXA+Xg
M72ocYvd/9wMp6poyQ9NmAL5proU9b+qWOFlv9WF4k9+WGjoTeUJMjMwqlfNzJgJhap6ag94Paoq
IfI5g3Oi6BsCDJ+lRzSj3AjO0D9a4fGShJYnG7gaM2Kvc6ozqElfy0kimLOpPctFD7bjR2GGGURW
lLr+dm0Xj3KhdiI9AF+sHzsajtTvpexuumVpl6Tp2ves9cce73bHvwnRxAVauH+Hwq5Cf92K74jl
k3uLjhSCfuBxRwvwTIhmyAMXkveT0BHt0ukRHIwdjXjmSuJuGSWDsAIcr5H2MsWJFAzayAJS7BPn
XxU/0LhPHBi9wdC3CR9WbxV/iEzdBTMUl7HmcogxorG/SKSBqacc855Mvas4xt2eZqU6f9Rx1x8F
+wSWDLsnFqzKYsDvjT+uFyxbQGa+MSLvwkmfHl8XWWnY8JOO2XXkaJETWl6W3tf4DlhrSKBpqlNB
GnYPea9enQFJQW5amVOrA4Set+KHR3BkHlTrQj7F97c+R2ATYOayvBXdVqyJOaTO7N9hMq2TzQRo
WpO/m6lLx1EGr8cEQdp3PpNqz6ca7hxJ3/BFOGItCMEnPVZUrs6YeFVDFlgcp4Nq3UfKtuw4ZV9P
asX4UPnL8TwNK0zUIf9w+JTorq92RSt8lrAv3Z8G4FAjEr9dOyYLUmbqnlb2QFU3VYTyD1CKymzR
QcA1L2+kHZvlROlrCOVdSYuexpfjW1FBjlvpt29NjZHHMmeeeHInrr4SYXEtmCy1AOoTsu/slN+X
WzZC810+TPL08xjRh+inbDEdBRxsypAIRgN2SP7I4JLBUnnihQVi8vwsfLDyckOE5uYw2TM3R8xo
XxcxTiI455h/x1R3DecNUuMvnpvkBpqck+OTYGGKLn9vKqCu54umEPJHSf6miLe9gtaDcTnst5j+
3/tc4J8KVKWscBEHtOCIG8PIcPKCxd5VjmJYzls7+JSe2Vbj/LpFE4XLzCWJuKgXHdp8+vMw2KSk
acOThG4GCNXByEv7RQgmAuJaAa1/GtlCrXTS9RytHeQsn4N5BdK/CsPP7PB0RWJipYbOMMSvBGaq
BY3yxQOGF3fjrKdOcmU1rri4hkm4LFOWbXA/uF43OztWgcCyhjBdouioQVvUfe1hivQ4sMHlY029
s2xnmmmp/Q/N/7W/xJsriG5oky+RQ7Hd2v4Wo90alzwVUmx3iSihp3ipdODIcPZYX5y+ui45Ag6p
PJV8SFoa5G6YAwyh2TC8WCMlMVcqihXUKvPOEsI1WtVEMnNfI19veLvBO85GXXXdnCALaCsxS9ed
ljxK05LCkZ2m7IUTtRVZ7Zz/dhXKglRSFNaFiDPZtj/Oek0rablkwgffcvNI9uwPAYWmXlEuAr/P
yqQQEMgeN+ZPxeEggPOtLoyKbHD4QvoHWK9SaX4GSondxpIMcKVrvxPBviMbWdmCEtQnEMLRTLwa
8FhnOXyYvG27o0IG1nF0FvUxtqx1Zy5flne25baL+hjRIvdO30ZLQH7yeso6qWKhy7BooNZijoL4
SY2nLpgg3YIGz4vzzAHpfFq8lG4yDZkOuZ75dX/ieBlh6SU0L7+rrnQD9Bl+OYrPGOlL/UmLO5mv
kueQYaHxFMHZzStxJ0vDSGo2cjv592NVCeSzErfqJrcC9LE0vnr8Vf2B0GPK3+xbu6wmoVx4o5c3
uVEIw3FU8qeChahP/41dbPTo/8O8Ldqh7sorjFWFlRyqr4FZcrORimTHKToRh8af37V86ofLBg7D
fiEzWMeiu1Y0iPTH6Enev1oK+kyIPi9yom5BxBdgs6DEstW7TsDXJmjgxmK56SqJR8mUDD120dmc
t642KPQnPsyHdm3uZpbjEnDbWemwCLdxAZQl4cxVxyyXx/BN9GMO0PSOxpFkaRVqJ6VGvagvLzBZ
S3KeUljzRYkSckShyZ2nEq3DxpbKVot8MVTzmGa0eJOCeS0RDKcOtVSniIlWku0umD9+kk0jUtm5
XyjcXxjBUTvkMx9/tdQnAw6aLSef3IrgayepWOJW49zay/ygu9SoT/EnUJSRYH/XHLrlCk/AZOTC
2mU0wTU57fGnBoTKTpzqkSBKPgIXJjd6Jj5+RjhM/q1cJT34igKjpeSaimin0yRckgQEqrTqM83S
e23iGm16YdTmzShviFn0dOOBWywYxsxpRkWewCflQs9Su7Af09TMhMnbUNibhXVAZ8M8ETlBU1fi
sGSgORPzj4iB8S6j20Nv7LyqTRkI5/YWt90RH6TwL5zOVYBGSiE83od2vnvsJxe2kb04NoRAgE0n
uBXkoUWxUUdCOg4B6donmySVIbL8hsf9rwDgPqlmLVXLJw92BpY4aEeMtMGXqGrNVOTWcWOtTZOB
tZSEOmXktP98xWT27XvGMOzdP5NEQmlplz5EpLTDoayn829VdvA17xpeHqI+Trc3aBQ5LzafLpiZ
8YG3It3h7kTtVTeFoJNnzPVTBlXaN5uKyHGepn5DBAYjmTaaeO5ZX+ZX7jm9wcFjLK7lq52Q/t1c
uztfRXsSt44jiipbDl34JE6hhBIAQF/M5jCNzC8FNg4wV/rOr2oi5s2U2r2OoiD19ug0OtjtcCYm
Y2DPXp9CuLuFDTIy9bCZb1fKgt3BlU84ujXsOEB/pT5VIAafkLZDsy2/EQqxSuM5mxVAlW+n7did
fDg6mLjGW2dnD5qcLIULDJ6dhIOwAKcrvHgd3m/yq8ZwXrVshve4LPgsw+pPA9U534KFt32H3CZA
nN3/bc8AxEz0BR9BZmkP4kmAFKSclbz0kmjJ9LkHj/UUTYDTqGQ68ctnTL4ZJODdfGCfWImyMQq8
MEEQTcwNkqZ/cT5I7tneOVdSXcLHk3gqfyPwnBXaV4sHXbafBbdiGd+kNuRHqdPQFYmTvU3wGhOD
rt8QNKMwDY6Vtra/KQ6yz4SEG6HM+SrfRa1EFSItSJ1PuES4f9D9XrMaD7T8iYGE5mmMq135QZHt
4/WLRRMsc/iSNwRMP5UYpcqOqrEHPBMLjUa3KVjroPE76fx4skIszkyYEkthP6874nOqCvlHxSFx
5mt9BP96+xSxEMOpUNTu+5aFQ1mK7tOkULsaun4VcOZ0CCcpmUPw0vr/vbjSJW8T3ddrPTlbMeva
4xfsq7OUHtqxaQQZfF+kXo8VeCWRqufznthkprDdUEKLDNawdIcizK53sDx/ieq788XN7eP7M4eq
yqascBKbgh2gJ4ta+a9KuMjs8t3BRmV5LcSMjK+/Z07fEKX3wdR0bFameuIN3qR5oOCIH5ymKNrv
qWjwr7OlDFLWVMB0vHx5kORKby4PvSekRkyoP4dHuAzvhVno4oRAOrVWehBdP+xJaHLkWrynkY2X
+/3LFDtRkC103AX7WGVTt8hKAl9Dj0y2VVGTxhyaP+TRCideUPtYZnorx2euvd61dC4SuxJudtzy
comqexD6QwmVgCgsZ3l4wReY3e8Y+qHw53QX0x5wgy89jtKxXrUutyxBtc6n1XCdMVbEeikPMYWW
kZOceU1Dx4NwxI8GlH9JNAAZi5BxESbLbFMZ+jxmtZBSxI6ncpPX4rjX/rpq+uqUbztDPd7B6HSw
jBkwaYrm6URULwcv333kNYisv9Yp49xXi0mPFqZoGnOy4RyIn9Kg30Ydo+WW+zSwTnjpQS6KjIpf
NmOjgrhUyAFwVH46uQcgL/Smg6mlw8G89keda5XUrBFM4DmbbEbxIXOQWfhtf12wbIx2CSdV+JCM
cWVUSZOJA719dBSo/MLj+5UDzgvALFqoVaFbmxXNmgZIpbokui/MUb/pClAyDni0DyExT7G3XMi6
FciRKEhq9Wtt4t/zb8JBWIY65bXfDDb4YEu/ICdzaOrdtIYBMmfkems9c+p/ZMSFXHmMDKSP9B5A
hBJe2CLeNB9hhAGtrGPYkarQy/6jfIw1zBSzSvO4cjDG7sD/t78zTaL0IuL0Fn/ldIR7XkWczz9E
7AZY4UuDtajYJaEMsuWoenEGGcqMN6oj6b5/C1jACDJUCyM9atvh6ceT82xWcKDsuSaed7pRlbxv
sM+m+xyISYai5QYR7j2CvZ0xr4b6hyJ91MB9roecUSQBtelwp60Eyvgdo02LgwmNIZPAzeLNXHpo
RSWs0286X5cEHj2KjoragGxTEAwyi/KMERRCZqbfN3A0CA5aUL6o+wzlp3uo7FS/rsgXBLxHMn3H
OBrLJUaMqWR//ep7PBWRSPjUdI7xx13JFKD4LHY0xZ9zSq9QdAbpN3XD4UEeTKBEf/WGyG8fNXDK
0vthaa3TDTI2WJ4WPBmgxC8QIzHw/5kzLiTgN7DrhTeUCrLgOVv5KHufTz5nAPnlRG5FGZI28I5s
f5flcndPGioAbswC4PEZ822ZIxdZeG4zXm1K8o+zvtR+IrsmgP5SHmUtCvqpPDgNxC7swoOWwcpo
5YpC+Dt1gwXSq3V4yCo+0oCOGtV4RLAfspSq7I+o8e1xzyzuW3Y647IG3Ake/J5Un+aWBaPsqNdY
vwHKZKErowCTjMxngdJ5of9gIhO49O2vXc5hvgpiXU4ACDDG2/hMyf2sNiXRmR9MNW8amG3YByPR
abQu2uZzbCRRhWGDU4gBWNVUVLIH3VP3Jk/sT6y1LkLG5xX2bEBiit/Tuk7iuGuOk21C+LIGalzA
nJ8Mk2ArFobx3dHYoqV6uuJU4m3UFK3jTfxt4cVjCAHGv1u7yt9whqzv59RJ2oy5YBADLJ+992/j
Yw8AN8Sr6lguqNiOb3gxa6Ldh/U68oVkPbV0qAMAq1pUrUeHFksmGdAXWmbdYIT7eu+5jTV4xCG8
5gx8oR0c4kGCt3ofaZtF0R65kSy1qKOIsJ/ryZxOZ9EtLcO+UwPYe6qFe3QP9IzsejFQyLukUgfN
bcyQXPvWPGnfYN93FTsThYxMon12xLchTMjQWsIux8lwQyJZy0JRyszOQZIJ92ZerJFC1wFcbRTr
9cgesGxONJ7/YaZYV0dktty0mZN9YXUB5s9dPALFhRzTr26Pq5xviQE507okyFtEf+DTTHzSw1QL
JHTkUDp+Mrb6Hdxb5qrf1627gnQ5PPwUDQneZZ+Ev8MYe8LL1h4ZAq30FbKpFlTukIgKriqMhDLC
UwGLcCg/Mio2DdfUy9X8uaFi987mViPkUm3mUzcCLn4WGMpkerY8mGQnoNtHAEiF/MQeYTwO15Kx
/oaui2/6KE2+F/tfy/YYJuCsqA3O+Rroc+KsK0Bawvgm5yjgc2qRy3iquCfkDWv6hOMfVdCrC9wl
GZ16Q0dYXS5qqE1sHUpXnA3uN+o/XjHD7LXJND9e2ztMnPJm5L+IknYY3UCjgQMh2WhKWH2sATyv
SZyFzNuPoW4qGAa1jnPOczF6NxASHNQyuToTW1dA9ELhnJSahe0cTV2VEnSxn1/K8llrq8m+CEy7
Sr0qNan/CQJSES9X588GVlOTLukryieENDufKmML5Joh1P5nZAInOERUxYv0RIl3RpcyD5ULGIrD
6LO76Kv/xuj5J8K+YOkHPN+ajgaMiTugGnDvnmXXDDngmigts2QnBAEAtRSbeEnCrHd2gbXYaXVY
1Dpk14eKnSbUzsTg1mdCDC0WL7dDVSwCtdIQN//mM0hosOM8Cp9+nuuBLDQ6hYOjYBfkojmmB7s9
Nw8XjGeWpBjfJWTLwTyQsjugpsjaY6OqfFnPjOpJQKaYLe8a3OVm5ueFzoz1bLaEXNI09Pi3Ry9Y
O+z4UZxIK8lSYlpVK8EitIkq+Jc01JOyUmClPS5kd08Ns3sMaM3yUPq0s7hfZXNn9dIgkiT8BJg6
5kma+0LYj0UAkJDGdUCUA25VhcZOreSyUBCMUo7fYWTvIleV9bwZep4DVNsMqB8vpuX6kFJaWKYd
85J3u2ixaTZnu76/9qcreRFl2sp1uNync14WQEe9VESp3Q2pX+Bwz8jkynhubS+eJ0tLII86H7y8
qMFI1oG72XUziSohodsOv+BXh9/RpmUUDwZpE+/K7xD+BhDpowEbUjgzHh+gqrCeGVBe7PGHnC1B
jLtFWUmwpvRYKVzguTvtzHEImsNHeNT6Jd9xozhj8Q9MKixMVYqCeHVa/I032evaQhDHVhlKSAcN
buPWNgMdCt//tjl4R1OWQAOhsKEZqTnYlRCcxCjMBN707kgjdmaRtZH4HfzAXqYJqmCoJkzROGqi
ebvJg6PAa4wY6Wkp/upbceJ+xI2xz+J5JQPz/q1h+4Kakx3ettWWsGct/gAMT9G3Vqu8jLOgorFq
VInvcRPG4D1wRiBCbO1YBlIUgiXoXsJHrCh1DnAlQH9Vsrw6IAPMV/tNanUpBTf/2+ztq1fjqoml
NHrVM2Wv3l9UKM1IA+svuUjRIFBG1+HITTnZYrfdfyji4ZyF16CGmLumDkVMOfAn/MHvQlqgdU8W
p1FW2V1NFcKVutGhqKHXMMcTmBbjjTg3pTXeyGiJtL4JV3O5T4VWzJzUfUmtqmqDN698rIuNpNL5
6TRqzcGrOmob6DQKYF1RCvXR9bFvfOjsOJA9qbpJNz8ZUq836IABuIqs3E8xUOQyYw+FIVTJqvZR
LocgPpuq5JLSGxIzTcqS0+gxdKZ7edeGGpQR+fVFKVH48068blO37ADf4MjKbfLV54tFgKSuWz8H
vjpu4uUnALbYjhAOxYIJefInCxXgNOfkjojoy2iquHPYDFcTyagUXSFeoCPVcWcMEuQW0nBfYuUx
64H0T+tf0TssHhblu2PWGqWSlN4QdYFaWOK385x8zVKbna0DzCSUWk8n7hFEnKKSasYJegoYmpn4
WmZfONVYjcJKhMT5hcYdi0xqbkQB8gGFlr3LS2BgLM3cd5/IiRyVY+Qd6d5+APlgI5DYpvuBd55s
KqKl5BWrAZpTaB/1YcKjJ2rSZtTa/V7kx62naQNDpihbdIa5Bjfng+c53CHwyW66b+V/CTvRCHEG
p2z0fNEYKJ1pPxmZ6pDKwb5utR7xjHrzjN1j1KBjgmVvybycK5RxAnQPTt2Fjij+RGIyYleIARik
qLn0DhY1V+w8oakbFRZOAHxVhEbkcHgIJoSBMc9CY2sYDr/THeueecjpIumcUMbYu4S8DGS6RdLN
3uTE4mxxH51O6qsqkurqa+VfYpug4uQatDFrxiAl1eWg3Z3vx1Tun9/krVHr+6JAARK/Hzk3epon
DOg6ivs3w91iuFk9RsZGVJG0HJXSULr+txb+b4fb6NMFFp6PRUkIFgkaYbFEgwETNZcMKpQNyFcr
Rx2m6rgbR2zxSPZO55xA3PJtCcbRdw3xQPXAS7QyU5ek+Ghoa+OJWDb/pPLO7CJzqFiSM12NRD/a
vQd7w47t+TdIhlMM/5jkWt0UawcMFIkfb/GGUz+DQi1JsUTVewum8NO5NsM9LhPHWbw7NuVisY0M
fSmUUjwzgu8mmTMR6SoM3at9vJQd2uesShlwDeGLxzkrVPW9zepmzW58qgAprELWZwoiHjL3QKMU
ejqH8OGkpv6S/21VLUK+OVoXcYG70hf1oAJYgEzx1cWV6O84I/ivgswOOYcQOhQkNnzcCbFnbr86
5zyz9fGurjTRqgrCuplM9kN6kdm9q/W8zF0TmNv590oj2MG9D9U7uNQ38DmwpCu4ILLRJTbQuzqF
5TIx6M3ZIAuYDzwdC+U3MdezCE0zT3EmhshWa08y19Jbrm+OiXzOFlmmdLaMXKEYTNPr3gZ4OhVc
Y6h2LIcCTo4djqEvZcwpwi+4/IvR6DVsgzi4WxeIx+XYGT6Sid3FSHD0/2gqZ29rRwQWVfynVCyE
3BtUZ7EvXWDOQtZZDiFVws4kr5lUUzyG5UUHWuIthB7Zdfh1+VdhCU2icEUQWETjlrYIob4AQu0a
JoDIMJNPaJApLzij+EP0zdYDzJ092xVbwrK0T+Ofv6n62/2XDk+NCTDgXKHKtwJ+ZztovaTLMShD
kQV9t9juuIqBpBONp8p+DSFDWNSsQ10vE8q7wOCMCWdFIvNa19jMcHQEzWDsfcnwXQ6zq2sc4i5H
G8VqZpt1MFdqzF2+O/BMCaFitdTasxAJWsYC0jvKeY+t0lwDKFfRQMqKwYbUgJqQOvJ1ttswdls2
1LDhKkZN3YG/I+280a/3TViEgEFbb66JzTiIbjBqwxtfkgHcF7xN1iy/RvjIxJeFh07wX/Yi65Dq
WWTYPFAeou0DieNucAmrqazwdbqQtDPzwuk8u/ONgwDynEn0KLzOakaHnOGpft9iPq4n0BFozBWK
9dFRQGE7vznijIYTebpTLxhs2/GyVcKDiZoBWAiIT0ssbDsbfPG+MiHW02Npj3U5UeFWlQ5TGVIp
EGu2Ic4Lk7EOZtmUJjGA1dRyZ2Jx63UPJzp/PMWukp1E8/AoM5n53v0XcJGzKd+sGi66n3/PnJIN
AfN6qxeD42V0ytF5bC9+xVmGXU17CXv5InUeFBq+5EGz3FWSKgDx3UA4L66a57SslgxOymllSvRK
qnmE8e5aF8vIJkbHnij30RPWgH2AslyG80sHs5ED9Ayr3c+D0t3zpi02s0zP4Lo/mXYT69Nhja6p
eOEUlWHqPr+YX5KyOzXUKBGfdKkTYBrWFDsiCNn/eFyGCXpecpS4icl+gelcpVz7xBZMiV+Het5n
Szs6+dXzT9YKy8vN+Pgl1RabAArQYoBdqrFQua8zRmfpxi2+UyrxMaRbpDTPY0aQ7O1SCtnArBpH
jhsZD3R3/MtzSbDgAfFuAkTNy5l8CBHpuWDhZBZgdGvCwZ3Bvawr3ydkvPGmSzwQTKHc93k9WMNK
gaG1aRLZAqN1r/XWHuEpW0EadwtgNz5k91ZWM1JgqP0rWeX2m8RY0fAz6/YJGIC18QAfbabcTOc/
mD9VvHfcf7jwLxmeNm+Keuwo/HDG4b5LcUZzAX02tQogGKkmU8kJOa6vNX6mSOpO36UgvlQUKhoC
cLOJvbjASQD5U+vsVMe/wg2Fi+M5ixJWjB+rvF23vzUOiks4uYySfdRE4FSx1WfCqKkr1ujfT5vr
MU3YZhAbuCQxt0ubCX3hbsuImK3Pwb97rAJyaIdkyZ1s7FkkuStG/xVF4SrbeeJUu2zRgkfjeJOk
ZNcHljxMyPeW+qHwsmXqu1ITg7x1jssFAlvreBJT6xOYeiCBKxbj3Sue90iEtCbW8CVt+4r+kcHe
FTQVrQKB2wwn/nYybI70TeRkaNOwONAwx6L5bF1HggR4R/gyCWzlLHvfCCQYK8z0uPdTQJUUinPQ
hfYSK24ZBT+V/zV4J0QqFP4lanwcB8/vcf3FvGxmr7fdZxfV9pn/Cb43gOlwPUMpVR2kK7KAKLjc
GPlfCEOyUZy4zGUUKJURgzPdErHaQHt54bDbkO6HBEf2zGDV5BfWhHl+0yXKgTsMlWNQGKftInaS
7q2D2n6xdYobQb3+H+TYFy2lrKjaRmK5IkfWhKFVQY4IxX8RXknmD5zwjLZWEtXJmDQzE37m431W
EacmHY7oZOI7Cy+6txAd6MX/ydnoSMol56yCZOYrZk2P6/RWEJ39T7iIyS5MDVw6Yds/OVUdfrNC
wClClH0AF30pNU3Kw8pwuGGdTdNUjTMMkOJoamYiNdifCrX0sj5Ccd/46/JVaKIr9OmxNXS22eDb
DVvSMTsyNdD4zXUbQB3qAcjlNjzqS4qfACaAj4/td0hFv7pC69lUVQeqtAzQogND2+4ZaCICLeQh
dT1wnide8ww4sPG763hiteWRUIlNRo2wbulf7B+H0c83Rkikik4GPJ/Mxo24F6LpYlp2Gh8qI8Eq
b7C9zQbDSbIBhWHeftviDQcav4kdO/mE+2TXs6eOYo1K4042cNdjo1k9t+mPSwaNxryrb3Vm7SPW
cBYfYs9oZ5qf9ur01UiVfNf3yR/O1vAjWzFKa9yHUCb8jPoPQt70yV+HafC2s1P0niOhKqKsE3aH
3cwhC0cB0qAkdaFWPbUhCgBm2roQlxNVAYZo/AwFtUmcG+XXKZMJb8MMxM89d8u9TegGSP8Gw56v
wHgXKIN5i0OT44nlbamtyZOmHNBNe9GEjXaXNzJqeKJ14EKuEJ+mP0M/JjoFW3LxiNvot3wCoIrC
Ij8xCg/z/GBSEbGf6vfIIAPENMBJqieYcdS6lkub5J9eoB81tad+I00+r0ygnvZO0hwTrKPTCuuG
zOeVJaldsjy3pib2Chju81Q74cPylOlEpU8N6wf5aAy0VuoEu+tlPsJ3kSDcKt2dwerLXgvY9BtY
sFYRyR7IYZ6c0ds3D4CUKZ6nyrSRXmBWLCrD+3Z3l1wAMrKquAOIz7D1VS6n1tSsBUtj2OhpmTuV
3xf3shdxFLiR1z7oPpqpOJnXufyadUg2eCgLcTiklNYHZY/rYhVPaVQl+aPmGJn0gycQhKBH8RjB
Q7JgMPcp/c2JwA4eO8RuvuJZqkpNW51lwAuaWYREjo8tML965KJWk7juxu2EOcag/J8WX/fuMy+n
n5ByZpLFX39sGMr72oF12swB3AzFsaMvPiC4lRsFaueHJtAKXDrHYxsgDxOUv/sy84rzA9HrEL+V
1vvoWRmt+7R6OvSb938jh+rgoLCBt8kfsFq6OKvsM+ia2YmaXqxXLRI3aMIwm+8xj639L9aFZQ22
h7X9BRRxYbWcF2h/L2C711uAnctrO1wFCE0umuPduTIua3FYB8MDNsHCRhQwVqcVaC23ydPgJZUF
iWH7+USkdvfo7li8S/e7c6dMUYrfbkCqwnMypIlI0GTRianA59ydQiUc9FEPp2ANBYmJI3wNXMn4
yzx99uotxjbYNxzqX8LYOtFgwErDeIGJyq7SEhltNgOmzivLBQvDP+oMs2XuyGO/8oIEay/4wK2g
y1+zN8gTnzQHY/PPmPxzYQ8l87hLHqf0DFU8NAyGgSCC+lqlwaWO8rZxOwPl7ebPhBnFfKPx1Cz3
+0TVYod6KJ23SFakoSEGfpz3BnnNq4PjyHi99TN8cA5Y+batasyqyKkNau8UYWS6vVeEjKk4UrBS
VtmubE12pTTzQBSz6KZNKx/G0xSuTRD8Kg8p9ulHCTRPGKYIin6rp0CyIfr62v4a9bVL0DIl8X5e
G6TZ3DoyuFdN8kP/aaZIAL3wmXSs6p35gFEOEAj0pzBb33CF6sZcdR0EJw3BkiHIGhsmhDyDLqE4
+kjXBu+rEbrX2DBg0cUjFWHfq5EaxAx6YcYl7oX+meORYu8P+WlC5DAJ68XoSjCf2N6711X3Alxu
sVBfu84NB/1Jif7F53qWmjHQMo8/sJsyry3Zhhio1q6hbM02j/qVsFIhTlAMiZqm3GVYEyL+FDTk
zW3JzYOw/dMve7B53yorsa+zlb9ver/JMc9W0cJK0B61biWL2OtjQDK4ZJ9i2P9zs0iOfJ5loOWb
P81U4upGiesBXiZpSsjgvgHaVTYLTKseq2XD3/9+uDMiT/C9ry3q9YLES80hU1C65fN8ZKGX1vBA
y4tm6SmdNoAG9YQVxFJgVR5KCCrQo0zRvt3KRuvbrZlA13fXIHlj66Qxkd4jV2lpOb1U1zqizFFu
mx44OB8M3/WH/6j9nZyGnnvE9CjhD4DIuQbAow+3dWy1bRii8MBCvxRc5H9+wRxBMNi25kM69Z5Q
zCvwRNWvj3lOTGc2htxG/3InivfCWDyABAkJY04z7wRU9eytPZ3bhjXn6UFkjnT/QL93GPR+t52k
GtiN3ENPvw11qhM+SWV2IiD4DJNHjk/7oph5zrGqeyzQtYuCF5m1LKTY0GGg6XydGMa5bFaGfBvc
QVJ+xi29twYCCg+FYOJATHt4lT9PiWF8ZVkMXmEyqi2uqAX2LDP4DhctO2x7FVxZPMyGSBfSDXYX
QQESWE2D8r17PsEztxmSVSXgN2L34AokjpEZ69wTAEZ/nN2pe1+KnW0iQcZWD7KgajaElfxzaBAq
fnN0rw86A4jf3+8oGIz5kq17dtqsZMxiTCRo7BMW+eQ/BjwT69/YWMI3ZewuykVsdXOJHuNDr0SW
dTK89+/h14k/4IDE4yyjKtn/7ywRdTRg2Gcgz7waWUkmLxUFnAyyNe6JVjQJAnaq+Ud/NpHIrfnL
lAgM/ItgOOz/DsBtJYI+HrBgF5NEo8DU7Az1jI3hocxP4FSMgXi4qdv9M5/Zw/3BKR7ouJy98H82
vS6ywqhn6tqHju0S/g4MtAKpETkfAgT40LuaDWjn+JoZ+fU7mYRQLOwvmtWSpkvjpOvQ5jHtOlTa
i2TUaYANkunzeEXBMmc3uBPlUf6LZYkV8X8v70DvP5vUoPoybXloMOKtm2X2OKzkhM0bENLeQvkJ
pA4laCIXG6LAo7WgcQfayCe4z0/70ptqzNu2OPFfX9JMZ3WyHKoOcAprJOEUl4vBsfKvqPum5FyT
x8FfDPH7/ouTheRuwNiofQy+eTJZOMS7XEI2XnKwLiirGRoCPTzH0BxYH+RL0olaVaeISZ0i1ejr
SVTxtrKQVDLi4F1Zu5oFM9exbsJuGDnmqtCqJFWbx4Ywha0ts3FEP0kO7elp/n/Sqb2SDbVgFgjD
ipbsPSdYIED/I/AEMbNPvFcM1g+fWL9Yssrs6Ib5BKC8TJVuKxXZoYyBn5eEh8/E6na2zqDCC7+X
huVUkNHgKZGWRgjGdjNZX1+061puZhjhbiVqGz2huE3dr/2Zbt7EDV7g2ecDsGRHRozNi5h+Fd7S
007nk8IpPCh/M1wSILGQzDpoWdwwGbT/3kltv4b1ZIlzz48Wm/wtFJQ4vYU9Pvy84BxRe1OHY4aa
KCI0EvX1DbUvDw0/2emSozxtPP6hZSx1LOuouPjR90m0ac8ubrxNwTxzKSgmxeJMI6X6yWhxDqUV
/k7XbriJOI0FpSNd+/jVk2uOaLvxyCVyBtrFgdXpgFuPyD6wbilm0FhV3qRR3GywrVuLET3a6Gdf
G14q0I+3Z8ELNDtvMRgYzLtzEmMmnio3G3Q+WkpCX6uwmzdYyrKYW45pfO5nMsR4XN3jl9iH4/Fz
Ec5s2GoVlLTa0hbfJSWs27xr9kykN/qmctSTLKHlN/V/fuLbors4Ai+90gefoJfWhr75CDG4HivT
5X9OQWU/HrUQb/0j49rsh9e5J/nXHvjf1Feo5SHbBopxxVsFt49XUysCkhD2he/kucGeMyWQXgD6
jhsMVwsCoJ5ibInC190RLqJErwv3XVhUK+DOGWDklJuN5QYDOeMZibe3s7sfSAIzELaeVi0aYVuj
Oqcfac7HiVICGQRsU08yzD4rACmH8O7RC5fXWgmfjBk0fCuvBIW5cwjvBFGQo7FJ79UlZiYZvizj
JT3N5zwLZ+85yrjtt9HfY4U6EaRZNUK37MDcP9zsyOMljd2ivF/dbVwcLT8y2mdPbEhjlEMPYlwb
0X1xbCMkDB22nnjI8D9J/0hE45auVgYaxyuYiYS1W5fZtty3smxhVgTjB8mD/zyLyqcbeAk75A3I
w9+ujuQoM+7cCrhZJ10VC4U4FE5CpFGhNbCWkIJ/vUp6q1lxhXsjhGN9NJuAbHw/AnHo9TRPv386
iR49lZ7dIEIRkbuIsH225WcVfDPBGX0x6ecWsD4J48pygyEWsMtaSpkX9DZDaeOl6lJnvnGsVBbZ
dphpXARf43GWhHJMcYvYP8Y/pAutPjb8+49kD2mvFx5BLa1zIv+TwuQMqraEDXGqvPt70Yv4K/12
47bgx9ZLfjNsQBdBAojEo+qTBgktiYzqAg4Ve7P+M+GJgb1TMDj9FKtnrSZ6uFtM1Ei1jorGIvTN
guDiwacfQ1dSUS5gnolGdpinL/E0akRVbsXxfCp7xzrit+BQsoHdie5mabcfGvqqqQN7l6exkFwc
dZOvh5DG+F/kzCOLxsc9p833KEJtMbRK3Msmg1C/RFVmB/w/PQxzByuNBDTlY3qw6N2qeh+TvRF+
Q7N6geKXH4vdz5OkhcevlVxEK1g4PqgtUDbsyaJfxgbRPHr4Vmpg2ShERov6FgjT7MAbOEbX3Ly5
vPvr4YskvGeCgTdkYwDp2tjWhXg1nc9eCZDcyhYt1PF0IGJIg9bMe53s3mIdXh+PfKm1xeSMO444
BOhUXHzaMbhRIjlbqKQeU/OehJD9zheNohk/dX/v8KXVxlulBi5KMh3HZMP+5E3YYqnIkhyOSw3z
udKFusde/dYUdioDNbFhAzFt4LOaa9mJhheIyPV3A8/ByAASB2cxUi/FW9F5WTXcGvCMozbe1VSY
KWKzaAT1+SuuWa0JOYUtaDsOagBv5rlCbYmNboNMPJj853uYVUce6CZdG9AnpTvXNs18SCcebULV
jG11QmpRRZn+LTyt/iCvsGZw55RlpySaNWfm1kgh3UOWg7S4shH91MPapfXSmCJ/L+QCa9DsgLZU
zPe2HJ1HxsqcypYrl0k6FWm2qXV8nyLvhSPO5Rv/H6Ucu8/Kju0V15RzP9EeZnc0uwO4IkCsIaD6
7LbkArCHKA3l/SBrfs6Kirx23EeThrEX9pXW1cLIGL/bJjJj+9aj0hHnxWnGpY6ESvq3LFwtLayG
W+AH9fE+hSntDq0wNwiwFhvM1hIydhPc5tqx5YRsyGAwaCQScfi6TYoMoT8dW4yupzL9ZyyxsXfb
0d/eD2tLljjt1oM1xlqDi4GmnS3xC2WZ03zql/OjlHmm/bCKho88lh7uZCDTxruIVe8psCJHHA66
QcYFLPWK6c2yAidWX8E6Ue/8Swx4ccGPhtJQbASYhPHwpi+lRV4R3VWTGxACT4w6OHCxNc0Jv7od
IbsDFI3FWgG0UdBehoFsj3kT3ClzQI2OfGrnFEf7pqGjKGp0pDRznkLq9OAWpPFn5wbjf9GeGnpx
f0AMImmChFyohuCM9/Gc+gBITvlZt/FLByK7WNQNA7ll4ara5Sk/eAVBXwwgK5MwSA65j2ax71qY
AJdDRYnfCdIMaGrm99QK5/25ctKnXYzPBlU7F9DOg36oEsIPfymfI5F2eUrm+18RwcTA0JahwzBT
9SxgpZdrdojaq/irVO0lS8u6NTfn8BVzkCtVNHPztWqu1fQNbqH81IwecJhzwSuMyggWZm3j4Blc
VGp6nPxrNlA6BY988RIvVnw7AQtdUiZoRWWR4Z1bY5joO9Oe9J4WAVvED6p6M2BrHk4J5zAnWvIh
/IKnA8saqIvazXKEkzHu3pKCw3xpuGNyf8/onV46mLeCg2plXKVQLMc6O6mgO02Epf5o9uJrjRJQ
82ldCrI2vhIz7udbzL3OoPXRzfAkyWS4BubjHvmDM13LnyBKeoYELzF83b9dXmqmt02SoP0MPzBR
M9dj0GBhLhY+Ilgh2qNb7sDYGuu+zh5u0/h+mLjB34ueGmVQf+QnOnJYagguBEzMefFMYV1+bTrn
wO7mzny5X5e23X+cvKOcNW5JtqmTWMst1Ue61++SaFxMe6gK0vzSpcl8Vuq35gIDvJ8MhMyDcWyo
j5GRgVtAeBeOuIXeCKRjsL5knQPvH2+w3QT8CG/MjhBioUMiGAzceEtW+bCIOfxFi5UKHalP+S56
ssW2Koqqg4/PizCrn1vHZkABKfVjAdNoElevEjk7uYuaYA5aBj0mwAy/Ha2IIhgb+MmeYg19p3mI
ZIQwcpYV26d2bpRRHCgX2Wd5H5bvvfdI7uvzfR8ohX+S4cLE2kyKNQ+t+Iffy/FSEMWgCcPt5ElK
ClvvpTuUdacXo7u0XVG70ki/T+P/sf+fqigPqlMyTW9Dgv8j2cqku6wcnMHGPOfkqTXOT/719E1L
azsasY/9uFbXux6mTnsPfkB4KNStuVsTThpu8pb6VNBxjHbX/sXqWahHI1Xr8XRDnmmaArbQuzlv
emZTjCAdb7mQn2oD8Tte+kRLQ9BEuVzahP1PERfgTdFFO5PLu7iWwZxGiLLgZKZqqJLuQL8V1NPv
h7d9Tz7+rIwabl1bm8+/1kreVDSyCgQVMSee4Ljd/hAiHd5qc5HtVaMlxI7pzUeT1ftSQyYd0Ux4
eq7tOgEjr7i9Tgg9zQR73ANpLD18gJEPO8WlMCUhiye3C32q8Ugq8VrAuxSz7fZ6qElDFI8wEdxa
KPnyCpqZpsaPFMhAaS7xXbKcof3ZI3oSup35Dj/3WePhJf/qLGCLBhBBGUId564+tgRm1vXq5juu
SCi+MAEmzf9SnxAcifwq6vIGG0cxpmVRwU2dwn8+X4q16IJPIyYcwS2U92u6pjvbvJ4a4AqCdXLN
oV0+o6kJa90PcV63oBz7ycrGyk1uWNiHUAAHcXBGlJ2bGZK8fm+UHO1M1Usgqwl8DP49N/812nX2
7eDa8rGin5n+BxPtDB8g97QMTTRocRc0TOQFRjPg5VcbRrbOhWxYWwruvyMHP7oEKcZXllmJG2/V
wH2AdAaU5K2E4WA/9Q4MBHrYW6qBYCqM63zZL0NquWXGT5c1Cszp8PeQstMKFHWyUe9Uzm6eZxEz
5L3CiDJcCGyEh9HSg3132BTq0+3FWLQ065BZqy1nbObiU7miDvezB5DgwkVZaDvW0k6Axvp8W9tZ
nYuFqGgV+OvlCsxItM5OKIFmznXzpuf5XVKfO71vELWjGfHM49Gbb/dU38rqSwHsPiJUBqbD7naO
vI2baVKBhJ7EKbEOeBYyco86vvlem60QnxfbAUNsqtx9A5A01W0/6q/pFs/T92qZhqb6fdUrOB0I
Po0qGw2cVkPPB66q6PpG87gw2X1Ta3gu7NAXRE7t4/2SRkRRmyZ6oTST6tdsQeF9FOtbbZRTDThn
7Ij42+Pr6O/mDajj+sGgTfIGNM9QJlE6cziTilw4k7pWnNRGqbV8m06MusOmeEYiOHBfs6f91Kl8
Ho9lxkACViaaWgMPplsrma750M/vJQ4H6mi3Ljv+q9BahouopGDpZ49ZRzk7fNwSjcKfX8/h64Qk
5G++N6JSw3kdC3SRTKDR4bs7cvmf2GoRUU9uUoFt/2/8My2We1pJjXvkuEcQ+Htt8spBSdiXUhVB
iKYdtSGGGCujXcQUEozSxIA4C7Kio7JTc9Lv8tRthGwFpxxc56tI391sdDHoIHIY0IfeNc+sH/iW
GEmhbsG9T9ucNeqW18Y/sj5RJHuR8rCqbYzhOr++EzDK0I0mOaJLeZx4w5Vk6d60MEpG478atZzZ
F7csMDAJ2/h2ardbuItDoc3YyKKsDu5PDfQTEcZmeFeQCrgZy0LeX6+yMd+LC4eOjmPxG0/PGoTP
3vVR3qzdbpxht6dfMmryEuu0hCQh2L2YwSqoa1Pu5VeYwHvmX+KCoUaYuRdqFwx6HeI0feApi/lK
n2QDxOsWBMelgEZpAXmPmvp0P9atMqRRCdLjhqOrGONIEtXyPJSQggrLC/hShxgdNviyyCDU8uk+
CZg5vAQcAM/Qrfqcxm8kZt8uc68sNZXSanvYlessYvM1DJcPyhH8YFGKAqki1JytHcDbyzdvQ59g
NgOE0MTIhbJEjXJQYhPesWz6kgKfvYoe64WFpbJmSZdhI4x0j2U/cErdkjlSEoHn77v3T5O7UVfC
Sluz9SzlTvKxOg2wGQP9I+iFNe/lna2auNhSXO/z6FBjVAhy4PP7qc5Jn5L+J4T5tsB27hhSCVd1
16hAu84vW/e8HuBCQyMcbupmhNlq1/jlAZCuFwyeqNQ3p9HymZHKV31sOBZe3duuyalzO3e2q+H5
KiCsMhKV1uHK0Ok0XdLqTocqez9XZbg8ThOO9NisAEVzG6XBB/6n+q6trtkgphidegVfIW4XxIjC
6erZ3gGWFu8d3c9sFyokoTzj4vuY6dKkofarrxW+C4uJ6WfXEc4UKPATYisrRT+6T5xuO2c5rJKI
+zV5lT0XrRRFDGkxHEiHvzcuAAU0ipwFia0WzgRJ32rSap0DzeGGpfPl2N78tJG1+PDvaXEUZ/wU
pBChjs5CpuApVFddSuPqw1e/KRdVg4m/e3bU8yPRCZUUz/haRr8b7i9AVm4p/ekDRaOh7PTzE/W5
YXTaDLcnVpR44zRhkBxPNbHPnmxRfP77DWY3nV3/2gBpNqMctFBbvNHrrYjvYK/EqSoSZEiNcHP1
9oofYZ7KVKOoB3N69Z66mlAl0FXWCozvkpoOlK8YvSHWSzNTgavBIxFURFrMP3o3nrs/DrDzTtgb
Tkfbfbj/QBDPZA6uPD9i18AgGFEhy53aikN6sS9jajtUzUg79qQq2Bo3neB+RvU5hzVkVarRQycC
PUKVqwIA5+5SY1HshVR2tF7GXRNePreQzff54SLn0SU78A+5bEEW0jeukkcBb9NcsUx5d4d7fQnH
4ff8OQ1t7ZYT9B3/uRVuoggJ6OA2IUl0B6FMJj3wl6uS75gacHG08vce1pL+X1J5gCAE+BEcGZra
P+68FVuZrCC8o86ZxDltha2xP87LV8fqrkLMVZx/kGIMNlqQBverPgjKFWgbQQsKxjza1kEFmFPG
Xh/VkQGThVeeKVctvZ/qG6qRtElch4di8g7yb4jxy6ACoZHs7AvzlLgBQrBWD/IA2g7d6AWlWXl5
+HT7UlMNejHVypu+TDKrQUUXXQpRCkO/5MfLH1r+7+2YP5nxwOO6P/z6GnOclv9L4z4vGPrsdeWi
XLaO/NMoocRD+u+giyRvLEFnph4+DzOf9gQvcZe8ApRDpeaUO3HWq00qo+GARRZBJ7DUkH5iXkQs
1PGuVVeJuyhV3qtiPlnrBGpq0G0gKsZsIVAUEpzT3yjTUwyefSNp6ttI4YKCUIzUYEGmCA31OnuD
Xh/XGTDL2oJc/VIgaECAwvULIpL9mEseeoX47Eklk61iZz01COvqMkW1zItgM03Czp8F02q2qCpx
u7xmmiqzvhsolumbSuIuGTHtd4MFd6HRIBBneJJNHn2ZRalFCCKuqiqlYIGYe2Qy+3B6Ay1Ym/0R
/k389Lkm10KRmoW5hQc1xtAl+Z7czhXoOK/mK3bVbcfUKz7SQfb6i6y9+B00nmS/bYMKKu7uwBJz
vTnNvAwCiIP/bfuOX20h95O+mAm9MSP9DH8HfnVnM7Yib/QG9cN1VF02XETsOX4KyhAshMjJXeUF
b6x7cDaCdXrHgs8ymkknKD6LpgXMDs/lBwEYy6DpLbP5E+DeKoTP829jLipICII6Xkcu1lOcNis5
b6IpL131uCxdsuZqTtbLCR9HZilUqSbWnB3/m4JmagB61p7lmcARUjUTWQcfHFOfEqGItb/kXFGq
WpABi2H0/uVaKMo/YiIaD9HfMmTkhZs7OPi1E3IKxKzhVBmsoNeISe1CPcrMIoG8i07JEiSwMxU/
Y4PR5MUva1v2s758dYt0wOBJgho42vJPBwGFUpURMGG4JiYoJW89Pw9hpYi2m2g851ut63SXdH/9
Cze6Hg95CRZphzPTGYraNYHbiO9ToOEWbQP5sSCSH+ns0Gfr7h3XsAl/qkS/rtyTD86X7OnT9VvF
Gk6AYcWtefClrnjn7f3cnLgFrYLTfdYdknComuF2pnpkdhYj2XD80jkh/VsfU1BoI6xuQf4sx33l
u5qb3JiIxrYSqdS/LMhk/oGD2yaeK9CBmuJ42Xj5qYxoE0ozq1K0rsq2xpT0g+cZRYpbRhCqEW4A
VFPIS5RErHLxzYAT8gGXIONw9TNOPar6SmBDNUss89XdFAgpdsdQ86UJk9xsa68/ip3UjfaFrhjQ
VWXrqVDyC5FKlyF77ANnbtfE+gzm70QVyZgZxqLm5gEMQJGqtei+X2flQSpW3wR14hLDvngUkoia
Qs9Ax1rP87yaE19xLSimy3tKwOosHG6NKNXL9hPoN6H5bW4EmFy2D65+z5tq+Wo4wvxJCBAttYDr
+1YyNe+WrAl1iXj7KttrYbbnHWiNTrkQPNlEEIqJJqzHU1RxUorY1iTGcTwTMmyuWreahMs/ZK/6
KgL+3Sz53ZazcRbrg4N33qSY678pjpPSuvwmwTtq5KLpwk1FDXahiaO0+U9cK5yLdlwBvdh/cnzr
7qFZpK1fn9tfylJVFgMi4wAbnZMtnIUI2ouwDl2WRbgeNqFUHGK/vk53uL9R6aeWqEmKJG2Wz6EH
1ZBffG1WMDjegiNHvYLRROl+xu6umQBcNEoEvKSI6HBQcjYPokkL79eVoMo+XJMqtpuJgZ7c724L
KFiUN/Wh/jHHJFPSWNKMhD/EcF/lmuuUA139dVDv8JCLyKRb8DRlNS18RfxF7yHed7EtH66H8Hqy
9QxwOky1Zfc5KLRnOsnUVvLshFJFhQwlC/pXunN7U2w1lEjXX4imIE/rxo7u2pMzATRb6WHbCQ9g
t6ugJwMArrDdu09zn6AHZ5sHUYQPTSGP4UvTJBSKo3qe2WKV5pDr5vAU52Trdt4dsFEfzHl6LLqY
K3RlgiVXJAV3UoUu0pkmjwAu4ULzkgf4KgkCr9Q757HBSNVDPKtuysOW8SIW6MLU+YPgtoI7KsUf
oVz2vw+/S54kjHbcw7HsBABigqdrxPDS9IOGY8z05YmD2j55AJvlTM+SwqAeA6NPUNqI20OjabDN
b+w6UNPl5m/tGJhyMu4BBtM9DTSDZBtdwsDQvtHpyr1ru63wAOO3u1CGC7UjTnRPvij3NZ/rwd2u
GN6+z3LgTzt/ZxT8qBPoQwUF0NR8LJNwCbrC1pw2fg8uUGRCBIamI2JFZ0h0yqKnMsrqUHmzxKBQ
CGwWZixhmy0WXPyUWlnvxNcSPDRFsFWaIrWBbnAuBKdO7Suebto3PvJAfqcYnwLi+ISbPoAJrNOu
+0s4/MElBFfGPrJMrMJwDITeP2xkf1nW64tWLRDI2qDI0gf4/CSg02HaKOQhb5raXo/Lz37wILT1
T3J/NB9ft0Zyn8qVA/cNp210hn5Y7HxCUMfxO2IdE/jRYxpFlD1LxyOxNQNXepCXnknFAS4jcGu6
PVSsGc56l9HNAW3xA0vru9/NiP+Cdf5RKqUvUBazNWUrpfOM0fDA4w+S/Qzc5hgQ0vFhSe28UcDt
3OUv+WvKbJH3prX4xO2Bqc65znI4MqHmf23EyWYw/RfmhdOOgyH9qXXxHdY27dJZWF5OIaS8YNLp
31Uu+DT3xY768rXlQVTVMI/De/Ie3GvjS7JYiL6LHdC2xx8G4XRESkHKbhBZMnDpEh9pVYHM/jx5
wkqqMettxFUVz5Y8QH7QigwhJZzhmnQPcoKTQo1xNfYLFjjhOezZoiQLYx4qvfU1coybWqAjK+bK
r5bwHFe1uNtPKb+E3UepgFqGSyafs+zuEpuJpeL/8J1UTMHaqaGK3SFyTXGvKjC0VbBPV5mKDDTo
j0Etf6vgsGanAiqpgQ/6Aet+3T3kvMosohdHCtWu5f+Oc987l1miYabjGCc0NknibZWts9WA5rPG
CUylrIWxbQ8I3HZhXBHnd9j6Zr7LdOvr6NccxHqSbWmYgTWSOJO5GTZeiCvlED7zJpFmmdvZ5uxp
zP9CKmTEH8KxwFiinvx3S/ndr3Fp07H0j1oj1jUpf3ukO+ygnAkI64WxLhAISyW5C+pYcSJ/Z5ba
6acwPrYfy2wuyvIXVrfBO53zx2aM+LoCL4YRHVC5/mFfHMIh35pXcC37TTHSk5k7KlYyg5MXnx9r
XAH1ItNR6t7Rz6gETz4GU6SKSC1P8FXWZpOCH112mWbCSl0J/sxKLOcWaIusmf3VfD8q277xE3kN
WpZNHIMR23klPtdwWcgfY0SWAMwATDcdWPAYhrWXXqAtBvpqVtXOE3ChMOHPipP5dbQ7faCUowmb
dfZu6pXQXSmLP+WhungUYQV+Eh8FtI3wkIkXtuK5b4WFVddNjBti3ghjXgSSlPW+PSHk2elSNv0y
FHAtNjJngNtEKI7aZL9grEkrBkIsgRNVvPvZBj4Zx1eqJIAYOAtKoEjEjHClB0YxHTOpPBURWsaU
O0xApN5F7qqlMlQW2QFQWzrec82LjMjBqwN95bgiywRpw1Hkqxfjw1fLa2BfCWF4U28zWVrr7REc
jdC7awxwym5KLhEm17gAe4f3eW5aCzzVFg3QwyeOmzzT36FTrHqor88z1kfIOe8Lq+v+U3aKpvrY
g9UK0UgaNboXIlZ8iXXbUzNaoedeH8DfHUUeE/VdwrEvFoOM/2T2BTYtFqtuhkIjlN2eZNmKBXrj
ksik0tp8D1cDV1QdUm7ereUjqvVLcXVuo1GKlByYf8Id59p32vXAgai3+W2s1fFeZWYpOIdOVQeL
q8/b81nXq28f0WnVVvZCqFpv0J6JI30fr6uJqbjnXlWjQTpCWbuwRbGLAYWpmFQdNvLB9d4H30wb
OsHRS9dJuu4s5aEkZtPp79GHBdeCWPvNdF+l0QgnzeEE39JcbdKk9Sc03sXKeYpSHvab/K5dwVVu
3jEUeksZnU1BTM++yrz1pmw17YiwVQEPPTxj9lWj9sr/gl56/mCNB6Nk/EHm27G05eqZZytMAhSG
+47AEegYK/AnMRpKMTdPRRwi2aALSbAE+SHvoXX8aa/Y2K5PRBnP4Ffs6fBpozkN78VtVOGQrjnF
3H3EevtfeJEN5J5wJnYm55F47kbPsnWr0ppplo6OIqreAB7SI5RQrlk2dehpXxXauUo5z5kLDzz6
NnNvTyI6atwLOrlWpmbf1VJmz+YZih4MtW5w48k2F/yoa1M9buODJDiBOnV/XqYfrQhL0R9dSmKy
0KmBmtnpROA3o0cbHG2NvBpcgcsP+UzLeHChHOxYfZkpviclW3CFv7u2kW4OMjpjWZh+sP+9YMKm
CfIxIMdEPVdD5ZftGZo+ppgIun1OcNwPkznSTObY77wmWK2bTSgYno9K3KoygIlb1hO+9T1AvKun
ykts471/v4NYZAC31CH99Ur0+CxsWFBkKWg3Mqn5JS/sfSQWxMts0ymMEM3L2l+0duQO0v+zU7X8
i4mAl+doLwzW1ctcIMVuT/NwAxVi+5Rf3+9YJlkUp5v7EbmEmsTXCUL0yHu1z6EZbT5i6VcOFiya
Ut65r3vhIPLs3ytJGB1EXv59TgyIHtg8JsnNwmX3w9hDXu5G1vt1WGmjvLLQfaAzeQ7CYnLsftSt
9lgraPgC+5RosEYP7FKtxQXItX/bUU9oWifCCmsSKaMt4Bd9X8UmY1w8Xv2T6PG20rNT7xUONNb1
pKEIwxzp0dviaRNZztLptUaSFSSi500w0ymH4CKeZvo+6AQAB4HGBefARC7/HoXNtiw7YUvKMwpN
97LSUz5PFfGSkO3q7ygS+m71idhcsh8gO0DBSjSRqKuYqxPazRVJs5rp0Dw3Rcndsx+lo9zz36Ka
rX7ozTEGDW4yXQLZq1gWbuDh/EmCZ50QzC9yacu+S5BghIu0/IcnRtdv+57C4KVR07IO5rb/6VkI
4h8IIZ6/f6aWm3s8rrMDKYExzEsiJBj2nJDcBS1pIjjbNB7rAQacJX4z6qkga6FxkcmkjSmIKDAH
0ECo9rTiDCYNyVGcS1DgxNmQytsvUobO0IK2xhJiHuLc9kTWNR9lgFAIJ0GogN4XAVNMbCCJH7g4
uRuGjTVXwnXulPbRh+r+6mLRvTiY9QpyswfnBHR7K49VBSNOf/BTluAu6PeFb+aUdHMs8aQJgVPL
bqfoMa9EG3mgeMGjsMqY1aYPm3kmEsf4hxtAMWD/ZU7OrpVOx68xfoCPyvzVGbhdOj+PA6MmR/V+
nGTyyP8wqHHoRdTYhgw/o4hVf6LHzodhQiOX4fnx89UnAzOqS/Kj66wHr0SiM8z/weQhmw3B7hBE
rOyAkjOkCaMia9uuX6t15JTd5x7/nICuqow/mtIzrcmWR/UDbZBPi/VSaxcjqXnoqBYOykkU10RA
PsQsDSSx7qxZyIg7NHxLtXPiKO54s6rYGPmDpbAsUC2Cf3JlYyNuIHXcM2SGEBWETg3QN23wFd3p
T35IRxkhK8fJqImNbnUXrMR1GQI6kkNB+KV0wT1UbQGoKXmnKfn6Fy1xdApMxwRnDEo8eGBRDmHl
u9Ihoo5l19RewwkAkh0F+dm2Y2s3WWZBFO8ZoRrXGuqp6mlkOp6bJ4xfOnTc07D0HnUUDicJRglN
wYVazQ0Oyx0IOF5ANVQVDGcVK9R35PE2miITPxnlJlsYnwZZLR+DHRoR5oFxsJtMI4JmgHeEKMPZ
K4xKsm4PLwhVtBZTIsMBdPnWQX5b9Sjuwe97Tm7rDgTzEZpKDCpsDcuoqDUGMaR5DYW0jXl+j35/
p2PoOb70hpa8GQFYOtNTlmC1WScpdgOVPQ9Kg5kRdfYu0zXO2nTy0LLzHjAyP8GzggH8bwD1czlf
nHURrFwH1ROIXhzQx7hUoudXm2NNTrii56srwX/aiwGXkcbCnYWPRVUqLq/YZx7gdWnbDZNljbdS
Ly4dIcpnhOfKXr9JXZpFK+4bKRQsZwcHvAX9Wp21rfjiJVV0vrdDML2YRRUaUIbfHlVCisJ48+Cf
en59w2Hmuw4XvxA0c05mUJOM2cRiS4glwmVBFCxa9XyJWsIZ1c+VdiQ55GFfmhUbmyjitAb/aR3a
16Ni591u85IssOUIXLm2DvGvLKZHhQOP3ogvzZ5WvtqoNUkr/AcUveQSgacFPKRM1WNfEcCN2B3Z
XwrjVE73yQl0vJ1/pi6YyzfLElgYnh2+e9vIVEsZkFQpAB5q+uinxLWeqOfAZrFPXmTHQWrja1b9
oZ90PpVdp+ZZwbQGwyvwSYLQ3Amo4YwqpiDJqeU0zKttaaF7U89FUOhXoUpBfRMY1Gyxp5FWlv0u
Vu9LM4wHr4aQ1IQ1ioDxxZ0/kXFRXgAupszleMTbodM2tLZwWCQSZVSMPFbCSrk1uu9Tw00aE/sD
jV4yj0lQa3N3+7D+yPL0BgSz65DAulRrTP4a0qTcEe2DyFfHzA1jdO0oEEXRuRN1/eA3RC0MbiS4
A1vAnb9Um4C78Nydy9M2qz5XkqxXdEJxw2b3M6QzBtprulPacdyohAwxUyjBtAG1wDAi0gegUv3h
zXsTy7QWhbj5O0/vgLp8u7Ggw/dQZy0cv7d60H4ExS6oQecyqhEoJwcljJDuIRmGElqHs1tiohZQ
Wq+jOgyWXyR6n4P5YygYdnTz2uVxsW3JCRLe4HF3TyAHE65m0XPL7eFoZhajrKu5lJabtzwiErUO
RARIlKUrK2X+UvdDWctNGe1eW/8+BY4wBZNFS/NwFLBqSa1kjQiChM+cf/LfhXhJ+r2k0cukLmeL
hNY+Bf+i4/Rf2phIefuQ4xpZHZXDLanRXTnxO+mK4NggVkGAer5F6TaHewwvQnthPbIFh57A5vwV
OG1Wedey+Yp6vcjuyxrP0NZbJXcQP1mB2e+9NWLrnLPyv4P6iyz9MnbViQO0xy/O75jhlhAlzVgq
C+YpW5qCOH9OZCYueBqLGICN9PaJ6VPuutNOR1v8GPohTQapOI2lmy6dLlZJg7LPpqIOmom/SPM7
RXhwbe9H5B2UIZ7udGbYxpVTwJyHYs6uks7dCexwRbwhj6TjdQ4vCxXfq0RN//HkoxAjf2CfsY5p
t9iPvMfOvGgdpYxqwwfsq3z+NgWAeBspyVX3s6yCU5aWcCn3g1+0LpE0y/8zrb8XqBLb9Qm5iFcG
emmEVIz9JGmXvNuPR0pQUDqdTpZiPsweysAmxYhHW/D75ky4uqD6A8QLOFnsEOm64aXrR8wtecm6
6htDg9jUx2PXQQDsrxv/0hmYGiqC3roxSsFFcwbi2sbmqV6feFZcXa6rAnbb32iqtBihfJn81RoU
G0FG/7Wcp+DP6Sq1pO9U1o9f3EsVRMHpTfCUbDJfd6ARD1IVULEO8Q2ZARnLI2eSvm5j+LEiTyGu
YJhja2H5/7/V21OcnE6HBfmCf1c3oHFBfTkDXU/e+osp3y2u4Vf9QgTvn667sUs7fOCEt0jD7vXN
O31iqhW87569CRf5Eoi5peUb0Ucjkp7gv60XMbW19Sapb0xs07aisiHuE/0XVpB1n5osrLetnWiB
oZV1sdcEZsKW4/MVwpLBy4UGfujfs+oO3xKF/eqIpPvkxWLPD0m3ydfCuJT9ftCpuUvzBZ+4d4uu
eu+i5gop+9ZT93D2bzWbe1d6G0tSymCO/PkeWXEOJghx4GAOMX3vcq5JaqmiEMBa/oXKHLB850uB
K8XXAkpg6mZxPYFoa1Lj4tCFaBqHZp05WYBjxF6gPAtfQNt2bDEj2439FOgDx6Llks6/KIRFpLGV
N7VxPptAl2uWGyfBxhx/TRDAxInF9mx4p4l5Iy+zdOaEoX6bmUtWIzky+xoi5/oJ54c7I+z4qRBH
T6Id7jpwyflyFbQI0fZQ01AfU39Oogrx4BdG8DEuj/ybf4FrckrbFA2oQx61fYP9dZsMnu71P9RH
/LIMzkgMOHhc63jFkMvzuq6vMm5Kb8ADTyB9gG0GBKQM8EDLvgLphtF6lcyzANc7zvXtTKP2fAKL
RrMjm0ZsAdwespV/3mP+cgQypON/Rw7qhEfr0n5ZuMMtkjQquyzhyfBxrCK7ikLcDJRceJXOVEqk
Nj1QOT6D8dhPZakdX9+9C/8J/FBeaRIFgAtsXU1AdgnNmFb5A2xyV62Cv5SHjK9pXIXObcPPJCQO
s2XdD2sEBMaSB3Zs2RFt74LgmT/5FwcIMoAaZqeMsoqp2fh8W1PMOv65gFdEz9JUxhcg2vOiv0lN
naZRPOhyb9WKwN9JtLYjvj1aTZLSGFEuVaD1kIEyp2ypTmwBeZKvpUUbfHXIIzFspqagGVamJ5pb
cPDzKxLYipkl2OZsaDXZ7rYrK5xf1ZHhfCPLrngpeYMsDBJdSAuUqqsEP1LosZvdS3wRBXnaIIy7
eq3Q9+hd8Becfg/SkKKU4afphRkiBKT9iv0inY9DKNX+HdUbI814eaC/ro6DrGmtqKh3EWn6m0FQ
nHoo8c8E53V8zKT9y3xToPhG9vam38e0myaVk5XXN5ocVgPQsiJRgAFrSUObJcV6YxJizGYHnGju
ujv8UnwuQElFmFfgeDkuBtTTCJYwLmgyPWom+Az6BjqkW3ydL6UyQE/qXb1iwnIk0hbI6dbgnvbu
ZccrQGy9ZIVFiOiLPvCl2CKc4LjrkNhGJtQfMaHFcF31uZlakO99lqzcHdx2JAJWrQLfRd9xXeAP
zkr4hR9LQjRFUwYhu+L6DtnM7kfeQIM3sjuFvqm+S7610KMex9FaEFRkrlwh+WqhdArUHY+YZvrT
nQEWco2zBoSysqdIw49E2qeEa70dcSlvgf//pR4keGTug1NOxP2eaZLRxDekOSqFyOCylN/s86ck
/zdCQvS3hhjPtA46i0YSKFza/a6b5K4oen7Vet6tKmx8vq/o1bxa1j2xiRkqGPbyiBAXcX4CFaLo
tP2zt7m0Z2/0cTT2B9ENYc4GIucTz2VKesYaCmzlclKppWQto9eE5cJ3uQ9RYI4IM6Wwn5xtpwKd
QfR4w8SLXjq39LW+TtQ+zt2Fo0Fc5H2644IjC5UKlOZILsTaYVNncxoVR/4E8grhJHKGq9K1zWUS
XSiZOVA6NWr7zKvs0qqUkNiET/jvYA4mOkknahTUpEZm9h4sXOjGWon7ALWAVQkM2MEm77naWjfw
suHRtJoskyGlHcdJA+8366vtqzOFc//9GpNGR3lCWw8nivKjmUSFDf1TK5JkA73jc5MracLt61Jk
YxWJNUlCtxKQaXJSTYb1ad9aPcDqG31JYMRCmoN4e5A0jUh0S6Gj785vsgiCxOGkVJErm7iJ7fWb
HAKrh4lUO2FnXi9yu89Eus0b2gUmA/AZJ6FXupI2tc0WdqOKbixNxZXTTiVzXmce/fPG+GFDQd6X
pQ0Vu72W5g4DVlTMp1+I7Xvew296VVjaLZFiXTVANqa9+2+3mkv0Ik0wejl81CnVtDLqccC6hieg
U1LOP9S7rDVcM2kUfWEiKQFLHiV5UtDB0VoizyHJy4+2K3a1aWQntahsKs6y5I+yJYgTcs40lF1T
tG6CA+g2ACL4p/J4FgW19px3FFKki1w9By25cRMr2WhTV/pGgRgV3vPZ4ljP9RNVyDbMk/ka+ssJ
QK/Zw1cGHjy6f8q9PkrRFTgCt9FEoBkg+zor6wm6jHn3eVnkvPaTRQ2TWHoaOvjvmpitHqEc+oks
ILwNmSli+8UL2TbS8NlBJVOTRyCN6MoKBKhT69Zxz/FH6rCm4mDJmmSdWdDO6wN1wUU9o3umDKUU
/QMtbKDeGPa1CxPHyZUU99vqFog/EdlcDdnSECq+2VRFYtJYYLC3z60ASQBxLjzxSuR3QM6tH68k
ClV3/+If9M1xWk+yx8+Xzih50CYoWVIQGEMpZSslSwpoN/3YQPWnnsWIKlk37QR1KcX5dE4uwB7+
/lRZL7Wm95WYqx+II/dqEAPK3Els9HlQx8CWthK+3aueJfgKtzZyAIggGLwVroWIqdSbHMwKaani
0XpsccsvuNrUHqJGvj7Tjk7DEozC6dLvWJZ1Hyg0tXiXCfIB1lfgdCh7Kpe3FSLErQpDelNJlFu2
v7Vqj3x/SM/SVETq9V6u65e2WcXuLARCun18zNagLFWeX8Cat29Hmri1LYCQ8fROL2g1DoXr+SGS
G0AK4U9oYvuU9FSg6X0qa38Sri2+2ZZWvUKYXx3Dad8FIsZPPmXlvDI6AKmgKFW3gVNk65hqrLxW
mjiLPRl0yXLBXTPJeBvaWBfEWHWLmSFpc//McREJcTcpO/LOPqSMT8b9g/Tqw7NIzsE2AykuEpfg
0PBYPB4GY7V5WsmIfDjs5VKLY979c/I/XoH+rjH7OLxoIFGWjiKK9kfxznkPkMzciDnGeFmCe/hA
/+NPg37vdfUyAXbLXx7EiPD8A9osSjFNvFPhrH76JZzp65khr9DXWERpunYDbG2RNm3YRaY0anXr
8nQ+X4Fmwh3TIc0yJKrygDRb2kRX/qe1Ta+dgfUJ1nysNXHUp8DWdvzyE81GqGJEO6m6wQ3OuLnD
g5oRy47hSr30ESGfqwt1N24wE0qqD8BNwWDQ1yYm/05n1NgkZhmKAXYlOvols/UZW95CbmZ7qBPB
8HRB6DiXBDpuznKnaPFctAavslcA9qWqQUOq6es3lY82IkzzESfsmpWsaemOjsdbeG5KJBjte121
+m5+pwpOEo2auSPPCcamJc9Dkc8495oGNi26s0TAvUtzJXuzBWsijgsrismuCVIA4A+4hPXxWS3E
Y30V+fYevdj6Bf5c3N2+K1orwH9iX2hADy4RU38LSlQLMXqsWx3NmmDfoWQ5hAYj0+CmkZdemlXQ
e3C9LdFwj9HrSYhZzaICo0vC9wuaxEky/PZOaxloJjPWXPT3E1+e83vfuPQYDSCMIiTkD4+p+ygG
abE01Bz9q/oViLNQ8NhKGCvlgdso2FW1EWauBCuNlcspS250EjM99J2ybeu+Zz2fb1S1SiZ89fp4
YodeAojOG8qqgXlQ2KMm/TxFUlbPyJeoPXMo/oVvdOorlC3rAujYrCYKfnmmqjpAhsvvO2y7sPz+
o09ImcMB/FEGnlNS/cZOd2KC4OmWvnm+4d/wM3nazri0Nc084FQE+c0i8Ws/G3LB/XPtAMVFGR8A
naCr2XRP7syThGGH+vff4i4QiLdyR3bKw8W0Vz5KDVeDLSTZYudf6QCc+yBpA35ne5lhgtRjWdby
kaYO7HdUkNOlR+36Z0mdn1CkaMi6xHoomD76wxpvFSdvMLSNXPJmMFJte92xmSbo/AvgA+hklpGq
NS3Dae1swzeSIwhTMDz/RQ7JNGU/pZx7pkyUDpLK73s8ggLOzuPyzluu/WVOFuLgLFbYT9ecP//L
2+hIm9M39t4cT3Q+jkU5+ElK5hxOHaA1Qn1ebaTwT88LSTcHRJNU9q2UJJv+PgavVyUROuLvoRlj
WNttDlYScGxOztbFvdRvEGQLBM4uKH6g0uvgRiVT42I3hE+zsHx8P11WVdPiFEBRs1hvAeM29W3N
4QlAD/50XtKCszXSz4EiZ0xKoPhZhiX/yc8gvERWuxus7lSZpJAi5+QCPFegrfu/Q100ViEKFEP5
79nw6vVjlbiwNmPhu3FAjOBOc1XfKyHuYP5ThSnwbVo768FJ717UCufJOyxk2vc88z0KedumS6vJ
UPHE8CmRS/oIWjWtN1zLT8KH/YkVW6Cq8n3rcxh63YAZJWRlqUfW+TCxy7+RGA5/lLcLjgrxciM/
klt03UgxqFNWU8yKdoCH3busWatWiBX3j0+wFoSMjCWcnsCNYX84tf64B+sRKhOzwNRyGvTzli1o
1BSN6kF+eJpCgNTI5zjiR7H2La+voVRTbguvnCysTu1p+twxFI/1oGk8YnUt1gRaC91VlQyyimLG
/KZmqwCMYhjUyC305ITH/lR2Ho+Xl6aVaOnLyPJ9vh1Jt1d/3o32MfN/3+aWBxLGyE5ZCJHnAh+p
lEFiCjLIzFtkNglC8JqnET4XTzZaBzzzPVm6ko1Uy+sodbz2+0edlbdy5S63wIGvCaakb4TJAG8u
SoULNmzk9hUxQD5d5G8ruqm+nu2ZmgYSA7TBSgi+c/jvvRbkpg1EsJWr0qzOaRcKRnm1/p+hMqYS
dgsG4nsQE8UCQMIOeRawmMr1oNOFM1cwOcLykyNsjkVdj92yfobAxV6TUmYc9b7inyYaYKuSCmA9
rYQWdskJWxiCCGeJgLxdkSocEk0cSWnDRYOIoCXAn/mUpBWYIluW2Y6if0bSOnRuHNXe015GhHmS
fN40l20b0BnwU2By5sNGtQfcEqpobUFRegJspcQJiLzJDuwLUHYQi6DyxKjhbM4yK/Bye+Aw/xGE
7OmpNNmzMLUPT3xEp7QG1OKd2akMU7qxO1ANqPGdY0tVjKeMOs34Bamfoj6jsX2y5fgS5rb/2XuA
/+t5KKeb5CrvzFDe22XW41LR7jt7xHKx2cFhxEdNocebx2b/b9VKb5U2QEd2mGGrecFpbV6qYXHB
hmqwosgnvHQE2jsA2vxMVeh3Ts1uwmd0y9lNw5/n7hXBLg7kenIa4zeOL2+2I4tZH8hF43GRPrvZ
eJ4X9zgcyjpwRlVYoRX4E4TRZB2LtfKRar6Xx2yCKNZCZjPiT+LpJ+m7l9fwdLBiv+QPEszZ8fwK
EtC9IKIMrk01cIXN4/CH6hcYhjP0V6t0kBt3V+Oqt8K3HGP+J9mFhdDPvgct1SzL9Zy4C60ibgJl
JSBXwEMf5eG6/29/bWXxF6oAThxEU65BSojCIPD4Q4FI5Txg3k738iOu43zkn0DFCub3J8Alvh4D
6hsY7NOU0YPJLa77C4fDQ5mBvcNZLrhS7As/dxpyTuOOdJ/rBiJ7ueyJ83fO/AvLyal0SOvbAgSm
8UgMNrLKHDg8rpXOIkhQcmTFqsICKB7yKgNECHLXW42QZ/l3DiVHjAeGeIPSx6lCIrXyqTNRi/j4
gjmVYIW1MbpN7w//BXgXIg3lYnzXp5cWhQqavBOx1D9UFdsraGYPyrO+lOEg6s9M2lKuUI3qYWnx
fHXOXdUa6BA6GZ5fkzbQR0/dd/7k/YhNZThRiTTATFFXO2EUMLONVc9LtXgCI2AFwZ1aQxmHbzuA
dE2TzTbF5VRGRn9hDevDpEittDN82IaG9JrjrtZpGFLz0FZfDPJFILtnqdwiP0a9YxNmB6A/DZRf
fasxzvaGPQQtckEGsk0n1OMnGjkUim2D73asNGxLmnaOp5dhTszz2BIXKxAHeGi6+Y0i7htf7eYg
Ou3Cr2qlroLnns0p0ENPK3L/gqvzEs7NzLb2G4hoB4bLS2Sa4Dj2zjPTwjO5wu8RGvXOCPPXj2bS
RMX8qa7147c5l+TB9Jbea1TyEqJLhZ3HM294fYFCetmSrcSDxcaImXila8TTFg1rOrhxOCLdNCM+
Ocv3nKnyf7GsDz6HmVM9TratqMU50XsNoPcu8mPCPUxkLHj/gNPVRzHwplICWm2m7WBAV5eFjSeV
yadD9gPzzA8GmJAwe3LPZMG/hiPRK0Yk96ovqaEqdQDcTDUf2RJ4Apu+0cfxujFArLejwkxzIw1o
1IbVZJ7L88FnDMqlczp9iBMeZOFTA2cpaD1r4oGfIZNaBmlan4jRn7trRRP4qSoHEXK0CIJP+s27
oBFbfGls7e3Qel5s345UvghXgoz+iR1+9xD3KWMm5cZ5bc2zBoLlcrowl70ho6yHbWdIEAa9AFGM
qTvDv/KbferUWzDlI8ulU+9wozxAnN6qzkFi2qsCHdpfI4Qw2KVihnql5x4oNU5dpgUxjtc4GqQa
NFOL+uj2O89rDehdbOIY1u6cR4oKYXyblljp+M0xLTo5iKvIfF+/QQRaY4AouzdzHXGCcyxBSE1M
XivU+RS1bDltlKLC34022iEZlyk7b2YPI+Zkgd0GoQcXK9AYG1t2nTU/36Y1oNOXKihZ4hbFfFpd
mWDZkV44tK0zTpdZPYtSFEJH+aCURNTpYNT/ciikoKXCE9O4aDY0XD0XB0DmJ1epdHIrx4SeCKSG
l/e1dFioQ99ofxrBWeZBg7A2NwnVG32wuYgonCnfr/F6vD2dY4hFGt86msdCNFb+uOTEO142SEWD
BWje52dM9EU0AOe3mtGcS5ojDemlfzQgwMMywtnrAaf5STNZipUvnDLB91SBny0A7HuMSBGljfuW
GdfZMFaDqQ4NqnHZvHkHh+icMoF/bV12duJSb54/qcjxGR1MrxhLebPiX3ZXOagkB+lET6X9l4XN
2xdh8U+i5Us0PEAVNwGg14HrTdnSXg/tzCbEWpbU87LNXNlRY8pyVpKbH/SGTZm6eceayKr5jBfL
yrZm+xDVVGn9Ak54QLIv3ZoPEEJCWkeC/3dxZg7idaVL8thrX9SC8xIYgQb6QO2SeweZuBMQOqrL
h/31mRntd7vBUDOS824QLE2gtWi+Nry6G+GemMfUNGv1iZREda+y2H899ZtVXk//DsoEMHQYrrFT
AqfHBFO8M1D8Ado29KDgbQ7cTNX9rJi/4U9eoBSoju5z1kTpp51WJUliTz2K5pmgS/jroJrYs9Hv
NE30IrO5k3LrdUgY4F4QrLc4StorI4JqfQCGT4MsgHOnolgwV17nHPp9ikb/IVO7/FXS0aeJBQnW
8yR+5IZmZ7ylXd5/GypsDnMZ/Rb1/jivl0qGV8iKuBQlQyVHSMgAJcz3Yezu1ZPJC/YFtymVsRW+
s+oJmTDsFz2me7sD9qpCO1e4gRQWnYVENb9ZGI5q02IVbk76zGAlgzTnT9ynONauZJXZsDrBzbeK
5vT+9IzOlycmLZAxHM4UY0wtyuxd21eiuU8h+1i6edrgTaHo/9Lof+m84GBfQng837twvEruSxXM
mQw5bOeZP0mNfcUjHJ+LZPJpsl4AlKYysISiNCfWmDK4SEGW433WUhNzs31XQBupZqO0Y1uxJ2vt
Gbgjv5OceDZKN0N+4YS7LMEteiSzURfkronh2ZEsPsgvrT91i6Lze6pyLsQIovSrlf68mAdltD5b
ZmaOB3NfGf1+jv8bWLDUO5YrY4Uyrzc9+C/IwltkLF5oEklixoVW9ahumMzA8yqeZpzFm35qqMtz
LipuHKK0uOmRQQHO6qLXkmN1NCv179XNLjp7r5JoG8X5ohwtKZ9Apedxq7Dhr+3bIjYW3vg5n9Dm
6uA9qLVdasoXKd+JlbiDY6+zOLPJld8iFcbJ+MxpS4DBnUL3l7UktV8pudNJXymUAOgomzMsJ84Q
v0uniBaxO2CvuJcKSTVoB0XyehgWtk1q8ma0EwwHxEs3KBvy8NsvUgJdZMYEfuPgse+/1SyW9EF6
rpYa0HKul7Eb0c7DzgcQqcs5BopeznMnD24G03xS86yUjW41rAp7ytROJWpXszTybKKc5Ec5l7de
aYOzJupTfkhTuXy2hghgxqR/njtXtMMBwWqIVZfiG5k7dBdKoLpvlNl+eDwpWy6svwUt/ja6ou0S
b6kTyk8mvoeohKraOkDiHMlUkYtbZ4CeaDBaIUak1MEw4lmtU+5hvwHW0T5/H3ZAtcQiN6P2AOsg
Mxj6Wy4oyFW1pQZEYKQ9y5lIUa2ivQoJwwqJhhfuJccUituY3ZQ0CG7NIPf9zypwfSL/vPnpOCpt
8UOL8/3ANXc6xpoEWCmv+S49pvfh7hhb576pqGxxJ4h0jM6gVLOXw5fzCcTCuT/97D3+Fm6IoaeE
42HZoYOqun8BmudLxchx/Mp789BkW/82i8Hm5TjH8zOeckfP6WZi1vEnS28iUQT4kzmlfbcx8L8Y
Jcn7BWsjQW8WjegrrZTQaXYEac4onn6RsW5yFqIKuUtQlt7KL2iA19JqnPJMUnCo/Rjq80qPIvIr
ZMgYbCcWQ4wXD4ml7rsAGtoJ+Fvya7HNVZGr7T1cEUi4+wNgzFZWG82BH87cMueYGqjxTGzz8VRB
PHyP19WqUGxaShzJUG/2VZUku+mEBSxgW1DPYYpOMBzc8Bqr4xjkbWGd3WeAgLH4jX8Dt4k1Olmd
Q3epr0/23Vr+2zr1ZQTIqoAV0HUVnC2Yl13IBsALD8q4UPTp+FCWC4fxDdIGoIkdEWthyDQRfEjh
6FAZbQKMUlzFrfTLv5WzSbf2cQ+ysIvnHcM43kJ1EiTUfFl1R5G2P9DnXNfEWRiUxg7qdWBogfUn
Kh1HkflxWGp2uPqxflDirt4sYRdoe2/1qIEtvZx38dwBHwxem8Fzu+iPjiPpkeYrs1Hcps7H98Oo
YLSkNLu6OwaQ7/TNkuUQdd9RHu/0PmI6NZaQ0Pn7eea2Dw/X2wxDiBYvLBEEFEWQ0ZvHXiy0nRcY
Nn0jssvierIztUJuDtvEfRVEZAmx+zRAFz/2pGjxrVlLxJSZNO5k6BDuN3eFzQ89TScSRld/22XY
lvxypvlME82mza5y1TO57dyKfNEd0LolmBNj8rrsGM3RZphaozX6y3tHkW4QIV4J3as6kDouJ84d
sivDDEqOZx2wx9dkpvX/jq0v7vMrbnw0xRCN/r1J5LQC66NWVvOCXKQWp3hSgZZMBYNfwM/yUm8l
CDra1BomeThC4fL4qI/AAHZzW5HGU+aKEbT/WuWTnjrB+PaexMYAu5Vzq4ySPuaz7KcI5Lot4OD8
mSGDi3rTJCtUxEqO/n3Br0/orJNSuT9iTPFxPtP0enl/bBcQwF9i4omC+AMg6DQpBFo0/BHMgz+w
KV4eRPIQbZjTZ8midWGDVfoNh03cb0sUcqS8xCOrVDZX0WuoSsINBsvAm6BLZjiVWwz0mGaFPoKh
6VdvTafT5nk+Rk5bNfUp8kJq/PTk9xi71oaVYrWyaKJ4jPM2tCpXEH6kI2QMMkX4PZp9Jph0EV1C
vF8O87MKJ30kh4i9Vm05q456L8EXfltkIOAutlF+9MiLIAkw1+8vo8lFmEvZvY83XVjb8WjPHanG
FU/MgrWedL5DumEWZSus4vCoBAkiVBqZ4MJ8+rCEZoGfN799ftl0RN/lOncjiPPWAUHC809y30SP
MNHsQCP7wQQ9AYTkWRzDeRxboGbci7d7/KnH96BGzntxb4RSEanajfsE+9bVC8sgV64WxmPAQS+S
58HKmM4062WOhVyzR6ajbol6SbDZxudoXhFIF66TlpBUVTHXPIjw/0HpTv8HSR+ln4/7UacCZSAE
fG5485Y4XHdqwzaMaAYf6MdkM14DEoi80AkKjBWJm1MbNI/4B6eV4Zal7D5mlankxIaxf1vFl5ef
Y4KkOG3wq77IviHLtAn0XS2Gz9A7G5Of6e6epJRlDvSRYXAREvR5LK0kKBBPTBAFL70fs0mzBT+U
0+Wjlc7LBdlIqs8gIcaDUDx51VcWzVAC44a0pvjKnf5dHS0nESSk7dxzr+BCLALRLvHaJNtwQysx
IRpMW8Ty+32h2us3MXoyl6Oy0SOEFVb8gF31jDCn84iblDyJRCY02ZXnSrgQhZNEkV8U+LeHV+yd
OR0GpcUBUHkwSm248bS4Ydskokk+EEeGYhBVL0SFdUfoWy/YuokqeTOPxhr4nmEBf1ku1yvDKBAY
/57qzsusFWqeff6/wmtdQy8y6HZ1yb0a9DirO9FhW8MaQdlwv8nXdMBp4cCxdHjjBXSwW9EF40bG
I69FWRgF18E6KT7+Dyr/joErTgOsWxHugAshQ8lamzn7GRPT8KHsQCnqNI34rHRnRZ+FoRAtbEtW
Qsbd8V1GcHyxZHx4peI54iGkwveGAbFv+AVNvFBYIHYueUTvlgFjdMCPkV2f31ZGDUOhG0IDmjPC
h+aaL4FdqwrHmXXBI9Ae5eBH69a6/nGfNTpSkQa2s3aoJiv7J2EruIZY8NYEia+TvWCA+io1khbi
do99bs0i19Ccb/ZdYv21unzP+vx17R/n1ln2bx9kVMT8ErOVOJQZFEDhs38mvOkdl20K/hXASdgT
2f+ExxcNKjwoakEXkepnJQ/jDGE9JXDk6EYGA7uzadmsZ9HXsDgWLWQPCqXMFL981S3PoFSw3BnC
u2+QGQtphEXNyA0kufE0iOfkj0LMzha4l7sFkgauqB8CKpR2ykCLMzhYJPnxY2vE2ORAedxqJe8Q
7T5KIXRyPj2jdMENa/ClM4fwn5ll5xzxjgeOznu576hGduD5Cob863AQt6cxu27jR4stoSX6jOwE
rQu4Rhio3voGwjF18x7xmQ+ZuVC+KRyn8IvYn8VtMOcU2et5msaeITC+hjNWITmFt4LrCToVz9la
r3vVGSE/OF8Q6zCFKcKNuQDeOB7BXOrAfKakR1tYRlU8pSyupU6FwgtxolGKX6dwHqz0WpOn8Iyz
2q/sTWO3h/h29xL9l1YIh8jmhgK628uiigHZaiaVhvki0E0/MWl/hsdFM8bYPs81HfBqf3JNQS/f
m/akGA7fOTMz5sNdiHZ/O8QE712opHgD5NXNdAH9w9pOgA3+uA5f58mpmdkwimY+odjAPPdv7Hcv
w0IiHhkKZgc3NhM1ieItfTxjI+kz32wZhB8SMaZzOEzRvemfDaj2YlmNK0SL/5fQoLh+vr8JzKxP
wgtQiH7sHJEpK92fCxe+Ux6OVelFCRFdO6TuxlJ0nK6cfi8o5ns6Ypfegu2/wprN0iiOVqAaCSCn
N4VqXFZFZdeejmmOWimT3IiJFzgtKczr5eqTw3JrFoPGXK2aoCPkH+ntyuh4mxdFX69Yem4kw3VO
8Avb411G++SVX2WQlrhU1RYO029qOCOVoH0EMyy1gLDot58suk6zKGplChtRSlOGcW8ibeA005Oa
U90nNUCkem4XwNIjzuaFzfpKpQF9bPdPOAHoO8sDokw+KOf5pNef1Ls610d97f3XFZAKsqi1Z0GJ
zU1uO0TE1Pw6ISpldXdMQKe1IKzHSmity8qdNkkua52lL6NDfd0tEF7fxlaoTRNiXgnNp1PjMbCz
QsjoPamCsHi4gsdd5IeCNcyuam/gETjOnLfODtIQy8JlQ5yBe/Vm9h4Y5mFV2gtI+ROqEUZaajb6
J/lMdZnnfQNQF818mM03u+XwxEXu9u8x6gMzSJJRoRyHqo4EbRhPWGXmEEAP1H5KJWScRn+dl2+Z
dYHdrIS/toIuMTOD8s2HPR3M3w5EQ1JblFnA3mO73htEmgyjvUHksqRd8w2BF0NF+DwiR+djjY3q
GCY+lhT32HpMmxgi+IRNjNVqFSoHrDAMy/LUrAyCbmctj8Jo9XVFt9vFlfthLJ6E1WDrpyyFotbY
F6kfnOW9xwWnAzeOguorDAeoj3a95QSuG+mQnEL1cqgihK2IwTvoSGSAXK/13n888U1piyW5h7KR
pfAh3LGJE0wRp+kY2H3EC49TlnqOaWms3aMRfkxm8JrECJan3IqcI+yzxiu+ahHcyWokE0MFzeym
d1s9xIm8o7BzxXsiUnR5lsHOtPAhkFS9F6TXadtvGexAyUA3utN0XMLTPIFwANxBP53N+g55tVEq
kl1ak8JxmQmF34WqpuxoOL1QYWQnm4D1xfq+dmwpKv2j9KbLc30XyTSzEmKJihtIeRldKpFxmiPE
Ro4cdZ79/7rRUQTYS1naF7tvh6r0QNl7spVQ/QYfi2zu1Krea1KrS22hl6L4oPuZkSvqtyXZid9d
vY1LCe0Ydok91DjU8Hx/jqzeh/xyFV5vev5xTBgL72NnIkg1lj8gX8qQtLroQdnp6nYDuIqpTBE6
NLyV3AyWUSpIsNWhHnvCINGQP1C4RAsnmJBncwp2xWHhgnm4bxsXnJAthr80KvlOSJ/pjmiAWrQn
dNBgov2kTj5WgQ6Ozj2kLbk6L8ol68t67Or/+W+BAWZlBcKgtSVmulVd9XThDHKDejXFaMHb92B6
7ulok5g1uKx11jUwGJgRzH6zTvnKWO2akD3za35b6kguSBAUufhKEVhoeH4YbMorMFOGvsROlO/U
Is6dqFLjN8XdJAWPM96E8z7ClB50WQHSvXN0mRSVt6c14frjb45/IwMeQkS+4ym5lZIJdFZu8o8p
8GlZEcnuP9c4/q6OVrILoH4Vv8JjDS6poRzoTplfLnUqw4gf99QrpI844jLlNRaoCSmJ8QHuThLM
I1l6CtGj/ackENpeMFQzJ0JR8utBVyYT529/tPY7Db1DT6Zh7oULDJUBO/EEKJsFCCqBFjvpYxP9
xj6OvXCqpO2BGFMRbhB6TzA18zhX55jqWYTOffo9GaOJLi5T3ANZMrV0N3dWoADYIQE7IPAThqVN
Rukj73d0IeSlChGzuRgwmVXrTx/vwOq1HGhj+9/YQ8w26Bs9HPwiIhQv7nKJNK3R40IlsfubLnOn
+h4H4PwUjvEi04nRVNLX7ycTNShbTcBtGYAZMaNHDL8y5hBo4GQEPrcgJpO0SBa2P10Gw+Wfymf4
HPJDqmiuU+4DmPA4c24QYVdBqvCVJpVPv37RxPzrtFCNXkeI31KjX5XoMcEZiSdRvpCXvtRUCcE0
5oLfKd7tZ0hnR86DdR/9soKCSeoRFB+RIxyYIQTSag/YeydxnmnyamZUAOZJZz2reYwQ8J2Y6AKd
RgJDZpg5u4UwD0RwhsrWjMY0EZoiu5OQENSrV1kOL7MdOQymjee+sckKfpHD3mr690hYqJVi653l
Y7/WFD5DH/QnAReMVcO2CZ3W6IYCWMGe89MwCbR811eXjVz5YHtKPv+2r5w7cgLKIml12gkIJ0gJ
hQlE2yLzOmd+FGVSmMyzO6SvtIsBAhOJ4b/OXOLZa9ah1vxbhkELymfq9EkdosfUR3SAucCvmfX/
tgNH8jnVAAOthQVV3gIJucHL9TNuyMgMZiOOyq+0yEIE8HSyAXdwRA8xCXnHsT33wBFrCusaZwOb
QgN87vUfM0qcybVRmmcvXJpYnKjlQGzt4iJaEYnw56pKZSK/Mu6/3d4KNPf+KdPKDEZVE6eMyVox
a5SzHEJ22vmeZqR3z6/b9sBOPIFQ21Jppz7ozCRq5A466NqkId9WuhAsNG0/03X/z9ZSbwhcTHAg
MtWJl0yn+NHvgBNdbo2xZToe7sOS7YRl6xeWJD3Xrtki7xT8APBuQaTxsSzkEDJcU7bVn2qfln5Z
W3HnLE9y7DaQMKkgLIAKZAbquk1BCZ2CnJSm0ssJ4eD9b3r3UCsc8+dWK6Nh+jkFUNzZaL8OYwVK
x7UWgcdslfQ6nVVgZaXUL2RLKk0FOzS2aHq/ftWEq/UhJv8zxPPoWSotu4EMEjkZfgLpmpxZ+OBK
vi3g/nRBwm8hG8hWs3UCjej8AbMj24IdluxjrnWeosfMNF+8gdckU3WW2dzD0bnrFk42QUcLpF/4
a+Tiz0XftQ14016/EGCp3BTmyOOxqHr3rniBIGQs+nvVacLCGCicfKBc8Sdd5DqKS6aI0bufolYi
WrwVzaO0PPJRfEa9kFnVu2ohBVlkyjT+iQ6BTw9+LeFlIHwqL+cgO0GjrTpts6G9etvmWH5Mgta3
GvymJFVBWjcO815dYShtXbW5V/b4dJX0VNhCIVnmusyfCwRVjrOta7iB47uSaOHjG9zFsVnzfllB
RtP+smTgg9hVwbjI7n+639j5UsCs0vaXgb7WfUAbSkEPposXU8LFH0lLwKCS3XaYN2R+EwD1hndD
KnUCkhHXS2PmeSrfAjA4cgGBBIHqdB5bep9ngJUjI6o4ZO/R0qb1uMjfXs7ljwuprQC56kpglqif
XKAwNNVCGoP+aq9CxBaPzxXZKTy9q9XXtYlc+oapA4vcGN0w0lRW3s8qWBsC2ZRWhPQAK9G+eXHk
jUQWUtYeiUTodMf73oM59OiAcwkCcZxW+x7xuGTNfKonxO6TLejY647MUBuX/Tu+W9X9BuBouRDv
WRUl88/XakNz6pyIQcwpr908AmxnIWzztCdolorAcV4FC/sHdvwAqw20vPi6Tbd1mOVNwycqxt9y
QCgIOG4YL71i/DzT/d+tf7SLzSdi46TBxw+AZTQ+nHLJJFwJ+DxIqyR6Dd5AdGbLBCMZJTyDl6OR
8D0N5XlgDtPmmc3H0E57PTesKvg2OStTzvuUeeTYYDlRq+w5nMsFRNl27yvU2IWpAqUA7MA2SXf4
ri+0SGVhnK8u0ozMk0LHPSFeLcSjv5rXI8yRsBIUSuSeV6nTRDXkZzwThuKaCuRnxa+wlLcUyCgH
2LwZGn36xhGcoNGKYpA76LlFi8shHJCehbj+SvDGB7ucrYrFXG6ZV5kfd4Vsc8cQ+lfWXlgoXFr/
EROyAWrP1td6eOEZcqbqNppIHy9YL+K900p6ToizeWR42VXOhiYN1nE+97Bw5oGSll2u2iiq0roo
+lW4fqbEbjG7leKjpqiD9kjg8MJttoVSGf7UhuSK+BG8PRWpFRopoxwbxNyO6TBfo3IfM+mbjfmf
vV/FWx5rwi2f/Z+XTNrycxvpKbQ0M3Nxa2yuMGz9NdC2U/RO/akntat/gNY5q8TtBgaUO5Fp1Cg8
raxOByALlOnCmkcdmQBsk8rFeWFDL63V7lLmH3HEPFoKBKTXQmqWnkc576gKOgreTDQjgdcqBpow
z4vkIb+LTuFlxdwaKjyCwsVHN7OJbu7p/AOjH3NuaqhAgfE3o1tetq0YRo3nK8QTIUboq0sBoTFt
nAPORCKHzz7ydQ/r/CvXIeZRTWzaAteBq5eRoctZi21H1FqFOI+LpWIlrnsbNtBfP2BcFjPbrDIr
uRsERmaQgUIZ0I7kkhbqeffPtf0a0GJEjcY72cHtYKz7IpYvEbh/crvqEFIzsGUPoKcX9GX2YY5H
oIkmQf6yQ1KAENSFksSNDgfpU7dFozDa2rqIuiApFa2smGumWZbto3PMHa9QC93r9LEmOPTlTW/h
zaHPp2VihtK6Autdmy13qUZAOZMzykPZ3QCEPRAcEY2OcKyHr1QRslQWNuULTNsjYO6PwYUkKLVX
+I1FsDCD2E7vqTTLtJrUhgd7o2TZIYlcWFgmnW39SuvTgqS8LMoBUU70PX5JvL5g/qivT/v/gGLr
bJdD+3XFxEDnBlmKIr82SRoNgiwESS+aPEFPAKQadkopW1dyXJrGjpu8BSPOtfM6ffhW9KEP28UB
0ND2SrJU65fKFUmMGd9ZpcDUt2XKkHGa9s7+u4UH0aOqskb8g0H+2z3ne7HmxIpVvgavRn41TsLH
htBRpe8n38SKhX5pOuqLctPnrQPxQ8EDSU2Kh8ZXAKnPeYXXbNMCmjOPq7SGQvq2JcdL8Et94LPf
hylZuiwiSmU8gSaKDjaMfBB8M6/C7IjOpylJ7CL6tso+wSSH6EMHozcAqVmR+lkzByq7sY8w301I
8+uS5ad7MlTlyN0qioJ11m+6/Pi/ynykSS+SgMfJWLlVHHKcpW68T+np3a/XCeHm6nb1zJZyPmMI
P9qcD1NGGHf/466vZm3tmTCZBhvPfPwSVRg08Ip/yMk37kTQwMLcX76hCKlE0Uc96f+kgeV6MqsI
XVeSWIAOe0wQ9RjIuO4qlFDvlC1ov8mBv0i+xHkJITUOPk1KuQgRfoO+Zc/bGBxZj2fLiLF6Ctym
+j9qJTQ5Zc8PQeTX7Rp4khHpe4jMPhEiau6eCERlc7nFWVGDmDdYBKNierHCYMvonK1hD7FlwNaY
HtQ22wTA2TzPxJlSA/O+n5lvAOIsguTmO2Sd675jYsWW5J+wuk/ywzDrVor/WngGR5qJbIJyde/L
3IsUCjhu7iSfD343+VSLOvIWnSsBXFhuRw60pgWnltLNFsQ66NZdZnG8f8I70jt6qLgwQQL0+Y07
+BZNFtmZ+EQhY61i0UH/HMSn7WtHl1Q8RIKzBLoFRbU3ni6npI2mETTXLt29xUK95FDpxj5nNZkA
bCD12DdpNO+qqZ15DX2qIWjXiEeuUvxI3w840TEgYLeKjkXPjNzGlhSmXm9b45f6rd9MqvQmqQXb
KCwUQdf5nrucNzJ+i9p0Mi8CAajun7DEhHd9vL5DEwK9TJIRsVNcLTrEyXSBdqHg09JFaTqx+WCQ
vFhicI4UyLSkowvWwkM8NqwRrm9zwFAnRneVLcn3Q0jShNiT+DHMh9nw25JevU5JAp1zssX7Abb0
YFOqkiTbPGRSMczGld4CdDeKbQvHMdPzBQsRKuvq01TVuWJ1YigW2UPXc6hWhK2yv83jrxA0CsEq
sSy6ULpybs5c7m/TCERpYZb2yZVYQ6CVqyx5Mf+w2RpowqGzFdzwSK7Y2ji7Zj09Bp+cv+czxTz+
+Ne+FLhlI3ncR9q04X8czkik8sj2LTVe5C6iG9Nr4tXOmF7qQXHtdLSJHHo/LaL9BjzXPsZMk31m
ZFcfPBMSRkgUd/rMsmru1IYCx4xoolQpSzXI51hCo/bGl1nZLVB1AGn4E2+Rkj2ZnOrn+I00tEqy
7qsE1q8lODZqAnE9nZ5xa2XNb25YDJ7pbJTyHmQcOwmKzvXO9dgIJdiSTClnSoFk7oR0BNSl/fJ0
WvwW1l/VEs9diewjxD2RxnDj+9TyrPL3FWCDmJQGZK4t9cKN2g5bVeGCEPorBbGx/exOOqBdhnxs
Yl4/QSHWiy3PxkrSx9MaIIwmVUpefd0knHDkHXld+g3e1Ic8q4SWqOxpakFulyT7n9FDlKCuWoQW
ZIQTnRzl8gnmly+KzRfU8UULkbqrC36H7gXCe0UfLO1eJR2qrOhg8MPc1pL1QCgU50TtuTYqZtu0
OBphfJGxmUf835WbaOndvDx+lUKF7BJ15zI+1/DMvWx2kIZcbCR++pfSqxuQmkLRZ1wQSqXJBT2I
nsDnzfYs3WQkCT460gIX4WvDrGNY7B6N3pSd9KQibE/ZCaTHwp4gbK3Qx+oBz5hEz+d2UyaUMZd2
wYh0dMOlGMpZm03rww0o+4j95IjskamXurU/giV/TkVqBHkytSU1t2GImBg6isEj/CJTQTs4vxQe
msek2vf4wB0c4pGUiW7y9taD6I0VVcmpg7LKfeI5A9UNxCJhX8PM1uJY4p3HllsmEPtYIRavp44S
92Z3KqfUmOVSdDwC3i02CuYylxA+3BhufNPtNvkTbLmXwdI7IPqAHnWR8MOUTVrG8KoJAHfL2n9U
htM6q1Gyu3O3bOrsL1EwDCr4PvJu/APmjpWxw+i/L1qth7I1YurH2b11UxkTsPdc87xgzsI6NOAv
79JC3w5fERUyVWimcl5xjlcPaBXdTzoUTYSFcqAEDDyOEc2FJ3OV4hOyqU3CRhZ8AYgsSCZg/YcY
brGAy1/Vd9AQVxDfXN3pYyXB2K9X6DoG/UghKeSTfA1irPbiocfVIXAa5WSEkxfKhZph5OiQgOwx
NB0A0mEr8Oc92uowuWPTyOq5TaT937N37uOa6wp9F32wVXn6BZHGJpQoUyF/um8TWhweaF2jpkdH
gynRQK5w0XDtnEjRAZFGJZD/9W8r96nmgPhucsrTJOWqEGwRMrF6Bg3FX9PhQt+3jP+lmHpnf2r/
KfK1ytTiiDUmdwSiS4KCGOyxWVWOXkCMkoXGL6aI1YRENcouOfhYQ8vSrbYnVCli3OJLdHmyT9MM
7Hcr5p8HouepXuSl9snmuZcyTVivwTay9EmkWrxjFDEoWcaUm3pVORknqSr0GG83npCKY2I69mxc
e3pu77ItTSXEZRJ8UmaqUZgttMPGswtRV4GhHVa8E0hzrQnTAnilHCGGq6whFFinOdQkKTSsWrTu
P+Gzuf239T03r5hmJF+cRObNmI/ndiGaBi9c6OTpfhJx7A3uXCTN4nbTaX/XtJz/u7N/o5p3lKay
lSBdtGnnLu0Adv3kMHpjbjRcHb/ENry0pyJO4x3fCWhj/8wrYQCt2775yMkMuDft88DoSgzgs0D0
vLUHeOcg7DNIqQTMR/zAF83Wxb++jUvXhVb6gt3lJZsdx3G/SxJbkkkG0HZgsQR06UqUSrW1Ypyq
r25B+mRRzqOAIVWhjR8QyLxI6l37QbsQmHvTtXVqSlvSkO05eC3+uVZHVB2pfENOORSf+M2V70eX
yWcYbk9Dq53qnzTt3qTV3KtMYHtWumRt4aCTMzw1SwbTG6HZwvpRDMRhH6u0sqn8VUVJkk5yxHDg
lF3n0AJ7hYXVgVI93iiF8THpEiTtJieSriV1sBdgxSZr2F9SYEyTTRaicN8JPHLUPYcVrYDYU7u/
Vs87ImJ6zWDLeIsfCcOWNOlSDel0NcFIojOKYLDSuGcLq7I0G28Zyxx8M+NDsrnHiGGu8dSp0XU/
RoN9aaxrLsTO1uzReM4mKwraARO4AMb62KRrWqy/8hhptbnktFjlL5Z9xf+Qda2dE2yUzPnaM0B5
Fj8YWkSV6kJJzlbiDXoP+NMIpwIkg33yEOtcAeH3jU5ckhBdrMrYbPp6TCxIujoF3odn4R6tAZ6+
zgJBj/V4AZ7M9/i8LkEoTXxEPIiTdc+PFdBI3hWrEz+GEmZK/Z3/bDPQFIvhoLahhMvoicNGaSa0
r3fyMHTHGlJ9Ypa+6SDr+HhpiTbjp/b0vY2YNI6H3oPdQ2Q7KfWgX/6EjBJFvSr3jexXSKF2pEG4
mZJnez/UjTMVvn7wzML8wbQ1qPl7P23nKQ/RT5qFOR3nHx5/D8ltAapdkBId7BYfbkdv3Oj71NzZ
PT0rvVRtYZCiZlZ5FPmthkw8L0aCUwKanU5JhR1IQPixbAJHm5qJJiZV91192+b5p0KK7SsCz4Qt
5xloPe7DleRh7mH8IVoRciiFgiOzGK/tHQkbGpVG/1UtOwLqANZjmtFEFn6KMKLPeXsEcZFQpN8a
K1H6uCGFnDC1Sn8OuCmKFIJrbeL6JLLRSg68JAthJi8bqnuQk61whausRg6iQuI6STGCd4zgV8iL
DwkH/vPDgzouKeOvXVdMiHygcbNQ8XvYbIIK9GhZQqHSsCMtcJha4DKy5yzijuJWLgkqkase2bXs
/1nuT77P9xeE3zL0Ckri6KV0Krcl77m7Lw1OfkPzANWc74CTHRlE9ci6SJaZAW3SxNLANkFZX1zo
/PZXiEhfdxlGDZBh5uStLXQo85enhSq4YetvHK4nS8pZsDqmyPb208iGFvl7pwzoFQiEzeO3EVj7
baZABF47qojzuRAYITv/P5rceNKYLeOHs7lrV620Zih5rGfJ/i2RHh1CnEPctEAPH8c/00VLwl4s
lW/Qfkvf7BJhyZo37MwIeNSkE3wsJWXE17WimywCNd2Ta5e+MGvz31VYgAJU5fAvrzoZigj72KE3
N7xTSrLDtWzGrdqpR/FuPfEZ0A3YxMmKqMpPWJzSsX4H+1U7WAr0ESSv0Mpq5eDdhIXTgmM3R6cC
c4Lq0tsXy1dn8VlSfuZYqVhGcn531tNgJWoODokxJfchqW2HWyFGJvWUihaIaFiJs24vS3ZstAjP
k9UNDXpTAKoC1lur/gQRigeFvDA2mvQDz2xyPaKUsofOS73UrEbJPqvqPVRJISCGbvNcml8FI067
XxwC2EoBrgFLjfGeSvBG1E3JSsZrsvdGj1R0yMFq4zIOGszOSpZjngiMOE89724ktZnQ5opft3J3
ZiXz8AtYxjiEeMEtVuJfa3bL44MVGx6XYuqYZ+MPwnzvH5C4NA12LqXqVpo/zLRmhc0SX5H+spTv
V7EzTBn9nzXLnngv32oxbTyD3y6X6cPBphdqJbaKkPvt0GLloHDWz5vRyvmQxsnJ8tozFGswyGxF
nPVqhK0JMsCQaq8whXXsdKI+dY/FsJlzN61JGmaSfFDZwQwx3Vn7/loA1zGI75QogRYHRU/HvaHS
Y66bKQuc0NDvBAXR9sHPAqOXMNGuhl1xLz64d4MvKmBoEzlMMura312JmBWFQouXIsx1/9iz+ZSS
SwQTFqRLrZM0bt+eJRnG7VSV2R054i0HULPbxjznPBtIBFkyNYAGfzNBP/EGVportEzlSGFil6im
HPRfyOtKjIcroQmjTSq4wOFn/bBkEA11PFParQpdZsEf4HFtBte7mGK9ASup/WH/aiUgeKx9+Rd4
czt2amJd4dVMWFn3HB0t78HHVtQadEkY4BHfVrgMQ61/f2OjXh+uhgtCxPNvQ96tSj6jXDWB3Dy2
qoHd1f0T3W0GBallwuY5p1/N64hXeKpr23VLfvZ5x6g9HJo2xQpbGz91WxFnCBZZeSsnuHgRlBsF
wgpQAA00dc7JRU0C1a42BHUkjj3OhPceOIBmsv8KI4d1cF4dCVqO0kRyWhN+m/vZ9ocx96kEhn46
rtkLfE1ZPa6r1E8g2xQK0iq9V40cdpXrbhG3Q45VaZ/XITJPey4AeHe6CWLEF6HgO4ZDaeOHO5Yw
2r2aP7s96kpoQcvWyFcp+Wfsww8BKvPjOjfffvK7OaWFfxcDEIpAdPh+UOH5SjDOtanwtZ/At7em
bjaTR0+Ow6hXnpqrcF6b2/QwLfiPdMQor9r/LNXOaSuvADnWOg6/jFMan3HoaCz/+yTy4Rob79JZ
JqwKE68djVGmoIdbXMIlODGfuKGQZUuuyNYYkdcLBb9qHdNgu9RhOnVpYQ/kOe1yc5991BvLPxiI
Akm+pg7O3o0K76a8P+R+4l0yHwd+njPl1E4WdYAVkuGPdcnP8ACbAKgTNsOcwuW3G8mDsvisKxwC
iVys/+dLHkEd4Pn8VyeyW5EZOx7z8Q2t1Y5hVHk+3FOS4HSIJS1LoEYj1PdxqgLpvP76jjBgH0yD
flRFzhPj3dykNHMPIGBy/T0g46YUv2qzlok6Y3reZvxSO6JqODug+dyg5RlT/MbGav5CCXYhlm4A
PccQoE8eONr23nUudKKxt1exwy8fC8DdYeQrT4DzLDMPCc80c16DVOzPHMEySfZmZYP5uD3ifHsH
XU6h2r8C48kBebbyP28UjuBF1CyYEqAEESisiqra8OF4GneWgomlhGGjM7IzEuGE830DiQ0YpYKU
Dp45sok7RrG5mfTbLKEuzRuoAMtH36uWDirnKXUbj8B8stPaJxkhghWYs60EIh9GOkVjrcAwvLUG
2xLGxmZkWMNMEbfgA31df5UHhVxWsBbpjqbmMmRw7DOwiuZtComoFnY0weJ54apIM7cIyarXCjD+
PIGcEuYO+8pisCbXdC0ea8IF0GKZt58VNkNh6l5eGRaQFmnD/dTSo/ooPftD0bXqgn9Md5h98Q3P
B+Lz6I4MjIs7ji0ykv0zm7sVkkIO5XjrtvPMSDFdGr+9IfT2rX5HQdDSDCy6qjxl4f5qar4eKZ7c
EnzddEDgq1ruxzGm+DWPPhhziguuFwAMlroRTS1ageBKVQWuum0Apv4Jy5TrajOpYu+hKCITbk7U
C84gCFvUxJHRuZKOGCN4yly+60gfX/rmnq3F4Lwa2WnDrf3wKWCP6l+htuWKW+BwHiADpEAtvQya
ioXfGbXjci9xJsxGpJ7ExF1DPd9R7bmx1y2w1OWpGZCiKbsaZK47siGm1yIdUgOGBSJK9rArGy1l
JZm8jz0uTdUg9lOSKDx+BVaDa08t2mA/HdDmyrqm4DE9IsdID4LOCwLetoaiNv/g3VRuWfeKMfxL
Lbm2+VhYWEe9n/WMG2ltGz4uclL4GT1XWPvDb6vgqLaggMbHmklbqDU/EaL2h3qTeLyeI7/q+UyF
A7/2ak4oF3nz1YZtu2rgg7K8pPDRz4zemnfbgfrShcggYBbo+d9stYPqUBUfWpvODeeLQxZjSs7t
1t+KA+WKvvLkfsV1+a+Covvu5PF5PJkuRJlPbRV4gXYnxi/HzgytTuMPw9DK5B6g4ffqpdI29cuF
DqvE0Ne5lGIUTX81Vhpe2r3VT6d0C1IpFapKDbbnO+UOn3ScWbFZFMSZ9qI3PbHx1HaS+2v9Hjz3
7Mp9B9sXJhBOHasTD4Pt8r9E9zBUCkZ+GF4FY9diUudNVkomjA6n1qKBDqNFhF5fyfvq6UvPdSLx
Jx6PyA76/1I2skqmRn1eZiFO22tScNAsU+PMkAJSzMxfh6FGKWmLC+ofjncn98NwG0TsMFZSbcdv
EvLKtsoeIorInp5BXWsPgIoWRe9GKSmB9EOTpfaj4UdQrIHMId0uC62/7fu11VddpPcjevT4o0Rr
iV3tIXI4w0Z+entdoVYUJeoeHd4RH4/yIvLmR8+BWe/3NOX12NHcHII/a63oxm25Hnr+gaVxfcXe
+6oGr5+MCdS9CpSI9JyIm3sfu0t0mwg6q7GF5ju5g2vCFH804pMxE/7UJ16SSEfR9Zcul5VYHRjs
JHhFgzB3c+5bA9Je77gierIw1G9qq3azSpxOOa2Zb4LQ2yZi3AmN7ipc3bMtCS19tAoxo9uTiIQD
6sDYn/xhnbgOxiunVqiq/islGEaOPtorvt1tx5WF6+p22Q98KRwjDKA+6y+WuEXWkuCdJKi522pQ
8zzmoikkzBfk+T3SQT1TgoEBCVDYA/m18q+kYAhbbUX0qVvIrP+cQnFt/Nd/yG9HTo1e0iN8pk4k
CwYeU+LsIXIFGy95t/nHLklrVuClb9eJqidlNedDgK2WRQflONDr29rPTS1BoH/YN/Q4cwiY/6fJ
sAEE4CxvsnvJjEi6ofAxK95eO4SKlMm1DEf377KFKOC+IueWC/SKhSZgCkl1FEaUA6Qeyi3/puq8
XmpWhizdLysC3rSeqegBfCB0jEtWVNKO+M//DXAhneSeLuwjDnMoETk53yvvaiGEuLCEejF+rB0L
yJXtSOzlX4ulnVgB9KJdU+kBSrKDw7LN83W0yZpniYOGLxdh+Q+S22AeqUeTW192n+MvfI58Vl6E
JJ6BpWUasvDmAn+6sZnvRamfavDe7nxNs64Oncn0KJf0EO7zdH40N3Zl/Dnhk76zZnc3AN8UWpTt
4WX7r4dhuOxLgyH98k1msmvFsC6peqpzTtF7KeHeisbRdW56coDAJimop1NEPRWL/ZShyV9S3oiP
0T6OGTFrU+fzAHHcsZGFfWjVKqj3MSMDbaI0JrDUjxKAER6T+h2Sy7HX0eSswXkMif7aDTNX9bSc
8tDmqnC9XWs6AozgpUptz/ZGIQ3+MdieT+OoZ6xovTwK6qhNgBRYJWHAVT2DdKh5Dzs7c0ai+8so
QWvsnhP1OEtL3y3ncUq4uXgTAzq/AEcemBSXUgbEHCW98h+ffNusOZl0AaIYvDCetW5JFEz2CQws
79K8w/JYD0ziRp9zyGXrWoekt+rGpdi9x2rdhmr3MXKJGd/3Wqb0l+o8jJsgB2cPshA00FqbgL3v
+KSoSgo5YykTpX6dCvUN2kiN81jSyeKewMJji47W/c4c+eMn2JLHHxr3tWX3XupdqjOc1GR3FdRQ
attwPZsVPaQ5SMF3UHrQBkLxIpsLSaR2EJvMScsII30b28x5l33J5K12VH5NnhUcSpLAEEcIyaWf
xgzKHkL3yFif1uw8rMksz1LwZroCqWpIDL49lcdeEgizr5BITHLboTLnsGX70XKi+1SpaARB5hRB
HNGJzPtbtR8p7/eHJHoOVwFBVnUG9SRv8MrsWaepi0v6NvTFMP6uoH5tz8ePBnPeD//IPhB+zXCl
cNwIEDFaUD/UnlUR/ehfPcBUvK/vo42jvBGj5WNZAUHaG7+ewIELnwDEAZbA8nNvNTu7XWK9AxFF
5KMphRgz/JAzL9p3RJsoLp7F6we0IBQjSkr8YLabb2vgpVhuFTYZd7JTlq+p1aoDBtoxU4HuXQXB
rHCdFlHxCTazObNseff43n9KUlNkQgk4gWWwFW+kZHAJCP7TWIS9ushsINDkOY1DLBQSdlOotVOY
OZKDqBJL04xvEMChaaxV+LdFM3Fx/Qo4EEntE8jT3FqmI/Bqffn4l9/UOXVz5r8SZtaJQiR+nhhI
lUXmwN02EOU8VOez7RA73Y6GDG6ZdN7jcuyoFLLufWPy3kjpU/CPrfGkrBH71fUYMLsQ/RLEeq5R
QBr1bhkdiRDlp7awvlEds4/g3qCzhvOqBw8ATMfg/796I68iOfK+s3ysBt6grbmAO8XiXXSvbt25
DdrBa5mtkmzJJRXhZlHZH4Yf+AtXVWDhs9MTaXCGXmn5NNhlQcCJm4ACuWoWG8T0pkG2hZlIcLtX
PxD/kaLTbCZYJRK22iQIc6S6J42cdkUlb0WlIxsxbfWjjCTt+k45k2Ndnwg+xyGqyRbTEYAm3zFr
0MHKsI9L+UmweXuXADedsKLQ7J3Gm+krVAEXkFErNsH2tmXXbTPDyjpUCtA5W3TX8JH6x8O+4mON
RpUJhWRpo9sqMQW0XeBB9+WxgyJB6ObQA5vGTW2S3+asNn1TI670TcoDiG0C9f0k3a9JZ1dbzrKp
Q/b3lXJG55yee51aReasw8llN6zpayqflOAmIKBhKavbttPtaFcIdKLxHhHoEvA2Q46smhj1Dspj
QImQASEVh+AaMwsjTpkGu5G3BYFMBTDkvmvznvBHIlSJZa4svX1rWg0PgRoqwcfvy6nIkIJ3QGwx
x4Vfx39Ev4yT8kmtsBwgTPFg2Svx2yqaHH9wEa3Z4/G2XA9y980RYhwdPJDUfpC3KnHHKmRymFQt
yM/yF14luqLhur6hHwUtJYTDkYdZRT6bb4/rJH4hxC+zrPdM6xHK7IH/N1TUHoc8VBi4T9Rrqhpk
aH9xerNjoj3bevHRSwz8vLmVpgFId8lopRTP/Cq0Cy+4wnf31r6svhTvdofxCQpKTKmM8pfcAqtP
l9XKEWbTRQEtYxWQZFMpCuX7HoLMyImPtFHKoht1+o6eed3L5A4PYuf41k6sndaFDr99W4R1qe2k
qqfSFs2ced9K7s/XypDRdvec4wn1xM6TjkCvdOy/dBvFK5kuwogeIbW8zrHLLiHiHKr3cbXGLNee
QK+soPcdPpC4+FPcYTCI26dTIvoCG4fbJDO8CkBsaXOhRe8iv+nkVgYvoEhWG2kyn1Fk5oYHWXSP
0gIzDtQHXSdueOiYmF/vFfyJsJHe1l1ZEp/hj18I5Ia4orIujc9vGmMNWNVVxvQuYuW3FuOtBtux
8qhD6c9Tzz8G+QTFe9s0K5Qth714GNU4T4TDJsTJ7giM4CR+x1vM+dHoYVMjYTdmZQaIUvO3aBpr
T4Jd7NGr0lIyh3Isr+djDmNWpK9/VcvBS+8ks8Xpj+DAr8xgWNSaC3Ape4dSeetPcGAgRkuBO6Hl
O2IRlAbJEm8PGPwgdNd2OWmSHkXF5i/pWxArzucxGA/pnpzxB8y1Mnvwa7/wM6DOqQM+9zZY9AEe
HRes/bUS2FoUPZ72U6wEYK5i1hFfe11zFAUzPlxJQPhnB/0ztLohmC8psam8J0WbuHHDhpq8ZqX/
c91Ib22dLAJmTvI3bwD7rAtzrRxy3s05JYgkogrV5b6p41uUw1dKv3Vb5v7FIc8EtcDbkbUag8Xl
wvbqPFLLKLthvwWtBtguRzvkGZ6j8qnKMZ5lOXeC8yiysOnkEcG1VfPdrtj4DBN65W/OjpONTRa0
69zcb0xdbPvHIyIkbvG97idh44zl6+Wtmj2SA2OUC3nlmwmhuDIGXMnyrgvd+BgHh3E6F4S905is
DK1Z4KRMWrTmtAjOooHTtDjjNCyd1ghHdBiKjl6zmJ8QhrrWb8H2WlC/x7WpYcWMFUfGhhziLntw
kAAJipV3Y2lxwdPXPAZXU9XBI372A7B9zY7DA7MJg5zTSpaC75ZEffnUCvy8dK8WeJ+RpeFKaKjz
Gno85hzRxTnxHPvJNaCmGx7ftb4ZigFpv6yQ/WSZqMmDoEDfHn0KeP51ji0n5KJk4CkAXF9aJalI
A/u3Nq+AxHnSSuyCHcne6PS8uwFAY+g7j0WdaVSBCx1aPVrsErOEi7SJMGV26B4Ac1MRCOn8CEuD
/SUY3LrtiqtIFD4whO50WoihKcDfsAcRUiU4EJE4//KeoSp4qZn7Fqz++IokSvEhbqdXQWbUwZN9
6DWgLwHUj5zRexFl42Zsbgo3joTGsM8nT8UijNa1VnVKyVX4KlPEtSIGy63nvvCYAiFYpqpEubR9
sG43/bl12ahEgM6ZTP3ygc0FIGtGAunFnyE472sH26hUPoROL6/p3IooD26vFMCqgi/0SP+j5CyP
R90iLEa3H0h4nRleDERNHlT+Fgs6Z61JQQXG63rJwvCjZNYoFDvp8t936ftQUx7/6BWpMW/S8rG2
JbRfL5FhkH9iJxKsHgaZyLRAEvdWwFAOD0VBiYxrarDvD+O7hy5ZpKY2JoJzbnuZ0C85zvlshMCM
9AlhXQJZvk3lt0OxopM0aOy6ZVxpdt83KUJIVjWllxlMu+/VehWynkdb+KmrXuDCM52fXn8cMyqk
lIQxygyzM5Ta77UeahfZ0tH98fT7SuBhAixpox/0+uZtYeeQQ0pNiaYukyNEh2nG9nVfR6+9TSbY
hTbIptphlkatov0cw3bEolI9Nza+2PUNMXGg6pv7nHB4lP09xjK1PlFDkHul0X1pR9L2PxSfaS+m
jkbDjsA9nP6+dMMrFmVnmkdXgwM6maF5/7t2atSbku9wnnMEfrekjuc8DWq1GsQimWCRV/G3VybO
besuQJjHMUfOnR516xi+77i4za0Ho8UZ8B4PO2H1r1b8BboUJ2xcUJ3Ax9MZfrt3Yn3eLy6eIAGO
BMicaBg2pEqRYX1grnSFM5z6oJyf4ybrdraMWTLt/1rTBCY2fZ4V7j73VVSIWX58ZYtmiAxzt8U5
kTUqgqgr31DcDHBdmBdM3BNMqM1suIeFmJPr5jpozE4vuRiHvbVL6WXVLzpws2pbeGZ2xP9OshMe
5GRWBrpr4wcVdv83dYO2M6n5O1jcHo1nkD27aGd/2KKdhFjKf/niWK4Kl4zusIXLy5C+T6lf+3CQ
l23eB5c1nUSpa2A9kZ6i/sayLVocG4FojfRXEgvhF3UhFjSZiTUzEh7f1fQSebyzQYTBCg553JeC
fVTX35y/bsq3HlVhmcYtewQj36HA6V7NovbF4P+e+jsu+jyNIHxyfhCbya2Re2FHHrZBJUWl+2He
eyrxbhf7/qVQLN7kDIrc/INQyd3dYPffwOcXy/+NEGTNBTA7KbFCD15EtsW901cxqxO4fTcnmHc8
Xg2s6aRDUksM9eK1EMIH/DHFcDC0CAM89qHDbewEdSnaRu1StnVXTkncpAsjMmfjLhQbmxzCLwMk
XCnRISL3GzY6zUAbXfZMeDREurEl7ycxPCelUDh5gjInC7uAGo10kMEbFwGERdSjcfNjOCXefDao
vfOSeRSHj4zPt5pJBq+bkf6eQXWLVI5KBm1vXPSLS3bj6lpIc95dvCvLwCfIzsroeHzDnzgh/q3m
k4GLcADAlxabqeWuaHNFrIxtXfyztOSCK73B0ysEnzaK/UmkWIgOFJ2eZZ9lLV/INQICN6bGuu6n
qmePU6vlazV2jTq02p4YDZkEgiPYWa1C/7h1dlosulYEDXyd+wdBtT5Pk8kChuQU9+2vlnoX9Esr
O/TgJZ6s3Th27tQeiYNdOq2SPF4Hnol/XhDzaMcUA6/H08hynZRZFV1uDgmefmDnAmDckDoJtYFS
gTkuIE+O8tc17ApKWn+0IY60vjkLhtIYFVZqdOfmUkFV4iV/sWPg17b1J72zUeBJCcDg79ulkPRB
tCB6GBtvqNN1M/KwJ+L8QKGhvM8OFjKzqnZoj9LLkD8iRYEiZnLsu8/BXcxrW5ukNEeLAvFZ5qX0
ua9vab+8Dfzup6BX5yFb2IRmVReLYFoLgWGhqZxvRa6TnDUMYlE1otbI0OllmQow3pSCr5Olsa9l
OooOym+S7gm1vhyq/6+O5VSkj5ExMIJtwW26twF487rUbaMVYjPb2S9LgoVGOlvnh4AT+MdXvkVC
HqZDV8rR8IIWc3gMLJQHaGjrBJfhUzoQJU0welIRaBCY+q7bRBy+oVs76+hukDplZ0kDg+I/qz1j
KOYwa8D53Istn7TlCEXiwjSrjOlUxELOYWpKxCWQDrowLs/9X1nlWvsOorJJDc98q0zzUevoVRTq
Xb/s1Rkm22j/I5FGcxCT89b8dMAKcD1nL2XSfXkhs2HyNhOzEg3FRfE2q0uP/cNvmvnnmm7BuOSu
5xSLR/ZAYNNMVbaZZbAw3idAW8bn7xF6UqyPLzRwKyP1TcirFyUlDvDnhC9AEasfyIVoziUOOmbO
8PyCnU1CVwxTiHrlwQQbac8/pemFooR/fPtAHv/m7xIx0X+cI7nOM20ZAnZ/F+tJbrcT30pJkfHN
0TIScjOwTww67rfibcFYx6c8+muB/9UBaWMklhXHI0MJN7XY1f6hkxS4umHlBtlgAjsvO5BqiXaJ
M0mOSDYasQFWixpAV7fKiwuK9mGhUpNJIsQlqjQ3fdijaVnpJjmCKnF6F82ax5ao7RyAQK3Xjzcq
JJ6Mx3/TXdEsOW8ThR8GbaONGJVfvA+WNuGDSTzCWVLcm1k7/lTlVrJd5nTTVnBEIVvSvMRmgp8I
J5b9jJbyvl/Qo9bPiHydK3gOSJXS5E2Flfwruo7PNh4p5JCPBchM/AtKnEVx6Q8M8zv0gk7g65QC
XpCb4NI4LLWNyGM+NOQO4efFe87vo/Ed2tg0lKWOKUOA8QQyapRH17ANQmahJ66uYwHsXIN3jfga
eYyK8vM+/6iGpdACdPawkvGehVUv8LUv8tyvI+MW4F/lfW4SnbghE85+q2HJnST7CnemGaSukwVJ
ZcQNjY4RMq4/q3nLN8rG8lHMPEyJ/ooGaHa8MS/+C0w5bi9hlF0u0fkPZ6Ge+7Lq3dCapaSmdpZY
7/oQs6EprhMhfxXFx0EnEMqVir6x+lT9opHep26orjTkPxS4VN836kchBIYBFBCmsVw1UhTC2sT6
7A+IFk1QMsv9YfWcGnoKDyFgcvK+Ifidrdpp9lbAlgry/dm7lTeZer0rzvcIRxWSkv+LrObix6VM
1NHm5Juprg5K0OdmpT7c2+KeK19d7jR57KBf8QeL+emH6gLE4GHaD8OE4tOHgOedt8EuFmt9d2v/
Bslet/VyAa3GHtXQYfDW5Nht4wi0ThlfF/noWbEPYJsL3YBgZ35c74MYPLusaefCOuvYXfGFUsL+
cqns4pnnCIPLEX/4E557EGWfVEqNA3bMAjoPYVxor7bZFyxBB6T3UJ5KyeYWpa9NrQMhGIC+U8+S
OcsNzG4PiOO+swVMO25QS1F5SBK8aH0U3FmR3mnMbmazvmm4RQqtukdY6xKYAfnt1fB84LbXyLpq
GdW85qiKjrXX0q/r3V9RcgU4VvkxDr52dCenqwZZf77Y3fkjUhSFx+21/aqs8AW8MbXAOvW4DXpg
BIQD1Ly7u8WPsKn/HxheFFSLithq+ms1FVOfj09tb4ns+fkQDrheKYSJA/YwhRF3c1BxsYoVn/qp
PFWJiH5xKQHluadtfMccnwgvsa6QMNFUKf/qdgfgGI/vHs3iP+RjK1Q1XAN65LDrSrnbeYOyLc6/
E5QtKV8bd4f12Ibkm+gkh4U5oltUaA2jkiXP8+FyM0nMX0ixD/EcX+YwXkaKGwhBPK7e2hJo7hUU
2Y2+VrrNn2txd0p2WI2feObjJy/TR6+Fchd511JDB8wV9VrLjvauZYURdF1Jaent5BBGXyUX9tow
g8ebqK8pCz4SVDTpsIc80cWgglE9D1jUaDBXQA9YOZvhY+HorIMRXWi81KRdXHTHFhqyCnR9H9RX
yxpr9kzNTrH4+nREw9ZmCrvoG7k+Ne/jtVANhiTk0h1tdMDckbDGgEcPsUamWSWNeKR8n3Y8CXhU
/jCok8ubnnmjIuY2ssNF9eMmSoEyK/fw5blSU4U0KMY5+Vb0mtwGs2m1WP/RKA6JlXJsBZYLMroG
gMKrKsDYU+VnhlROmXA7P9JympuRdByfOtKzFFkGKZ+DucYKpAR0mq2m87zgPJRnzI+wn//0gYiz
7pl9ku6w0tIe7nVO7RPm5g+pGFeSaXmjFrrgqRRfknjGI6WDPNNwLkUxcm+rAOLyh654X+j2Qm3/
BSzP+GkrzL+I7yBwkv1JMtxupQSDYG5+nXLiSkSuaFkjgnfJUzn67eq/bXQzcfpeYq/0vuV0h5yX
Jy2x7y6+8cHF8d5C8ZuWaaQLok35PrUXmBw1qC/wZzzDPvtwNGZZjNWK/xQ0vTSbQr93kyE7dffy
2bKGUcBKsU0Nz4phRS+U8ycQwAy/syvHHgGuKHrHBKW+Hzn90xljxXv8eu1NJRymPty1m90yNpjS
uvhniY0hkkfnfi6dIukxsv4dvzq8xrQpjKnrcR/itcKX/BFOb8ixZLHqJzmKZ1jkS90UCaLJknzP
TqDjMWI4nmNWGPcJkapa1nrYc/kw5jYLgylfLf/UMpYD9uUnout9vRfwmgpR75AVLn6Z3oGG2l8z
LX4oBKvZl0ql1dd2I2OA4xtpiuiXVnfmkpMTQzBKTP6uWn3IwFGfb+XjsCJbn8kTm5Ve24XfniBx
9YP46udwd1kPz0sg0dqILey+aNjmPIJm/HXCjcuBZI9W6YRLySQiEe494tBeLZzgnxgCKVNEpajg
XbfRUTbnc4FV7jzH2ZMOlBrdc18I6g+vVbKYCNF6EslyX2rtEjJ+kNno3dgA3fkt+MiBdqHmHLuj
wvMz5rbDmXNkeQB37zjdWUxp0+0KXy1HEwhi640nDV8ClUD/mi7cu0UKLVJGIa/B4gG0Dt44TXWD
t0q4h5nfCB+FdNwYltxq3xJjpJpWgvbWUOZbFY1IXLhsAWMfZr5isttxzvIsC+A5j5FVUJ4FU6ja
PQoj/grejIHNCPAucva82B6BmVwPmgch21rP7BqiDjQf53YLSArBoNxXAwdYKp6OZvfuvZAdmkLO
dzrSeAgPMce/L40CZA0yPgkXDxdaDiuPhpBYsIKLxX51f7tZHsS2VPmKIWTUKQ9qUaEYQ43p8S/q
+DZt7Gxy/K5mTVrFcuvXzGotLGrTX+ph4Y+SQ5Fh/GYUB2Sk4+ZSURk/QZm8oC7Sr5TdkOKYix5v
MjbnNG3ptSCPL07XfFWfVs5yLAC8QrdnifMCnix9mXq2xJJg9i7e2zSibNBIItSbkQxPvSIteee2
BM613E1Vi3YDSuAN2Bh8pWWK/rEZsb+uDubqBKeFD7JIAMNbfYqudQQONexY2lEJ2t3aKe2qzoqp
e09EQ0HwNaUdr0BA4il5/ZjwNEnCiSXqxbsShmXvZcuAG5XNzea9Vh0uaEkcGMhKtO3VOhTxZFcd
zgHU30CAhcwtc/2ThlXG2lC1DI10vb5mwGkGnj6y762ULBE8Swrx613MaSMPGbLjGefrj+AOnAu/
L+0kE/N7QpsEfmbBmG82jKjhsf+GP5aWguTQH7hO6QlPQ+7GB/suQc3jFmEA+ksSwPdxNKOJb9KH
wuYIQ6sambBPspAMGprErzF2I0rOQOcot21H+XvzhSpS3p5YCS6YR61n9s4FHKHHF8z/IUtUE4FQ
wdk9tB5XvUREgEsLv25GvUp/IQPELHiXuaqMo5YDN4BQbLXeuV/ePW4hsbSuoHV2ekfjYbV86KUp
NSKLcg4mQnOyikbQ4IKOSV5LF8nDJgBj1BoQP+W38ezOKO74RIJmcdbytigxUceHjUXntPLcExML
BJWHAuhm7ThCApzo4KjS0x6/l1JkviEd83lUlz+T2BXrvzihp/dXsn+KBH1fM/AVNO5XUh+Ibg7D
PuFz/9GTOYrYtfWArBRhwS3acWHiDm0g5PXWb7AzZgOmSkbDoD4HvGJpwWiqjAwzO7Yn+rqnWDLv
NThH36Vi5rs0vrRrp/0BExGhSkQFrQnGUAE81nnI59bKL/dTmlHodkHzdeF0mADgSRWFRpqVHegJ
amnqIzwu2Wa22MMeqhWqU4UVV2bAe+CvyTjDlXXxjpN6+Z4k5gqUwKImWi33YLTJGWIoyvnlL/Kz
jvXAN+KUMk6DmAhvYJOsxW+7s2GsCDvTVp2yFEZ5bTFQiL9KoH4VJGRDFKT/iOnlNWrPYWnZpP23
HrFXpJeFLZG6S/XnwJ2JI6pO5XnbeVrLVEv3VAeUYh/IZVGpSCm9ZIlHAiroj+/KnObKJtkEkCdw
mF8R+QqhUQVFDcDn4bDW5HFSJ2/O1WIu8tS/4kx8FmjuJ29CL4Zo3AFJn3uQi9E1lqSW5O2AbfAf
BfPVHVeERncAoQekW2e7XiFAZfraRjpEV6PebUbMAusPjiR/MnhH+5SnZYMuhkfwSz2ogPouTacg
ttzTdjfw3CzZTSAg26uc4ZyPRwm3HzB+f5/2z+5t1vPFReWQdRPLE84vaO5Q5/Tyg9S/PdrF3U55
adrnTh+CsjY8MVC35Tau0jsZ4QuKuNJGEd68u9RkyuOB3P+/3dL9FlgauudR4Fxm8+g0C5K0EvAi
KNQ4cM/ESJKqLDyw95s3ahWuxWxJRgp4aQ+wbbPHK3Z0VAjuyZygKKEmeyHEEJ8J3Oz33sGaXlQU
qkfo2BP+lkCXREelbJmhtrZeF1c5IuXMcRY02803pogZK1mh/HkwDDlpMDPrw8HsJO/ddKxskw6b
8GgqDCVVWDCJQ4X2Vy5Po7oWQPupilR19rCQkYnHX4CQkMZ66zEMN9y/F8GuJUnobFm7VaZKWbWv
krRSRZhriBDPv36HOeg8IRdEzlWk86amKwF1H7klL4q0GgS0U0yZz0tUsewtUK5fTKPKGyhJn+LR
hnnhRwS/pw4JnDJW81p0gDY/WLyXsJWVz23CmfLcMxZH6fXQfGFwcNL1ll35zS7P2SDEGQ7/Bpbp
RnZFpq+vnCxqtGmlQaEHpvgCQDfkHsRex5SnWK0ViLgjktAQZbCpl3y6m3hIZ+Lvufem43vWnZWI
6f3BPOi9h75PiLXov0VRapov3Hdm9amp2fUwFEEw15kA/pweLrppMgUCfIRHZVcu/OYKZ7GAc4L6
wvL9j4/1wpB+UnxMPs2V3scmG4k+6O6zWNx4V/a8hL6DDp55Jzg66z6Vql3pK6laUhv0Zu+kg6AI
7QPJnxqEMifmHyz/873DLDhtYihJS4uHEjDr5q479ePSRzVemlMK7tCuDdE4j9IgHjQQAJ0lvm8B
qqjrSPm1yZCOI1g3TSWpTWCTudjcRyR/Upssr0CmFCsNrYzApoKcv5m5dvFET/K2raH8EbiX5DXi
h8XalVYT8n7dMg/++G5tZKfhq9u3yyRMB87qClkyoJS3gHNTcsECA8rupB3AjeJHopdDcbuXu5X/
Ml7CLxhnUq3ePGLk86UGI3FfcRgeTh8qJ20SPeefcLJHd0H/4Zo9ubzwjG6BKTB2LrEB4tUSPrKM
hGMg8BuiTzVtF7/3WgvdHtz+Na9bkrb+c5Dx8GL9tGrrrfS972R1n8f0ddlvmqI1VGImipnFQzww
GrGIOZ12RljFUxWZphwaJjhpz8GxeMGsKrJZjcWPaexvtLT4DUKfrN+niHgGEvwyptLbQ6etXtVo
x9/Mlrvb6Za85CL3dtC5ArBAORKNTG4YGCyE+Bffk4A6jzOmauYlOC3TvDeHOvF+y0EJ+tW5H2U+
V0ITkY+p0QyQ6NYT2m2NF8hn+84hzW6neWqFur9AmhfmMzqlFvjA6TRnGVKsclE9/pPMXwSCw3hJ
sGTYHiAJ1rUKnjQlta7m/A3G+asydL7A4It4R4UkoipJiV8rzeUr8JTbJs/PUzM7XZ+yXVFoIrpP
cHRYNgO3294uDQs9F376ORNAJtivpBYlaZAIlkwnd5vYP3tqxFm24jWjjdBuLQqHXemBOB7SAejP
a2G6p6I9jYu0kmnswiZxRB9tsnfeTGwHZoTPJtA0yd0iFqKfrSnMH5SqUyraEhknRh3khoDyK1BP
UtWbvdpxx1BA/VoWmS7RkZv0X1c/n2tGExmW+ERrXWEx2EIxJy/EU9VOn/1VGx2NQU1paP1A92us
O7ivfPnd3YDX3kjZoiyW6RiTIjSDVLdzywcPOVFFQc0GPi29m/a1zrgNpz92L9CTKwKUZTIvD2v0
y6mpigDysy1dnGriOaWTH7MCCBi9Cfk57CRUzQnnZU2FDvRYEq3OH23d6FF2av6gmsitsP433T5W
C1TklAWJbTP5MrPsbDhVbBnsNrrZuOuDBIXF5bp4eQxVo1Vt6ZnM/I06nfsoSbNvQ9XeY10bIV1U
UwzRXB5Lu0o/B/4vDjNxHLULgGDq2rPl+POztCbw3HWbFTPXxotE+gSSJeDWePVWrXYAWqezps08
BDHBbpDogDtQjFtYxS7SHca6TC7r9qrTfhrlddvZ+P7+4bf+mfo01iEB5DbKhcoDasClezSY/q0b
neTnYE/yvN/PV7OVnkIjRBr56pD6sSaYxFxGkLOWNFZEOtWWN2a9o2g2ggLeCvmX82x3jrv8c5RI
Y15SDhrynCQof3JXHo9NvUJxONUK/czIWZxgAd8S8uetnpR+D4OK3WeZMfRzJsG7dKu26J2qea93
LCyLewq5XwRTg0ljKNvQalQE71fk8Qywon1Y6mnoRlBjdl04uquS3MkECXew+RnCgIQfrPxbtZSE
Soih/CIFji4y0H58btPrR4z1yirm1CFPVI/5S3jD5CYNq+vcvBFoHBWm2GsR3tFag0l4SprIKKXN
aDIQyDssQlvrlb2TbjdlWrAxNM0Hvw3Y0Utjt0b80rxRtUrV7osIlewoLb4w5cIOVhbyU/hqSs6f
8YjTQqPwBphh+46nqQjKPE9e5mnK2nBGJDelJrUzpb/1iN8XC+937MgSjbhW0Bh6uY2DCf5/yx6T
Dn7nBJr49xg0KTwT7MeJUtmMth259G9liGod+KRRZztt3jY2A1JGkafAqNHUKIWdj2Z+obzdQT/Z
OsTFvW7eELMFLANNbhKQmVvCzVjrlADQvt5fAWHICw8NjKeKP73AkQtxVR5hvx58kzVPdMW9DMvH
vildKswFw/7hcMsDvpGrt9DlgEB9BGYyw9BOdLjTZSD7WAU/2XfV2Q8WfTKJ2Nrklk9Sz2IRcZyY
VOSe2yBWUCqyBbBjyvqzqhfSIUunZIQabE1sNYc8wmIfXEjO91M6AtNmTtu+ipYhw61YbdN9AVHw
KwAglW+3xoYqWcBC/VwR9fY/MVYuU70I73khrZJ37n5qAiIGxqGV2EJtJXGfZCCBVLLumWIOieFH
O34D3HThM9aBPIChCA/BcKJ9be7otbFrCrIiRkgBZx8zwl3KgF7irb4GqL81StWceAUrlxncJSbn
KFvIByvO21Ux8Miks9Xn85HWBOHw3/tAHoH2AtujYvpUSm4LtfqYOf1rAk4khaTmz5IV9IhKX4VU
KugZbpusqD8Fkh3X8iv00sHAMMw5g7MklwZVgiWFaU8aMkUjnVJE9yx6FNMpFqn8tEoBl/zHYT7e
5NH+gQj2WUreg1AZBE2Lj6SezPpSsYF/1PBExJBPl53CMPpcx9f50lkJ0SEyadgxUgeLXSZe4LWP
FmmPK8YDivqXVnT1NgoDgBfR9Qq8nQCEz4M16hSxVixBNzYOyK2Re3Kn7c4LPfttu5WB32ifiQD2
u5MN6r5aHIhb0N0BSkbtlt2nu7wCAsfiH+kfGV/7ax0nLAeJcQUEEzuXKxG6cSX/8XlFY3v1h2DV
gQNzEqyqPJG2wqOC0ykhXr76lrb/d7Bv3zVW3LHKfyk0psKazgb1cglZCW7eg7990OpEnOIVBGWI
vHYbVDc+9wgX9uSvDnRMvdXFssdJ5qgpHoTK7W9cly1DE3YLDYtJBy+q639qHUhMa3God1tl5XTD
D3xkarKudCX15mhCmimgOqe43kWP1obA5fLEJrf9TaxjMFdDgPLkK2nDqwu9nmh606H8kAIZYpo5
oYDwNm0Tkket6yWyMdIhxNKyeITH8yl9BHIR0jq+UWEKrNXp0/mQE0lAov/qG/eUTQfdD0/bUqM9
THiFPj1cm57nYojgKl1Jz+UDCpgIPZ2bHdrqrZc++EIqPhg265VWjaX4OUSW5GdsKLvby0tCQRiM
L6rz/CLoJCEP2zSLPdzn7nxDFNz0oazkOtIhV9uDclE7JQgW9tvkDL2MMKRNcgKk+b0b7Tfq1zF3
8Ah//RVqVVNX+5iuwaPfl/Ud9UDNSFYfOCuXqVmMLT6RhBePkeneEpfQpwykf+khAkPKZfDAuiHF
vRA6b8hIwvnbFAW20/ANpRnfatr5Hl2yQ6djZ2FEvpmd7bT58gZ8u20+II/rlJL5fQXLUqwgUl1a
7VJ4IV6hPP0s3FWg0wsWTcRWwoyavrr+Tl+DyuYUbOKQN3vRO30L/hbPqeABv6L9Eq32RWSZU+Vi
a2xaVK2ESEGs5dkrbLRDe5pRVsayZO/ZDmQw88MlsC+0DIDvhFusyE90ymXw7ZuY0gwMLOY2Om4r
ALhTMuR+PnrVunnQYDHIuRta1my/JcsQgzdBUEUYSDTpkefmTBEnX835XUw/7KoAvrtC4DPQGG3C
12ZL2TRxDS45Atm++U7cJX1RTxGQYqwDhkPAaQir1rHsl2/IuFgJvFl3+/oq6QH4gEui1hPn/pSc
S0+8CcvCR7ZpM7Pqpu2/k9SPdrIiMAgluJXuqxBFySf/Lg7QninnlmL6mx2YiqWZAhR83n8QnTUg
iUFRd6/rtsY88i9OfJ6SkikjEz8zc07azHwXE2J9u5/m6j3CkK0XzxtaXqGkabfVF+GxO70snRQ9
L7BlG5PvilBPikqyviAJsGu1Lw/JoHGLrHxY87Zwdgud47iYNQNReL99XNs63NCjRbk7GQehegRc
LJqVLVGc8vLczNjR+GB3In4jbcWXZUdOFXbppHShtoGyRfCp2J+/n47tzNezniSYRCyw0rDF/sk7
a0Mt9CdNTe4xsAPsn4fuQa1LZYZ0BtK7vUqI76olG90gi9UFPUBrHsAle8NreFzpTnVcWRK2a4eq
KkByBkra6HFL6jWF4vAaIuppVb5ztlwN71Ux/7jgj7bH1w5z/Chgo5OMkDc9Kc1c691HjFxOCJf9
OGAZ2LznSTs3OA+tqiYhZCjasz0PSc8vM/oYTa1/6SiNKsjT6p4qA4FVk5hybX495ym8gWLYPGbb
q0cGh5TyY9i86vVrIBECi/aHitsTxlrJ+yXCm2Gb+y9+enkALRp4Ju3jpsAMoTyLXtyw9gJLinWs
F2nhecXajcbX381CKHH1yxcwa6cVP5xHT3dlhSAAzfT4yj+3L9iEmS2mIgsDCAmciBXehsP5vGNd
r/HvhdZQgFuSfJiwWH8sTIxkAJRCc1OKVo6sZ5fOuwJiuxp3+nT3prNYEOnE5OogG/J5yOFg6W1k
+6LnWjGHWaRzIZvbJpk0upXIRrwyK1XE7Yv4mmZWRmpX+2c6ZCMK0VkXTIFvalK2iS7gkKKxtNZD
hzrpxbXsgQvmFDPdulaZ9ysBWJnsQgXJ4qqGH/347GkM3IXp4zZhBEFtUbIx42zqd8acqa7cRCsU
SazcSF8cWGhYpcXwhtAAj2ijK2i0pvI1xo69s2CKJ9Cg8AeiBAGDdOqJT9JkmqyUH5SscDpXsahh
/b0pQWYvPBM3QYVaos25D9MADsNCVMF5uhHgH1W8WZ7/oAp/Is/9COCogRJSdueVZsK9zCHuEBpU
EIgkjfYW6esdIcKH5hAF7ONlHzMMJtmbV/fcoGW+CoXsgb2916LZeemCgziTviz5s8txLOuMXpt6
fMgKoslC1wNobYI0QPptGOFqv/3t93heOVPwfO35MY41+dqW3z+Wuug1vBHiKVAJ8IImRFCWP1Lq
z6AK38yAn1k0E5uZrThehtKj2wjKSCqPyGq8WpslvQ6u++xtl5dWQrj2Qx9EE89+tx1aq0PjVMhh
f89nZ0zLWoZifOOpEqRxScDWFKHpoPpA2Q+jNm+bNoWgL/rrWwJI6pFKcMMml2N1NLYNlU4sMMfO
fthJdA7bHkmHXK12lNetybWmjnQ5dMw1I8EmqdW7w5HVwzeu3vPrOn6SSn2gTf4mM5SeSoBP+C+L
0xgIm+6QsWSw3gtFEhDAC5blUpCsPIWxBt7dKpwdguVeUk4haw1UKhZGYcIOpRHzniGfEVntpRPu
LKrI50RR3GhXV7SdchgYaCstHBimP+Te+GYBJBR5O7JN76VIE0R7mFPBgSMWJoHARnbFjmI5AES1
lBh5GFaHCeSmsKvR4pa+0/pLWD9O+ylbSOrYQDOCw4e7PiNOQL23A4cauiwNu2dAJTbz4WGqNJER
3IAK+GORPwPcvPxvocZAnw5zacRzLyh1PwNh+tjKt2+DiTMpDer6UQ8CHrvdRtMziegSbBtyZFnQ
uoVekETEdEL5KGy+j0Xebcd8yzg71UoCt2bt3v36JHDUTIFOiG99Qkt4GzSrgrSeFml0wRc56rr3
8azTj03QIBNfre9QD/XgTLxYHNx1uvH47SS/dkNQuu3HiBu+a8WgcduBGfOEEXBMPgOfOc8fwsTT
1CvdvuuLFOCHoSfl9gEyfY9AouB33JxnhTlpYaNNRAMdMn+DfdwEnz1ORUZfQNVD68zCxe8CMEAD
26RlXrT8J/Ia7UfDYl/QxIAU/jt3ZoPa+RroSNR+5TGXR8qjdkKHmE7239QQsbxMdZ8geYjYAwZL
eAVo9CNQ2jY31qqOGeeD+xus/oVMT2+73LD84+XYHeWl92PER9f4qoz+kaVBU4SwouSi+XF0XAXU
F9tTLDXOJyKhidpmSIeMcsS7g4glOtnBB09BGl5bDYuuJIaF9VmKIoL3PpIrJahiFFTh+s64giMl
fDXTR52z6zDh6KbD0v/qMNczNqOkkheXPBbnMq9mABGRalzBfiyAFB2atw1JwfdCEfEjv4Q7dPAJ
l6OgPRyy97Yg05uKb9Ea474ky4BmxIaePQWEl7Y+16sr//Ko+/nyur0c04WJJ11YsXfVibgA7Cs8
kZ6jTQNUspuwzajpXbDhB1gR0JGj3lhgvfwQLNmXmUydPX7w5otshwTRjPiw6li2vpTznwnl2spx
2nbPeut2wrVbNcGB44kpCJK3naAycy+Drd/l/ICzDXFwR1bw7gK2RP7LWHk1+bsbVfijyotdwWpF
9a1kJwYtoqpxnq9++eCvVLhJkMgvt143O+FxlDr39rhliGEUIMrgYHu/kAQS4EsiBdB5SShKSSi8
svuU9IDhDHtmPUoy4vLUSFpk3vsZQkoXIrRRoqQO379C741mZczgNHkJ3IQQR1mEJNHZbFa711Up
wrB7TnyIFRkVshfMkL9GBqnYCuis6o8oQfhPlAqd+nOc2/0um54YH2VTxczrHtLH6RwUEzPOqpAt
8tQeg8mOyCLp5SwLCZUy5X+jo2/U+Tu8hphViESTcJD0NkWf965u8c6gxbtevh5XWwj6AE5yM/Da
FI7ja2lpjF2QTELcWP+sVHb2lz858W3MMyikE2gMLep0UpHujDpPj2X++DmZ8blBda2gTRlEDQWu
YY1TIBggtRN+thPckgv1N2BTTy1u/n8ZC53QCiK/gxY7RHBRVr2e/JHK/eqUrxj/pxCQWwQMD937
1XlsqvWpEoQFyOPB6ej2+nks0qLlXfUwsuIpUgFO8WqRUhTZ6r/Q/BzBeyIPai7SRIzkPc8IkppC
+lKV7VyTkvQuNsEd0IK5+atGSY1Vd3Jdw6YN4JWeRN28KG1w5sbjIz7Uhp+rGZHz9NK5pdEAvHgD
T5wcareVn2HNkr5kLd8pVdl0i17J+G4jCkguazGEwQN6j2Zyuz2/HO9BQF/zWNWGJBIlLkD8N40h
oZ1DdNloEnVsgSzO3PMJ5hxhztva6PQn9MYZm2Cz4nI4mtks80Pm/DqTD2Uio6t+LcBMnoUXexGx
rWcTGmVFk7ZSf1A/iR/o85huUudcR5514UTxNDwtHGzlWAvljzBvpzWk+UYg/6dNuFOGQHG/VCLU
KRsQtnyCCOUJWvuPpaXD1d8h+OiJtZBVafltTs1Pjz3V0If0abB580xTIynMkSzvstLiHmyIwpRN
xjYz9quSCuivQnq3fwSsOz3g95WVHS5d9nv0+04UAhJyWtBT/JG3kmPmhC8qQhuEzT8uEakL7tMh
tG2ZwJOfQI0EgLfbQKb7VlvPaA6E0eI7hLuShi0JbwxdfRFTnzLdWBZ0EnUQseCCWXF+9qTVkSNi
ZQpM8yxWKhDkNoc8yEg9QktqDcKdoc0+XFTZwsFX4WevIBpuZWkMbu6QYqbePO0gIH/YePqkvsBe
+m/BuUwM92RmeT4crmQXxaXDwQEZUbrxKseVs+ffqsGE2aLv8Xn8KmtO+ylDvh50EXprmbcH/eHF
LEqs2QrFHzKDIdhi380EVUbolifWb/wuU7m0DVWob9gr9BckhMRkavlKxspaO9j05EoK4HmhlOhA
Vrfrpk29cJt22Cddcs0nGf2D/+/gvFebf7SysEwDVgoSj294Ef9JnR9Ihpjq+hLaGMfq41LP5TWA
9/OtCAh1r/UqSTd7DANRdix2nUA1qSf1WhhP2AGztT8vCUy0MD9+CCnoJRc7y5H+5A8kUepTfqC8
tt0m9fLP1PR+pg2mSuyGuQxpRhRYZxOEfa+jDcF7o/QA3tfMtkmpGNa4m4XmygZuV7uS78yqnaCx
hUQBiiiYnnVOo7IORxY2NeLh4cZvJpyC+4gA6l0LeIDQ2ahp+Rs5OjHKPSgngja9KxMkIPpKBgA0
xcBD1iSvrgYcfH1KA0hRKjjQvdD19XnYA3mJl3EGnUpahFQWQdL9lnrAUehvzIdkZ7//uU7mAJUV
G0dZwMgYTSC8PdpRX2RmFIUL+YZTu70p2F9jMvx5vE1+vWzcyuesmDwexKBG3kO0F5w93tkI04k4
a0yScyWSnnyj0CosZymDij0QjCb6p61+dMa6EaX+OJCKipsaJglU7cwX7e93dnlQbgwZx+BXkc+M
YEMoC2JSmSwd10uqKh3p1cT5yuoLrkMZ0GBOX78ow2kV9MWY2xZPaAHr+bhQgw7hZNhG+Fm7dxL0
qNVxtA2T0BCoYVqti2HNNc1elHupz4R3zHR52KgDh6B88LvL6gYNdK3mfsku6UswMl3KQjRqsKKC
8CUqt+J2fYhwlbEsN8+gQT7QO0mGykCMGioNJESUvoMU0rLw7cLb+DtfGxy7LF7/C8RIm59a88pz
bY0kQwbHXHGASB44bASQYtxNP2/h3qprCHbKLxmzScZiaHGZ9nctsXi0FK0iwpXHreYr8BXeRIIR
TcYuu8SRqGBawntE5KoncwA78BB6IsxtUstoG85sn/eNgwgl40xjhS0Lo/MY/ELtoGFIfwIFlsMA
XaV20aVwcYjtjTmZdaS4SGTm4iVYjoaIUlFcSsfOqNB3M/1DLEj/bLfiavD9Sm81nkllkMlryx0Y
Ld8jtPSLnReu9unWHPbkXEfUTuqzoeE0mtbZI4rxV7j7DxlHcAcQ9xd6eR3rj7zOU3yc1/gkh1Yf
wowsfH3rkYf3WyVSXiEtZ9yBgvBpHHQ8SvPJe9y5AZsxwRufA12Cq+oBHtiPLoUSQeRtzF5bp4W2
QeFsS6+Awp1D42QBpmx9t/CRj7571Q8qtMX6BR93tTjWKo2hXxMax5mG5fRT9dbAITZmolZ3pVeu
dmXettb+1n4FNKaer2bHRrFuKdlfeVW96xweKj6nHxz6wrO24GmxtZdxVtTxKq4YjvrwepEBAzWH
mOHkyNbTsBhBCc4jF3oW7t4/tWPR3VRYLHgJavKNhwSK8ECgYhZG0wJtCDnR2bXVYqyxsXLARqZd
B4GP6gDQL9LvL4DPO9ajIQMv21HQarCy1uwN4DWvpLTqKg1o47fNnazYUSsaVm3d3CoW66zKMxza
0UMnWASB29iH/4CVOk748UkKp+R4ToY6KpAvzF1Xcmzdav/eMwNcgmOUAYsW5eyugj9G5uFwOOmW
0M+CdHAEcMUp94VuL8tay2KXHVNNZUwD0gygLF3bf/oy14sZ+G+ABKPp6ej3z+lGuYsQeN9hTPAC
LQKrkPaUKYcexoFtkBHKbYlK8FnSV8PG5go2YFpyClXVAUAGk8WtNiOQamgPEhtRytqRf7EnJNdx
6DEnvf+c4USXCPNo8CyD1KarHfMGJH7iUWogbMt1RHDVEfUJMM1xVWye86wJ19KW0gUGwXfQyNAa
Xxh7b6vmTGcXjhH2anQhOjeQXKpVTLMpuoiKNQ142xnNNvMiARd+AhFPrujdLxv/CPYq9RixEoDZ
5w1envtkB81Jl3AV8pLmEvD8mZPEk41/q7O2Q0IsK4ll6AohkGqCjPSwWf4660l/IGGQuwP/9eA/
XSA0DNy5+G4fyDIpw5pAdNyPq31aE+kYva7BHtvVLy58cClY/I4tWCf6G6ECYjenlBWtx5aliH8s
wG2tfHfzanztPYfgPyYSgxDfcDNLHkQ/qaZB+NmD+JKMZrZM5xFoOAOQznpl8uAsvK+Rky/WmsUm
hnAWyFkPMj0+TRPKAX4dWycsOZL69nscj82imO5kmP4NZTxxCmh43DmkY7XfWDH253IUuEoTETnH
JZMM1P2jjP2DZU2Hxz42Y5gJf8QhLu1CQG9SHAUUCWHIYNqlhzyt92TiiOLupnoUpS+SJycsq1pN
c/WIaFPHKQHHlYNJh9Hbi+s8jdL+0O/RaRyU8Wob8FEfyrpVsbdnCktxWXQJ9B0JahO9lAXK5+OP
IRp41Ie735kDasKSTeH82mOgsGM2xa/z317oeVSAw/bz/gqd30biNHD4phtRz2ePC2QwWoSniBs3
JSN0zCt43Fr/cpYRcanQwStHVRKTFfQjWyIk4iMB63WAGKyFHlU/cGyrcoikM4nEl+CnNtdVyFMw
VWoqauxX9lw7QJzkRkVEDKwqriw6YlR424suOb0PNZPBiEaOckbE6++7BK/qoDT4utTrDSRyrd+A
9syjl5pNrX8zdSlSN2jXJEfbcnxF9MDmkSlKZL6T02rVg45mGY+yf1Jy7K0VYfwWeRys+sZnm6AM
OSX1RtN8ul5Dfs0T1FPNBePC18cJAwGlP60sc8rcjyaBvnBfJyvMJcOzEYm9cZ6iLVjfR9fBetZ/
8VLSNCidNz36vj58zbdRuz1VKGg1iTkgTiLMxjdb4FQ8fs2ERY81yzHtYYJIAuHgXtRbKh1E+q5f
sBhzkVXL4XcDjz42n9CjuE+YPclJxvr24vZ+BE8t6JJj4pZbnULcosNhNhxZBRRv1cKBYdXDZv2Y
GLwMFP73boTeZ/5nkW6b+YrLRwe6Ld9hJsP9SCNdsOJK75oQZdRVhHR071yJQEZlm6dnJOntlNwP
peEPxIRYPjtUWqsN/IwVQGANqKVgvq5ubF8ng+1befEKnrbAptpxHKPIh594+5jQyRqWNgKdDBBl
Yz0Rcmugm0SFQdOBcCEh8lLz3Fr3G6xqsGgEDoFfighxT2cQyVbplXuVP2oeB8LdQ9gguGb80rMf
RkR9VtdElJX2PDBIZGLHVXiI8Sr960ev/ggVpdJVuVcvltCsjWUepzCBd3jtRg4ZN6azFrVeaSQj
QMJSOluvTHaq2dey8DBEXYyW4U+02rHzzKYrut9fdrf/Ef9gJYvhcmfR42S8KLsiCn4J9aleKStJ
5yyJw66N78D4dTdVREZSQdDsl1T7YXVCticE0uDDheFfNWRCN7y+qmLI59BEmhMPLhFu7+sYgzLs
dVtL8l71UzVeRT1VKWbVtsJFi6n+mDClArjznXneInIkdm2uo9Y/6cxMwRf+GmkNsvT3m0L3GDWX
LtaCl8ebmcW5kA/jO290kYz/zmssG/uLc8C26V46GHp3iB8u4cb6OYD3oPsox1oQcv7qMjFE2pOC
6KlywBXamhwIxfsw8Zz4buL7omWGmddxS09YD7kWKiG9tT6l6TD5Xqrv+pIBBWG2QtIY+qPACebc
04dJyXo3DRirL6Cze9aB8KquuYybCXhsCW0fY7/A6lrmCJIvrBWewXpHd60HwPI5XUJzaBOYVaxK
UzvMD2X9GhZ5uncSjA0HqPRXBJrllavsrGm5YSrxFxKZ1CSjs90j80uu+mPMYAmpSLTnrPVfOWrz
hmsTqUH+i0mSKehpXFubiZjxQtnKTu+Fq2hwyWfQ2OzLmJuLZ4E0i7/F/rdVqwrxCI34eI/F8tPg
KwaSldUHIC91STjSePqS8NG4mYeklRLUM1B13L7hGePIG6SrvC0SzcS2VroFdQr5lMhajJnpjNq5
pqHfIKBt3EQC6tCsXtglSfGK+Kn6MkB1o+EQRFoCk4UByYFQAFR1O2SVsiyX7cw5dwA3S8Z0zII6
Ru46BJg/yEidBEcDq7w+CcYOj5QsAeXIC1PIJiK1HL3mRUs2Pay1AgOgqONTSEdjrR0jIfy5SmL2
kQmI/zgFjXT4q8SIhuJJ8cNg+A8dFseCFjIpQ7m1fgE3BSlrPjpJ/N+PacCbd2z7sArpgYXsqCVO
xFO+q660UjdLoJk6gyLOU9Nn1zDNwSh6OsvcfIEAIvu+v0AVgsErRzAG4+6G5S56aZl653bX1LfM
hLliLo3zGMzK7Fj1bKD+iT4mzkIYsMRGkFIRx8NsZQmldPvcRoSLHVNMHOXNWVW6+KdjkK/LD+al
5zonl1i1azKX9jc2EjkD2SxR7fU64StA8F0bbB3Qk/lv2Bj16dQrdQT7d/Jnka3mvBR5U87ubsoj
vErKy5/rJ0wcxN5j888x4mQ+/7IdfTqxAzSOJ8QH4B3uW9b7BXUOSDebUqzm5/TQHPrxG2yVK3XR
+Alfp9FqEOWNnMlEUjsm7ZkVmNvElPRcPNmrGKzs3bBYEWhjS69pazQT4ajDX4eiIojSSE7KjpK0
cYIkzjQ2MT6fDT4ZGbRGrf5BDI3rLlghHzGnQOjwzDc1WkifWQjN0vJ1SR32uofyTFwMLt1INxPz
uOI32jL+xdNmBzNKF0uE4NoUnQPHYs3kNmIbMoccjf0xPga/rnNNzyIwmI53awINhrdTj0EwGsoA
Fx/cn3lNhzAhTbkkPPJeZMKKwi6MbUzuJ8lifBash9Q6zPP3M97RH36kQi3G3D+rUV7ri6XxfaXf
SHE68dxhDX/uuHsucegqsh8mkcUmd7StrrJJSIzLJ3DpQOrzpyWFX0flQY6muuZLqUg2iEtc1/St
746qnUavL9QTDucUAJSb0Omhu6XS+klFYUX28OUTBDvCt4cFcIkx/YICkZuyl+XFBitUaqfP1/ky
uN2auv5J4kIdpDt4nSnE6TbJRYauCaB5NOKCCqntuOpycxUZ3W08wzGuSlN36vanGBZNXHzY+Z+g
Qd3qiHmwzl+/RVExQfng4PwBuPXzEAAlFqMqQwe+mvIVoRm3hBgk52gsCryQeO/vkixYH1sLinhi
l4Q79ilqn3r7UK6my9L3Pwq4bGIbLvTRD+PbtjoCCi6j5UUdSsq0KG/PiX/k9xAME0gAaiWd2pvU
IlvaYBAAUmtKnGPsPElvIKSC4be1DQv+X4i+PDG+jPQ/SXjWj5rUi+LmOMN1qG323tPhpIxBLrdw
+rkVJqqr04O4wenhR52qXw0wAwOWpUKcrAvB9nwUXvIPmJGfmZbxyzXvoVmPf+TLwattFW17j0Is
Ehw4qHiWXuOUCV4T69O0FX0Hzv0ucVe8ZsVxrBC6LKNv+IlvZ1ZDct/x0kBMbWpAbFEJuSuK7gMY
WRovlmmT2ROZ+f566NGDI2bwmaRiJ1iPrpIng4nlMAMX7SFMGpamrmJ7oDTVMKWnmWMgv3hqW0gb
p4EBBMoaJuBoR30qHyedKdqB7niPsyoeBNaW+3h9fzx7JI2EQnPm30yWeIpZ2Wak0vUBluIO5OAv
8eIX9PHIvklbqNPrOQuV3xrOhnBdEqNVeD3A170r/U9OIwjedOBnBxYtEABRQAwam5LmA2madAu2
yZThKQ9gjVKFdNe/28z3SCuChdf8RKlPVYCYZ03flU3h50Vb/Girhd8W5KlqcU8I4I7Umnb+8mLC
vrVZae11G/fpYv3VryKPthK1tLbdkzKMAIaGOA4x8GbR9e9AZbOFbKd266DIuXv98/LA2LW2mbiX
gZZM2OwwhiGTxQMSOPGzdGEDcCACdS5VyhIz6fp2zJJjk7kJxxQf4QKyJJyAbvtv9DLkAvTZxFJh
NNp7dgWM/cysnGUP+7s2XsFmblp8YPwP48Tf/ip6h8TL5eF5aWA14uNAKuWuMh+e4u5NCLv+qLyw
lpWn8ZV/T2ciuZlI6PcxUK4CJJ2HPlBxWypMxIuSau5NGbs5r5Dd5NDiEmr/kvgjczsQ/Dg4mKcM
hkSUCo7CyuwUDSsYo7X5DyFwheDFu+Y9CxKBuD2CFutid6IkVRwMHSOuZZw7pPnOyeFxrEB+AYt7
i4ehmCnmjJI775Vr3VaLYa7eRMyF6RvrzlC2s9Emsiwatv6AltXNrJYN8mHY8Gv6gk5R2hfCaQ67
2gvasJq4RcwSfGvRfcnyLubyVEaBepnLNlb1MBkCTK7crTS6j51+9Zf7O/Ker6EdnD9R3G9Sb+3J
ojluApqPnVwHZWECt3LKYuQbMEz6NADeljCL0ijBZvoaHv3ls9SuxdeXku6PzpGudlAV1rqYZwCV
bIton4uC5ClOcVB3IwuhCyT+SmZNgZBYzvx6smE1WwtwCJF5YaruxK1scm5CtPGf9HSHcHQuUKpg
36m6UlR8Xa2IexMO3TWq5b72z4ETvWT8TJJ69RB6iWO+ep6q9V/DY5jUAEJaxmV/CvQNDtUg1ZvH
bCiR0p0KG/z1Ii15ymeRlotoY54GaNFfTmDELuAvihf+AfXxOgTexgeSyqZ3ACjnGoTMo6vLUXuY
q8PlEl5RFHJiz5DUUD90cI1mUgsuwE8boLWuFKxgODSsxPvB/7ggCvUu9N0we1VT5kMYBlAS4cjQ
PIrfDasaoUD01y02Srjui/ezcM9CCaFE6IISzNyIryVJgBgh2FQM09jX8fVZPpOXThQ2tu+uPELo
9tylmznJJxEE/2vZ9MUUS+zWt8nUayRgjK98WoVtReGVP7sj7xvw0RWlmzbE1h2sY1ax6OcYg6MT
KjXqOfrEPgMw19go4pPpKqsa5PmqamaWUNPUxslX8y4znSkm3tzom1S20bTmhMLoBprL0d5id8gP
1GiaFuX4q5UC0kQKAVR2qyBXtiFNlyF6T7DZfeoB+HaM6H27/uT3Jskl29XxKybPIOfp8184xI2r
qBHuJ6KciDc12TRaPGN+ga5866jB4AC+5apJPYol0kKUk8EcXRc71B4ghcMjGKv6eFXt28Pqq3Nu
0amgYvnIRHotiZce4ycF3eAReCZibZdoBCLJemhXzD5i0Qah8a9mmcjtXAKQbGKjZ6Ap/m62pjJx
EUMXlVcWeiN76CyZdfNOL6faycfrVdtXI37W1mxI6Ni3SNXe1rJf1QZarv3AQkXHy5EBQrg/WMjV
7dCI6SqLtzG67Dx3JMHL480rRfDbOM0R1egqxnddrE7YeNNv1lszaQAg46SzS2miB8DQHd/oHZUN
mUuyNylxyk84gZLs78lkHIqi71hjRPFLl7cBkSWiWsA1rfKfYCCTN5Dj41ue/KAXB5m0eVUddU2K
t3oqTDhNppi/4hCsKi4YeOqAziyDY5SaYcgg5Bz6CXSrhHxBjB5+0VCX3LyH+N6C13MwZHLH9Ljv
urEALfvPhm93a3dXL8pMo+7z33BeqWvM2EYCyNgDHPGCz0dRzHiLAaSgGEUOcQfod+E0Wo2rwx8z
OMTlO2yZwr+DGbzFRLGIlta9f35iqNLdHKcx7YcYvhhfYHxOR4lOKxkz2WqRNcI/+s7BXwrx4gjg
rbOz+CMXczS0xm2cRnow5V2xu+GYTCu3xSM+lGPl9Is2gIOk1CE6M+T2oMUpy7wuwbzwsDQzd4iN
vYpeZYEtIxEYDte9+1h2vpFfWoKX4Ch0U08AYJskQYKnjdZAKZ8KJOXzrA4ZbasyKfCQJ9nBrB8q
xTC+a81MC5nuqheGED7FmGl6H6SvcXAgAiRxxtZe9bT3KdHEZaZTrIX/ea1HLiW2vmPyDklRpq64
Bhq5LsfSTSHkzz7tBoOIRdBDKfy1P2+jSJooFP3fgNvJ58ZZX9euTdHBi9wULO+zI2HKeUxQ8PSq
uNsVziuFdlXvipoVDKP8eV1AstwTWseSplCj9mv9NcXeqq+RNMReJ6K+Q1UC8S1/BTCO3nsq+JDY
mZxDVLXiTYkkcoikU5RhYkR10u37Cg2ZLG0QpF6ey2MoN3Zl+2scPStFb/ZEu8AD/ihtFGrhCHsL
aQpoUtv7vGfdrinVNJTDU34xVgNmV36V5mGdM4Q+KLpN+UNIngmg9rRChfeYv81+WfDpf+wE35K9
IF7j593UwAubs7BKpO153IKLwDKdS46GAZGG3TXP+vyvfHBX7r9SCAppaIKUcZ9Fcq6kKSNEOX3G
kelUQLy0iGC9ZbvV2K6QmXMf/drF5DuCS542dImSEvOe9eooOATGOoj1komF/beT46UOGiM2ydCn
4++wJM2bY9lcftvJG0ng6EgGCpQtI7RS74WSbBqwsvuhncaBRcHMXLTafrNX6T9bboYO16TuW2P/
0BgvDHX5kXDBNVTbwsbLAkRmYR9VxDiHyvQlJ/xDXBiPjueMt7hJ4ZU61LO69g/x3x5jEL8snLkK
pRndyB4f/Q5Tzo0KGUOQ+e8h0LgMqKvRjNkDahiJn9OkTPfnrHHyGwtNdNaZudLGkvZJ1AnvBOvk
jZIS6qaABRuiJsXp3ogauxTmQN6rpu3ASpFcZF4ZoAfBugSacX6Idc2FhlpzBMPVQEuc9KBbZ+iw
lJbCdCSygCSRF3jjsckhOCqFGWVrYbYWcajXnV/xgiceFAdjSwgqstS/vkKBoQWYSIOLAB0cJrwu
e83yjWz3/hTtaF29ukQNiu6j9f/xioO03dxdVhnwySUWZ4FeXc6BJ2WmVE13S2z5sTp63PaCmQHe
I9HEzWCC1qM5fC8CLeNRLrWR6DNmIQflelR/KrOXlqo6lZOXOYeuJhsfWj5/m6PR/XSD1T1tkjSW
9/1+oLzIdvHD5dQcsMpzlESAv+sXapB/BAXpFgeV5zk59lZJzlUy3TaXDm/eYmmqwP8vBqfS5pCg
JVJHOmNpNpJCFSkG9/DGOl9DkP9zuYsyG3drN5Oiw8iOVlPMIMppj4W4Fs/m/dB8K7oiHNiR4hvy
KSij4wllKfnTXnZaYi7hg3po4I2tf81l3uR29DB0bYKk8Apog3n6Vy1nL0SzVLDkllryMPc0lGUy
epgVpQHZxhgnZOuEPHnwGMGzbJWNBCYzNV/L8Liuzz6DNnf0LXPt4ABX/pjQTbGquKRj2qIQ6O0K
NDbN7Z/Oa6u97eaytz5ig+XMYgQLPUbKrEp4LTWu1cpARNVmjUhv0rFg9G7ZvruSIp6v/zxGSmJW
r/+6CRrHMm73DFl9BHRWMj0zOWV2G3G3PC8wv81e0kUw78rSPwnOEfqVoNdrdzbwv2mDCVQln2E7
6ho4RM0s1pJL7+FeFkLtN75PacSqN2FBD5GfmT6d28rQ05MsHoJ5LKNR8PZaI/EN44+YQBULsRpL
tUoBH9yWiiFf2Js6FZ26IYZRjJQMiyjKqLPRQqiEadqdNVEiobCMVO1irdHC3oNRWoWb1GsDKK97
WAvijKcOhKhk7mZOL4YAlTNM7BzyTQinlSvvtB33IkwQDMHfl+rXnLSahAodq9X4qLVopeMryyLW
XSAqgu/lHNXKisUyPO62+FcX8/SnzEsgzVk+o5LHn81sCgn5F08bxjXeTu6Awv4aPcRUdCSujaYv
6WLFiCLNmtZ5LkSZNPsp91Wt83BdsQZlkmrU86vQhrs4ENqZ7YPSuT/EJ1+hKmfiKjQ92rGEvjEo
KQTEdKeorXO2PkFSyJ+X9WB0/jitaWE7P5c+v01kuXO9A2I1RcymKmYW79aA23dFZJIQI+hpJ8a0
dBpGesH0Jm/MneVmAk/Jn7vtW2w/CQzepD0ZmEQGK5HPRzlZnseDsZojRuVHR7SJ+CmDj0Ux4uOT
wP1Rkzc3SWene3BN8HXIYS13EQtKPidYVuC7p5lS0rI+PMwHSbJNfcrLSm5wUepTF7PG7I+xlDmk
Uyf6TkfiarYemhMoOAye+GEQS54apBrycczoAaHowd5CFHv7K140lUQhv3LRrqGrV+qmRhxPEiro
Fb4HdOeWvaeLsegFZ69SqC1JUhC6qwhaqri3mttW4ctW97siOyl9KZU1DMMhVw65OM/X9weAyw1L
qGHrzdrpw9TW7MBMpaXBoCsRxLuPkITrWIWEIJIJrqPXjNhRdIET2R/Lh58etKoCJDfYs/ZaZA1b
CuQLzjgRfHQNp5fU8D0ERjh1aHMAF1n7VYEblWVi8zblJOhyI9hPHjWAT2gZxP0LazJfK1L4uXaK
p9TDjDarDmZd1mAuuhYhfV5t2pkN+MwIgYepw1s8eTcZ4XeZuYm0ymcHOs6FieDDD15J1jVeepIu
XXZGz2Ik5hN4ClYEa+SzAIStNVx/66hYEslD6WEVr7jNlojOjJcj89AxaTJGaCFZCsj9XhzUfv+1
rrZ3Qq6hKBcyszOKzr+aVUy71xJCP0aONKfNwcOD4y95dH+cwvIbwgvbFBHB98oF4/glMqDnICsi
ZO8dkVNhK5xCn7MqDBT/rlr6DBC9WaGPJGb5QbKyt52RPomq2M8OAmSTRI8lusTdSg4TnsWenv0S
IDXwjN0YAGktWFufG33HpxgRXf+h2TLakLTQFGSQkxIQg+fYS2ZPNqJG3M3RX/JrAY0TQnl1onCp
hHGkCWZxBmZMAJl4Nxjske6trVicygflw8xE0DI/TGyDUmYLio+8+zPa5pwf426+LH7xi+qtfUko
XfWZe2RE/EH0mdMCuV/3tY759yuUyvzHnUyVgCuk9EBC+NHBXCdJcMFMhSPCGIGNeb2yCE2v6MUC
U1g53rcerShL8FdaxA/irJCT8tmThGsOU0h/pI5G1/M0UYF9ASvuBQzY9PWV36k/i89mg8YXtVxv
6bbUL8NR1Oi98Pt/0ZIeCh5CobS94bAa1n/tEx00QZUim4ctPjB6k++AAe1hizYbRlqns7ayfedh
PSX1EjgbS3fJFOyTJPegb6vDPbL2c9ZeKw2Gj2A7Ql/ULs8MuRKLj3ifHTyPTIh3ccNGN/uirnsm
e2xGniHl1/UN74kJgDuTLBqxP/vUQC4IAbHbBVtmLc1nWqTui0PrdFukN7AiC+S/gS6ra4x36gwg
t2YXAkmR1PTFM9gj9axAqCdALWMAWBVWUHOnHZpFh1ymRnOOYn6gB9vN47bUXgco6S4wQQHekRGi
4kCSmu1+lg9ZLC2uIG9iE+ZFyQPsFHo2YtUTeiIeoIWYRrllT63Cusr4K3RlDOUg/zNaeEBCDBld
2h8faUfK+OpIyeDIPpNZNBMwzHERAoBu/IbDYKUeNd2AJARXiKREdLcQXxuNAoCWRKOrVofpE8XF
aZN7MtK7qa8AN86HKVXr7QBk3E9BLd21WeGcEvpAnBRoNPY0QPjwgKHjjNLBQo/Xpap+FsKJNn9J
g7nig6lduZiJXjHNzE96M+i0SciSZRnbcrj+s/6KPZsfETqzICWniBvxdQxDMsGRJQlPPsci9NsY
WrntDIF5r4FLSutfagb/FeZ8LLzamoSV9ttbCqr8v3EBGfWZZb5RMl+BKueLuSuAAyw4YcF2RABq
nubapooVChhC/ocKaUvDk8363U5+j4Aa9GB9winqqWze2FBhl+/DG+FUGvmkyylCvGFmxyzZSFED
SUnR8s6zmK9GaRCV1jNIRwak8C+H8EwYVQKN03f7m9FVksbfTWHRbnomAuH9XafXWNYkqOty2pDT
y6Fp9D1ox2HnVbrnLG7QjfowAQqWkRblsDjo0+Cm4kVU1YG1xC1cavv7NR+kyK6kkQkyweZdFBEK
a9BniHrAlDSN6++Hj/MkOeKpvUwCjIJlI90yUnNYehw2lCm/du6F8dHmJxmyHxpMseerkRGLJBja
VnngwGZYmOSglYMTC1PKy711vz/N7MD7cOcRp/+YETY+dwSERUv3zjvV1K4rAagVc2923qHt0GtL
ociET5vqwRQ2aKdloE9hmDTNiaRx83x+Pq1LJz4naFNUL53/nKV6wwjTkMPAp80mpEGQOszPv1nh
7xB3JP5Nnp2b2YgCGWrERDCvUGwmaIlQe2DnfxsJ+qpoEcWK8Ys4Qx0RrIw0GKaO+LM1TbJux/E8
vh3adnfH3ZeXuC2UXD03UWRoYt6tG65ri4o2QR38uLBaCV6YOaNLmOGFeqTFiJRQ5DGECJnLzTTt
j9cCAPQWlslaCJ31118q+2Fwet31EN1TbDolOGIB2b05Tdx0BYd+Gi46fOYobUNCHBdhSBD49kqT
Bze5xkT9xiva3hCZc6zlgdMBxNPl9qYuE3B5IPog/Gm6pGAFE4eDAQI1bxedrAfClkqBngbdZdr3
hAtfGhRTr9LcMwoTL9SI90eJ4ALAO1vzDcGY2P9XOjd8ZqrQmUZT+IVQVrGZ6gkN2vRLUWMxWSBi
/EW1lG5fSXxN5ttz9qnMPfa7DmPy+BUx22RwTxRLbkx96957dRDCulnEIvRp/ArDw1pWMJxxt0uS
pdd0zZ0WTxisi4XGeyhzBPqpScv6sUaLHolg9qjjDKEQyK2HHXn8EadRTGJpt0yUHmxtD4Dd5lri
itwEi9RC2g8Ff58GNjN4NKUmEsrSPC33fXW0mAPHe6e8BdJ4cPUhdhz+3ON4xaPtBfyiG9d21C/l
1zRxB3kyPpociEhZAxosBSN2dhJpZccmSl3PFjTpSkKlcVvsBoTSxo7eWYkpX+WIdygwQcaVtoky
dkei96VOcF17Fx3PeHzFMgc9omRDBM/SQKNUGgpedH8cSjRz7RqCp+FBv0WEt3KQFz+KzDR8YILt
aNHnHeHlNBnvuKg0ocIIpJGGCy2XYijIIhmVmpw8+e0oJi0M32O6EAYEnDOS4iuf8ArUxOf/SMP8
MFebJtoOjHjn5AD0vPkr6y2HPIhuwkiRwOzWuEClmJQaLmWl71pUY0RI6SM0aU6jv7HXUOo0Abcn
Gmv4uw39hWIe+fGpCVWSS2qmv3rr9pUx3b6Gc+6bA9GjRqGIMgkGOFfJKPqfI7Ld46S9y0DZqM6X
qbyhhVeKiY+841Djt3tUmb0AtNIc8nuC4m+IyC7PTPfY/6Zqrq1wI3uYkavuUXifb1jNVTSPxBFL
UJUukRyDWhfJaJ+E8Ip+tGZz8Sc6oYbyNQKxlSQTJvLjy+ZKZSBsElofu5gzIyrJBWcjwiNRSAqL
A0wrWmh0S5nmpeI3+FvoXffuufgo2d4d9pIz4TWiJmsavft6PuKkaBhwZcZt9E09h+MwRM2t6MIo
+1DPtO4NlAUwAiQxCWaV/jH3icEjmfYmHDiNiudpm+7PSQNeKo+4ex+sgGFrQZ9bLmV/4Q50Tihu
mkOwwut6amXqKtDMfCcVFx2lb1OkTJUK9CNABJ4czqKTYNkWluv8tUAumCcTGekHa7n+FMtMP93E
vpccFxMAnZZVY+sobr1ROcOQvxCHVyvad7rmPeGfGDW/j4yKLZh3yI+rtfyYDn/2l5MKpSF5DuJ+
jBcDiEYnAj9aE6Fprk2y40sMoiwQn2oX3ZwshxKUKyj4bFAqGATeiDhiw9K6qvjtqhBO91q8x0NV
DWO0Lntbh65H4+Dic36AMsnWUHS3uDX3mZPbhwN/uhQlfy760mteiNxHK5Mc1OxkB76Z0GuwffXX
ecv/yNp6UvNKh4p4VbbB8NvP1vLAyXl5JQgxHD6RZnsigEg90viAv4m5XzYfJs3rnN3E2JxDK2Pb
HfrckaJHRmOOr21j3nD1Z+y3rsYhDFQuSkw3uUKrG+uOT63CuABHPXsamPvkJ1VvGUll8Sna4fl9
L4+jf47sm/ZGGP+kC6T88aC/epzUi69Gu9Ld7zB1B7hdxlG4ThJZTeMmTovcC34FYp/N1Md/T51H
H4458EiuZDsXSnYZ125J+mO6JsIe81hV+/+Pz9wQmDw5alH2NwDqIltCxFn6htDvfO6PNDgMrzqg
KueA9z0tqaEIA47UXQjyJ0Gmikl5jKRdpuXVlVx4/BQx7fyMit/JPoskhlNohfnmhr3DXpxFX6gB
na/UQEp9kEyIcByUM5qU+vd0rbwVSG1GyDvtmsMxSTJgt5o09rQEWGoRYY9VYuIXrhZMDE5MMTdy
vkEQKvqsVQK6O9EQAW9ycEmcrofLWjqiW99pPCEguIaMv4nUXK+gI2NtgcCCufiI+KIZWlqBXRuk
1X0dx31+/hiM3/bBQcfL3TU1ongZHieKC7r93gZEzKejJZ1VFybK5mBT+/GTZBulA+a7AGOfx1Zi
AYLdsjOXhm2qChCCe0m9KUQD1GyDuliAGQZ7cKY9DIjdPRSW0psVS7r8NzIfgYTm7q4rZtn10OiJ
piQ9omhOYDntzOuRv/Bw2hENWFkY8+jFKAqEJdxcbpFBt59n9jYOY2FHh2RInk6jgVoNbm+RWQPu
csCAFPc/MNzF6ra9zi6gqb6Oi2Faqj/OEtPeoWGr2cVfLQ9AFEqKAmIiKfJyGb6NT1Qok+jK8Z6L
3B8YcaYW3uZhdyjWa/06QoSX5i6kt4nIgnTl0KhDBo4jDcJ5YuRQIvK86RKn17Cof6Mt9eDwAmXX
D2LwxHtF+CKn8J/ovwLM4a9GLwGr25WsN+tHHML2/c2e5oDrCemCYBqO8fHGEc4CesnB4WZpyRzN
zkm8kZj13nbgGZ7hO853xWXS4B77PKi9Q2nqslzrNaHHgQnCHy6M6IaeXl/XCbsl0RGsnOXTjiYL
us51ptMS4jGGLGwAnB6/81d4L7KlbbWE+yAhUT+/zY0p3NJL3L+zJI1qX0yDGbP4nUGccdHaJVYn
+z7bBFXDsINgLkjA8K/SllRQUKwKbZEl6jWQ70dsvNx86kcSumeE3SX/VOaMQ/ljOfThq1MtjYUI
bABZX+LKRJnxUml9XOeyPMXz0FL6/3hmRLFhvNX2G0+UAN87eVXmp3aHXDJSO2u5fehYCULpxa0r
Zv/OXrfn/YL70lyX3K74tScA5MprScwh313N7EZ6tTBmW7y8ptoYDRCxUX7TMPQkZ6RfM9cI9Ik1
OEaNxyz71zJd3Ef1qLwdhGKMCj6J7DeLZMHWUPr4Ywft4vZgsKoy1FnocwjfF6x7aQzUD9Naza3S
Lskp2e+k25X0dY4a1WGAm4yFsQ6Dpv99HuG3GoGzzFIuTu7NNvShOjZHL09Cq0NeJIotYUk5jCFn
iTUmavWIP+HmxpGdvN5hjhmi60eus74nLTWaxkQgP1GEcNNr64cEK5zW7QHuCzwrIbaDmBUQVGIE
UVHKk+LnN7d8MKiuhHd6hMKluGuOsKb2jNsjQBzmMADBgx54baYCsSEOlZDeHDfsQqi0mtSzDxO/
LqLywCeO2HISvJQ44Pbp8BV5sXDDSpGWXHD2S7jqxDHubBvGK7czqxTxfR6wsi4jCdRKxlnS55kI
GgFI4vKiTfyQea0luPGkfszdZKspjSHgFcH+Cft2O4dpa7WhERaVAuN/9EIZlsyu9neCKHACJCGC
8cWMKLPlaLF9dN68UCqL6fRv6N+OCUye0GCIKTJg/ex0U1tuyq8RhHfNC0gMkUOJm4ZFLg0MoqZm
CxgFbmyYO4axnhf3pI6EhtjT0Zm6jD9AfR13kKn85KKwZwLPTyunqkkXX+EYH519zc85fQEkXjja
xziKy5SBUosC/OizKl4KnO9Cuxu0YrIrNt9PBNSzXQs33WreNDslzydj5Hrg+gqLlcNkPfavjjOB
BIY6k2bXwyTP6ASbeVD/xF8WIiDqqMTpnIBjZxjzIkFWB5wV4TmmCQlRSYc9eUMvvZiz7lyo76lk
QQpfvEk5QisDW+7s4Gm/xun9QZypHnvJFly/TIHCaHaLYO7wR44ZoUGJFKqxpkZvb549dtmyP+mE
r909L5ReQExgsz9bHhGZilwWQLtt2wRqjobVeKef+CshHmq4YEzjHh9l+q50c2J8T5UYUGNyhyuL
1dPQLPNy7KQ6nQr1EXN27fQpXwzuUUBeRPrFr+nAWC1H3qfukd1JqFvL6PeL8EGmPfGOCiEn+zuH
7kYyMv5KHsAiXbSNOAd4cmqqjrlk9B9R9ld/G4hh59hRbwapoCFfyHhov2bAYkIqjMZG+w+GHDFR
2GjK/+HYYqX/vegffN+USbUR7qVD//s1MatoH4M1u/H9G3sXHbrGggvPY4e0P4ivsQm1JvyhVNcs
5t5zLvjyzSIKatNd51g77S+sO5qMn3v5doHxHpa9f+82BoohKwXbyr7S38gHZzAi6z/Uvtu6iZHH
R1FuGKesghPnWb9kHXO+remLmLiaknE5JEtP2CKJbEciRrz1BAAD8lzR/d3r0DA85Nv3HG23ayRD
LVFOfVbl9YMyYnCTPC696g0E9o5mFSzHhEwq9ZHk7g3y9DtYawfQfUwHjLbnCpNK3IguLj/fW8bB
x9FsPdUPZLz7/hTFvnYBgQvVQP0OKYuVYdi7R3B1OXSE5kP5ufnQFZ7kFnXbOJizryBGmomPBl2y
p4L2PWlgMLgqe3tPkQOZBX+Z/Qi2bI7QcmXxMq25d0Z9hFDCdlfuKoOXliK4rty4F2SUK/3MlZZz
du/TZSEG0VyaHxHgdLf0GlyhrLTat7ckTNgER8OL01r97dAMN/yOkt4+HWEqaAEqirGXwfMqjQQA
g9Nci0OCqdIueqQiLZmrKHCpH7ufwBdv8wPXQq+bCrItjK8fmOWTcp214aw63553TkRX+cTVdJ6n
sOLdqawcV1Fuzv7GuK4m/sVI2KcufpPFaU8CsgGehZOYNrIDKQmEHCOLD31n64/9HWPRt52TXj4Z
TGDY6EYxBYU9EQDBvTdbQ4TUE1xyJ/2aMb4lDgXLTqlX8drZCT1htTGVd2TSFogElV0fgAqT6PMr
42f6Ew+ZgbfB1ejVYTTh60XeJcJdP0L0pEiSRrKFpuHN4/RFg5yp5tOG+BQuh+aJCCchWf7s5s2u
iU1IGOrUdseacEx2HW4tU6NfKQPf+12qOA8QeIzUlM2MlRgN68le08z4ikM+00edDcCexENwAVK8
VbCBMpspQ/btIRTu9gIoqGdigc6fawtjKrb8C7FkPFnsmwW0xyvf0PumoQJ3ttARGDktR3xfGX8d
1Y8TuGAVkqvjQofWvrOxZ5Ver4rNxyTRbeeFdY6s6MbCZPiGTWud/7HRAlSUCt6Nek2np/zASZ3o
v7nrUK3d+zNESzHCJogGnUXj/0PW+SfJsUKyYOWogUJUC4zZ4p9dUj73+RPZvlQ3ApXAIzCrpA/Q
wYFXvbqADgunVTwhno+cX2d+AW32/E7U3tfEQmQrpLB36FkC6PdPNIZuW3TCqdZxW6bCq35uV0Hr
uG1JbFZMP7i8XGpFuwbdNvKxIDK+nWCjEUm6V8TbZbjnc5hlZLAaOA1GhWD5ZvKFpGzhw9MIqd7t
ESoJgJAW6V874EtdTr5oS6lD38Ral9gjZ9/mmOtvB0/5N1v1Mqa0JRA+BPvjae++BEcJPjb2jJge
NggnqFwUAPGpLOuFvYHyYQUWEGvHoperBv4iskY6fXCGJCRd+/J/auSlOz9oZumLUkQEYg90/xwT
rYAY+KN/izs7cCTYFKnuZ2Lyuj2IgRWix8X+fzO6jIadnhm74O0z8jbboI6KkoYWBV5uoWFEVgEx
r0Z0FFfoOtSktl+obZaRlalwWpyC9PK6+/7DNSTCQEYB4v0XiJyfJ4YlbTMfMB7aZ6m12gSZrCfn
LbfHdnYUlEwL5O+gJXZMePme75XSOBjybIE0dZkBJpnjEbAdijr0MWEsULig9YmHpRroXJPMOcjO
tg6sVxZ7TyoWOSMh8w2IMdSrA0pRi/3qDhttkanX9fBNqbYGg1ZP99yMrBb2TTE3xg1F3asf3egF
z7GMyyK9aZokyJB8tJUYVAZ2I3Ih9YF6/4pTXIakBOG0GIAWSwHNGPIqEZQXlVG4YmoDk0fADqP1
CCZj9ajW8NbRKvvq+SnNZuuxRz9rO/Q7vUAbzRvbINFoShPisQNd0QmwiiGWu2eci4kQXZ6O1BeW
oL6UXqdVb6CDUBVD8JP9zGp8iL9rqw5W3zjvZ0orFSuEc5OeNaJNrQV0FzAKy0rJS/6kPV+tRHlr
ZKxUEVnEp4onuaHbnPksPEicM06Imd83XThejlPl/bp+g0ia3yrvcHBTty49HiYnHi5HdEkOIoHL
aA0Dt3o+qt0d3n8yTzTx4etGaGfzwlkHCvnxRNaHG2K3LbtaKAbHJRfbk2NnTM07mvpdP/4j/ujY
Py5D+AbeFE4d3fajcZruWMELvz8E3Tbw42+oIyrsFqFBlQun9cvERXJkokeImGnwXx0MyRfCuorX
p2/L6CX7qAoOkIdYHGQ4McumH/NZtdkEvYSUb35Eco3wMXVXGMCJTFm3TI3djoxK45gkZMKdntoq
bTPz7BrRHfxYpw2Z4Ksipm4d2CGQ0yv58lzSnlfY1XCbmYAtIpWIykGDEYtOjDCRQEKg83o9Pwbd
DwT2lESpVUKop3egOnQd4gQBNpB+ZjLKbEvxxXckNUNW0Xmuz5Ofr56dsFcu+6HsOtltoMnH1Uwv
u8KlRC131B1bcMgWRu2XDcCHs6BK3uo9NBKgk4T6Uak1gjNQWCjvERAkg2KL4TJIe9dtd4QkOMiD
g8ZSXWxvhh+Stk5RVeFex+E5o4twDGZ3F/xPYULJEsTbDAnAyvgieaV23JwrCk5hLZ1fyp6YqojT
+SPEq1vR+zJ26L9ciUqPsvsU1Qzp9mUrgIXhV8xn2qp1pJ9FButT+sRuMyW+uzz8F/TXEHpobVed
wXySWlilDo0WZ0kZGUo3af0O0O3DxBKDiKRfnWG6Ii0gOkObQW5BQIm3qJboxIUX7ynfK/Bgsq6F
9MpRDyXOVaAxnSU5qNzHlBl5rIDTBjh7fckhPmNePcvILx4VYNzVski7TD8Z+8EER5GYa/bnhU8M
eIXoza0Rv0685Ngjg0w7vA1h1y9VEd02cMp9fCj06VQ7JClUFD7ubWzL06b+w1BgHlYRCAzBO97C
YhVKEMPJfzYQJLWg/S+dpD36TAW/OMqrQlEcgFVILVGt8a3nQbhkmoI+2mxWEIfXw1M5VMimFm56
RYtcx9pJnwlHtONaFcO1Uf8Z6HpfBPP/RyU0qkmcOy0/uf8Doclfjh1UC8Y2fW5QC5NYC5YvMvZM
dTeXfX6rEEBtd0jSrYvuUjCnjc56KdEGknQUFBar1DWJkwLpno2udJajlCB5hCmWaoRCug3ZC5gq
21glvot8cN/3TwIpm3nYv0yDzmwE38j+9ZlzWDq9RUhCOb8XEUBCeKgO4n9WzYdQOds6ay6Xx6+i
q3bvlt/8MuSF0WQbDQFvDNEJuanT92u3W4nAJ+92hTFUetxuMOj42kp3Gd5d41Mz4YphV9eJZefr
CMONkVjTdBYwDHuG4F7TMeiqWIuW8f0b1IpK/a2iIKpf5vMklJcGrolTmSax04KTUItGvg2aAeTt
Shu5oI/7GOlX2AQvA6zexlZiTpId4L6T1HQBf+XL/V/YMcGuwwHvr1RgMpoDhLusYqJJAQu33w4b
+eyeehZrj5Mg2QwuCeMZ7lxjyrlW875hUkafXGH/HsXNArYEh2dP7yRL3ij7jIWlbwfCKOk16/vv
q/IDkEgCggrY3uXF3jVdR+KLdpqmvwgv0m1kXDkUfMnwDNmB+kO3PxqdR1QvaXWYWHJjQCBxL+7V
Tm9T8LMy1qKl8h1iaslkqSAcxV86q2hAcOKC4GI8zoOuRiLW4mby3gPyRfQZJp+SbZxkdSBBr2U3
0VqWBfaXCwlo+8xcp8KAGDYcVsI34pJfKBEvYPl2ntR5eX0w5Qd9aRuIsTPSdA9yw7ZJc0p6+npK
04Qeh4jeihGMWmdZpc62emDo924ZDr2dNZgSmNtAOf4pM0qJiAbtsqYYhguwfqO6sSFnRWx/MSKt
FuMp5tW3qM/wqeEATaKqPsYGWDgQRfHo4PORZR32IktReRP2PMABtlWJg4R6NUyE68P1yWqAQRcf
/3K5uVmI9ccqS+TyXA3tvFPXAUrpYqszmfstv7yNC9v+G9ijPl9VXBYE/i5nBP3lQDMmZw2v5q3G
oBe3qNMtosx+5kP3j3iCAUDG00iJ6NMpSS7Oms+jCEK0Ot16l1weraIDc/rO5wNTXqLxzoOilFZ8
ecAkTdbPBVXD1U/fMl0hs77ExPxwgI7BQzIcEWSj2CuDboNCwuIgLc/6mFrsPEtJ/jOZ/UDgQCgS
e3k85+OFCOKuAm8XCunh/JyInToSZ1OfS2wNSAmCZbq9La+1MDv5YxuXkgFsPgg3qwaHFOlNd5tX
GHjYYFuolVrOD50AbIpiD/Eoqyx2ZY8Kej6GCdpe0YlX8xMSHwIwMp1vfdeqXZiGKkqZdtjlpYko
AwGmC1UjB12IUGTM12ycWM2t1HtpTIYDXySUbLE4+ta5l9ZfxE8UBT345ZSx5fawDCTUzYqsL8cQ
mhtlybmY38ceSrSF8q+lUlm5DVeEvovXgpt3+VXvqJFe8hPnUVJ7jeuY46n8D7t58IDeHgNYfxkh
Q/q1rJ4ZiXO3YsLW6pfTru+9p0PD9fmxYbrbm32txCgYhQx+nJwpqxvYEw4ZWuk1vW+G0XjUtrAU
u9t7bHSqsVx8KaZs/iyKHVdvqzrQG6jTuBAuX+UOnnou76pAXyii9dwISMtICrNoz/WuIAOS4BQg
WKIk9nKI0vei6Pscr1IwndvBt6U+g7u0rSm5kIGAf2Xpc6TFGNLqwHporrsAikDHvM0vEAaMPyPr
cSRK2lWumpPX8ga5KrtXmqJVdMvgdOLGM06JYM8L5uJwxgdBwG//4MRM9kgcZ4sQCodTNqc+LJLm
i1/t7QrspFsXt4AJisezxOYLNYZ/CoLjKhmZAKPlUeYkXDFkjYu1cPDqhbXwepwDnMMgF85TzKMx
6GezzaiQJPdDz9QquqaM/d30KhPwKAWrG3Xb9fCItomEysYiLSez28mMWuV5QnuBJvzOXmlZpQdy
VAPDCVuFmA2tAHjMMEyuZuqb0xhJVAVyb651seZqt0VZZV1i/2rfYWkTWWyTF+MNKkfgdtBlrQ52
HBgFqqAisDhv+xdXU/T95oA8BiZllYNKTJiq3XBu7WidURwKEbdehqpjZoP7lanFm+7mIjm4CkqR
XDBSx2TRHu3urwJNLIGBLIXozGCsk9kJhdpGzpWVb0+hEgQvmFxfubK3qwLA+i/tKm+JQUJGMxSB
ana4LZANTGSzDUW/mM5LQKU38PZHayueyQyqpN0eEmU4SDTEZD8VCIDm0YwVbdVoTWDYtptaOWYq
vBvhPiN0ymAjj4QweVYE49B+z46KIh05oXAnud8roGzi98EYyo8oga7b3R3P35YN9Is2xYd6nUvB
f8j4aCo//8gV0FvS/QWJZJXZPuO4ISykGCfI//0GrTQFN3yb3bZWK8lL4+KEUD/BSO1FsfT62gMI
WzxRWa76N/sFwVorJlcLoqk5EiMQQUzukKFVWoDrKvHjUly5UECi6MoYZnypisiZfsVJa3z5K4/o
fvyaDIO3wpYG6XzsiUHcf+67TSAoVvA+r64h58TqjUOjqiVPX2eGDYhGxkZEsI37p5rZqhyKEMif
vDvnRrdNkoFNhXPWwiY/rDz04NuoEpYwHqZhLzD7oahhkM9Tj/F4jVvjf1F15Wg3FUrR1Vsq72Cc
F3LvHQe1xccaCeZO1LuVd7AK6+aXdEDHOe0UC5Ozwiu6IUP0meWqQG9JpBif7Xwxhr58Aj2PyXcv
lnr3E/hFa6Ua8CdwGKGok87TQZ+8tL7zE2C/e70r107pinHPJWeOfJp4njuHBL5GfIHel9WqS7De
IDpFgsBtq7s0sSVoWpv+gKko3PfBjCN+KZClJNzjoADEwfTDlH8LO5siKrCSk+Q4uUnIWVKKf/mz
pzD9keup6gyRojI8wHoUWhOxTWtNyTPLj5vR8Dyix/6GsflIYBvVPjg+KTouYcEX7nMFkCHoXKQE
u3uj38VH4W4PtWDRi0d8vwddwn449cZOj4npOiTZ56ISgVb2uul3/6tOfsGNNWR3bMqeA6V05cL0
20wV6thHgb4k6B+sG9qHEEz6Iy6fknzT6Tm4ZiR0UKg/aEUHhSFL7GXBPjNNq/BKixraPPBAQ2qN
QgapnoFdRC3zrMStbrkgRMEwFkdpQu5aoj77UyI7/C0VE38xyLbcxsfBgOlSg0zH5Z0RXx3I5WD/
cZFpMMzlJNl+p/0BfjwGDhpva54SmnFAOgBXlXIPWwxAyoY5gmHmMXv6cMX1qyWsygTA8zkS+lWA
lHZ/tTsMk/mT2U/dxJfim5cJ5tM6+YyUQXCc3/KzCBzGpD31/1fG7Adkf4fzQ3ZM/gJ3Ioo+Fn3U
XRAXDyJWPEut0qOpfGYhC4aw4uCz74sxohh5Nig3OXbTg5WPqf79iBOYoyQBQcVhq4j/i07pTu07
rRZEETiMiqNicZByX+dDztw/qD2C/BzBVmD2YnjdGLzNbxFVuFUjdi7R+fbAfqKLKcwRF1WVbg9j
xIs/iNibrEKmIFh7AryP2DR8UXecWwGI9gaNevvlgYecPzDuzXBewnuo1lEC0Hd48XK3Ttb0QYT2
Dtf1VN6h5s17+oeWbZhX93HGUsQ0hlo/LcdQ5xsvYcN0dxDNyVn6t6E5QEXX2OKy078KLg6mZ3FJ
NiA1PkZRMSFqsHopi5+iU5yFq1FP2IDAgLA+Y8FtgK2tEF6B90HaZhS4Mf5/TlzVjBZ5EN328pn4
/nI2LmO1nEWp6RrqfeFQAnkSLJeGSHQy99a+F7rkoMS7HTd10Udp+p852vDcp/i+BVXas4o/6Tfj
j9roPI8G+LnIhPkr5YQFBAVyDbZXd+/GFGoiOLJZ/eZsBNiepAowg4HPNep1QopxLpdn8QJvQx1y
fRFiPXldr1FJkAFphb2sNhsvfZy9RNQSX0KgUbc2XU7KuCGM1daTq7rSgzMa6IytBy1S8MGNpJiW
1retLsYU9lOPYopd3t15m7nH/K6zL1lrj6JXzvYOr9gb09DtQmaIveixgZrLODFXrRwmw/C0aGwD
oGUi0yIfJMYiUvesupQxaMEaM8zImQpHFKYn9Dg785OOn1xB+mwKRrDAK3PdmLJKMTGfcQPa5dw8
Ju+wJ+X646Hu9IUb79dnsjh8eonCTd48FG2AJRgqfrFRC5iwCW2cFrlb3f+x/4jupQTMABywXTgh
fk9oqdNd7BA8tWexxlK0G7gJY+L/kOu5ntWPhk2QAorLX8FrDG7Edvs2hpW9QUq8p0Jl6owwpGud
XLHiDck+uf0u9BR2Jvpo35+8rRhyiSeGFp31vaUgkn6R3pDF/XqTVX0HgF0uqqvOwumcrWEnSZiW
2wyMtO+NF+hanJOEBEIYeNPZIfC3H32rtAHp7MzApQ0BivrpA87J4q3WPdfLIXaWh/mcQTZBZVCX
311UUoM3Tt08Bfk8dsWy3AabvxQAa44yU7lePXGbVZSqChHpZ5Kxp8pEofc1cD3DYQFSn0nca+4f
Lrrf5GWBHeK1VD5L8xTd6kZ76fBalVwumQexkO2bMMfV8E9ZaNBaOIbgBbmBsrh3GFy95nKiIufb
NDlEyfOA1jM4E27FMPpnR1iAmisOz5kQgypJJgou6PtZfl8bJMGtASp9+graeckUUOq8BlISxIn3
qRfmWMnWBwX7Xf/Jb3bp9sLFGNJLmKo53hPBsdknMf9TryI1EpIz+8G6LGc2ko4e5/nHtvLK82k9
q8MNBk6Sc3wuwnxwXHrscwsUNcCW8ktMmkuWOV9xTjSwHLHpjABgfMpj54BhbVAB/uqGR52z2Bts
Yok6F8TDrLdlVuzdwfyHZUY1VXFjCw9TelMdz+sBc5ofQfhupoXkgMW+PkzrtT3xdWw7Y0kzCOBP
uCQs7L5xsJLrO4AfDQ5oF5lUR/0eBnejgcgarqmLHssM7RczQaxkHmNvh5ay/Sn6QWU2BPUnE6Lk
4mw857MvD1y4BwVM7miaL0jjnOf7iUo0SwSgAydnHthlvHSnP94EkPZV4bwHXJBegTWknVBrlXo1
pS9dHMW/0cO+9+ExpM3ceHIBWzsFTADAjTOm43XBWpH60boEhkSE1GIQswG4ggHWccG65YG25X8T
SpkIXjKxoK7OYFNLHyavthL6C5wUPaVWAW7PFY955NYVzyggXB7HhDGMaZpCf0OwURpl9xR08E3v
zYcgyNUPRFg4nErbLdBLW6eqt+GX0rO6UqP21bsw6UWZZ5mM1+WJuS04YRFerpMgXIk6nkuPzyIb
oXldPd8taWtEdi4iK46QJz3EFcAqvh9fC0XmArwa+QgI7lVMw+prYk3voo4vPxjyegr3fR/WNnf5
8TRR1Dmx+6it3NiR5fPGwoo/v9gxKsMaMnXuUzMQQFktuyTvCoHStxUD7Mh/0r9Pd1K0kC/6emXW
obKOaPc3HON4BXjNSfc8wPwdjK3cbIRZr8ltWY1ErkU7NiP22G1IOB+PXanZuwozkSDdf5/p9DOB
6yFBal1hAbfW6fKY2A+rstExSRbjggFfczUZtFkYV0jeCRf8Rw0wn6mDQCdBsJuAsSaDdz3srQjV
WIQ+Mlsx7qOQQKYCbCVuqJk7Kbpzh7VVSWmUjT5J0l2vQpbDkk8Yh6camVRWtl7G6g/qbzszKJWL
hOSikuY4ZkcP3HMrp2dADuedLLqMqvvcuwk7Wc91dypaVNjXCbhg5cbF7oL1YtbEuF1gPPH+legw
7XJh4HmXxpLmmnhr37xqaYLnzinpFVSd+qBosg3EXyrGQZJ2cIkbkiz9gmqJ6AB25UE0eqkFPFDu
TMrrLIUt1AydbQ36ehWxxtCYqlixPJUgxLNtIAUyGtzDhD1KW5qvuipZ7DT6wSD7UR6C19/mJTD6
u2fTGO6cfKV/oty/BhQjjdfFJwPUCf99EGoJNm34Bh6oVAGtPhYj2bqyy7cn71c0IS397R/F7ONH
NgPlnDP9yCkutCiVDw3np0mVt8CrbWPWHKmgId/IehINgKy/lV0r5w8BkrStf+w0GQgd3Z8A4fCQ
nUYVMRtZAZXVrne61fGPhB0SSrPBzxnnxlkFVWxpaxXjdexJRzrLCS9AS9myv1zD/E1k2+O5wjue
dg3/20uDXKzUkQOchdxaw+jsGz5k8Lrrg2vKigxkX7tJz5hypO9sA3Py3JkKAheMLdCMSWdjPQ+t
zUTgBisbcCHJzeTmnWbdVi4t7MYuab+tu5F8Ojuv8RSc8Xt0ORHtR4aHP0quSZDFZtIexQGhmzB/
wtdOo/uZbOfuE5QavzZmuPRlmJMq2cJ7w2U9Kbj1vDRIV8hiPPCl5bWoMnJypHLEJJKKXDYHKDgp
dJexsfxdejkK+zzjACxBC3qXsZBaQ+Hl5cu2F5GpwAgjv93g55/G/zzGsRPP6EVCK6WIUPbHuL4m
5P+znHEkD9Em0nCQzOWheXQjmgX+q/gK+GMOeHUlk+MKRMqjRfyAX3QeLwQO+vvU9ynCuwiEAQ0g
gLZIOybS8lIZOvRGcoP3k/N0n3D0pPojKXwQvPE+M/kvZxUyj1ihvjtC6R1z7XoFma2yrUm3nk04
aInB/6QCru8MH/oJ1OnpF+dRlo6dN/u5yaSAT55H7XEbnGeKUsxTZ5pcm6KpxdFPsdUaPTWamUD3
93/66/s9hEU03nXSUQb13Cq1kydbkUK583kHSNjXG5TgO6EqmOcUXoHxSOGtxVKkGCDAdfg0nIFH
X/Ek2xTCVKAmT0TAi9Wx8EdrrYaCtYaJBMT8fk+XRh1wfTopNTvJ69C34ePA09oqYDvOJdIMza23
ruP6uVZrANPCvt6dtJqy5OVifTOjy43QFsVk1BTSflGke694hsKqaFrJnuzWkou7MLYfMli+71LQ
nn//uzmeFsJ2SLRUohYgvdqUn+JvZ1/x7bGpn6UKkiwUV0wytZq+EHl0ZD+ds19/kOkYuGKA1+zP
fBSUKJmNMJKbXzaFu1shHMBzbmplrJZSfIvP9BJhHWDUmLOIi/TUziBWVE1UeiPdXz7tGmRqsK8r
Gf+2DSGIMIFdbdtpzKQY+vXmJ08+diXPl9687xuYrM28W8hdv53AprnqZJ7oKWk7aKSKwgLRN66f
fqPQrA7QloBaNxQFGdyy4DfuIL7gu1El8qSgOcRIyTTsiG5zxzWWpE75kWEXBMfJXK80t6fxtENm
6tzol7TvRfDi9XrbD6Gb9P1xKRYU8nOrn9mNt9l3ouGD9/GeJs0binLsqXymlsxw8rAzgwAHR+hi
39sKBqKl6ZmvhYXu6usIxiV8sTGCqV95dzm3e5Pkkhusur6J0RoL712R3Dvl7h4xAepvry0UKsjl
zLVDWd5hl89DjBKRiw9G7q7CHpy2a6FryuS6gPFSh8uheyX+aV17f65xx/XnzEq9dW1zlu2MwyyK
hPyh/jdf9BKSbWnoiPlbJGJWbYrMGJ2PSr7kfhTsz6DNLEZuEjlP8F5PRt/EQA1dw8vdU0BwAJJg
bxOscpP7AwGoqnsm5UeJ4Nqj9IBL6NPpQU2c9tK7/rKicC0bcFvzDhlVZeKOmLkz6ZiZ/+vsV9RX
msVbWgUFDqHwisBb6l0r9m0o5N6NLQJka9gVCA71GBbYH+KnaSLUEZ6+Q7A6bHCALIXmthePvYhK
NJ8eVVMJIIJTtdNwypWM7xdbPmMJOB6KwvxsYWcMm7Ax3X/HmhBJtXdtVHzcES+40XfLzoPk/64E
jQ6R40C4rifgPMyX/egxj1NKMflsJqA/1lMwHsaRUzEjj8o42JUcLL+6Hvsc9AIM+q3Dm6KfT+aG
b2Qbt9ThIc4heSPN6KG8ewDxP6RXb27ChPQQk4PqsKWX3VR9beht2CGYh1/AzKP4nTuJotAbAf4C
jEYveQ9FeKclLlsVIf32OF9i383Zqb/L1AfI6oCLd4Mch/ZoSSPLeZ1XzQC47BAi5KyEPQV4lw8d
FDldq3Ke8CH2d1j54pbcLaloZIf9C1xD2L+ikvCinjCBPHP2jo8FbndtGBj2XvEAAAG3Bx+m77oV
kFy25ZlDW9PtCiL8AXd0c69jTWDhoxRVnuDhRYuxQGCBqxR7eTd5ocpBJpxZJMm/oi/yxhKh/Xkw
3cfLo8UTwZEqQ750elf9f/JPZOxt3pqXf6vkBjkXnkzQKXbDaAqJdPem0oV61bcDSjT1sKCTX4cW
aUXAaCQ/1wdEkYHASmfcrzQTg+teBbupjUpJZ5Q3r4t3FP9YddoRSifDsAVzUhLoh3zbUsXZoDZo
4hsoKQ1yscm1TMvWxfTPY4NMyYCArQNSF0HI+UZMnCPCMyE97XESvdlWU4Q3oiUdggwU/1uLM0Q0
0mBFVNEO6gvv6nz6ZNXizea7708PhpQ44UiWE7eV1Fgs/SblTPG5K1eURHHs8rE0/rtoGd/4Y5vq
+NWiyTgKCsKQsGM5GfeTyYZQG533YWNVor9qM8S+9ZuXkCbLL/Pt+b/YVv8OcZ9HPklvGWUEGRVj
vKgTav9F3EGHsgdAkVIzgQ08e4sCDxy4np/JYIAvTaZbtRcInfygeOOJSew6b3xFKxXOnrOxWEE/
wzo2TabjvZBsmeGTAD32UTnWd8HskEPeJcVDh6BzgMtA3H/Nzs2ZcAlh5HrZfrgOOs4sNCdAWxRh
gHLFYA7gQyQkLukMO+CRKoxTLEUc9b6jz55sNyvz2YPD6vry0CnMlY+nty4LnbN6zUwLw73UKw2A
T8AfoABFH3nKEPrKZdvApDUFdcFEteflEaNzM8YZpAwIA5op3dOJkYalij7lMaJnOfzn6CnyU4TJ
U51RYgKOVg63k94MJMTEKcNXiOH4dD1ZpZ9+w3p95wvflHafeVZQPkNQPoqbLr9gVmsa6289/H+y
cfBJklPH6SdbTJsvho6MnraZUs6koz5fYxs1Rj9/BDE8RWni6il1CDNTzohxQYSFQaDQYikJ1B3S
9zS5seMRJW8xG91KTdyJKPKXHLa26t8e/niEyz89nPUZfzNO+cn5BmvjBjJYnj4KuqRj0g7UgNCN
4ysKn4HvuYKarTEeSsgkHHXR/7dEHffSOrq9MVAC3E68qmf1IQ63PIVmCwUv/FOWEZDHEb+H2SQz
ic6Nsm5qogJ2FvCU+4WODqPn7zBvHBi6G4EC9ShWDNIWjWrMc3Ow+GvojsQ38BOhZ7knhP4jwSBF
3tTzYq6dkh0W9Qeq5wKayU6rlTCtC7aZGfrHWL/4a98kXWwVOysIGW708KEDfwWRKM2cXsK/kQk0
5rULUWYr4mg4g79Rfbl4RyqsYtnpTXGI/Sfay3IHAM8xbtNBo8a7f4ZyDAVJWMLo7ZBNgg0eftNy
fjz7HttC8oh6r+Mx/aQoG2nuzUr5/Mo1cyxkpKpt4BLDTVsjc25MYNPZfm9qBvl8pOmr0azj+cnE
oKQJphV24lyjPSH8CJIGFbTAfJOiNn7CAnps6Ep/joqUTpdwfA0vPdWPEfYuA58AHyVDq65XwTKm
ilECuwnQCIsnSUkh1RT/Mk1uozQhk0DSwyIYWn+dfbCYlh8WtqdMezJ0A8FdP/A+MtleY47zqlO8
qONjCGkeyNG9Rpr2BQUFC/7A6uxBVbL1T/pLuI9BDPXa3O/hb5/LasBaeIusiPEk5cU0MHSCZhNz
ApBuHrjaaRHpxXFa6RXguskr0SDew7QTcSp8H0MABRzjDm9JY7WxSGBUI6InxICY1CLOrmcRgpxN
Nc/1D54f02GyOz+9taTApO57ec/VoDGxbdVr53IqVtF0FIaCSSHRl9Os04P3stbVCtaMiUPAq/Zg
t7vByekwzm/kLtRfwPEEbMatgbgDY2kAxKa2xazuc3vxnmQkm6Rdf/BkpNE8NlqaNkpXUNRGMb6C
iXcGFkPHOU8NdIGLHCYMR+LPumChCNuWIICqGuiPuM/tCifDPG70OMHsemEVXUVf5xucDoJdnOvC
HXpjD2Kk1/pJBcXDUQhQhVIIJJuXD2ZYs5cIg9vJIaRDdiG2V+xh/kgykdvMJrzD5pLQbt0PNcpn
07yeJklbwmyd81cvrUR3n2HWFHlCa8ksb3feVKZGPhL9LldSQ7g0Gvcc9EWEhNLlDrQxWwhQyFaF
DsXOqH/Mu9rD8dUQYO095g545EjymvZ60REnkd87IfZ6vYyjhVJvY2iN545peLYxX5CjAJGkc8a4
Pzu65EYg/N4hh54C9VRvIaK1xEFzwZBvFNrgilVbiMYIHD3Fj6afz8WT6JYGKqCW4zMXfHt8bJ2A
NaKWP9nwpZs+zZtPSDF4cqWXCVJdQrq1BnsmmpkYkSoRtJfDPB2aoqZt8yH/IVrR+KOr2gUzFL3n
IWagdF9sol/J8sG+OI+7zEjLuo6qyfoxCFP9Z14UA3GGRW+tau2+znJ/6LfjVeOxshDg1xGWm4Bp
Pc5oA2VHpI74Fnxz/Lcfm+Sc/4db4xR0HLTWZl4Ep00IpfCNnPGmz8LatY+P2Megb8QTYy2236CM
DxsX5D8vnvCJWIQE9DwSBZYyAGS1HKV5ALVtHPIkIsIiitc4pLe6RDTw/x8jsOYVZ9nzu652wUi0
7YsEeTPVELK6Wuw9gzWRCLa1ILzymhNEr4QCIy6ZHHCCLSGUYARcY4qfR4LZdmfBrj/FFSqLxFZ2
yxsQtN1kFCjnsA7uidCQzQgCOBOtyVI0uyd/3n6EawDATVxZocQZb5d/56NDg4iY1rWi54kRa8G1
CXQON8SL7VBbVsAaAjPLpQDzcyAloCUctuUBfAJzX0G7i+BKdDy+JaqeSY2LidtWmeAGrbhaBxP/
eymp7OBYeC3DPc/VztCHN17UK+vCkjVx+MmZvsnrTwsxuEpQtqHjoSCgAMJ08LDxZdqVLlZ0oFIK
hFxqJ/NwHi4YeaqC9ZrPSmNu2/osxNZatRmtT65/yWf2JEuH8McnksLpwWp1ocN0LgvJY2HWU/Pb
qs0S9W4l1FKJ6niwll03p465MpzYeO3ie6DIJiD9qMdRS4lxToCowPKeuBbeLbXg2NWVrNS8R1D5
ZAEV1GGoGwuhpknX71fxIslscGp+3pdk+o688FwMxpp7W059S64Fb8Yc2Ghn0vlvT0ExtCTcdjst
uJi59OIePO1NpVlbHkKfeDggcHDgWi6qkpZGu1EZEEWkTOdcas7PwZJqApAe+o2Qj2rFjOAcvsU0
77bFu32IqQ2lRqvVce8QAJRhuOQHzTTkP1V7Uu6ESQJ26NyeHFUc6CmeGOn3hTENIrUMwymtoQwG
OYFFOU9JhG2aw7hV3ZvqfR2Y+6EOcBM1sb1yrIos1oSWiuDLFirzWnRHON2cawwbVhR39/9ULHa/
TF1EduKdEKO2IPMMp/riX3qeplXZt9OPHqrW+kMVs9hSiQoiByzTQwB2Mp1VzcK+pAmHEG281xKT
5DeFiX64TfLhvjVTGmEwwZIJ1L0ZVRu0PauyHQYsuedoXtuyYre1Vkv1g4nyL7FM7pYWH46SVxcl
AEW82e4U8tmDKMhsYn8VRQqmTn3Wmf135Uaea/0ud+1XsQHtQpzu7LbHed3RL1uyA41YxuCSgzys
Fr6wyyx+LoGe6wmJSBqUJ7YH5YMzr1MYdGyH8mPyV99rlvv5636Tbmk6lxy9gdBoyTzxWOJ8RPQl
TcfWwavBXTnepYpYnytmrHOF/gRer01Vl/7L1vJYRjQUII6P6aI5nAU9RgPdF3sz+U/3ZfuW9xYa
Bwy0gqml0kwQlOcY4xf7QGQZVgp8bT1zQaDAboJeBG9eP8VkTFynkijGPflFVQN9Mk15n3lnpBG0
Ks0rvwNvFMdNNiBfsrOq4nBNDFNC3ADW+HA7+S3BU1X3eOYMy2dCT9ukXWvhUO6iMh7PDpJPw+AP
qxcYDbKNwrEQjQHlBqDR13LJp1Yeoy6+h7beSYFxv5+eLetovx1g5Vuf4TTj6BwDrJN+TJ8Z+9ro
Ysr8PMke8dR90sWq/im3h06I/yJArp6ThUkR8mAdfpcxxyogf8CzOgTmBMrl2+zFkEeEFEWHYkzj
540DP6n4eIorzLsfobH7k1WH1V8dR5Qcq2ExFjLTvfKFbyZg8V4t+1LsqZiKrod3s8SKitpBFEYV
nkuSSI4zMqMCDTTidKWd9gdOP+V1cEbgg10HevQrntjBzM70v6MvYG1MDfoZTWWP74k6UuSHfxbp
PCnUhT6BuyNlVCOHSBb2DMZXcVNCjB1UU3xFHG7wp9MlhAJt/i7oXp2Vl0Mt3vu4Jh379Z0Kdnve
LLr+woUzfK/TjGvy6lxlsOg03+FQlA9199X2T/r8yRQ8ScbpA+iqQmPTETrEhgxJYNhnwYbqOPDG
15v1awYQm1HyxacxQO8wh1cKSVWftZiVbCO0S/Dzn2pREJDQqSJ2qgiU/DR/fv/mQWdfywBxbHQ0
MRrklfSbuNlGLk79LqGtJpAdfM4YtzHeRvGgzSmuXwYUGpicVRGmlGuRcmwX9ns+JlUOrwLipY0Y
3TIquWI/GOWem4+elwCzUx2k2+4Jd5Y7VBlvm37pjZbhzOTovkAc+cMHlCyaNpxRdKgBbPkfPL3R
hSPNHpOKNllLZwzd/pkt97Nhf0wGRXNEX1eA0BwuLp+7gIubjn8MZBcQgtPlmjN8wLycm6vTAgUW
3/ClnY+L6NGC4960M8yOogGBMsId7vZoYqHymuyoDENQX0PjXbQ6A0iYmUja6V7kYUxm3RBce7zh
rGBwLd7o0pWQUDYlONmFRMHAxTZwoCZZz5T/iKUhnHYI2RtwzMFubZscGtZ2vsl/ghhpEPbsbsT8
7nHnT7YqvnT9Inu9ctyIBLXtWN0jI1JnvWWQmbizMzJO5q9QQ/chgmfDsmItQ0A+yaiNS+ytN79p
ol38o+4pkXcy/8F+qfx44UUrzClF6ZkNFtHxe+6WHh1MrpkTliJ6Au6ikn7VQnhS/Bb+bfUqvcZA
BPdQEZkdVoCGNqbmsFwbRcCdmGVDorX/HePHQVOIRpBl9uT+PMrbn/zXIpJBEF4h6UyO+p6k0mm7
Jdg5VYXaHlrTef8mHwmXrYbEeONPX6JPSmVxwtzYJXpI8GOvi8pLEfKp57jIbMvHyqNwC7ZE2fR1
m2zjYWWKaNNpiqJy1D4xB16NVWUbKGYOCy+BTfm1KLexmZIpb2Ck9W87x6Ww+lE47viTFmN0qklA
CM4yo8T/AHeJ2yHC8+pGkRJuUD96/eZE58yIYvNzEICMefiBPjFZ9RdPhQw7pVOT6KOcNUTg9BXS
yTx73klivB6h4A9QdWidq2/J7ZRA+bPtkG0pfcT/4Ak07RtLYkIjojYcNYbnSe0S3aim2tjlvOjf
AXOLEVwTo5w987udfR1bdph/Usbb1ipUpgLQ1sbCi2vVIrweaKCcRKNGN5+LwVw9+dFH31B6B3rF
J2PmSpeZOE7dMOMz8kl11yMeRNUHvq7lmXgmE65L+xZyg+ioiOm8V9yyyaExNuAToRGipo4tIS97
tfQhG9C62A/WdNe4iwwsbE8bxvQ1J6rQIITlEkOx0o6pvUoEzPjULEJehjvuD1JXG/qvdxb9ZmRp
hBy4OQdcyj6cN+IIzvt9mdNGfZb01UVZbYlUCqizml3yQ2QNHvgiqq5Ig4aurBQBQs70Ow8KsiJx
xEU6VcFQRwHAM3Wg6Z0Cl287mImQNu6dIDgsCl52g2i/Pzj32j9xEAudq7OMHbyClh1sdD0iBqXQ
LhZf1oX20wOGDI5Oid9m8qLfSMygplmoTxNJ0zKOQm50R9Kr6to+uxMxV0o6sJGFE4Ei2bGQGQru
yA151PLzAYbbJq8xCgivQFRRvzPH6tKJ59jl5IqJk/O3qjdYx7e6ikXDqy0S2ed+PHG6lTRr6qDK
r1PvE+9jnikgNkXGduoZX1zq8VMBaC4bRowHyWwv3tF1OLLObVXMSoAJCRqa0gSGhTPdBowV1/qi
lswsbpRtzyVJbJiXnn/wgDuB85pRYtTgIMCc4BOYtU3e/YX8h3j/e6kEt5Rc8vVMGLhBbW+1CYQd
HZuT2zFXvoogL8Chbm/4/ls41dawepUDIodHDK/0b1dQWfgzBlgwzh03VjMloBAktUKjwkncflDy
ZuXENKHMorV+GQUJjid3WvSOO0HVi3pOYA761NwujpC3XbXX6jgFhoTu4RzghtGKvbrzSH1YKgoT
JaUMCbXTVRpjTLqw9/LrPQAVkOBMyayH4u2zgl9Tr6CO2gmaHnDEXD/tsZnPWKHnnp6MKxGijygz
enblnSblvAxwDQ3Tn/wXCro2HOOxCrw4qnMdWCFutzFh6sesfI9q4H8sTI1oVMRQrV/nudWe3DMK
/Mf8WZN30V5eEsk0AIiaksafwPnKQf/+UJk0MUHt/0lYVHgr71rEYGlb21qEisnivQLf2dbD8PEt
9z0G5kaZdEtWlHViaYiU6noo6JJdJO0Pt1J6gFHweDjZIWwtptQwAD+r2NEyPG4J08v5prHSlzh2
9kD+Rrwbqa1sOEeQaF0+jpWEdzTQOmyhY3F6EUAGKw4e/JZ+3nEV8UjFUu5ImAOMITnk8piJyAo3
7MZ7Z6qkdn9ZdhVWjmPeKlyRGeD7998cXE/vwBezxBOVzKbh4C1rrJA/n6ddBs3PlAhSvKjDWfkU
ATqXlJHHKpGk1tGEiG1/2KrtHKtxaqjHqkPj6UrBpPRhxUSyCxwbbMCGd326yPHiKSqDLVPpeUlD
hCTnxemDQ3jsskdPRb1hy4H1DIXCKgHpE7T98Wc/9kUr6gxlZc8N6N/IhkgQpnFZUY66N2tBqnHJ
lJwCQrPbhM/8QBhkSh7ZlGUQ/tgI3ZPuqImVkGRDf4I9rPSz2ETS3vz5Lj38RCsyJFJ4iiEiq+xV
CTNXYYjf6XCBMW44Fp6ZdfUJxFb8pT1nrg5pdajMnnimyZjkzMh31L/kYiLVnqowwfDp5CU3FB4/
USm5FWPUGq6ujdphVomV3DlpKZwFhmGNorjQuPwTxXEAD+ajIVd6yukHLKD98h5UDagU5W5+unQg
RooF+gmBOMRtjuls5WdVJnu7xiiAZ7vK7prqU182So1c4O7p7KCWOSALlFUJ8SVyvT4Nrj33xoXD
6Rqd3S+gHALpAmCDMyVTFdPMYLJaApSqy6GnC63qc8hPE9/POVgerBDnXpwFWnd6jefupIkVFb+Y
ujPdqR++pMOSyB+gsVGO1uPcoKve47y1VqjsaikMI4nmF2lIW/mna7SkidX+k26IB+64qk0vvnbw
ntuZ27IUv7wXb7yf4xkCqYYSMgBFCfqu0NvRKhZweGNhDWpvB1zEmL0CuN+Oyu3NsTix8BNyaC8d
aZXHoy/THSHp2czus/jHp1eSsYSrX2Rl35khYdloW9RsVaBa0NfxVAIA7srUXezTNpMlxK0FvFn6
k4DmJXOzBUG6V1NcTTLoSDrLLJriQih7AvtQRFvJfX/Noa1ngHvrvdtWZCOWvIzZ+pmHYvBHfJXB
ylmU/qixLO56dieMhzvALIOjOc4Lky5PG3DuB6qf+NrkGt3EIVUaUGuFXUK0f9qDOYqYOl+7Zf13
U+Dllen2zsRNdd4hNXdGyOWRV1iwqhSFI5daDQot3qWNyaGBUmwL18/6DCY7G9sR5W04HFwa+3Jf
pmG7PEQbvIlbuF5Tq6oGlzZXVM97T5sDqmKHW5y/jWkz+n9eCKvE64Xw3IiGLRYyQrxd0OUam9HF
83dNKegOfiP3+fzSlbYqIr1+NnAnPSJYe1AGz074hpAHhK8sz+u2VvilYzJ8fAyW0JG4KYvLy1gs
tLjQ6KFk9UMS8n7LR7jjV3bPJezHG79Vm75pZeVGZEcswEtEd5fYWr3YV854EpF2Rc511c446VSc
LllUh6XLBP4fR+XwfSkuJIrrpzhhGId7HvReeXafzGLHMsipFUtN2kk3Z5q5GgcdEZssVotNRLqN
d+FsTZPTlaiwKwVzUawGojSIMJP+r9OHkouAO1G6MubwoEjw1OED+eIcWCqjaS0sjsPcojWentMN
duW76KHe+G3P5rnhAMCK+IsQ+kMIp3wrD8rp96n3J90dOCMi7jQo9VyxJTQdlj/5p+xdjuehKS2l
VvtjPfRL8fc1Kc0ym/xZ72UnYctoUmpnTpiqk6G762viwnaWQ2/JlppyVMytrAUMhcmooaiMVHPq
Xoj4DKmeonboENrrJTwv9U2FvT6ZL/OUf6UGI2LItMh18wNCVpQhOnuBHhFF5hK09vi4IT6TUCN0
QhR+VCigMX2ippJ+M0gvQjuDZnzPXGzp1gnT/zf5BxhHVq9Oppl/krUlQBQ/g1iZEfOIERtboF/l
JxVriFCaLB0ux558mkIH37+xkLEqXBmHpHh3z7PPKvyQkFp+19sx58KYed0Z8oVhmmJ+wWdlcu9r
Y9PjHtSCb/YuNB8W3sX8RCwaMsyuT7ZxhzRuHkHJxCBmYCbXKn8DEySZP56v+Ycc9Suzp8zRQUIC
x0C0gjX4gbb4Jx/X9lnYtNkIuWhv7xMCWePlMkKAkEZOVPAO+2uZH4V1UXXCrUFfwSCDyI00Ag83
s8JO9tMQ3LhXEgCrbu1x3fb0+A4DzEfQ5mvvlOkyJGl8b8p8GgIsvjPjp5tIWf+9iiiBOIhKWPI4
iS0hQWztBXuPDAlFquusdUVUFpq98fL9GWqiMiiuq+irf2pFU1rVu9XB2ckbJbUTSyTNoms0/haT
JtwhBqOVE4LGdttMUpCTZuWwK7Kivm+7RsgTWNKn6M0BccXFYRa9H6VfNKxmp36uKvVV9Y8UcAJD
gjWD1cy1jl+utbjOkhKvaRxFyRhM2algj0pVh+g6DHGxmH7JgzdqsWcMFV3VZSCHF8LoXJHTTEKt
9BrnQV0gMNUFokEuExs0mRz7KEIX107Zh0AzvBCwWY+lUVmd1b6rBv+D/H2cBf5UmNK/WQGAsrlM
QBwwodzwYI2f1nSsmeAeNcWWrYta+qsla9s5ruYF80N3FJqruoFVRHndoHNiaaxDyHUPvlRvxjBQ
X5nGy4q29sDJ5pvZhkIrPQYfD1fCbw5Fyoi54/EoNMKp3MKHoQOkm6p2MCwwgHXCdIYCKPjbe42F
LfF6DOklWnSVmoe6q6BKLwIUhrFqS63bEQDV+3IB1QKC0BP0UZzvXvWy2Y+hO4CQ4VpHO1le52G5
C8+4gkjeGrwwjC0FW1ckXWyVz+HAnJLVUWR1a5iJlEaEgw5+Yd170tz/nKGDASDd22h08ENqz0mn
KKxL0+kkkgsL+tFtcZwAaB0DyhJKqZtT4pH2rI+D1pS0r0zquJeqL4+0oLnpyVUYecfyfAe5eiTV
RKXqKTrC9EB2X7hDy8mQyD+32KDoHAAc1lz7v3bz0VW60ka7vxJwlztTCSqE27iui9sH8SwbO7fO
BWaRGvWleRQctQ8FfZJLhWtveItV2o3oG2BdCk9z0N7YTFxFQ69ijvcqit7+QSwVG6xzjgPjfeBf
vak+khLvS++UPZ+q4z9WnRebkl2UG/qIRsrMNPEEHBT7zUHwjau8z6PeJ36PyxYFqO3FZFbzvn6c
pn+1bKgvcNVvebuNKyGEpDYovnRHcOJudZQOhiMtKr0DDlvfY1Q6cYhqyLN+TDNMtz78FHiL/WtS
bP7xnopz+6B6QprziQ53yTPoOj0btu35hTdvP6N/cq1HsHP13bHoB79s8r69d0Ae6guJsu8vVAxR
nbVPu/1IqQUDcXEihUCVOP/AIgfV2tDdrfbkISMZFua7255BH+CNqLEev5ejUpjk3NwFApinER7S
nFPDc3Kh3hg0jZg+PhznS2mvaeVU4KaoyXeouJ/VT40RssLYVDGmfUFjoxZvTrBiJmGZlmyskDJv
ECBgbRbrevmpx0bApxQNOrhg0PU7fNJeRNqJ0ZQEHyhsVgRGEwEQ5vNlWyB2WdA9QoKuJbT1401H
1ZvfLx51owR/PFD5yYExL7+/3YCVOITiy5V+E3fTj8FnK1pIXKp5SSLpub7Aw01rJ9obLlsDruvt
BPAx8JQOgjKB87X9BSP0CCF00ockyDsL2HLN0yXaHhY8JsRLCtb5e23NNY2gg0tmJE+mYKhIs+hF
NjBmezQHA3gLLlJwZTbaZD6baYxE8gJMVInPGBAYzEL2zjhFIgUpvxxI4lUygWb9LnSOpgQf5nHh
cbTwiQ2e9IrxMTyRLhpoe13GTQr69TuPcPODgchoIabV4hIhSRbN/n0B2q77VydNx/fDauqf3o8W
CBoZ3IhaxA7X327Mm6KbVmc7hVywavzaSEEKYt7VsIXTUfwv3tV04Hj63XPQcstwTxcjqrqLDl3K
aGBM8olqg3DJyZOS6yyvXHjTZwTMFNdXyZd54xMAUPvyPZY6/K7HtTNZYj2HLvfPB19U2/Zm5uvI
+fAyOon7GfcAe7DX11R+sXLj7RhQHQUg+lSZskPh9m7pnCt9bdF4OQebc32N7J8SB7djmv2XDu46
0/xOlbbzefXwKG+b2N2zBM+3J+PCCOnYh79ualeklCw38BvKFsCoeKyJ9XRVWpUNoOoYkcW8l7hg
R+ht4qtQ6I7464N/WdeKAsR0Knjms/MCWcNzMbSlJhzcLnkGh9cCCusdtDkgW8Pa/lmpDWwfuXjV
WoUXxVa/GcgDuxK57PyrVamybHZUhkcybcDaAaYpbenEqSiX4BaJUOceqiErN9NNKxOVXGzbOAKU
UavGE41Stt+MvzMy005mS+D1LPyo624U/QM/soTWlZJUGK9RPBf4u3aYh9q8z5wnuibruCDZfjPT
7SPN6UPKZ3GOkNS0aPljkrnPWyTF+jtwFEozpTFc59PjX89yGH4MfwEaTZJrJ2mvflWIZeKSW52j
WVj2ZugJy9M5uW3MWhfEuT2YX5m/5N75wL3/I6xx6yv9Ks5SR9ORf7sC2VyQmykiLr8GYWYQIUhC
ZjDa4CilIf2kaSMBuLAvnoPa0D0KyXcu4BVDv/S0hxjhFbOXl42qol4guHgrBjiD58NN7R0ER4w4
My1NDc2D3DfATE5PwMiYIxrOHyB3AjUav/kdPY6Ndng61Kbqj08K/Gh/4GQLvv0q26i3kAFXsbQK
XGqnxDfbty42Z/cmlnDURK82bloE9Oq2O/+E532q1LG5cdMpUJU207v+vEVtZ5d0Qmvl5yYHnETb
b4oUCByGrrqpRAX5voSEwkhW57hGiKtxWQO2f2ULjWVQih/xEXXPZ+noWNGrABIhrzMNXKKiAU83
Xbn/gRmd1kVbgIOhk+2Mvkua4U6d1kEHxW9BuFfwX6TEYhNrzySoIexrRlJabe9A+Gt2dGIyaXt8
7heaAxETJ4ts0LGmo625Hh8jb5aSmgRjQH29rJEKCIoscdhMNMeF/D8LKFSRJiv4478kZ7Hvsydp
w720pmH2/fB+Jy/6MeCfd0gvfzInPkf/eKYcj1YB0CwUuZxW9XDJVDkspmYiLskYwU0L6iz+gM2J
biC693n+LdQ30FHKmLNIX2jcOlOxGfkp/yf8jnzhJTsLvU6jWadn7WsPe//UJaVdYLrq6AQ6rlcv
Bh/+njVYfUhpa7XEMbLztZ89aGyyzNtXnV0Ubia0qvZoYE87mOUKMgyfuDeT6VoNYVvCvZU6gYXx
S1M8VMasRq+rgMtcd7WWAUp30ZzNtpzbb4z9gyT+QIVvmwxqwW/jwNNJuG6ebiEYGI10n7nwGIZY
fIVzgRTrxUX5BNHwtjt60w0c4e6nfpz3+f/HUySbmOooZnJk1vc5Pf/9943sMB2ZR6sduz0prjvI
kfRGTJqL7AZ/DmHaTa7HDv9Qhr6CiqMn/3mt+YVWrK+09Sk98Xqd5t5a4/wOAb5i7q19XPlZadAv
+TRBhYz6BXDLQSnyuZLhWzofVQ8SPGBxr1NQUAadBTx64OoXxBIrDlOalbZXmQgmP53s7CkVqJIl
Gq2VGqoQQDQ0gBwRLM+Sm2fMMIhA0zKoi0HfJsz8DueuV69ssQg5Maadc5pTGeGTdORS4PzUz/Z0
tmOqEqgNkNEoCFM2KsHGMuPVPeMdM8E3QJzEJ+WdT+zB2PDFu9AjngI+HaOGAvoZLfFYzt599QS7
7Rvb+LsftlcSOnHi4+eb6ytM0Dos6Wz2K0Znvt9gszxhtLLUEaTRGT82lvqg1iFxlqeH0MZnqLoJ
7oAD1+uIkMgiCf2CsUd3a4IUQ1pSX9g0Pi1AO7HdiEDq5bJLKPYXpY8bQT86YfolyqgN55jeJ356
cE87XXRgDUoYc0jDP63VulBCRAAJK3CCm4GZMIIjCEhGJQL5ZLrwd+AFG1v5vCVpfDzgLyK7LNoi
TIgGehr23MzeNvcUlh2KapaPO9zeKkvtbEPV/444jQ2uzbSlZFT38VrV92t19DSYxMsbzT9Hpqc+
N9Ig+MFhWzase0PmwYtL57RqMK7bDqpjEnNVoMMMfKN4P5iSWqATx3Y/AuIEbLFOhzlcTiZHAjDS
5GMo4ln1SOu4EbKvxisa+cMVs2vjLndjsoQcBbF5IuxoNFu2nFJa1EldNk+eieECyKY5/c++2ZkO
p63QAWV26LwN+57rgoFxmUADxMD6VZ4BEGTAWPjpAUms6R6V6m/yFtl4nHsqnznU/b316JSo3uKZ
HrRWlV+DPqgl65bdVgXEivZfi9Kj4h+nN0AkjKs9qob8O2PNjDNtATXAVhFCnE3DR/b7t+aPVenG
gRxO54aWyxETpqaY3CBwoVL9m+uYDaa7O5GjDzW+xPRg8qmCpERkbkZg+LmqRd2XekyJpm3ILPvw
2tf2qV1RrjH1AO2pB3fotf6yk2bfsI1iixdiUFS2tveO0xTKQuoYN7F9/e0s2nwSOFZ+0Zo7CUYo
RHvZQH3k7fa6Wq/UkXAkVhnr2rp0F0nCVwqsqDPsYaBDc9G2aIbfoHutlea012Jt3OcxQmak+bJ6
MVhz0b7nkKQ//6BDtgX7/fK2BBSRBkrcZ9ryW8xTs7t/kRqh0WtiMmoipEehn03RsJXKe0KFK9Fs
Amyj2rXFSZVeaTBVUsUHhvLVENw3tqgubb8gg4yoYOiWosiMz9Az8ss36405ew8YVR4Yqg1U41jx
wUq+gRILUXg9CPER0/uTRHn0sWqvM5jMJyhlXy3/uHsT+Z4Hui7Bae40J0xPYpr3Kx+zzp9V0p5A
tQzmjjK/qagt9IEmqDPy3M1lGVQ+1NzMIhl4eKfvDZcvxQsMhMKEFW8s8P6yK5jLgVKGuB54URD3
ImGH34l+sgqS3PZHA/T4SmQjiq1evgneOQOubffT89eyo88MqizzMgwr9Dyai9+GhABUhicAYs6u
5zdSbHPfH/ol0lbjm0r0b7nQS6n01fnkpsXUeNn0peCVfIKgSg/zcLjv35MnqeLh8n97Cs5SZegf
qny8FOW+Bk9kQ3StMXlzztK0UfmR9khNFKo+M1PMQDwp3EPbg8li9oPqzROztBN0WLurlFotElTN
3q0p8Prl+xcuTueT+crkxSNIQqDUPGsk610yKP2gh+J2qPTqyGrzLQO9f9zQlonxaTlNW0sBNEfT
U6HZWgJhNLdmAvfb3uQiUOyP8GmtgO7tbe8Sk5kQ6skn55YYkhix+32fLsKpDW6F+sTuY+Hy7tWo
nDwTtu0Hy4/iXPlHygrHFTNFymN1qF+kFnMebnlJqk0hE3nEEq5d5rtoCB860ecpwjrhP1ZFs+uI
nAlqMYCEYMWbxM6j+hCr7EisPFwlWkqJGoKjC4VaharDLVDf8AbDGgm3986clExdyUIeHBe7ok6/
cuj4na/e4oedAmHgY+st/c/zz9xgJkIpibZN1euJhBqE6uwpyBVvmr2EoKhNecp/JR5E+YYX8gDZ
nqvUgqAZDkkr5z55SBNktqR+OSUsq/2FqU39At3vjpmjvWjrEry0UR2NWilr58QXF1B56BZC37iW
wCtHITItedcpIxuF59TW10csX164Z5Q3V5iLoO8VPkEvUeLArO8wJXWTzcDSZ69JkHXxE8gHZCaG
0oqw1BNVK/+tDY/KRIKXRPghFWJ8/fVeiPg0Q5X8sbg3OIuHwkCo5LBmPku9Dveg+HK1AlXeuGDZ
pGHcquQzOgLtc837l3JbQld6rYJ52t89kRZqLV34vY8JMUcpmgiKOS+dk8cYH/v/BWTxPT4gwdsX
nfA5PBU2R0TIbnTbiL2EzxtxYUWiqJbtn4/4qJsmdieEghW6lWPRo8DafoBoTXjEIFlxASpglbW1
XWne0cv8erTH/AcTi2S4L8/vEMtyPorrbvOGgwtSGCec12IpBwUfQa8AaEi0SqClUhgG2/Phgp32
YtnMdh7fUha4zz8qlE5wrODikgyX6TlAe3M8RTn+bW2Gs8ne8gm0K6BQdnHMgFSOZ3WQ6lg0QGze
SAfVflmmEZ0Y33jlIKuZ18FzPQm/MejogiTw8N6Xn/DC4rGPHibQFqYVPu57mCAVTpJcNlpUjgkw
nApqOq/OHp34XECAyv5dsLPHI+rzZ9aGxzngJP7gIyR2vmKdGv4+Hz2rMeWEbbebPKC1OEbL5LCi
84wMWfZBc66yIbBrKnq40eFRuiOlz0C5Rqf4KiTrJEiOwgGOcYsMoDmrXyvHHIu/2F77p7DiI/4P
UoRGE20Gv2zcyTJuz//GY2CmroY7cBdgwfmxSolH0WmoeQxvHMvdVp1DEpr+18zDjSVXAB3Z5xFd
CrGSFElxoWG6uNvdi/Il16UJcIyO8sCA4G7SYdlJZKj+XcqSPhkWolthwWT3AAZzFcwQ+FneLRr8
45aOXnwqO0+O9xC4na9vvkQaNsg7s2RGZ5CvIrI/2pRLn+kUQAVw5acUl2GBqfBZEwwRE+cPkxRW
+/itVlRR0ripjbNj+zs/bG999mnHGzztUVQGKrvbnlUruD/myuXREIzurYymF+iBCZyY2VNkiEgI
sd39lPd2s7iOf6KQ2EMMcbmAgeHOBOvkgIe5i5A3DDRrJTkEXRT9a4UiPeJl1w/6I6+T/aR6f16G
AxwzSEXexMIa2twnEcsZkUBfGg1II8vEW0dKFvxcSVabvX+dmqAjSYxbFOYfOvsqqGhNjf0BK1xN
8ow1ktXKPdJUd3FrSxOtNamGolPX2YBLHyGutUKs97YnDXRzYXb1hx9ZPG+kzxJpRFOrKuQ6fK3J
/RC3mkDebTTKOqRXJZq7CwIv+ghX/R7TBoBkRALYZBMaTI5SIrBycMSDDBx/vqReZsZaAK+M+bXd
fhkJmjnkJ8DqhmfJnWHJKcsJTDaKkDddl2jU/zb0KmjPWTwiWT7kIJYbkVtDmBhnJyDH01XRabDn
LmwWPNmqBaIwm0O1O8iiD+Zgibp2d5Ty8YfelMxtV/kps+9U4JqhST8FUsSFfz6EBYctkyODezWw
42Ccr+X/xnSpXzZ5j5uox6i5faXYXhBqUCtdeT07K6QHZj6q+Pw8zhLex7pOMUTUackojkAN82Up
At47L8E40O6qciy2pfdiSJiZd7kNo8/rGW68Wo0UQOxAedMzR5DK8Tbpvix0SJQ5l4OKPCJY4L7l
ArAyghfl+uZPixGB0DgAoCHfMSbDqdMLaV9F3P+ysSaTaLWslF7LjY1M2OpETgi0aIUvNlWbIGXb
Fv6cdkWAOi0HdYfAJg5SRJbcuhiCsPamCVLnHQykrb3ODH7zh07PdjqAYdp1hG7LDoAGRBovogDU
2oSXZq8Ubny4ApNznWgfGM65TVHe/SPPSs7nQWF8M1BRLynXqZ9oVkJeortRrKBMXWx+RWrDCGqJ
wWUxwng6K8G4pFyIBQodVYg6mRnR2kpSvXK+kqIX/IXut2jkwdU5JAkeT9TBWOa53JEcAsH85GJu
7OV2AvBNtB9nnotIklpCYsgYPkTdOkaiYWr5CdGpUiLZB2ZLMamF46M50TArPzoUvzpdERdHVPle
urXE5x010CnxoZB0RxrnX6efVz55i6PVJ4TD8n30RjbIQ9/3cr3KaqalHwqXcgPp0yNv5YdNSq73
W3fQJnlOCFcCUJsbz3cIU3hp3MBlD7vLXCIn+E9NRfDPgJcUr65md2lL/0wylK7Um5SjXU+YUtA4
gQDY6cbdHjs9FC3PedVdLxwqzhEl+o5RgZJN4f99AEn9k9/88zGMpuh9I+5wt+K7nEF6WkXTUdes
Oetdz9Vss8dwX9+hZj21T+Cj2/+Lm7+nMttjg/sTWpofYL4OacaDblDBGlumg6TH++Gfl+wUXBHu
EIC4Q6oa8vrDjZE6CcUR1NQNlikWEAPPWwSGAxujpxHOZO1uWt/Xlw25HENJxLqi8B8cXLyAc1i5
izEHYueX/hblK/UDSKEYuz1UeJQFDphxYyhl/nN8DRwfrv8fP7VrEOIhYxfh2icD3OK93RLU0X31
rAVpQnRS5+TPZUIBpIhmTAdm469ZWmxGJwxIkaWUiAZEiE6qUQMpSROZFC6nPmwI2CCL4V9IZQCA
pjHvsmEiNSqnTNxVBDZlhIKJKdbPK3mYxxB6BqRCEV8lAxBwt+eA0dRybld3LDpuJ9NZU6lLdr5W
5yvfLNi95Y+qMA6cmOvZw+NPcxjbaI1fNEpIP3dg9+3e9DHTSpOn1AgfV2ytcIIe4hSIyyy1Le4R
mFPK/kAc8hn4TanXwFZaUW0hjAIeO8grYiuAe8Sydi7Lyzl2anjV03wl0l+e0bbSDOa+w9B/tcMl
jboU6UlLt+q1mxCeDgemrFSINIRSLmAMeZvd2dg+tZyC3f1gBmWZYjQi0+P/WXzn+ap3MmLXl14b
5dZ0NqDZYhcOReVo8xs2c2LxtdMS5TcZ3bdpbpH3k+c/tJpCD5JWarhjU24wlbBvjI8irhwOoe/u
Vkr5p1anKIyTVWFz5w/Y4vS74m70Wq+oiTSxDonFiGqVr8+Rjn7UBCNcHId/R1iQ1Y+GAGIxPlTk
uliPORMYHVjbK7szINVOVU6WYQiQG+7PE7uH65ESP0w61GtG8ziB8JJma2VExTLufngMaWeL6Wfe
7N84yAgOU/13j72PbyWF6Yb+OXIjAJyJOD08fp3abwnpnncQ4wyHKs59ZnfY8kBycYZ3fj5Hkru8
N4Ke6Pm7D0sffrEVARgN8QgvGVvDYDmBpk5etL4HpgtVLXsI+bImpVpBqun6gsJ0he8cZ9ScTii8
n4Hkp4FTC83bDRkb3sDcervz2ksZZnAgN4gl7pOyCK3PeuAy4LtZJ5A34DGQ1qIBWmuuBXcgDtA2
XikfKV5kY2y1KrSKnPMubBPCzXvsc4EEbO2CQHrsSOB0J0PGmlh9LmXBZ+U9DJD3CrXswwmx3CsK
qcycZgfFIadUF24TBpSFDrTX8gDA15Q+gvdEuxr6uCpCoK5Gs7Yp5itQaceubm54+Ojw2YhL5Wn3
20BbK3yCkNGDI2OM2dVeLEoYXGJ2w2v7U709U6F8xJxykWuvT7eqo1d7jVc57QvKakIVM6gOeuKe
pK3rW/KjS4M6MYPjrshji1vSbJ3EWsrI2AO1qaqgxJC7rEG/QGSIQ3E1G0Gxu1su54dG3Ub7bQ8h
dcL43s73yBjSdxZBRCujflN5UhbdPNA0qkaP0IvsGoxqqf2KxtZHz84FtIYq+3H4otULkjFumT++
CwjASk7lN5dEliXK61YbUqPyEN39w9gffCXPOHznn2JVCl3IdkBxbU6vzMeCIINYDwGgaq0rv6QM
fIyfCBkEPW7YIcgqw/qye9VUVQysYFD3EZACBM8foCAGUVWkzV5fY/VHHgL7HngkcSfAAwSCQJqW
Jk5H+CdPa0oDS1ZgqMl4q3/cCKvXD3wwCFI/Tm+0DENj0UKtM0CfdOBpMexBj31p+LIVf84r4ka0
Udt1J2cv9eb8dhth0q0lMArsJMQQxBG7eqDbLXjxdmq7VjB8mGBV76Pt94V0v2amurPh2fGDSLoy
52KG8StwZFKJOUGr6UYEhtmu2ti+4FQyFj/p7IDAUCO5JoBhwAPZ2raBRhpkr8x1J1X9pj419Vmx
eZ6C0yUr14kuQ0oRDYFwrPHzIPvoCuue3/vMLiuU8YJNeho8/7lnTvK1Ys2Uug0XNNRlBXAZJH6S
nn6EN3/rre/+ZZLMLG5sBKXi1ptV3fBkUmWK8ZmR2FOni+oGkrwiqXiW1EA7mLOK47OLQesCHzOH
qPqeylPWLXjlzCEwQoK/1OjmajuVjcU9r3S4hSaEI38yxQAOtve8P3KatEk8bOyFOGBniT1T5dgF
GwuPCaIFdu1YquFTPluRSFMkL9SjQ0fOAfArxXERlBB6J6B0jf1noBlbvXCs5svbiUcgrcErFGih
HmniKBc5U5yxTV2DhVmZmyxvk1ArpkozgKqkyszOQ7tSuDWVHuFjRiV1bzPiMdA9xqGCAawAsnpy
KH1GdP/1P05200b2ZA9sCq/kfSdESuWetm9GEyvvgLRONvBxCeteLYTIRhcNU+ZJHE3h5Y6qqQZP
aoBAQpfrEwVUfhOnOldKDqRu2Z1hj79DDjCZy/oxZqEw1qP8uMGGy/UQU7UJPFCh2Li/paOIMSOm
DUcFnmt9q2Fx1rtTVTB9t61Jwlu96ExH55YgCPA06YIiLfGD9wGL7uA0HoUOHHFw+DRZp12E9HYL
oWj2j+hqLio9hxeH6YouzNy0wd2l8ziOEAOACmU65reHG+x6JebMWNn4uDIGZEnatwAhMoki28SO
upN9tI6//daR1vENyWQgjr17BtGy4HnChwT7Og+/yevnlQiBw8w29ETVgW+BpOsbH4bTiWJT4F6L
unLjSWWqFz/Yfch6XQoFi1Bju7D5sXmSfM9aY4TnUNoCL5ToNLYB/p1NBT6+2J4yZ/dbL94+haoT
XU15ZsaK4/Jl6C8zfgZhAF3bp6RhnNuwJ9A/DGpMJlJtnqZ67e9yVUkgNGHAx1AkbvDojd0lW9Tm
VUSUCkU0t8ykc5364XtEoNZTdqOsTr8tyGPFvXlT+DI9bYF135iEksXcG09e32Uw3lAiOQDqYxBu
Idj8AOSA5hSul/75BU8M0b478576fOI4Q40hNTpGtOJqX6SRi94ODyWWs3VnDbiZ1aeu+3pJ1lab
lbccRLKkCsppdFZlpI4YiLmEL7grwPInnz/o5mrD6UDlz4ckgroqMhBeyPcz18c9SHAGoW/DoEEf
MNbV3lq6kCgXsFDsIYcm8FR2AWeQKgtNh7jFpwLVerEU11YIFqVHnNgjJCayCTJOLh7cDJhfmGrw
fiI1RQDUMt9YbtLO9EVRtz3yF3IrcKYgeTBxuZq7HurYU78qb5ftMMymF13IPlBZzTqCkrwznVXd
0z7qr7dlCZzpu59jLb8mPuCw+qR/gzYeOa8cy2/KZaT08OHNuJUoQbF5njlMWSsrTKcMX1fanOv4
MHPW93Bh8md81OEWyVkEdxfO5h2o5x2qzDivFF+XEOlYqtiSjdHtZh9uGlwLzXax0PFjf9iGlBOL
cmGiKtsKcJcviaME3y5N0QmjRSTd+T1fhBI/2fxmm6C6D84lEvyIWqifGI+m2ik50SOME6h6K0fs
XkPejGDqL/XviTQdmpSiTzkofBXLHWdojtHIKoRPcGu5JF0T6K8PLuGMgfxGPB7NouYoVgLvpm4r
0lQYX0L90QFF2jAg7KEHqbVgGdrmPZe5WdPhXn/q1st9jCBmiZw4EnbJYObizlO/o3ZsxE1EPWKT
w/8pCAfilklbeEoUMXLS5HhcrHy/qQZNHtPe+5NDddFpOsvRZC4HiWX/pm8qy/8LdtAe2d4LlHt+
3TB5/WhaEdeF6sgSQwoeNsKUUbY5OxlNfEDO3KR1pXbhAdaT4Aa2KVkGqgZikm5Sfl9e3Z9ERRwa
p7NMbKlTUFYZbXzK2dLDV4IL8BdRWTcHLRYvFPot4klKY/7xIi1crDf2TPtiXNy3fSDLwPLSL4Gp
F2vMGTNByWuNZm6PcR7OwQ0mEDrjK12kQc9RHBPHp6bx7rfnPbkbc+mlY7zF544z+enIaSSQQ6Gj
TaLwyMgMfbh4NM8USpZ+gtvMonpB2MxDrmpv1sG8Cc0TQSvX4e/zbwzLvba6DPOXBDwO6A0C5uIZ
b/jtoPJ5vXu9HSXYYLk5cZud7rBSLT3LMFz2aru1Juhp1ib6nzl18lmPYnzD9ppqh1ryZBaKZ6CX
vgr0qSA5bLQa3Ytr7Ou/RlX8fD+XBDC1gajHcwfzi6FhRrvBNs4EnICyX0mA6SHpMMjyshi4d6HU
1maW/NHHKwrC1CoMXQSPu87+h2LAIM/OC0tvZ6Kl1LaIJi5nXDfD5oyJ9I0RRWc6lEw4NBQ2EFpm
K6W1yMr34hsK/BAHcBym0HLI9eU0xI8B2gmYvnqRH7pXk1lSaY29rQ/AzpkqIbNhqHIviXL9H8K+
DGC/Ok5DL2l1Zo0ci5P0o8kFbvekfdrxev89udch7JmorUmnZrYvk5mCxTJE29E3PWP6vl3zd+Be
0QUeOsRirbRVBbQT6UYWR5Tu4+u0K69ln+D6sXubY6kl3w5oT6is5m3xCFc9dPUgn5bFS0/ouKtQ
j9bs2CvGeQuxn408sppL7OR2fG9tl4sxw5I74f/QT1N2F3q89K3XoMdTd/0htoh6AQ8ypB+YsM/t
5d9w0/vbOzyRxIV/eAB15LKrxljqS1RKU3SuBA/l4BQmfuk40sNZ5OppdmUYLs0pSauUgnrZGJZS
z1vWaH3yCwdFJuI8Npakcw6Hs+zdWCPZafttQAPQ6f5lHrXYBgIAsPCcYUjLiNiinAltVV7I/niD
jr76Acx+fPmu/dKYktjxP++V75XEX9wft4CMhslhqLyvVWKtxa8yn3suihPXxiFcUaca7b+pVO1M
PALGXM7g13KjXN9ro33z+pxgQs+ydS1+Ea3r3Yi7MbdvL1Ubj8hFi1++yfyGBlxybqLdrbwDdOrK
KVtqm+M8z2iJF0+No8m3XMOVLaQHBTpbkRCRa75ucDmyY2Wy1SKR+xhfFZ+vkC+KZsiitbtQDCr3
YEP8abVnOqHWC4DRxzxKJHqjqYz3krQMsl7QCdFMMeiQ/XSfGq45hbmm+lSbP0zz/u1XyGHUK8ut
dxYjV9OZkXye9vbfDiG2TI1bsqOZFdHo8pS/Sds/Iq5DkK3wIiW5Ztqw5c3KbUtnqrbKMdFx4rdH
FGZu3Q00gOPViMAlv6MoUEsHH+cdkueFOUciJgPMd3iShNYDf/krOSk4ex4fyUOLLve6WxzpCLaJ
FzuJ/pVGsPbAYoI0nNRH78x+GyV98mlStaBL2B2YGotxvEk+kYqnRoAuNNyF7yuiM679hI624M63
Dg7jlPIjZzeK10GipNE0zvqaRZDEBXZohZT+8o+o8NxMpPOufMb5hy+q5RcH2uPVkxNRfyEeBJxw
yOiKfbYO/JGeYmkbRlJs92G8pDHwW2EzRdgwABL/37yYyWq+KjIehoHXoSWj5qJYv0YNMGOUBcWa
KjICp7hFDTYlL1gkcsYOELvF+jGR9mVTpKIvkOJqcAxvZmWq2hYjKdngNBWqezahJKlHRGDWpuTs
UijL66neMy96DRF3VhTLWX18Emej2icAwhfCNmoSuX3XFQh2VBOJN0N4yQgByHKaRqE0IeIIEUDg
jpcof+on8kLWAFOXUhlGsefqvtcLO28i4w/7OPsYr/0lKYCMWfEeW++viwwXumUNrtljnBzy1iQI
jm/tFtH1TbkiVH/rynkavi27iQqQS3BIWfH/SeGj3uxLb/ajRMhTRlSUjuBAv2AdtieKeri8BEyP
18uwtHYwT77HM1Wju80Od8YaBcoldzdliNcffrTptmgcHEfMMz9G13uVvLiZ58qfVQL/MDSpepao
yhzcxGem7jNM2rK9tst2H0POzSMV5zL1g2HgvTQe0St9ak15X6ajSRAwqr49Yjgc//tAqP+G++ta
rCPA9PdNsof0hxfQQOCE7T89IBXWM+QqGSKRVXPebdDqeSFy3cCxG4j0m70LZb80JQnGPnFyTjOS
THoYuedmi+UgE7sab9ZZm5xqzVj4zjx54Ny7ZzB6Dnzg2llJY1nLQQjIyZuoih+LLiq2ledFsAsF
XPZP0UpZwrEZkO3/lOn23mDoDPnyKGc4kerK0nQGVMh9lCDcjVMCRQ+gDis+pJ/lhbez9fqX17fo
r3PRyNJKzhs4GmdvgMEywuoNfc6Z7qOjnkTxMtrQ02Jawr7IKoY4DSVxQBOuSXAyluIijQKUxta6
bPI2aksXTa6cm3tvut9A+Itfwc/sAkXV29XMHwgWtDalkF1xajocSeaBt/Np7oElh5t5hnfxW5PP
cINWQ9yQ7ebY06eUdTc0DQlklXobsqbAIeM5KipW6MXxKe13DhmUxEnOvS/VhmGNjJe/yUhwv6X1
QbRvii8sRrhZuUVi+/Jm001FYUiiWMcxIzMUNKNnP/gF2ahsCUVqs5GvgV8DzqLByZZd+CCxjCNz
DQSEN3sMEC9nqAnHTig4rmF4AlRKScBlAklfdEuKshDGuu0qcV39+V0iaK1PUR4GvrchkQ9LzDtb
WbadfRwi/qhGXKRqjmOBSdiNRl76DuVcRJ6/3w+8UWU7ecIBAu8Yx6t5ereMAlhaOvsUD9bRh2yZ
c7xEPVTfsXdC81NE8ZX9bYJAzfxdX1qACPI4Xk/7ZpWiaBzzfqc7HmI+Ue1dIgcJgoXWVB6rEO0J
Q4WMsODAtZQHFxB7CxqqB974Sg2pLCcbnZQs1j8+Wiy0+UTwgVqOJJKWM3gBCGpcbPvOl1bALRVp
rewYiYCkvkerjsM8ZGc/aNGGvRmeJ25ueGTNolZVgmc622V29/ph6Klosl7slqxHLpfOpZo/d8TN
jWyflSWlTNWFDiVHIFZ9LacLIZ47GRw+OnGv2w1XclJg3GvQLuVlBLRTXI50GP5JcpDbqgOQC4xv
68tif+lEKjitwCjqnT5RukW8zs6PRQlk6Lm1IW4utoKg2yar4CaNUHljZeHsmLVeib6NwX+4M6qG
BVkbKE1xH20b5Tm8OD4byaPUI7eIRMWgBC4DDv5j+ALk4iUqZhJyBilQwDhV/g9qvzJgPS7ioyRD
S7844lwKctoN4cbjABNt6HinUuMyPYGEbdVR/k6x/xXaQsdBrm1Lz5/BJeqSdsuu21D89evbGAfC
LK69KfsHEurgKrJis8HcKxrUvPR0oafE4VrCb5LVJTUUqTyRNVLaPcDqtH9AHiaKN0KhC2ZPz6wc
1Q7nePSmE6fWCpRS6MNw+gbdfr2q+A7JTgMz1GUHTlFZVyR3pps4450gODYNDbGjGl6taE7P7TA7
fmVsclXs/t8y48Xr5ySnWYd7Ui1izrGbo7PbFDvpJ2QlBPMBO9ls0ybQ35s/qsyNdt06S1zaOGED
N0O33DK6o7IStiNNFVWHRAQ+DR/RSuU/JKHhMEgr7LIKJyw+UM3kXr2rahw3B7icA45s4g9GkLGI
w3Hhrd78715uK+oZhAmuHtv9A4+OoP4OEMOrvAAD+hhWULHsy8qKxrQke+MVjHMSAzUcowO5dnGX
eMs92rmLojrBIFjQOF5KpsVLu+F+rR6B/0PJvsMhLhvcfRfSB0YEZVRRKTDS1TsDt37urJqIt5Ib
VgLEC8pH9Mop60iqHuheYXk6+jvK+tzlfLWcLEeUMEIXyEDd8BpYa8AdoP84TsKe1FLZhtvjCJ78
8XqjUj28UnDgJ6lzbLoBQjCT7LGt/jfY+rb0cASR9FRwXGKJMO2tq/xq7PblGAYjHYQXFL/xxHPv
RgOD6fTGr+KSeGvU3XnwmEoVEWidaTKruCE5Addw6C41BrQ7O+xICv5fDx7XkpzyGIXimar7G8qj
HyYUcqEMWTqaY1w/ovwoMn+FoMLUV11aeUOgyD6IDXEOedcqYsNlIS7W+oVfaA4x62u+rIR7qLtt
uvLzNLQBCT8r+cBizhvflGUmMSSwHEPpWGEy3sDjOKCgXWmomrv+qHbGXYSdtuknAmEwF6iC8czS
Uiiz6V4AWvBe+CgMjVHuI5rwHFvIcj3y4MbRNr2Hhk/AQYpa2LsPGx1Ra3r+J8lpl503hhEXAFvV
OuQT/fmH5xcE5FaBqGJwtW11k5srHf9IlD0Dq2nQoFfG3mkY284bHBi/xT6n7OlV0uEGfOyYKnyJ
l9ZSHulEpz8I/nLjLwyLkTBjfywIHnGtrON9MMGb1HJGKKKc3H9UiIdXUUUNkdR9/8pET7+drMZT
Peq5Y9U7dewkOgUO1EZxG+QytfpcmCpHiP7otQ5KQPSA0bmQ7va5qEVd+JX0W//HtBKKnBZTXceG
GibhSncEYyH4dB2bQeiz6dLImoin58AZCgHfDYvc8IePs64E6yFu/E63dWcygoe6vUEkNDGbyIWx
LcISQYwGbMzqKBS2LKO/f11VgntXW0r3wVH+/qqb7V6iL6N91epDpevOkPOUM6JYTNE82hvKVo9d
Uy0pWm0knrYwDkjqEUWM4hUkvF0S6Tp84JxicB+8WvfxXvWebPYHM1EJtbnWTzqEigucAbmFViMo
3JyHb5wJAnu+BjN9Km5VWKB4kx8c8mXFMFzK3Ndq6ru7XbzS65SZOnw6AYoAJJke5LVPxsMmzkaB
W2b2d1Ev4C06WWes7hAwt/wI1Z1+kPwiaMrNWxddtyI81JXclLrBSCLPWJSLya/qz8UV6cXiHLai
+5hUw+y7Lt2YZizbO8gyNEC0OB2fK/HYPNCWqw1ZIsNM/9m4TnlChrN8zIO+YMXeztq2P/0jQqX+
ujaCXGGzI+nP8Eoogz8N06oWC+jN20OmIK3bpaSYuVgehHwuXo+2DuYrp3bo4/qv1CGtljJlk5mW
lvmAL8HZ1zFte+pirSUyf1GtLNTiGuEgCsNJBVlz2iDiZ6B7NBSe5fBtiRK9hd4Dzn/wq02ONH8q
Ql7FiWu0OU1lLx4lxXrv010PmNbJQT3srk0cSMZyR8AxwjLbXySwHZYDF8JtKKsBnJcsaV2l26xV
eqMG4D6M+lGFBnMeob+P1rjOork/awP5Bz1O+Vl3W47vB5NhQgL3m1ZOeCkW/GdMxX6AbsrX6tkt
ek10SSsSH/ys/WqlaeohC5vonch+Hmia8z9hn2o/1bqtjDahqUDJAyntAAg8/9m8DQBUw0gVNssZ
Vg0SQK+t4eJPUw9fHnCTqEkJjmznqP0yTNp7nrv9eGL1ok/02KPw8HZ8xdXlq6VL+fwwCngeDgGC
XKkpK09ZlPNZVT9MlBC0f4E1hspQm99ljbjR6ZKZWKyeoeGCTu0i+LK9/izXouZFgXldfm9jz4g4
Ussf1q3RWhKq5kx1WvVZLrUWbsGP61X4cZZyEMwP0piZgbPQT/I6FnCugTgL2aykT1h+NuLqbX6/
tNwLYom5vEiTHgosDB7KFHq5BQWJwfBTRjSbWCgPX+c45NGiug++lOB94/Lc7dz4lRNnSkvHPluo
LDLhnWAPtgZhdA8LkkK0GbyuW096CPMVt/FTfuJzCiuomADwyKuUihGJ2lrDJ4loL5yXDPcVHfq6
/ks5tT+NWUYrf9kXr+Efj0oEZ4afiJOmRPqWWfX+JQqK1IWAaLKZfKSeeogvJDsm6mLm0Yta106i
j2toJ7ENmYQAWLZmJuT4VGtXQIZQrYJVbz15S6Q3Em4F8Arun52n3Rn0Y0aoNTFc/3DmgAsSnfHQ
lBw2mSS0FGJVGSKBm+LpgDExZBIk/g8fZcrIyHFHgz4qF1jHBgiJxkuYYAhWKxik89rtdNL+cclb
42FZQhskKCW6Is4V4oVzSghMMu7tPKAs9iQDDmuZZ6V9BdsE5NLzcdLbSEJ3BsA8Hxzp2Sf3qLAr
uuEjUKAUOBExlqxc678Jv2AeOG7XeNRxASeOm5VNT45eDeAWJavLTRth0ecMmze/bQQvTmW0eOCG
U0ag1cQv7Q54/4lsVAFndztvIhRMCFQjs/YmU3paiCbZPvpnR4GTwF2/9fCHTFHz/mRLB8fwnVCZ
k1qR2/D27Sh27YnNBcptiSW723K/vLOx2gT8zYd23mS8ZEnTIVBAZ7XrfoPRtdB7B70wb7pT+eTT
tTGbEcl/St/t3/NEDvNagmIF/5Vx1FfYL1yFLTAAxT4THLBoin8jAa6EaJiuH50sXBAVS6T8IqUT
9nuoGeGpU2IgS5a8LL5LLVdyTkRFWnk4v3a8Cc3Vm6bgM3akCamE+G0xRFJVs+z6ods9O3oK7DRq
ttLpq0Fc+iPbBKUOEWSxf9bViDx1RXZyJR1UTSVlf43oD52rWjKV/SsKDbFzWQmytLV8FUR/p8Dv
3Rv5DZuQvtpwXnRi6YP2o6jrF4InkShOhryE40HbzT4gCtN3P11vmogrb0YOHeIrYpKdiEJLhhrV
C7kSpc2xj6mHayNZbr929wsI3AIpht0NL+QNZlGxHunSVFLPIrw7sEPSgbkkWRRDkI7327GXaDeX
Hukvyk6ljWbusNmogb1cYVrcHB8I8k4B8HB1EDguNJkZipo2e8EgNj2vSxBJJT/XWV3JQKtdIKNs
dCHNKa6i4swd/K88MwQm0lBurUOEU107IQJIPF/CnKo5a+J4uN/YtHRTOyKclxLQjxavsG+ArQZd
EQQZCvEuBGZkcCKkSBvndiJfchYS+YK43xVF1HH41o+ObBzirq6udXzsIsHUgiAnESpGOKpcfx60
dBrM5Ihq+a8Q0FnBFZt6ddv+oPXIfEqL9dfNJSO0A5XK1Yz2Yq7GkNuo4RRh+lppdDBF+WgZDtYp
xcmYan6P92tooSJU/m6rKf8b6WC70qWoU+fp7oQ8i2NibxPj3Wa9cvzg/PPYE7t1VT4JRUrM7Svs
3xCn1wV83xsw7LeCBx3ed9RBoFFpBQkLXa2TJyZ/xNjExcVmqKdwm2Rcnwr0UPVvH8rdVbx7K7QF
0BW1vouXnpYY5RkNgHiEFXbat6Xk1Q+4Z+B8hKKdopHZ4ox+1c12LaE+Ac7aZVhVyZbFxsqzeWVO
NjPkaZee0WICbunSvCzh3menl3nuT6zkofdzXYt0JX05/kBR50ngliI+x+Awqe4gc4CZu2SM7NG/
LdPEybRnv8NKqHcvWzQ41NGj4SY0E5TtxF2Q/jP6B/If689ehRzEiaVbuAgpjHyODIpVvxZfU++i
ZqIDqJpv2wXOHR7jJzkZ4snoSItXBuLXgPOR3+03aI3AiXe0wnyKLid5rEo0MI4RVq0Cz9PeHrvP
3Bf9FmlXxEr0pq13LrgcI2lg+RqrbrAFv45AWFbFDry0SkioXs4yTatek2enIjWr9t2eUJ6U9OIM
hKuIpl6ldCCx4aeLj++PerkvzUmIPgsHO1KTUBCS+LrSIYJn/Of+IfAUzFhyHAORcSzkDz7/tiIu
479jtEVhiPJphetiYe1JN8AqrT9sn+Q6snP22PbZ0M/nB5FGtOFggBYvMkGLDhOnGzDm2Fmw0dLO
dJeOAOdtx4mazAop2xzLiFcGUE2mdOGHXtup7mYCqNoCgHns0ByVqHkAYF6yFQh2K12PyFn6aUnR
QEMZEqy75lra3ji4lhIofeWvNOr3+tAnVQlLduOYQjoGiHtyiYup5yNCCeyrzm2n7wJrv8btgNxR
PMxirpuUeN1gBg9cxs82f+WKfdNDVZ1wzsbHfYd0iRDSwSTcjo4UunaLkEaa9YtAo0qaC1p5KYnq
8rEIvNw8torSBNHyco9563BvVzrqgRXOUyM4yJLTS5WwsgwjQfQK1/IvSJIshXk+mTaCClxEfete
ArK1WjndFm83Wq49rbWqTOJcdX1fxBQ6krLTAHOnh4l7RNv9oRmasidn2DujY82GRKk38xlxgftw
TasKkYmvH7Fxe5IyXifYUSHGX5sMrDxx4MTJOMoH6A41CU/lmPhW3uATwqd9I4tBYaxLIeHih4SP
kE2AHr82DNoiVQCY1geXG1czR9V+12khnYMVEcBe16GMVNSH5oiKmL/SLpYokn+6DGcZ6kC8Ch1f
Uq8ivHIgzDFtXj7kPkInMOY8sDecC0BXm4t9WArFUoV3gBp54xCq1AkyKNme6rArks/3vivV3XIR
t7hJ/AQ03OygODdGcFmVORA2kvICL+6k/vg/bbdzf9YMxsVx+uHm/BVF6azk3JNhJWg9651BjsVd
EfMud7YGDqIzMk82on4rrFhFY63SU1Kk6oJ4Nn/DH3K1Zrwc5pE4trekZN8R5gfapFSdj3dnV4Uo
7AHs17j5/ta/jeGkJyHeoEIrj4XGIg49kIKewUsQJBAvLY+ODozy3BSl4Kkn9nNgFRpmMB3RwZrK
ee44MeZ1nBnJx1VpjDwVnH7dJxp2qIlISaX/jSdOy7kDif5emg/iBRW9getZrDRtUV7rG9HyqL9o
46rsfWq8bqcqbU9JvQ88JCCx5v9mGcqecnp1pQqOOW7pir9rvrSCMq9Y+SNEzaBvue7jAB7IGeXL
weEmKBmB0cLOug/J90sJu4Vy0h6GXkiNa3Y5EjFLggoCi1tseREviAxJ52OeMdR1dY4ISZvklv8g
LITmqKrmS4ULbR1go3elI1wCtHjOUZV1eRE1et0WXufkLQCFcqnGgHkw0VKasiVjXqaWEzRzc9cL
jS8Lzhms29Sq7GyBR4JNjoz9Ds5OSaiqRMatEiU0ZOLX76zwzIYXuuNgtBOkyEnQfLiFTZ2iorno
vy3egX/0OU34J9eRZhvhzglyrnDao6UGoZhwn/nd+i1grbHS5OwPQjjVBNweTUgBW8JgwrbRFypL
H5XMM5AYLrFzX40B/MyEiSBlvTt8BOK6uhjPcc7pYaythBpOafbOxX2dBdLcnRONaTSZ7q+TnaGR
0N9NebizH2U92ORsxTUYMHnS0oU049+m8nDLJc+Ngo4m4iLz060LTIPs5AX0FHxDUKwvPqSe7YSW
yngXfFSTpvEAs3ybNIKQRNCkedsOp5Ubsol8gZa5RAVrG2uVXbCYz08lBPs1a+OzMN+8/4qrmnBE
Gde636JPZ0FI462fubfD+qzvHhytL06WFblSlL+Q8IhkwmY4oGEtpobhLv6Sgbrcx39lEYwv53dP
mIo2bIoGViG/Y/6DOaWgHMARDdW/iuNCOUbWyoBpZaM7EJoEg4oKJV/M/1CBFcJBU/87EYUTc9O3
rP2fHKwcmt9i8nJ9FT6cxhKUpr7GgjxllR0WMCJSVTKgEtC7YgFRjOxY2ct+ho9GQ5pawcsiNCKa
a32qdjJRTlMRhqaVNqCMiyyhFkPET+B7gTL1dIBquew142lLfOLkydtO15fWsSjCefmvlcBl4IoV
Frh1yGKM5OnMTPhu1xFSyxbLZOpWNSBwrhGNzuIFe2am8CtGthbaJ16iHrWU2LT/ty3HxNMBuq1L
9f4LsdMrH1GaiKDyN2d8l30JbYht+R748tIXJ61JQRItddnh4chMpc2Ovbtyxd4Wp9UDbQDx6pMl
62wWO95tml2B0xQly5qUZJyeCStqZzU4ERXx1A9WKO8VPbEsGT11S4ldb9lFuvjd5GIwvmfNyill
8FMIGV2dQYxenVWzMa2VPmR1bqwz1bENvG0CVw3uKKzIP0L4dNBBCT+Gae6LWIZy9BAlT9BImsQm
+GHbi/gof7qxXwYH2y+MFF2IKAwJHUQH1c/Tm593G4GTf5idudc0RE7b/IEJP52jj2udir/fj2Hz
taTqRWXeACUSdPwpt+s6wFi9lkBLARva6SdK+L69Y7RSKTn/FOpIyzN3je0qvPy4m6xq9tD/cZVU
gzJX/9KVslX5NM5QfMKBgyFmww8vmmx7gXJ6q75EM63OsV9Dgp3u8mkX62OajLeOeOGN0QVWu8Rq
ZoCIs+C5NyJwyonCiRvrUud1qF8m3Uqeq3QqNavdZIkcMVKi+N1cBhlPvOn8mErdP1fultGOHb1C
Z9Hr99NqD02jDHd0qawoYtYIMNSblUyzV6LX+FtKcbokocTHAAthDu1Tl1fTvt1y7Ovvz5nIIUfl
bD9EKmnbYSOloaz5demu4yB9r/BsGAbQjIxj8O+TluRB4+5huEllj2whRWqLoFDusqSULmauIyqh
5gE7TJTp92X0WNzOym5vUFrdXw4lZxjGVlroA3UO9vJXpCXUZ0WoLoseH6BfXv0C2WTfl9wTmHgg
4dpr7sCkOqrs4+R2Zy+Hbj9CR/nvMNdW0D8zYjp4n+tzGIMz+ZA9hKpJYwVXaCcXjkHRyruzpQ6g
Mc+ELqgiFuX5UJsVRnLoC923NxeCni4R4ue061JWasSNSszyfrBMaWA0MnvSV7Ic5f1SF2aK3Xpm
jVlYyuYIpHVjxXJneWoo5W+tCyoiafQWro5OZ10ZedN2TIJ3eFJb6krypwiZP5XXbcH2/2ZYq3Hj
7c3SgIwH2xeEXBU1SqOAiqhcl5F0Mu5i97ZvpfM/syftv09Gg8weRQX1O07W+cmrt0l+aLd+siX5
4XJQ9DbHPiLMWHwNg2nbkgzosw/7XKBggblLefx50vq0CWC5dj+baB9y3SHnFXu0PPX6qHn6/OV7
SI9p+2apfZA1ACehMZIeTsuFfOcfTq0rjopqwHJXsO6oE2P6f65b74VWqxcwf+dLv8UmmdWkH7jk
ko/vB7MI/folZZ9T0gu7zfcm45+yeRRUFn8E357HVUBOCz2W8EkzFEdDH9uB+L9qUuVc8GE17jXt
2/tnjp/PHYPlGqXCqfQ6na8Xxpse+WI+EgQ/3eGese0ziN77mF0KQSUca2gNqRM7W1YnpDOKsBO7
IVGbwwoAvfLHjQcHSGew2PhDozqiuLEEaVKqxy2SnEI2kJkxTa0anszO1Ltg4MilIVowCj2bZx9/
EClTom1iN/S/XTp40M6hKgaM6myTp4A77nE4U0VpJQDBZ90RU6yXRZwHQYdK26Imi9C7zc3GeUe9
ka9yM0qGdX+rhChvGBa/mN5/xD5LCRR91sn88FeH4YyUF7jc3prok0blSycDPzPMKxuoqD4qGMfS
ADEfL8f/b80jicW2c0rqjdsU75saNnRloLVqXiTZk6Po1LDPACSHKneyocglJZQKiX3eOZ8h1q9b
o0CTcJ9o3uFmWwcxGn8NRfkbJfdgFACnyAi4WqHqKL7klYOzwr9K/9wYZ6O7wLmeRLYh92N2F+Zb
iI+5xXZnRhiLeygCfGTm+4fNrkPAzyNYKTOgRUHoBjecX1e3jg4EloDhHRKQ8X4DFKknabcYbeh/
MGqQBVrFley4/ooIv8hGA/YkZgGZOxMMmegvq5Xwq3j5sjzr8JpMyRj6UhKiPLHEY+ej10qY+V/o
fb3Z97T7hftJFM3uIEfbbsDFKMbKLqPLB951BLCNUgtizA/1EJXQsNyrtauvjK1M5YFlv1sUr1Qb
SsWZVjSLM7VjJ8vft4Fi1fplXOrjdJi/y9ANzPXRMf0VrJqglT39jXtpALVLZAjP1zDqV4VtK5Ti
dgGplcp8hJxuiqiPgJy4cPW/oIsyOJf448OMvX2VNw3iXppEopaUARzLR1CIQ7KWyVefrM12EVe/
qAf9y8qC87J7kGBPgBW0EEV8PPrKeAvfxWlZl+5HScIwtwe0YbEhPsF5rjK2tcA4x4QxQQeAgvze
4kQ9qCg/ef8wXWSAD2JnW6Ft+SWoTucttoTLczdjATl1hvkbfnYtOpv5LBqm1RFv7Pe2wViPtxhS
6BV31cbZuOHZ60XG8EkAbGb23nkKt9uYqD2nRy03fUWbidk9K7zaueIZF4F4XzNHmPmbQr4dbYpd
vlBVEJ3qXN8YT1OGCO5Y8CuhEzAXvU3TET/9RCMrBFWDTLN4HG6pbVRs9ot31J0tOGpCp9j846TH
MLV0IeO6U4E1iYIQFuRptu3qAOE78FevHHx8SGM4bpkQhLmKlMh4gH4Yre8d7X9M46fLD2EX0bKS
tyY6WljNlkTly+TkEbXjo6lIXCHHLXxmzgwD86KrkLyenS3sfwVOpbekPLgvaZdq7R/nA4iG6zGc
kBdI96G6DgmP6ei5o/LwYVs+QSRh8P+dnh7UTEr0Pazh76d0wWm0Vq/VMY+ojtMEnKSyj368WgbW
3wNWjKW59pnr1FQxAMiXtf/U5haC3X/6K9OPXRxvTxuFoA0ppLWPXaxKP0c2+lJwkVp0jIPp3fX7
dglfs9cf3K1SX3lkoD7NkIC6f+jvIwrxmZy5MbErtuFAUCr2q7OdKMql5eAN1nf09WT+tK0FZrkQ
fKAZ0vwMNtK635lOiMxhre9G3xJ/KKR9M+2mNNwJmQLvXmboKJpShy0xnLNkTAgkNEF6xBrVmTc4
jvrmYSU25Jitj4ttze4GFDVk9ttKHVthXLvVzoZzxjVB8XCbQRwTzQ2fNCA4AsVKVSGq993YaFID
bUyT7pXkPlXThbZ+sq+ur2ci7ceh4tU5aqmV83Si+0KM9bZjXT013+1/WOQl7qQS46+1PN5qaZBm
s93a/NxEARQ7Bkczgrub+py32GTDq4kJx1CltJOoogxtHmN0Vs5DA3/xuZtnmKGfuIKbjJx7Q+03
vTOKdD9NQ2okJapTmHYmX4BuupIPPeNVRJeH+SFlB5ykvrA/+boMFXaJYIA/ACX3ajN1Gw62pTTa
OKSpezsXUr5gySllOmXXn3CaZYf72FcqJOLSYYKOh0jVSfQGS9DV/kvAgUgK3JQta4HTDFZ+z8tC
URKE/RVF9t6IOrm2ak9x7Z8N0sZ7dtW+xhT2mds2/HlE/aOqSRC4/SlEcUz00ZZi/b2KFOw2Cj2x
bNOg1Msl7BIb0LYG/Al7foOnEr9J8MqR1Y44DvHJGM78cQr9ONfBIsVqtJhoSg9ii3QTckG4zgX3
1S5IP5vwVCSHqZNw2KGPR1ed9EljZrbvXhCNvim+nttNckO0en9JnWqqOTli24t6qor3n4Cb9aP8
7Cpd4bcuXSGjo5VOa+z5B0Jb43fK/RiIPePwDGtGGP6huV7le6tQfSCWwDGrGP+AUkHBKX8qfnHc
SFJCQFusLitvtk2ieAUZ8DBugWEPVnXJHwFlKJHwLKGxV5isQBE/flv3o3DdSwVdk6rBDbdh5iJP
NcjAM54ifjHhdSlTLbgVvcfF3IvZrvBogVTMti2vG+3+xE66ZTiZeRtVjS61VzJ2RWboc+LJAQni
MZsNnyPhf1t0gFKAAaZSToF+JbRYHglHypsddbdxGB+jAV2QH5vKP6y3TdcFfZYWCIk+cyd31MV/
dk6gctDTA0PtIQTs4SL51G65l2tuhp/3lBzgm/fdhqWxHg0OCQPleTbiu3jlWQqjq0Zb0GhAClzR
uqq7FfqC0FvBYBbRToXqkC8eZ2EvBEKDdRpM8Oyn7ICzKiclWwTXmA4vlrm6eyYZHO4OcbCmq6XW
Xym4rbXshxEiC+oBvEJHzwTCwILHLJzK0uAW/wJhIOn8UVTen2dEGSjYMeQxUd7zO3aYS13CUpX1
iB6CgbQtDyDxWBB5TvAE9XxQOYvCnCFsvkxGBD6hzvQQz057PMm8wqL7jj0dIhLoYN+zQ+Q1z+1v
bJ+gnYx1hrZMRupXnBmQGoDmFPQ4z1sWEHE1tqzeJgL9wS15MhyhsblMVIPdEKvHIgUJQq8yvlKR
IO1kjvEbehHlvdxDZs+m2znVMf0o1OV/nwrnSTi+KsdhdLEktsgA4knEEtHdhR3eQV+ewVs52mk5
+mW5rpOWPscYCTP9nE/a/FM+rUzAJZkxnM2lGLavnwilRdZMQKwISqibCmrNogatKTG7I/kHc1qm
r9pgX5myIQRBe3QozaOIUGqjQFlKfdthk2c27K7HaGs3eDpyX2NE1oG4fnPgDy+zAezGrnRt2uzp
VsedboqvDdqcHjuIkY1CHNAFg2FapeqISjSA3jZTmEP6SQSCliKOJ+YZZ4q3L4uQ3am4Vw6syHYG
HeJ1ybM212SogGDZYKssuZLCxANJso7hrlXsuV403nGiKi9TEFDE5UA/J5BCY+BmpAK3o8DGcIBn
qZ649mmjQMwgsw8eD5CHMGdLW+9LzUCPA8BQv3lQ0w7dzyHlN6Gdp70qp2COl7UrGa0WrVEhIj8K
e+D3hJ4wJLiLIZXGuKbb624HETXywXct/aLoNaGiVzndVm7trk9l9FdCDSc2NHaUBlwHoGOyIYUC
Yo7+t+OyHvgdqdCFz+4pX1qnzW1Ia1wn3s4yMlOOHA2drocVNJJVhGXurdqSKP8fz8wXOqs5WES+
Z47bXAAJqMbR82/3mmWwcf77XiITTsXjM//pJ47YoFinGHP7EQpJoUTOVOkszfMCyAjWMwgXu3d4
rIkr4D/Vx9ZIP0Mp6CM0hbQZOC7sGknTpzO84axQp0LRyekB60vayPnA9/yynDvCThq9LlsKdcyE
Q9oJanjz2b965pKaccGvLVKYtjoUXhCoYqFTP0rOEbgzeeCkjd7mWXyySm+MGOXqUm6DcYmAYjvB
2e9ftyYiBxXF4NErN6MLq4rp8jFkm1Py/lpvy5TKAhEVA94L/ubiChFo5f8Q4Cc9GQ3nMDbthjOL
ciZh89WmvIwv43J2Yc+5bx77ApSi2nL6FlBG+GmAGKsxd0i9bwcC5PahtdIbGJCdRI1+b8IxkKS3
KssawWK87ubzwB05/S8FqYiN+cpjBI2MAd29ZhvqCsJmkHtDQx4Db68l4BNaXdZEuT40up20YC2o
rIioL/wLferswWWPnlT2mo7vbfftRL1NTOhEuGc2fZZEALaVdOmXnL3p1PSYxES0a1W55ge6k0oB
BvhNIjjq7Dx17BlH2ZmhVPQMm4OzCpoTyx7GI1qgYh/6kjJnYn7Nvdmwpyh/Tyhw58uk34mOZxQP
amd6DyFPUd3gtlfkvAqHGANgm7n6RBb0veQl1LSgjGkWp0gvroGaHIu+TRNsfncQ6L/48o4K0EnD
ZT3QOH12q1NWJyvm0+rUPB7pt6TicsGqbNLAKVMSyxp3+R24J9iX1pEdCY/AT8+klJ9mAKF8LuKx
qGjvhZtuHa6u5L7Kxu5UW6gni8tfwRzceWz0AUmWaYRXU+ImtpO8LdAMG/u4g6bA4iMdyYPEdwer
rqKbS4/XVFScvHKQUWoQQaFG1K9jW0G0iC8gRfG1HOfDbwqwkF2GatyrHJBh1apvLsUj9pwdqIXm
KLC9yhhPzdsK/LYJAAG/z22Rx+9QLSTsdpd51KjH6eqSIb1P3J1RnffhFUTFVIcqhB2/sdjqbMBx
LPByDMl9vF7jAQ30/9SUGtG9nZL1lJuIALLXWt0=
`protect end_protected
