-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nT4Wi4unC/EguiyUvoIrMBD7YYW6VjaqnLI97RDup61Y6m+2GHEr1aB7XZKO15eOZhZ2hA0sgeLO
N5KXmcahS+PMnV7rVpzsfRink3RCFiYN1iYWRu6loVOHmjYLBx6qOiVMgI9LyEVhbSheu6r/q+/A
DnNip1vd8VQJZph6QA7yFddSlqfiSFQM1BUS9LtBuzfKCyxz+dNbrMouU+AToOSYHItfm+0Q5vgM
+r3QEm4e5Ui9QYjBOSXoy2Ir+NiSzUvtUbJWF92kEgW+Ux/uvi4iewuj1M8i4IP4rmmnDEG+P/cT
Ro7hFNb2/+7aabzyadF7c7jYgr/NsvKUJ0UoVg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
imlzzwzVHW+6kMhOpWl7HsnK/UtLfXCl2FmTPqpNb222RPjoDA09imd2AyVZlViKKm8E79GTR8lA
0jWhEVi95xlyL/glIJc32vkwSR8IlpU5TRPfUTk1qfLoXImjsJ0w6Z8s1EtjbjD91w6E22TfT4l/
HUk5KUYEZwmCIoCvhEEYjt6WwYm5q4UZ7iUz04ukO02gQviACRxAaQSoAwl9wzFEZl8WrLQdSePh
kt8kSvHD50TYre2PBKKWo+eW4YOGUeXyP5Uf2yuB9GvEsn1Qfpx4/O6QMrjH5m2rER+KqdcILIF0
GZX+OlTxC5gZhi5VSdhzJB2Rl74nUPvPrQkSc3uBaQXpyvslXO5xUsQ4Di9Ds9JBBqJwMoedtint
3TbTs7ZLTq8+NbokGEvtwP1BKSwaGrabSG8U8uXOFF7E0T9aOcd4ctOV/crX7Yfb4sgw8/M0KeQz
ZV5zJxKHnWm8au7YifAjZ3oN3VxOouG0JPZtEfT88a8ZmU4jrRPLR5LtwlO/2/pGVB8rLPqhy9K/
L548pu1lsTtMmrSsAsvILl4yMItmpCIuzVBjkndn8Vkn6iVG7qPocGGcVOgT42s7L/FEVHwiemsM
MFFyYQtl/qdl41iuWzKU9SZocm9XGskwkv/s5ITfypXfbKNApsvKdDarcrELsithZfm6CjGxr76Y
u6oi6w2ux4Ock7MbBOC9quBWkcgBduJpVg5OeCQqAFEdDY/P80xPrxu8y47H/Hg9TjJ19ixSms9+
f8ZLnoGa08jSZz3U3kFp05ASsvFCzJIPIMCSC+HjstXbyygwmk31WVWOBWy/8OLQsgofBv802EDj
tqtNMTJjVaYzYaGW4snrhJuLVG2uckm+suhkfyoCDofufOoMTZQqsBfj159Q0/MCUmQiaaMIlnTg
LJO9mb7DD4ByR25r/fBi113t1s3v9xMVOAYpe4A8QAG/t5vxb/Px3wVLwUkTi2lzljs4bUo6HcOh
1LSUTeEYlBG94fIMCqIu+Rw6/1qqAT5UIFR67TSxHufj2/do5K1l9gdoO8zHZRQo0VceyvakaEv2
R0U75tRpniZQdMBiw1BW8908QT534rVE6IKYO7BAaDUNYOdTkO4c6KnnsCMXY+BCNfAavSm9XLo5
TjAZ3XUAMAZnw0wvRtfKcIslevUymwbq2AbSS+e80tV4ySh1HTp5b6+9wNbiF8wb7nalR1zKsqA1
2g+hipznjXkoRUZr0Tee66faPQ44im/V89BuPj+zSnWwvBrT9xvlAoY96nJRr128aPlfB3tLEfQU
WdISdsSw9v3aQjK53LEfg+bmHEJ9fEo3lJNKfzD7xZJO451j/eHvQ4UdGe7KvclI9kwcCkKF02Uh
lKWLDg/Sq3c64v2BrGBiPRSxdPhZSOPIZ5ZJNPyxygzuMl270Fmn6NUkdMdufYRY1+NqE+KkOhSd
J/CmEdNprmMwc3A2xdyo8/cZfdPnvDw+5nFwb3dv1PVfMH1abjEKcu7I2iEXDu6BAxJT+hD86xKf
iUBN7g0xg/eN8MH9dIKtLj754rabaUcwMDOg7ZMq15H13KLi2/yb9xbfdS8rjgysJbKM0CDOqUko
IrBQhsJweiyt7lATUKtgzMYLvWQrtZjIA5cQUMnoKyNSvrB/VxlHXVpM50L9fqPZIXTR9E9DHxxR
TutQecCOA99kogadc3cPPGnRL/8Pg50CxxZENtTDTAXJE0JxN+N1VWwhW5L+L1/aQ3VAJHyPbtln
v8bfH6yVSyp8twXQfHvERt3yMJbFTsk1CJUnzBZap1jCu+rGJ0yArioGmtgBxFhkt/qAAKWSnHqo
rA5c0Ou87AscA9iLv1jLtmZYHYX4OhyrlX/MpQ60W4Jwp5ysMs64r7h7bfXPLgbT1yKpgaTOdXb2
gcuWA4mRlGQ85OULdaYR15qVmppQDzyiyP87L3KjWeJfPG7NBV5+RNt6kqHTaHVKLFL72t8hnRR1
5vlD8CRTSaru/p3fLiI08rZVbPaT4BV0J9cxf9S06Uu1+pJTFZzBQKSukyUFm8wD70v+FuVdnedW
p/RGO+wMX1slBAUWkrbxHBT7HOBEwrZivCcqVw5lmE9s6DBqokgqoeNA97ke35hxX83uM6JF43pd
sZNPjbRVOVd+ugbpGh6uVaRxAkYCWA0oGRoIJIoO0ZmDwNm1uzWhZX36qID1Y1Pcn+BOTA9rxE1G
SMhMiWY8uShUi1fNQcVnw2gXQqEBmRJsxdAc/tDzx5FI8KTfQMJDaNls47ZfUuXy0aLjCVGNw3lo
W9jBN15GcnNuky4PHioiVVcjEIVIPbbOiobKr/dEl2CQMabodQVoygvo2/EJ6w7YLzOEzp7rDOXz
LRz+/lrlF+Z5uLSzL4oGgf1vZFM/YKCf8ItComUkR/wTzkIYiQMzSHGrHHEBme832rfQ1wmMVcAe
CgBEZViYLF4Slj5unvazJg+kKOsGQPUWmJrIi0IPEt1EzEDxSQigNLL2w4RurU82aWj0vKPdCACJ
pv2YewCQqFzL0NkWYsTHjNPNr1Cx4hGMVCpBno6gY4aIxDAdyX/lvvm978j6ePMAJi+BcSbhXsHQ
jHSRAsjjC2rQsIBv/WU725e3hnvcGpH9lNRjRXJTmwngfGVpv8IeWr/Al+jztY0wWykWVLla9IeX
Eh/QZNU41ohuW9TYhCFrrAbM0xNr9bAhvZQLcPZPX1fndbC2KO6tGH/V9YvwXtd8WSHGiLjIZcDN
dYOcngpQw5F9Y0PKYHXqFIxq4pUj/IhlBC2ddj4czi0ehOhJuCtOsc5XVekJAHgq9wSLPaZgJKUd
7JB37i5G5JaXgEszITgPkyzdHest6USULFC1NIt1oLSR/PXSJoKN0hxDSNSJze7qmyoFLo/2lUQo
AayNR3wE9FiLqLe9ZoMv6w/uj9Ard58v8XMsSf4m79r7l1VHxisq6zV7RN6qHbAnTCBUXJFmOyjF
FlXJ695JsLnkNtce++tpzxqMbsRKpRLuEer/ilCizUa8Mc3UjC82b6/6rvN5pemtQBN+EtPYoW+i
L//vJij0+96vb+2jHtebThAakclOyw1fAbEUR6XGtKvbU6P7apOMPbi0Y+BynRJhSaRAXtjHTx8T
ZSWbzLgZV6E0rQAmv0E7z/AFtYi/6bMC78uG5qfLY4thTCfA+NEDStnO5ObhdIVD8oWBYQpHp9DB
2HX26qs2LCxHgaVZB0iGN1uniTQ6DmXB7pV12zb1BtPqn8WKibHQ2nAoUkErcf1ruWlVbjO7EqaQ
V39tREw3eCQ2n+PuALiwpywTX2DWlIgSoI0cu7vdeZWE1eD2Wl3FF7UJOxIBMzfLnpKxfxzjo6XD
eEJzBD51NAnRVIra+yed/lFu8pVixrXL+tVWJP0RspIqrSQtbnOnRiU28WUtYIEWJXqpwwCerOVf
KW31fpliO73e22DpTGWra+3Lj8fjydJQ8WF/n8DHjsqo5e0dFXss7LPybmMN/bIAkVkg88nx8aJK
/q8+WOkTWN3G4F2EpT8XumaTC6xi7aXpFyJ4KkUgpy3cG3xowDtWyMuFolrTrqOb3JO0Rn6FQd0y
hmaIncfp7PwEPCejAR9d9GJcHsOY5Wzu54O572pkmvkpCkvhgWuxe1Iv2gyTjfzFyP73Qy/TRLpo
SEbf3A2gb6RTQa9FZ8HPa/WRj0fjF2Rsj8ePAogPSkFN3MLZ4C+Y9HgHCnc33ktHa8cUoErmmMav
QKw5eBF4pDwYZce6aHMkF0VgST4LeuLNIUoRd1pu4LO0zEg1r4TZGoiTRGCW+pv8PyD8GWdq5tHM
oBbZfZd0SsXzsXgQMBCep2C73vyg+dUBllItWasXYsUei97jhhTN14KYOfitBaEEpAIe30yJVr8m
4paGpA4Lko3SeL9WWERsW8edpT7cgWEJc7kEamB6T4WQXocpVi+EHl4QXNtu2XwgUB6YZTkEqbUn
3kDX5smoCL1u57AT4hXMyKxhJDeK10PfntNtQQX7urMBHSIE6PJMvADSsNjleH7PK/wShaJfE5ut
U6mSLMRWMuKXjbd4Mhxym08bOgS8DQKFDwk2EJxRIPCDuPD0zQgDMb+i+wRG4xigne1ZU9GZC+zp
SPBv7IYkOInbi9tEIqUdTX25e4s/LYBfmjvCKcaoFz4REV2t+uPqAR8uqIuLRRufCCqoVNcSfxiD
g0QTgFLBWGy97vRoN0a7kXEBhgTMHkx0XrTQMF6g/nuYGjA1QEseBTOuOq3X9Qx06glDr2zZ4it9
jNTnd4zlJSEkOqeSmdmkdOznJFgeJUsADBSFR/zRiMcCCkaAXVgEU31eyQ0F3Hlj5FzVvKB2r7jG
JKGIec+fnzzc/uEGmzG4wLmzJ0P8iPuHa+BLzy2UPtZVQnfrIgLtmB7dSI9wAvLlH0TC64wiZhO2
v/zWN0aL+snw9+Gth8fT79J4x7kgY7KV3zGNTqlm973YObpndIHK9UFZEyFM3WDwldPtb6wrfFHr
iolETqGXRUBZSMpWfQkAzD4ILhBPUrhlGG5tcxTkM7XuhsKOCjbMzzy8GBhpB7dZ+F1BwffQ05++
ajR98bPsQhtRcDYlvpF1ASW0pBa29Li6Gfm30xP+uTyT9fVZOnAPgqyC66bDFqlsqY0dupdVLkWf
d8cjQ9AwnkGJl0M3sm14InZQaGdJR/uwn4xPWvYWdB1OlV19BnE4hrw/WVoIcv1LyGW9F72C8IuX
P1PemL9lAPw7OmSgC4Vu4yO0z5y4NbtpfSIicyzpM9Iyg6XYq5ZfmMWOFBozt1xDCJtpq6N6VLJp
y0CdwdOMatH8Dsp0uDCAnEpaX9BpCz+G6TIv+eePhOG5sA9G0CWmXddItHWPqEWnL/+gKBLOt28s
WdM5IB0h8IAEeQxHwBX6fMO2cTGuMGexqb5aO2zd+qVC9/cNBfPXPbaJNYCf31fo4+jLwgdlr8JJ
oLX3v5QTQzw1IqhxxJHuuCjN7oGT77Ma3ufjlbpGSZuzdnlDg/KX1U148an11yNUp02Isu3P5MT1
Xa4/xgpGeUK8JxkTuxKe2VvsZkLCp07Pj4QQJ/QSYt6GTRu6r3+GBOFdAILnzzBk69Z+6Guttssz
XHoRCirj8Geat3nmHgOGMnFwKfb8lyaMcb07AsIlkNgRqU9gAVYmTIWQzT8s9qxepzwtAuWEvWGG
L+kwq0z3HBG1eWfo/RikqSLYsR+azQ2skgjO6pKYF51fyF0i9kMcdT0dIc6SoHNvUZt9+vot2d5W
zqyd9hlAmryzLJUVpJkTVdsgCTeb6+t8kG2Sfq0AVgNyZChwnzPMOWiOchZFdKcbgjKX9TIC2gDt
LWloIeyT4lcVQjM+AMmzFMfvS/Db2kFhlWgwW0LW1HRsyLVh0UrRH+4TUCnEVvnXnHFG4kz8x3e+
/AIssrnT9qdYrine0CTk6tHs5UvX5mAxwnLNqgRVQBc5VYTM6UJVGWZrsc83UfgGnL1FeF/cTzrZ
d8lAPC4CtE81y/dbvcb1zhHWstZMwOl83WO1Uhum7BBlK6Q8XEa4F5jOFonL0WFkh2xOcWfpq7Pt
l18liabTvr2a3q8NhO+9iOvt480WwI+5faoEuEVXGSixD35+eYV3AfB7pWZvV0FiKpFX713AbJCX
Zl1gi2bd4COBv6BeCWj7SnEqw+4bximqiPAMXRWsoZx2FY73+6u4krpuUtYKVdWltFhK1Z6n/Q27
8kSm3fdzD1JY7wavk7hpHEPfBFzNzYnoqggSkiPi3shVTEhD+VeaBxKsGHYel5/g/AO+mrjarX/X
8HPI9HbCkrQmGVitvRGi7usH+euLVCNNMz/Pefn4758e2ay9m0iFY6R11Kr6zW3w3zfPcb7XtInK
g2PPVBRH3aS37WBjtMCaZHCIzHEB6Iyb2EaHWRBvdZ+xVPLivT1Wvjt8yISNk+GFv9jWca7WxA8f
37+xLTn/b6NhVo+wW0r4nULVjEc0Y7UMcX2b9xalSkW85NlZqLIkG+b7sLWBK8COkXWn0CHckOpU
wOe+Eoc11rtvlcCH+X0iKUsWS7HI2Dk4aU0rmXV0vNZ79IfN+7ftzxjgiPIkdeQ6fi73K0T8a3mp
aAAEil7/pk62zGQkrv9bo8JVezbpvNeS/pJXVU0kZIuieWq/8iGL6dDsKBtuKVWJzA3sYPbySKp9
zahubijPATsZuF8RNnzVy0gOWNV4wJjpM5EeqSVC7qmGhcipK+28RpCBZyWeWspWWbGQCnmRew==
`protect end_protected
