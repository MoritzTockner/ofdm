-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
w8mgBdqGY1hp5ZKy30mB+5dXgrPIuNEpdP1gwJ6WJgaDUIXJoIEF6xn67eKfwnG8jIB4c+LisLsy
Do3icbBsPnQyiJgdz4lR2KY9CQSj3yFjPYHlU5LK4jtkijajWWKU+2ME9pwPLrS+31v3zpUO3neb
Nx3JcYXNRl+5QnJ4D5YfmiLwxacauyuSfIu4ieaFug3lY9JxvRoF6a1zvpVELnRGhkK0Jjc4LdFP
PenYEgaC9jb7s4z6gV2to/2DaLjY8yRK4nt1a5WUHy0VGOIK9LcetJFpnCQMNP51/duaVgwh0GZf
U7i+REoeZOvmoZ0RK282wJ0rBj1UCRvHSFptkQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
1TVMNWzQuxwKxXxl+JraCxGA0XVKlh1kAwsHzMpXMr48L0UNYRFZi26PDP+8lfQ5edNi2a7ZpNvK
q4/ajGQIcl2UD+u241zrOQeJYWBZRxP5SMn0DaZwm8hVCAPTepHvvzeSUp2GoRTC7NZkaOMZPWAM
gYb3q8rVa19EH93m9/GGpKMy+nIXsyuZ9lgiLxFqWml7h4tg2dwlM99zB1FNVLPfq0W/8t/ghr46
EH7pXgS48ggj0ge649S1v0U/u3YAsqwXyiLKVDsGl8PGsMJ23UYhjvSC4/TCx19k44YkAfAdvLKA
s3iF8NlwOst/Azmr2C66rZpIdE2x9ZvLEBy+7oFiiQYEboaXDmw7iRIeXEF88KKoSej5DmCAhf5S
5b14QCjSRRSDo8AOELuPo+JHUCZFLvJoiSLSogvR/aBb6V3Owbl0Mx3PcuX7ZN/EAjD1KC/blG0p
/v1vklIm+vih+T7BriGA6bJ+SUc1+Xtpv+nzD2NDkooduguCLS1pmxk9i1KehBf9ndCahmuft8Db
nSm0X12M/n+yQsUI77aLxy0NovTKVHn8z5/qZlcYanrYyQks2KJ8ewgbeIHM1+gfrbAKyhjDOLS+
Z268Osiy/N3KRwpmp2W3O1Yr5ofbx9oH2OKvnVTVMOrXs0JIgeDGTSIWbtPYX40b2kXLBYGOQIMe
F58gPI/Lfy952cZzcTTgiBcjzgSklZGuEtdap+3Vrt9kq5B+aOXuC03Zy7PtxwsF8DfLcByMjkGD
g2UNe7TgsgZDq27wdwqxIUC4gMwPXQctVoiZl2hM4IndueXJqjrP5lxAe0b0vOQhzWPF7v5qcJne
+jPWZkZwR/MKMenFCsJg2f39KQXTnO0v2npvVRAy8uFSzwrg4uKmy2BeL27feLr0RW1Ygp7Hv1yA
9NKmLsUz23eSfrx1wiRc8dsP20+d85uiLHvUSGrEcQubzeUTbcNNZTSpahQjX2sWZ2kSSDZS5UVP
Zd1T1H4DC5xVyHeBRSQEyAta0uaNrVpJnrJWu9+pHja+xgyRPU7bUG3ieugCohoPJ4Tc48ghpH21
YNTM3YvPIs84bAqHlZ+LfxbDF2EGrzQfAby4SS3GIiZRkTq8oLE+PNv3mDi/ZizjKwQuPcCWOvUk
6BkDe2dXs2JjE3kqSd08RUQoNBOzR0Sp44U0a03frbNaycEHI5zDawrplu3Zl82hK4TLIL1uG+R0
X1D4XpBFmBoSfimgjldCsaiYV9kEx1BYbB48++ytTFuVvpxR5wGdylsE4hq8y/KzCDfBK9HWE8Pc
SCjI0Rvl8j5/enaGj70IGRDjwm2/WKlWb83VQIvC6ZQV3S/yX/fKSii6YqA9CBb7+ziT8PG+U++F
OZF/9bBgl0hBZ8oPEWA1O+SpPOie9yGn3B/OjnDMK7l/9TQPdaTprFnggr8mBZoUqWKb4QBiTbQG
hjjnGLELsrZjmU4O5uEDscW990MLNR0jpfeVmhyNxotfEGF9L8ooqXEw33lHVZSmZe7iWSIRRO7K
ebwA7iWWWkoyLlU3uTeKhn5pz3JHbdpkwDfWyxzoosllPAK2dgk2A4+zseoy2AAiRJQD7a5ASrlt
0vHaFs/Z3jdnByDxOdpIYl0CuPvOgs0GKULDv06crbzpCh3eoXB7+Dyaq0g6sCCim+CPxZLmYGVA
nHsxkgUPFFtjr4jDSAx9qf0uGwqTLI94lx1upWzo3wWW+pPe63SmNYJ4vNOzBWpWwZla/2lCXbJR
T5+HfpcAKCBBpUFeIWTzowZl5zK6ChMrNLV/tDYiKn+Cb8iDpSll591AY2U8Sh1BBANajApjwhPN
Lj0Ra2/R8dk8p7jYY8PcvCr0k4rYxs/yFt8LA7gE5aZdoVjCJrNxN1ji40h0UY82rux1TjpPz0Hg
+eaJ39uh4jw8S6YsFPUSrzsfSkuxgm6VIGpnenyA+iVfNezzpr0Fzb6iSEiZMO9TWt+6o7LsgEG7
d2IfUIGyTJpDAa1GDBQefDxFZfhF6td61EjFl9M1EF+dTRRVu7wMBon/bdHYNRo0RYr3Hif9q1LP
e9xjDUzRYOU3LRTelcjYz4Kq/Z8ilPLnxbKx8mMASeLCAnywDhxBFRsl+HpZblIAZ4CuX7iytK5U
RfEcqwR7Nxx2tmEKFkYNe8xaPNGniYHkOY/ByCA1z2pXffuIF7KsVM+Bju1dyqgo5og4UabH57yj
V2/oJVjO8L+CRqTuF/Z6y7MEtmYlCk/MYaSPzYHjchw2CRsBuXiB9nw9neXPmJ1mIO+goVKEadot
SdOfUtq5AyI9726ISMEOgF81p3LyXqaXKeu+etB5c3zorghs4a69eG/az2soFvDGoeKn8sGpLN4X
kj6fSKX+BAgx8GFfW+6QoQazwwtRgM44I0tAXGH/UwCPUahZabdtC1W1O59p+UREmI7vobwDJeb4
sH6+JijZrKIkJJpKH5e4PTlng34xl+NlnJvIvGFFcqBf2tydUM25HnoTnWKHozWXJClV+dKDkpgT
aw8N0/3+/KzzbqOoY2n5orZ8s9TX6CHqQfnWmkMbLFtrKfHof73iBVAkWZfhUF6CiPE/lVHk0wbS
VTlWyifKyFTXbWPSU9dliD+qKiba4rZomqitQzeO8T6XVgjCdm4ZRqplSyH0uTuLmabd9J9t4cFB
0MMj440ZUujBtvJn+vc7OhWk/UxcTVe5e+9SVugXCemVPB7267fcshxhkd4draYCeF2Xfo/u49fh
N5AIRR4oAJdi1jNVPMstsg/f8XiXxokgALlcbiJFl4MHoYl3dIs0cAVMD5WdzFO5nj79EyXJh5zq
m4I/3uq8aGNyVm01Zcc9oeovaGT5tMqL0IcPZU/tz+AsuDWPAmtU+8GpTrj4+soBFQ+lrpwUKrLr
yFj9S5Sn3akSiUni7ZVrTpPCL7XeI9PIvaK/bTjRGowAWTdLwPa6BnaMx77raUydq7+k7Y9N+Pw3
pyMpOgKjs8ofMTGmFSOsKHAUdR5C0MmjWTdJF+7yzJ19mPgfOIS/Oz0bPI8uogabZjIl15kKlb2V
/WIN4V562uAGI9p/rXxNpx4jtFmm65D+2TywHNA3xZGcxrzUoNLuMRCKZL7jAmug5VvCnKitFwkK
Mpq7zjpnBbpKQvPGe3mr4cVYy5OZXi9aqXaldt9wbyhkZYYMJLQJbsv2OYtEmsSHwzm+oIMKUh3m
tffS/P8JXwleeNWlBxllUIv4Z2nkVGf76QYaQVwk7enu4hIVq4H2EQOwak7n9w051pVISPIRiOcu
tCdK3X1Gltyb++U3O4IrMQ5+/EnqF4lRfWX6JmUsTaFwDO6BtwnYb8un4Jq34lM4fF8E+j2fo1e8
i1QNo9lH7hI7yFs6cJFfFfoeOPjElIiz40JAjoSgGdkw33WWQ0YWPfp3Ix/UQJrIwf1q6miPNNho
YyJCxdvKeR1a2fFcz4lMNVWWDNzqRDKqKqgg+TdNB/CEqRHltyIruSZNX8ZLWBHBxDYZ25Et4jWS
FzjvNezuBHKPnDbuO/x8X+wxIb7KZq9RX0X0xEGf4TR+b68Byklv+wEwkvqeMLhFHVLRBwTTzg6F
6qoJK2ELglbhrBBhZR76wMuyTtc5P3/7jqf2S7t5BJBSqzxWLmZJ/RwitA4r4IH8RSno8wU4VDM4
SCq6tje+Gk1DGIB/BM6TMCgAGCdnV+ZWjelMVEXHYvxz1/9cPx94Ok9IBgS6MFXM6hztgQks1MKv
09zRbQsd4sMPjlZdKxKHjsuJpTBhdS38vzO/V++NnySR0cJdXyy1o0Pb975kYBCDspAEddX+QD+t
CHowRhwoaoQgJ89EvBN6WjjUW6D1+hOqHQYRiEwXuZnzq1psg6/jhzQHCzshzCvLKb31S2er46Xs
1BVxWzOlBCiJyaYN7QHF0N/oPzvyMMpfm/VESUcXbVv9fVsGlJYrKszHsx5002nE2fBqdZ+z8rH6
nzegXSTrKytIcYhD2PAGtzcPs+E2dOVyZgfAIEQTGWCr7Bg3HYNkAbty21Mi9WNTwdQDJ65GOeZx
5kKGoKnHZAiSN081LJvCvIsumNv0vlh5jmlYiRl4DV364n1WUahzT87Du4u6kaWC2BObpDw2jLkT
U0EmmkGWYxgoLDan9QG/XXWm/7RNcklc4W1KHtYFEebgT8zlMfeJ5DpuLQBwwGtqtgOeoOS07cxa
/kwBFTB7E/HO9ClxX/hwrd/EHLMMxqfQ2QaO3G1cVuQPSB4PG0m4p3Tt2xBUr0G2zPCfZCLnDADk
pZDuPfWfuZC1X3tg9KAnMJy5LlvOAKBdZ3vfg1XMHRKWIP1ehemdmiZB33hJmsKEzX4seHK1VKpI
8XsAKgnxCurN93CvzxWbBoLfMfeQId4DnbTT+fnKMML4A8Gm6QnlQFOZfJo+AEzZLbQQCFVsXJNs
Fy50czJGh/C+JSPcwMZvI5rJncR++5ojD3WLCN9QoLU41yD7SvDYU5wHe0ONei86qkF6XWDd7ua1
QkhZG/P2Ad+bU+CYEJWB0/HgJz3RtKO2FaHpk7cp3gAlpfjExJA8LIuYe7UHDNREQVC42kdY6FyM
kTcS7O9o2WpQnIdy+RqvC9R+T1ELNWSB9VdciShQuYFPa0n3PYWhqv855rfyCZpuVkLtaN5ALs61
DzFWQyCfWKiJLz+NCER6lhwLhYKKTuybKTeBiXjDQ+Gq67jMokaZJQmO9+IL+FAY6FN5gWiPQfuX
kv463mauSaiJ5MR8ui8om7DWLpCgVYJV9uuLp6mTjTLwcwDmWxVpWJiT/YjWT/bEiUSXgAVGbiRY
X3/icTrVTbJN7/4QzAr0AFIXphrkWaamsutnnnSVa+Yb/hfbPJX5Clshep/lzAvG1klQ9aa7x7jX
Wyj7swRC1T5ptcgKu8NtRvre/1X8mAAlD59aYFpJmu8hvKHFz2iDxw6IX2b9I6JEOjzFpz1y7H+C
AmjT2BFXLK4ZXwD8lHZhMgWWfZXLR4FS40VatSS4PWnVfNMT/84Cpoun+cP62AIaKI4QFvz6cKNz
ZIQ+N4lmwAWrleYl5K8jFBSqZc47jJfoCoAE5MtRuzmG9CUFCPBV5JbtF1j2oA+QO8mA+Ndk2V6/
AhaLC3Cbbi30NhO0vpnD60lw31+AIG0dpVCgeUfRpT9rkZJ36QLrxnuVmEUwFO3sQeeYqffAiRNB
hEsB9PStY+K78UqYcGpLfSPxioIlg/8Qb0rO64WtlLvt7qiAuMyO3YQBOmKyTkpSnaRvTkq1pZZt
UY4/C1pJhecRiNy1q8G9l3A81/UwEyiAsfbtTTbTNZMFAT9CZftdx7niazZ4REh/QqpJdvk1+NMM
mAfHaYuPptL8s5K+y4uKCWm912KNfRG4bB8lFUMxImcn8l7PwjtbQKi1dN8rs9Jy82uCN5gjW7J2
6owmCRSB+dA+i47IKMKg/1XIZTodya9Ux/OAGiAMiPC4XuAlxjbVBGqKzRXr2ECqx4V9CRPHkUOO
nia4lCZgFO0LsolcOPAyxkHoyfdFXE3qE0cEyYRM1fH1iZGpOyheRyBhpJmaLPy5o6YoB/Nnvo5J
QnI8q8Ve9EvYu5OsQybDpIPcQ+4zfZmHfrgF2wU01mnCTKm0JZWqj0sd6BHJJSWOgrvIF2jJgpMk
irBZKl9K3JRdRRBKE2ZNu1t37WYifeEjAmKtH6FDzqHIBhXXTJFxcKYQsWP/UyrjC/nEkAX+6Guh
nPE8UPYDiNDT+cC5YxeV3WY6ajFGz7apKF9KA1Mo463v9wfeinvp+ybIKlZvkjChKmxK/WTHHw9l
ZI44+7PugX6N5Ue4eRm+2PM8BTId0b5v1p0+dPm283KPyLEwpEtVKQZN6YfVTmz7/i0AnQtOU9Pn
Ozogrg3xgwuh85Ug0OJDEWcMj3wKRMbJYZEGX7amtPabI4ZmD/ihg7pCJp9Uxdt+QY2pJ49WsUUW
ZR9pjHsUAmMK+Ix58xe0jt8MKoQE2YI9xxM6Z/GMe8V5Jc9HFWmGcLNMT1R8gEPXpamP735SoPGS
79szTK5wIA70ul8soX2zWsQt4bV6Ka54kK35Y6lmCvGygZ+UExZgEl2XB21D/cCiWuYdkW9RDKw9
CpCDJArkH6v3aubI3+bzR6MjSHL3U/mrXcYI0r6Hy+CTf/qhFzeMc5zuW1nLoTzYXAvIq3b+xtfT
Zjj0MVwioUBhJ0Ng+ESyv05ZwU+7NWfH7sPVX3+aAnV6Kcs7UmfYPghzoKfvVi9rEjvCeSvXl+Vh
izt9gB71FJqsxTBm/Iwv5J1HGoohdDMm2ILF2WmnGIRmiyOosariljrfXIoxgOv+WAChECz8Am1b
HcQXzVKywHhLdgmvLdu+JV9yUtjSIKQpXaP1+Hve5Gq0lvQ7FuSuVWW4hECOSaNx9pLNzxz46a7R
Ih2Si6BiKulwRulMrx5UubEHWw19r4B4+xEJ/nvmxic5bxg9sZ+MhkCs7TyAZHZzFgZ73kLkTx9k
wGjjSCcEgjGRbK6Dtgz0hBAL6gZwZGYiZnGTLZPZJMHHPKramloSXJX1EpoFZrRsKIxPZ/5XnXUu
DWTIG9b3elsprb/8wD6HI2ikZPJrGdadMJKqN589EXz5iGkYxv0CdFcdeZgr8o769o+MjrrdP1Hu
jwzF1sAjIsrYK9uUs4UvesKWCdk/HZXJCM4lffc+dcl/2gzkKmeU0d2XDt4+TvPFa3pqyvYxpWYd
kEBRieKFK/P620ZxtcK/RAu4ghAHVuwrRX5Z/Wly9h4FjMDzKK1T8Hv+ikpbk2zPSWSEx2g4p+77
pDDt2JjWRmzV4ZrJZ8/0tBiXV7Uzfs0YTXuoXv+Z9vsk6rYFNdRj2s2fn9YEK+C25QPs/adeKZk9
k77biddNyEOZGt9Q/C4802XlxsefKJHy6yD6se55Jdzv/x5Kl7JO7gnJjcR+kEzGRQzyj+rouGhy
GPobC750w3o4P7FDwislTN9FjOz7xznDMNgbfPsF81Js54eQWDtynfxeWowS/k+F7Vwkm/x8oPia
9movbJT17x0USun6tivwwDDpP1HygzDKODNdTUadXg8+Gb8IQHvd6QqeV1zp0cND0HAS9hrO67Lf
JXZ+SJn30iyQSmPhjBkutyITAk6CJc8hsWxtxO5pM4yXDhzOIsNGNIFuCwMbSRUA5zWaQc08hyn3
YYrCIj9tRvAfSAkFuDd/QalOF+yVVvZ3p7QhFx2q25PGVLqzWVqKNkfM4Lq6OJKYL7HrjHlbD+Lm
kh8F8lN2iRZakK/ZK3NDqfhNjwO8cHvfAkq4GEuoTGZOl0fEm0S79visTEBO1hqP9rYYNhi7AX/s
wl5hxqTApUNpyVo5e/Z5vBav2S3CNUSi0VykqO/pTVSGZcSqiwvRluVH9mxlq/wYQ2d+GWt29Hmh
4PHWUAQq/A676DnGOO52rxtOgfINWX/7B/6TmRKdbx7WbQJXjy9+AIj5G+Nhn1h9GnHP3YPl1Ujl
5Fpunx4jI0EpTIfeF+1vC8l5IhdLnLs6iMdfh3VcumEp6vVAJkz6NOyk0ne7EkzcFdynC1LlEJ2+
zNC6frsRONL3OSvExJJdiboFJ5OwNGU/KZ/zY9ObI3K+Qxt0/VUqq09lX+UZOBjimhcmw0C1iIj0
EkZRL5RCwrUre3/nTWZFIxxq6IEc2AQJDCjT2uqElA4Bb7+2nnJ0V5lmzyNVEx8EqSL9tjCHlS6U
+q38KrAki+x4S6sZIiqul73wXOeSqVVmFlzMxk4xZxVRioTo8Xw6vSqhKkztMfczSsyKIg9sycoq
K/aCMbj1OcEbqCi2ZVjrF1XcgN3bD9464vZ7XNdI8JC7KZ5xSrWau+zhICe/lcyLbr7V7KzO4Tfz
f+1lUgRt7ao4vMOxndA04lSDCxViIyWfuigVg8f9lUxLdFgTAp31aBRg6LRSjwVq+8YE2Z2gYCcs
rYWe3xM9eCfJqSEj+WRqrqdYf4FMMUem9gHZrWEENnODxF2MBVJB38KqvYGGPiQ3jiaK3awcZMHl
PD8L+txVuA9yJkNz4R5520Bi0lcQ1LoQzKbkBOGkyT8hscQydBXf87w+k1OSGbPNvipxyyXO1HfU
l6vkL1GBQ56dZtLfeO7ri2VnHnHmwCSFdnJRDfoiiX4rn5pTdHRZ3MyH5o9aj8YC9YYD5qEgMWIm
9CdmHbn2vnHtdMnNGZ8q3qu0v1XZLJbK7U/I++u31Rl9YXscXpV9ZuK+hRpGw0nEmvsJ1rMiG8+k
i9e60+3UADFPOWXzJdSeBW9JAS4q423nprQ98/5I8iqwuK6pLa8nOUIW7RNMVvfnf9iX1nWNKJyG
TOrvTLLlHEWhnfuspwBkh33OaO7veoTcPQ5KKtD8fN/GSIqulaVIljp69bUpTgqGEtptAd/1zu6o
WAmMk2diBytmdOASeOZSsiBal8SgIsc9qPo9S8HOuxTMWVZjGFpj0Qr+r6Dut2fsc3S95CeNDpLJ
RKCdFGgSktNeDdXvrcSVrN0S79mn3f8qTaxI+cUHlfJdZOmc5wgFS/1WcDgz+fnXLhraoUoNsbeb
b9CX2rnkfov23Or+fBjzZLT0JqG63JVxepI/hiIG5sjhD4NdGR3Ou8LNQACNKkRGapc+d0Bbb4DM
pJDa7F8tas27uVxYGuvOuv5wW/GOy128nbXOc/kV/WldWJasRxxzGbayKGD2NxO1UK8XAeNOgezQ
KyZMBnABOnIrmG3hDa4AD/t+HRpuVk/+3BboSdSPpNZu1AwZ2SA0EGXGbyfzI8QqvIRckMCTFruE
RTbzHUloEHt0MLDcKS4JUtXx+BrjEONyjLGZTuw1qLP+fBvuhDoqLgtD6BxWbUprpz4jGM6JKAcu
1MWxuxZz30F2uq0gSm/ye8qtz6BnmkCg2xIP9hz8KQPwkE9Tp99eOxEeIffKztzNq47xm2W0KKmm
vT0yuFw6pFj7fi0lioEj/29DY2TS9BNvQorh30rni/xJs1v1ea0PWZTrPraOF4e+paRUu63Nm30N
ozNSmhDQfYV8kxJRn+wPrR6RWz8GFpEZVx3QCr/uGfRHMu23cxnVqTsFfB9MNgSU0dEc10Edlin3
c6K8zOjYSeLBDm4Qz3B3fgVph6RBkIi0OeMeMPLZxH9FCQWfSnHKrRbtRQnPKAzbk7JOn3NBV/ra
WbotwiDY6fvtFkgv+W9IlFgXgzuhwA0lXhLU2hPiQ0EAyRBd2SoyySuE6lF0xgNiajjBk8xR7sx5
AE03z8HMZZyhWaKfYbdpg1mkCoSKe/I5zDvsYecyZKO4APPv5klNxelQ5LOXfngcMVr7H7iQTIQn
9oOsi63XZl8OD/GyWt74Pj9wiogXx9WRSNEhnQGJ/S5xrBpm5lAxHz+/nhI4DbFmhfmveWU4EDxC
EoPeD8Adh7mMuEB7jh1g277of+8v0QBHqb4MQQI2Ohk4znyVsS8ViNxgnr46kAYkp79TJiJPL91V
frqCvEsb4GTo2vVtoUOKuoDAfQBeUuX/kUHCOK4BJmFFZWPK7+2ekTvNpQe0SyijXS+VHZyDKock
9+L1mZ0wKR/kx7BvvialqhbODIQAxpS16vo2wELGNY27dnmlVIZqsP55H8tFh7bN41yEOW30HOJF
jGaE3yzncZlRa3BqnY96av803DQY51tL8SBUDRuRHX0QrWEn8+rhczjh72sUwcgQ7sQrGMoc1kNQ
q17n7IdisMAPnspoV2wUJyoirwu6KgVWl9+lTLIEhSlzL4/IqcjRpDcDGkcU7gISbpz125DUEoct
5cpY/AJhi4dh39nWDoPIW0zTkgHEtvI69O8fst+D6tw5i5427GOCzJ4818yd+qD1Zh5c616DmNLf
2ocFuET9UvxKvNphZYVUvjDc6HmPKTU0ACowsKQolrcdNI8HcXRmUHODMqLH780GJk5p6eo+MAdr
D5B1GLe38MWPlEmX1+O5DKdfztoVE6i6myTXJQ+Qvu2hS8oMn/Easc9cTaAQgqT2ZqlC2DgH5Ljt
kfL/pb+mmpID6qCo8gTx6//Q8sOhlV6IhsXLR4ZkQ9aMW2liDhwms/s+pUFII3DHxY+a5Y89PBzH
uP/clpaiX3wH3PlFfPLgoV2//AgL1XefCr7S4eMUOl88uAyMWzrwyZgGw+JjM7zAOl/BOADOCLXL
UDGIK3yBErefYJGKFNq2tnhKtPSEaj+1HM/6QLjdOcc+G+rIoQCthQSdzdzYXH7zgNjCPkaGVm1v
Kmuk3Cm+ZdA4J6gNivCishn5XOjhb/g5FDVgSMGxYP/mEJybFjHQZP4xj4PpWP7Rpg/0M9xcNuT2
fOXXtjmNXPTZtB+O0h7FHSrCi/npZhPfTajx6hsoYjAY8+kweXhL2kRa9Jd1Dz/8RreebG3EE9F6
3Px0GyCQ93Supo2fvRaE8k6PN7oUJxBYAnrHM86nIvDjEdhQtGwJuNh3B589JrN8ZUlp65VGA2lQ
e56FBmbMZdcuMM9ADGmJjDWjImZCYjg/6CKZhlZav1qKSyl93yWVwKOKUbvvhuXFVCDMCFJOeE49
ahZwzNrb2Qql7Mk2iTSK/ulKupD1CFb5gZpPrLOECsyFHyAnR+/oj6KKHd3JXGfdfOuI85rSmFC2
u6q91hVV6qQORXx5vugwLvf3eO+xmDW9futYOBsaezayW15BLm9GW1Hurb4LOgbK1sbGhx1btHZi
Did5b8mnft4yddO4V/swUPAKzteverAIKF06ogW6BOp5UnIn2NuLiempwLTqqBJGdHHajtNtNvUs
2j1yIYDDV4D9YnZnbx+iL0TkHUz8U3dparc32NHIZpDCqOGmLAf/XJnKEfoA/w1KUtS/HflzKEFZ
6yzaRmCPFD3WXtPZDR2MUZYlqV+KcbjpEdu6JKhIFtzKOICThCJfAOlOuIaWEmTmw1AQnMmAaJyV
InKF3+o4ptlAq1xyFxIHt6edgQKhNH8sua3WHjLZtSOjvB1dm1DHDfA2oE/m7F66zP42FC9B6sLQ
DfgJb7y7r/DaZ/iWMKv47DouxCgJGu5+dEjvVDOEgbrzZRXcl/6SoVRv9mPrGZmPDkIFYcFqOM3q
rR72bXQiuNsqLn6n8YTxuzJ9gbFcA6T7hrOSP/2kOyl/g4P3sregsOa7DJbbAufEmZC8rI68IvN/
ktfWvaP7zUC9kVat7PqsepCXhu3gCIHaspYAvtTJDnpXJpDT+bBtFD3KIl6s4oFOlwMpYlUgmJiU
x6buIsIZNEtSNgMz15tAIlAblYUzt985nUx7CoVvMuocs+nu/ZbKPpeYCypvg/BlPFaEOa5xIFyW
xs1L62S8jbhrYTK6HWznAQIPn6QgAoZehYlfGo51UT0AI2H5EyY8ZarTC3AE82slVvQQCay5tKQG
KTTky9v1SXdRQUdh12vNrEM7Esk/rOIcdXckv7sP1y1JczoxgWRxhtipmwVNlB0rJgrZkoKmZ1m1
TtFMBDdQ5qqyVAy+K4MFgs/haH++aLfZzkdV5lHT7n8YFtu0QCej+UvJ/exiqjM5IKOCQy3HUBIR
aTd9oSimktJF7pX/jSF21+7kqatdpMr3ylozKCPpKlTrWcsjXEhzm5AxwRS+cWnIem7SHlB46tho
t4vrn66MjUrfr2auFHKjCXWOnfsmbzFzAzJsgbXpiOwzmEk/DRY4w0gODQXYvup5lxCQLdfqZaEU
RLZLnasONLx4TyY2lqxshcp02Miz3wt5ev/1WhhcVLkDE2CBEz6xBT5bRigicclK3ulHHiSem8kn
cMSaH3gXAbrEhyQiUKuvKN64UPfIUBq1qlkn+c3Bf6PL+gd0L5Km3e+Ya5iJDrP2U1k58KBlxfWO
Xr48gUFg5n0cNa9zM+Wyfjydqj7iMNfKNWBFgjkR1UT63KTQ/M8umu2dCx1jAAksw+KV8N7AsUzw
9JzHz6I1ITCLuiRZuCI/5O7lSoa9yjjeBcPhJuPQFW7HgAjv6pkqycycAGgMle4pMS9sV4jvt7Hj
Dg7Q9xF+5cXW+fGz7jC6iZSiur9RHv5O5qo0UshjO3OdDk/awOS25560EMydyG9R6KBbhV1+KI8K
b4RCOzgPF1dBatTNZshqIzCKNZHChWAu0SGHDHlJ7dzvEa3vdsosTSajQKCTsujolbk15sWl/YdB
R+kIaANyJpBFCoSlXlZbhy1d86NVDEGlIKmO6dMqfgryp2Hj3ECuWpS3JP4pdLx5N7uj6jADf8Ej
4YDLCHhb4GmaswGJdy9Ggp/XxqWWQtE/eGiuwMNAjQOYXjPzqfMP347dqOkNcXoQeqWKJ+eCcPxO
O97kiCIRg3s05DsKuHdFgaKaKZQee/8fl8Hjk6Y90gnH0VQA1UpRPm+MO+jL38O5fY7FoSNe5i3x
UHFpulttQFZlzZVhmHwZNhcUvDbbS7E4T993Y9pnFWUVHRAPdiCbCIIMK9kmA5cfOevB78aI/XYn
zZnoAsoqr/JNNwnVC+zIB7akH8tdHurVuv+hPsD9vhNemJtFdg8dY47jXDoHFL3h2hgihxHX7Tf7
cMnHfcGwXgISKy7E9D5FaNlfw529KYMYfP9/hNQ0VmtwsiteFlrv5F/PGImgko/mQ0zMYdb+y/96
hzVC5Gb1huS9Pqegg1dGiMt0IpnppkzGB2ny624glvHi5z//yZeQIodAhbPT2qvAAmg7Kiv4Cobw
R4hnVsMhXOFENt0fhl+uG59vaCC9ibRLpvbhwGxgcS/M1EpWL9KdOGK79izHEMG1sLWk057vm1Mw
61AVMsMW416mcLHzyLlrPdO7duVT2DYPcLi6yWa7FnlZUQapCpCyKRHRZf092dyHpsmHtgY16b+Y
Ue2rupsu4SRmpgAaUWVAqzsPiyPmCRovCaMNo5oPCHl18qUIJG5Ldh2UISH34NGFNKGrCJqmZ+3y
WWLE0CHqlzvw2PqAK0Jw5y87+mqaG/7zInbzN2RjATQZ2OPiYjd64suWUQw4SXfxcPymeXCLja9f
8W3bS8VofkonKHfYfjBCIEM6XQLk+M7BVGSJdrvX5l3V3EYxvKz7rAJaHPmQv9IByVGCcSmNy5B/
qm+vgzil967U65LEMJjmt68AWcWg81DIjEQiHKJSs2QqBDcIrMmRPp+VGbjf2tet6pqWTgQppg2Y
3SPeQD//2wq2fbAurynP07P77P/FeajmeR/XUMBqYnrIroFnthABNbiXqu7+uu7larXUznPmqGZP
zt+Nt8tfvOc+6hJ4XE8jOA4cYmTcnGQdGhEo20ZeepQ84IcmyCDHNrr6UReor9eqYtBBlgWzd5lK
n/eUXiTkUxZsHCm4QHG4tSVv/XpSS65q0zC3GcCyV3+3tmj8JjL2V1ZRPV0S0jxRrrcCFxInj2r3
SGgyn+jzEPCTPzJG/FqOL8KVMgJT+MKaAQA5Mqlggc8q2t1hkkAxTyBot38oZjOIq0doUjwfHvBT
Sp2hcDhh2tysrJAniU0y2IzixGsqMfevrEjrBafSaNLuedM3hEPrsJLasF063wMSqQQNsyzEWmJO
euZkw2tK5XduAkrJtFhPQatpYrFCwwHEA63tfgQxwkHN4t6rxmLZb1fH3PJCJF2N+IeUdmRNaPfv
3xaULMJnOnhMet4HB7QcF1VrwyXdvPX85aEvYdcfLGn9OMOmgL6DdzdOWGZSbP19uS2pIY7nZTwY
8r/UhIxrutQgVkhMwwSDSTdLlbrFlSuKkifGvtwC+RyYQlUbgszDP2Dt+g4P8zqZ4cleyP43GO85
DreYavTfPSITXS5qOZ1WGJSilG2HZDRnf/YmHW4N4BipMpBUKXI3z95nNfRrzhkRwOCroJspdUp5
L92BboPaS+Kc7ko+0Ers43MsX8ajIvjFi5GzcwEZlyh0TpZw7NWvvJgfSZoO9Mz05EdeMfeJqo6a
ORappziQpFC9VVIMneTN3m1UfsvwfFrUeX+H9q8mYXTkLMnXpEuNQtsgUkaA6mimoNWQ60qSchzZ
d3byvBVwhDgeLooqiPcFlLQyRZXcjclxCM/eX6wJPf2TRPwTXIWeRL4sBjqnHWnm9W6lTKXOMI2i
7OUJ4/pazI02SAZ19w3fCrtEIsTZsp5yShbK2YFjwILxGB5MsnJEa2iboEpoUa1CwN++58Y62F59
UP9jACYc79FSsrpyZ40U9zensi8xI86oqfQKcBN3AjkqE7PNfyAj/ILk6eeZRVQeQIsaQtPAxfQ4
/tAOxbdQfub+8gRz0OnEx7qK/QQGuTpZRtSNv9ynWnfgGgp12uTX4A2nH7lQzVApe9xBm/s7p8Wh
BGXZ+/BdbknsMT7P0v8LNoD+3OhtXxfhdLst8fN1n4nBw7JuJklUBruXEZ5f615h0Uh9jp73RxlC
cTlD8Rtlfb2P15SbtVwJiopzQ943pVSSnVu7mjRO1E52VW1t3Ejemb6O6ZZ3qVIrZpyxGXT/StF4
vAP9le7UwIisDVMDklcog+0j25GgZ5tJax132Dlh0VH76YCu6A7wm8Z3ROBo4WJaRgwBr9WU1SFW
RrUkpHBgzTaNr0c4mqwRqB7FV/yHrlx3DkwaCd/jiOYmpN8XqvQ7M5DkMN1zTQoW5gYj20dvpuYr
E8CQQMRqSM5YCvCG+lYAnO7B5gGYzqq+Rt6jgiJ+6UKy1NkarjoksuBaIHWs5wPMQ/PoMag1Fs3E
/1Z6Zeei7EJL8bNftdR8/VnIby1I7R7z2G2Kyh3xUxdV6M3ArxOWkjOWYsEY7ns9hs1sMrF+RFOA
0nQ87HcwjoB8SObwz2ZtofD0gFwKsmQhc5ucDJsQdPtZGWoagALLxXwmopHHYnKji5Kwiy64DWoJ
2lP9eMWUF4/uZUbiE+XKn5xH4ry6UtrLJLX3omg8KxTu/S3hfcQeDctvgbKVh0l3tVQcXjOm7d5U
06PWaklQNsFQtJ0bXGfg/HnwqjOiAwWBTFne1NKRUK7c2k8p+uiSI+il7uvlNm3L/t+7haxr6XrX
ooj2KPmuGSiNq6IpGPU2zkJtYiuVLnhv8YzJexOnZpDD8wzGhcj92u7GuT0yedQnl09nqEwZ0SkT
PC4C1FgCybhwiYI4aYjGU20S6oq3ZWxkRZvalPFHtCL4aBPIlzwHB+fDxqDzvGg/LSn1eMPJnzk3
VdMszMEmMgIJmNsOwQmIsw58KC0BJGnnb5rAyfzlMsAFMqeATxOaxcjPFWjkTvMaYOs6kT9MIhnl
3/J40epU8Bda2hoGkOOsngKEnXRYmO+h/UAOPSzwCYwDBjLFbK2SGY8ccd50+VD327yYFnG4aVyh
UjN4eNzcceXnMTqEYtsQN2Cf0boeVFD7aZ/a+kKAaDwlKwoz1O51e437Wzq2nZrKv1I1AaN/IJk7
JMqIzeH7sOzhstbwS2KJ3SOwX9NB1rbB5PeYb+pcDqLAnsCILvHmOhBHa+DTMIr6OejKMlgP1Y2+
2SZ3/Dn5rMjXpBAKwaEOofE8BqBkKvU9AH+llyrbXMTY+Ptsqr3vKBpGNWO9K45IuIFa8/ccYbx+
an4TAol0FYXoEZJhf/zHFqVSKcyoC2XtOFvtj7VLzvRu2zdsdaM650MQDVcvAUeaUqChJk1W0Q7Z
jP4T1NOAFeAvo4B0M8ysNForhkPBk+mjeLbE67vTsihxDryfHW9XxCk3VhjofFLcJdkzkYQwvk+a
8hrUWxnsguvx3pApsScXgxpFhdToeEQL9bw6/t/yAMnICrtQgXBtfClO/J8L5b9xc9lnQpeP6OFc
00p42S/Vn42x1ghWRHQi6SQyFeovy1RZNQb/TSW+w8AbFQO+Rgeim/R546qClgncTRiL5FgvDLVE
q17ckBDTqiwJ1tsm+trnjYvxGlw7MNqw52rWFky8ZX6lZ3i91zso3OTQ/0nhrrJ0fN3eyhmiLAcm
PZDqKCfUTyTU40qqYmbQJkMLmIRaU/jkETJj1WweZbgV79y6+kQlZUNPXRnpZcXmtbm7jOze1n92
MgQCgFWX6lUsy6YAFdpGHVTdjY0g17vZbkKRPoBgj9wip92ATdWtXjHA6rZGjBuaF5NYip2TW6Wi
uwpaKL6kZR+X6pWQ+DIUaQPGpZF7hvudqoxMp4kKY59NIeGsx4uTH98e461VPpDDgkktIu7ZZXP9
8bMwFHDBTSw2adM8FItHo3LDoCRknNo1G7hwRORgz8s8Eq3OKo9xbq9RleILkWp22ohUlDUzCzIm
AhAUZbTQXMJFehGLG6ffVRXyPMpa3AHY5YSXqcmoPDt+CTv3ObWfR2NypJSecQ95KZvimTVSvBm8
QVfSDhCBLNMUTr8ilnV2w7wMcSpi/psFxkzfZp0/KdxHC1vWA/w/AC2oZFuHTyd1zOCjjBwX7RMh
af8FzPLcGf++LaJzfp0M4+dKQAJjbNJXdWz8lPUpt72mjeLNtJJVCAXLwunaSA3WB70ppibBAFpk
cnM7RnnudUBqCoSQFJ6qYHOwu5+3/+ZGZgos49Ki5HKdej5jLXHKJjLnpw7F43WS6awjobpOQDM6
2/xfD1vfl52/RwfuGVnXFtPdcfljqocEdoiHPQJx9Og7GVzwNrq7qMi6jS5dijQH3GlYnp2uZ9CG
yVxwPJrsxmr99SMfqUXbC2k+iOKHpZT7wIaZ+fRo7X6pxNMx8/et/Xfi8BhRIJ3eFVEAi54y8PyK
qIT5ZkPX5vTHrm8KxkmLllGPYkWxf2ZDSaI1asTiErlqSxj+8WEJvo6mwh8qDS3TvAIy8r8sWabh
RK/a8ct5qB6FPGm0XOJVV7fStq0obZL52MMK5TNX366MagXmtc688IGw2gMfpCKUgFM1PzmVo9/A
39AxzKvHXMcaALTIHgqvaGRjCEP2/IIHblT52rkqKscj/fxq0/gE8eIAVGI5qLEyP8Iaqhdn5LDv
aVRCfs/k6o8sARtUuKGemFFgddV1u8YdmCrlGSXE8Xufe/tAKkVvWiUHWc0Ux9cCo/04uZsaTyqL
HKKh9ngDppMIGVBuMWL4bKv5D2YOfr4iTZYG8P2t1+A9veaBcRpQRWgvsey3CBrllYVr65rrn/QU
ANrsIIsWp6oaKRSVnyxRG/bFOIsuaPuTmV55F6joPbpB9eQ3YftXod2FWZWyiLL3YyStgengG1nC
x0C/TEBvZicpfOfhyz8fhgpYsF5Bj1pibRfWQQ2SbiSKgJu0Yg8fk17yf/3Sih3A5wZOxTi2na0/
cmSHLGRfwthw/cOqzo0VOXEwuGZIwkFTPo+opkTObJa6qi6xBhyL15Ppr/0SNppCgPdQZ2a41ymw
OUmdKK29JcqSe5X28vuEYbtdAphx/KpeKQOIJ6sgPEZi6gkYZKo0RGwWyiTIFRSiFLD3YcD7MkVV
sIVaA5ee1CbKMMBElwOpSk024fNv
`protect end_protected
