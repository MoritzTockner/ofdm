-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XvXwk2tGSaP3Q/XPwVaydqlPrQ4u73hoTr+wqagtSTrg/3IeS3SDd8wkReOcXiiRAtmuqzQSyJNG
Wm8l859tJVLKkLe9277er0+/jvAnDTrMtaPF0/it9jzOq1/LytLOC85xLOw7rQEC9e4lRJtddqIT
0Bq9y/YiUI3ti8oBj1y5PD2EC1exMNqkO3M0KWLcQ1qwFFDaUGkGf1/1cFqfyw3vhq2j7ELE8znw
4wkf19fi2FiSarU1xoZn68meABVlT3Qbjq4jwtN+9cV/kKEZgP+bYzlPvxEH4PgaPB12IMvn7SWF
7M7RW1D0U87yr3w0+cG1NltSdF1b3TOtgK8dwg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
OMSekN7TvoJr6zQ9k0koGSAXNr93D/MkorC6IFFYmDmvZynCceS1tgh4Tq5jdMs4A51TmcdJvcTe
E6YO2g8Cp5ZjPLGx7rw/rFNehtqrX6Xq4WXT07qjfQxFMEvfujtXbw6/Hx3C4eNS9F5kqjW+5INl
MDhdAMcYiDm4GSL9nCHsAnvyRkFJWuHdXOGW+dxxsgosjuPYaQbzxTupySta/XMhrYVraQ5lscqf
9oqQ26PJ8R5xgbEy9J1dSw620gQDGp9lN+x8RYWTnEfBaBdRbgfIwGf6ZbhX2EFzc1T1lLl+GzPA
1LtTR1IcTYyfaGBP5eBCdGS9FZLMcroYdU7qum/BAmIxx41rS2LHqkJ8xVgPOL+wr/XCJn+XhMMR
6IkEdM99hcah7CposPrY8ZQAl7wgnrWzS3XVpH4YEMsh+ebRqkZkKGRAwQPf8ZOXOY/PsplZG8Sk
LIy6NmAmiB4wciXV0TfGHyF3mQgKiVkuPqn0eXFDIYYD0puAUZuVOgGjXGhuWsCq6aicDUliUwkL
MDHoeblQlEK2idpPbyqgqjmvDNoZGMYbVFcHEoOy+op+p/3F/HKTVt8tn4bxttODeMOIliJ5P0bA
jCVQtLGIiCjbE3z3ndWGo4YCcrSzZv5DmU5Wpt+2ci0sAOuH762ZVFhJppGpE7/a0xpGVDxZwlE0
QeSdIBR4RGqtLqxc1vX53b+Z8dADOwB8oovTddB54jxaRhF/2PzP9zr2CudEMxb9teX7zGrXRhcK
qbYNYtQlGDk1ER+zeXhUoh0i4N0CuZ3fqxohseC+9Y8t53wseGgqIZMgD+LzUw51t/YE0n0WRQVA
ZiZ5M7iaAg4fT8y1hSFHrfsRFdXy7YyizBKKDJlw3+yRAuxVnOhnirG+GCl9uQLqjjyf9p1i+cJJ
Ui4720N9ebQnAy+WDxQguSJPtW1x1El1BpOitOw2OaN8sz+8bGpJpHqjFjOllUXUT3L+V7DMna9w
gchfpwfhu+7rNIvsy16tduyXx/oRkx6FCVzekdl7zgwjcYmldKwrmWfn4IvAcmfnohZMvqGyKZS/
1zdJJwEZ0EPS6JXYG3pGdJ3Gc/QafYd1RRiPLalj4gvoi5ZQJ5vLBvTRS9hxk9SdD3+GMnYvB5EK
m6HviClVNhzoUIGIhMyUbInXuBxP9yXDNOrqiwOD0qLkFMfsJn7QUvYBJLMiQEb/yYduMhhE1eiO
ALdMJd8Mx9YK3U6wr5HknaCpjBkeOvRNUftrObk4eJG2C1brHmI5Q6TjgJZM0C0S2sWLI6sTmnNW
GyVbNUrlT81u13vD1UZ9CoN75B8F4fKjIMFZ9ZfoBxcZRYIPJn8zwRw7frwQRi7O+L+tMlV7gOUP
OKkyMKszJJ8XJdYIyov4pwh0J3nfpdqyHZILH7dA+DARpWFpi0+CTz/2CqIau+0dXhJk9bUznM5n
8X5x06VScaKtrgONHQE4MlRo3asrVZISC88oyxqzjWOHsyxO3SLGwbAXjzEtDTaNKuCZQfms0M9R
HMvHOd10dDw0NaP76Pj9umFykJunpSKtj+BtXUJ94hOyOr6RLrwb3vg0vVYBHBR0tlZLLQgaVy7B
wQCTUZt3FH0icL4zyndYe4DEZP65DbLT5RQSnzGkFO0AIFfKFqz7/LQvAFrWn9+CRXc8zy/nC+Y9
o4pcPPR4F8DSrVk2ZAWttTCS4ooo5TrSbusQ773qugnaY1+8WOa/H9a57PFARgQDfpGssyZ60nr1
l4TRmyJ+Wd8UCdUOr9xZS6xxRtJd1Pu2CZYdEpCX1ykZ1hoGPCwn5EQsAahTXpvrW4Rm19UFz1QO
+sbumyxV7ZeHxyTTOf9czMKwgVFK4FH5WdcJvqQTOIjgHoBVevRTGoLipKFdYndqwk+rgxIwNzlp
7w/TBD10CHrJfhHbvYm2/58ZXkvewhhjh7h/qPLNoH/MHkMfgeSbhyXsacJwdqZbSKgjGrv3AqXH
FoPvJVOCRZ0DMywKkE1UY2QtX6w2zj0vvY4Mr/EI8jLkVrqLQxJqSMMb213qG7/KeweYSNNHlH9e
JftD0IPQBsuz05Jpv4PZ2lS8/57rh73/G0AzFn7H8hlDd/1OLa2fULyWKENHXf55XiWf2fPa89Po
NPYUeTEsoR0FzmAgb5S3TYTSgd5G0UEJWGtZbSCPg7DBf4RmG6mFoW+p/CwGkKD0I0V/xHD7CbcX
xSnHBvyKXLXvgfdMMgtU9nVfjNu0ja6hTfDUzHpLYv4zqFNU/eEFn0LzCZ21XAp04B7eTqcEiAkD
ZYXxk2oQsZzLq3Usu57sFNgzsc/2q/+2AOTsP6L0luiCqhePBFGDjZ5nmAHSkpg20PTEMvTqftOt
ixgx3fk+fXb+7AK6XPx95qrJtPA42fnicwB62aeOFn0+OA7Kvp0I2pIvkcnh6uzdMYKeQ2Ntq43f
NDsahx3HVZBfvnsGNR4ADZb2tU1QSU4ngms9vj4pIxxn2PF9FE7rwD9SqM05sRHDMHU1Ztv/sIi6
Og9d4KpRMwLM7Aoy3/qQXfZvACDmxTPnMjNDXiJbJtvNQRuPkW5bB0oUFhRYHHROE3yRWV1kZ8YV
g3FRjD5oszpUG5wju+cmeKOFO6jOAG/SZzIfVf+PGml6FrDRhj2PL72y4B6yBwC0suyq9G4NJQkj
llElomC0sZu/tG5oXoSGHlkVf5zGE08gjamw52rvCLdsf/C2Iy8sgLJgavqAD37bMiM4xjuAaebX
d+RxkaEecBTxCHbpNLzVn5B11TqNZESj2IxQfqrcUoIie8laY8GyMjT0G7QGbr0R1FD6RehIAQWR
3rBnrZjdZ7E4HMRJeD74Pi1RrD8UjCeTrdKGdcCa+RnR82sEhAjwi2MkWuodQjtL7NchCHDrWl6O
Ie9RttgXzUz4ADCHVCOcxuV+lKfw6ZCO884EItao+O50gvS52pCGeWpaQEVLOasltO2zASySFwFN
ACoDQ01GsG5Ij7WFP7Hj204uaJRZt+13qjUSw1ll4c8hsIgcF56F0FKPvE7rKs/5U3FeBjcusdqi
RNfkAfleEhW9i91UldTBcZOr8vknqnRQhaJWoj9NNKW5xdYP537Zg94fq61tdxzjKjrZdR46v7pr
qkm1oZ+4rFJo8hyyx4AbX0tBKfq7cc8IanqFgAN2qDM7UdEC+EjnuJyaB84Xwm9fIxaSEiFKgpQL
9kWrjlvJHn4sQSkVTJhRexZZ9bfCga2XSAkdBte4E1U0R+qzzdfuMNUEqgpACfwG9izfuXMJEaO9
hlJgVjtgkX3sPU97jzr0PS8VyyqLIM457uLIdHqGjVCwjiUvUnXkO7IUrgBMdQlkx4agQWKoor0l
UcJNjeJfUc8JpWz8DW+YV2L7t89BGNTRSR+XZZqyZ4I/wmQXaeOtMuM+6U/e+w9wj5gNgl0M/E9c
EtU/ICM43NodGs7SuYHnwXvJgKW/W9XJwLHmF3xuZ3AMgB3Yor+lIrmvT4fAgZLbt9ZOcyfcknsC
8kq+xzxG3L0PQRJkKSq78V9tZjplWlPOhlQkNVPNpvzixSZAI7Auap5O1yTS/QlfJgQ7oEZQAIgc
bwVdG1tkeMXZMYg0H5o5pUTurknWmiZB3g49bQ8CCnt2VmIMSybuxNpP268dEBxLcjn6c5RSWqiE
tUGILvGoogZ3T6Ja3Ic4aAuBynpkOl8AHOs6A0QAFP4ixHoXj/D4pPEDi/8u2mkIodlM3gVfq+3D
NW5PMh4i7ka+4lw+/6LpWQdwOnahNQFY2BRrpeMQUl+518i5+6+lDEcjve5jcJNZzxRRbfm+KJpP
S+sD8a7ATr0cntLaaWfd395xC3IqXEGBY539usBPiALfJssu7+Xt559ThBIvGRG2LGsj8R60y2B4
mm31hf/eLLwlBb9pLmBGPsCzpivKrBvw0UTjBviWpHrb2ENmEI5Dxo3hDd+2OmeKD8BofLptysPy
E8GD9Exyy+v/FjiZiAxJJ/Qf0XhqBBJDVaSwt1lzQr3Nb3OvFl52CTJ9lIuZ+e3EBJTcgvZTmUDH
7ppEtM7TfGyImDXlHA4XOnhi3ZA5ZqHbj+MeQo+rEr8QwHZwZh/5fmW9XTrVrx/GjoGe26alksyU
c4BnFei1NZZuhCsMmcheS/6Y8AVaPMgiznMXa8qbnZcZ5LxHD9Jnu1uvkf6CEvrThq4Pe3834rDR
/8Sn0513BvNCEh7ip/21q1Ga/eOS0C9QMy45Myey0gFnYblm0svbXMhoEpcHbn/FVNRCLHuiNXAv
cb8sJcDqNRmEDboYVz3rFCs08w8jqjY3Z/PjxBqftBlhNFYF4UqEWEzpp03ck6xpRmHUo9CTVkhS
swCkk4vMEvzNSv+0RoTNtZwf/2v29xHeqEJbR4WXMok+Pg5KGg383UGrQD0cR7ZSnC/9lh+fo5j5
4d2J7dKB88qqP6Go1UHHLccwCMk2c9KQWJFgmL1L+6ZNHK7T9oeoxd/GaLicBNDAzeyuGYbxqctc
MOazZFpQgq/IZGMv1C2gLR2N5L1lFECQISCCU4i7QrEwVP75WJOcDtA+2IoXjQ+UndYSzauXp4UF
Hj90sHiuaBmboW1X1FKiQ+D5AJgBjUayo++GdELC2NQK+YuMjooyofVTHyghr0br2VtcP+B7WBFw
ATMctwRbzJ2pAqUiT0GOvDFT6t8Z4OG4hFg1eYpwQf3m6M/2tL8RbkjZGTsyR8JDQcRZK23MMhdv
cwrrTTk66zcjV0AXD+3j+rAulemGC2ep1pc0h76LCQYA3nGeKe8Gt3MkA2ktyF95DpqKUMZvFFtJ
0aG4xHSLEtRtcdzog5Z1Fbqng+mnlhWp8wZ62h9p5ztR78ZwU4KLbsXvw9l19xdkP12/73P3lC2/
G2oebbMm04JrmWvXldPV1lVy0u6DZnyhgRQsvDrGulXEnVaYr8zwZ5bvh3KxIhKytZpoiUY46ivY
VvvCko3ephCRjPb2yah6sHY/Oi/SIpusmEbQ2ET0Spf6/LcD3fj0Es+0ASpNHWaVuklQ2Ud3BOfG
xA4OX8lglFOq0H4DH8GKr1IvQurUaF+mO0E8ooDaNWvw/6qwreUlyp+4MnX4W1XMTkLOZ4KAmIMo
mP5QUM66JNH+nP18Dbw2NEgV+GqlBFLEKL4dYYdwKWiB5Moz6RNLltxyJmDBOyVhfIbVq2Hc/8vH
lvc38N5VoRQ5tQbg858MfPnyTkON3vFjA3WbLsMlQRwDp7jfW2gI+T3+mSL1u0evh6cNpxAiShsX
Z/JTc7i4a+62VXtowj30xNfGct82V0MRv03VxB7GYQz5/PC4kFHO27R2xD61c4PO61GDgM/co0ee
M1OI7f+d2SdnbZ0b+hKYoTjBKue79niC1xcZ+L+SYBiOPMsQgbsxJuLEiabtoRsQCUbin116CZBf
s42uLB7o+EDHJ0F0+L9uHLf38VEsZ/ZE6nql8pDkr0Hi2mU7q1GVftukCiYqVqjv58IOanHEia0p
tz140MkFru0fbqLNzqUdgMOfsGvE4wx1P5YT1kxKDETqj8MMDuLWec1BYFJtMP+V4PCz8/TA/0CN
HrH0+yLH14WIqxIzw31EmYjRgL8RQ6NuyB/Oy9hwni3f2IT2uvYcXM1fO2h/igpUl017qg0BONB8
ohgcw+/h6RYslwuno5S9Mgo6g5Y4PFKrsWuxqOHeB4BqYdpHN+ny+iYrMYevm9t6GyD5PH1vzaBJ
XM7/593zt+Tuc/Neio2ZeYJGDca0NIqqPMiqmsWSexxLbyrLW7Iq8i2Mu/dY76wmFTxubt/yQgVT
R8LMhi08/Q+Reyw6XqyWvCe2cUICRfK2QLgr8b2rUfLXD5qQX4cGKKSBiffA5RRugjEdE9H7Znon
Ttf7aW8qzMOcoa4rqbx1LzqJm7YJV9qfR8ZXrUyS72vxzjUERyd9a0EIhOSUs6x7pMb+8GRZ5bTw
bdMbtWgq5e4936P3xdKIfNP9O3RZariNXlqMDc1dlwZ8vpPZYeToni5bCjTpiXjWhL+Qu13HhGzC
QEIxuAe/aymvS4z53wil6RnUQ66tiPADD6hEOZzyosLJ7y13oXEioLb8Is9/w4G580vsFBNu4Ayl
+gqM63Md3QOnb35qP/gTVhaW+D1ewgKOvLEb87HbDmF7gu7N8DpWmw+TdzzbelFqn51JYoXrissc
7Jn0QX7M/dsC0iXTv32OiTlVl2BRZBCmtyzFNCONjcH88K/gcHVUL1SaGibi61Wxri4N1rB5yhrM
5BJOudkZnuZp+N0eOtB7QDyruvC22hEizhy0ZWyj6Yy6cQpQvVaMJjnYEtrgfa58vd4alVNm7laW
hrT3HFReKECx7xvQWjLikYGnH09txpWnKgxXwy2Gr3jO2sBtmLm+kXI8g7ZWrtdFE1wCc+k7qooU
xL7aW3P8lSNBUQ2UQFApTppWjHgzRqgEhW9gfgSwrdtDObL3hn/WZN4y98Wp9Y8uyHmaugltQpig
HTQRwosO0CSuWfuocu9QR2KY5X9V0AoZ50xxK5PmurZfJ5z1MoggHD/sEgo12CBY6w8dJRvhq3ch
YVXM/aK3nA62hrsJIVBIY+MF+6kZV8xkCYv4GJtFq5q/SEitryc/r3tm7NZTGdmvowqmGY7WbieY
XdF6QQmXjb5YB5HVwgYSUj7vd95zALVEQK/FDOZs7d/HhAtLFsoNDUv6Wlu178AIMNOMT1BqW/fd
uA4QqJvsk5v7YDKCKp5ODTPSyoY0NJ+XLa0tYPQr1kI4G9Bf3F7528O9eH2LZIGY8GmJI59bDbW4
9lAZPMXiz4VveR3SNU5GwzLMafIHHZOlPqBN5Ca6BcpLV2nHcG6Set19rvqFSP3ri95idyPI6umT
t4EPOwiMEhaaEzd/yyHQJ8DttxIpDWkQMAHFxAnBl+SKX7kZFerQhHZen7EliGz9YUOWsmqXJXTi
P4vOlEZX1JrhGC9MEQ1FTmIVJ0bO7ImE1A5m8ze46vLVBr+vDcBuQ/IEIc/WqQJhTesiaijcdpR9
vlHBhwXtBtfEbWSSG5VKSoCGHdoePiEFS+glUPaSgtxIq2Ha3YIl48DUmxBRH8aOhrcfW20hgqup
6Nx4toX4yghKnLx2drvUor3TAj4wQ/7t2DVX76yGs5qxxJQkuK7ZSzyRqgOHvoh51szYOH8TAN9E
ryxvWJLOrwPByMTzJ8dgsnwKdI8HNVrfY/uNVGbuZv5csZSikUTc3P988T0MCVvrZm+fZ31ipt5q
R06msx4VVxdGZu/jUVxvhs/5ve7/llymcqkExuQUXOGkxJsOU63hr2q9wVfeqvhcIybh+YXn/lYR
eZUXe5mLl2ZV4SlWe06JvZ6Grp9v0nwz00umAC3ExkNYZJE6WciH0c8+82o2EiN7r7zjzKUrg1qg
sEvijCZ9beMbwDCDFNOtZTXZLHtRe21fQu3VZJE1q7CWgaHAtaTZVe0iMd9LyVnAXpneTJy2wUAw
OOdqVC0mKO+cckqujK3YRcqIgMvtfE2t1epWU2nI4CzSrTwQO3QvI68rIHihJmbiQIqvsBJIlKAM
lGJoku7J0qnU9uSctAytDcXftHs/P/WEorGNoRuP4r1H1M6Z+nuOpTYxDDcNp6JKMhwoHNyJ6QXD
lgU2YNX1GGPo9fq6N8aArOkbV0OcHPHEh27MY0TTD3o0pey99/+jZXeHOs6zajfTXrZW2NFWA8NQ
NLiYnjh1mpkw+pINPeQs7xEfYLkoIV85HXKN7QDxdqqSMFGKRy+TdmZ6MC1tDg/N7+w98hOqL4PM
rxmK8hqnRUMdXe53LkaO21LBQOucbBHtD4rtEFWWOxp0K1VEYPsGBw1WcUeAZcLjUYMtBPiQBR/V
mmkcIVEv5UL4+d2YSKFQpIWx0ZsIroyEjT+lAIEPe+8hyRgFHgvkxHMC98VAxFm0/CJd6q2sVZg5
IniAAQ6pzdXwXvku61svC805BGvzU2+PFO3pn/wv5nP5anJXmkc5srjSAsP+3z25VTuAP7hk+cFm
MRJ1aq24DcBzr2jaqaYItFXQyGw7LJQ3hWpXmwWzbe7xFS5hA/3YxAjNluRy0ZRGuO17LLnRuSdw
q/7s6dZILmmiN/DvBBmhTblNHyV8Gn4q16tNhB2ojGx/8WYQA/b97mgwf+c00ux1Ngxfy7m2yX9H
ZBoOui8XWPF7wmZ+U7/FOkoO4+rO0M+IeSFM6TxrmEdHbmYd7atXHQwSFnyONvzQuAe/z65WJlaD
VJNXkBf+f8ZcTurj7a/9cm7bNoftHSnzNljWGG2bnL5/tBhQTZbVeYVKUPPO253I69vcQkh+U0Vl
Zae+CGY7SlKJpyr9d9XRGalqvujoYi0DtiF/3TtFgy1ozkaY20ZH3o+iit3+1dSXnNMi46wejvR8
1S9Vm/TXKusXJAQ/5KFjXDfhi2KcBVApps5vQxWBdyTy4BQtD334+wixI/pe5xFQTGC++jJlJVHP
axgdh51q2nqaH5UhIS74zBLK9rjUMu9FaW+hhWAXf3N10FZYSRxSFD7Qp8OGLq0VXz2RQgblKD93
ERylDYNP6pXCRe6FoQ3vRIwAqigsWXNyDl5LMLvMJ8BQIbYYKvxs/wIFBsxs2pkKb4McVz2RSJpn
NevMGYv9KdP/7yllyW5Fku7WpgJSJXcLONPDflXcaztkSvScqKLE62S+Kg6xiON8VTMTZ+707KI8
mH2xCFuIG8oUT6QtvZrSYQRrFn009Fzudi2r73RObzWz4cZR/u0D01o2cxxI9lHBfKMJQinjq5yv
WqwCIGUcbCmRO4yTLl1+pIsl5hGjQzCgXBfOOtn5zP4jQog1y8VpXaPSyz5enf2QaU0dBVW37ti4
7wSOfKORnoWj6GNnaoEbt+ovdOakxhwonkY3wAINkm7m/B4eNnoxa2KvXkR6K62/IxzmIqr3hBOR
V5U/b7qLZE1wuwZeIJyZOAU37YuP9uSc9IwdzNQycTpr6H5OIxk8OYr5YwOTCxK8qSzKaAwRdY9w
v4r1mMiydN+am3n3IIXdhr7WfZffr2nL/wIlTuQnDKlPLZdZO/ivRZdt+szqcX3wKh0WxtuZhdfy
XvECvjRw8uie6vvqR7BcTHr5q4BqezqEDT+ViJwQor9FCyF2wVl3QhUqUmkwqsa2jIVZ4ceqib0h
/sVDsGlJa0YxIApRdDOXX/8ThQKjNFGfu2NYlKnYxbGEOKmIWSxdUW3H2+XvMw5p7LTIfwzPjxwx
JVV4uavQrU8gaWGM14S2ojgyH7NsKTsumOBgpjBbPB2R0/iY1f+6iBs8tITPtU5fdZTJBh54n33H
4pssF+NXN1k96ZcqM82WIZbuX2PvYJuXwIzl0w4ZTmEJnfgbJMNk3aGx/T8d1VjFKRFlrGoCBk6U
WIFcx92ExnkJ57ifHWhqYrJigSrFUb1wdJJV6O/ppcSYQ39a1t6iKMe+UmqT1TqhqHDNSBMVFWz4
mMqsYWgCtf58nyRfoUiSM9jPDSpw0qj4SrgeaB1mCGfPMFZHG8tbyOtPA8/YJ6O5d1OfnYqMJfnM
I1igUEwAeRiDMjdI6R7TbSxOOMq0WJjj8TKGprXs5f7nyoDpnFDPbQRhnzEdNCFYTpSfG7YxIqjM
q0lF7TCZt/MkYiHKfRC4N7JPzjH4TPYBwDX8pJOfZkMOuPh0sxzAgkESvKammsl+XWPW3L0Uzuj0
VlJ7skL7ZDVrOkoh2QjTUDWJ3zejLEDW11kNmxLIgzlNnGyWlb4u3gArmqPWv/It5w8esJ8982sQ
FpTQQu8uQPfI7UwoNZoaEeK1ktkXmu8aCnGVJngRtGehqDt9apHYY9egjRLl2fb9CubcpKuzSHXD
pkimKgRZOm9dff6VTBKsoNOGf8tXTY90a0HQBarK9TMyvicMmELHUGAjN08/raQYB7/LclDr5u+D
S4OsOYDJX5aL+GjM6WNf1X3qrWaYGtceZHqdZiduOmGilMx2lNUN9NUVA1YPdeYo0cwelTPbprYE
UXjDOXAavPDuIHmCgqrFhTnZ5rp7bVnEpPzPxLU92pqnxIX5EsYjSCydxTnGD3YzlPToprrA/6LB
Fom7jDG1x/MPmtzYizwwOovbSGhAX/x4abB73LlgWhZiBaShZ4TSRTNLj/1kYsYBLGCQtTfLvVfo
I+AQ7+V/3Yk2P9wCp2MvFfDDDsD9ZbR5GKhWyGgQXeZluMZDLLdfvLI8JoG+o55pK++zpo/Ix04H
nufdCtonGc5wwprBneDULnRPMtqTLLyylNt44rypIO+eeZDp2hQv7pPCHYtAbQMIFiEoNGaYFi3t
zkvzCu5Bw1CuVKuBCo2Zh4P2OttsTGx/mk8BtbLRhnz48f054Ahxc7UiZQOEu5n73iAPxedcmSaK
V7jNFsnAElzFgbm4UmSSJitBlVj4C2XfavxhksD5JamQHMYsb5LKHnu5HjDpK/VYB2X2TridGPYm
PMEEJpl5iYmg3qVvYsznE8LHEehdXLEbrZzXp6QJ8pSHl3+jFajcmwXDxYtle6fwAWTGzfh1CgqU
z2aZd5MmbQtw2ndh27dbqG3u73GYYzuwWojI+jvmHnbbaRS31YUDw/7pau9qKn8oxBUZ/FHX6VCf
KBWY50lacKMRl29YyO+7R2ickejHjdpEeecbfto/22yI0ciUbVOtkY69vNFwpBwqdeb0YmnOnmqy
vKJar4hfNi0jHPHJDGtsoa0HMKTZV9nXaFjjrM3vertbgi3CbG4SFni/AVgMbozLmH9Ht0gJl6Vc
7GiumdwKW+MmSRG19GFLaSiLb44fLOgzOYeJ5icRJFhrmiAp+ZNlKhQD0cYrvhBQExIx2XbkS3iC
6rfAQGRuRuxUTpHNP7Y/l1bGyVzETVnkbBTndNiHPTA0hreRC5b5xpMqT9NOqzNDZolIx8QKrq2b
+Fpvy/C3AnIz4xRJB0QHZhEK4IfPQVHqE9XwRb8I+0OV/8b/k1F6QJsl0+UqMh1elmroZ/u4zgM6
33e/5x+HY4/wPo6xE3bdST8FFHSl3dBGrRFNkteRZklBbmq6cjJqp8vPx25/9UAmOKYU/SYk0ZTT
BPLPMLU50z036CrDiAsVzbDFsbXtwzMKm9DcIR6NiJ59MwEe2+XOf3knPupeM0qZE13JyBvCjnD3
5M7cPw+P+FfdJzpPrcOrtYSf5REUl/HsyzGYy1o5nXqR3XockVGJWYn6tUhcO01g/KqsEYLaqp08
xmtsorOFLJbeFb+zgjW95EWKIiy+bejlJewSXIWvzd+yEFkevl8BLaAI/x6MdvbG+6f0BFuvdpH+
lS+Qnojx1rdtH1/FTUMTucuQrCslr9UR2Bg2GqI3yRvQG1bbz2TSZeqAzCspcXiGapdfcgeZ8y6Y
zq3dhsET2VbRf0lhscakJVMBzZ6Dx3D1yyAWeWklQIT14MdVJM2VplQixZXCDn2ZRRFbZx1Rd5C4
45G1J7eaWsP2q7YnYocPXaFRwlOqgv6FnvM2yZUTgPWazgoN9Cwhg6ZO1GNEbY9oC2iTTi06bVXt
ovaDmZ6YZ3Qgui2/Wg4IAY65YBdgzN6xf0m6UpOalz+gSt1fR07qKFgie8/uOX+3cOFWznfVEdgh
BCfg/yMiAQA8se9C5oxTuzo8QZ6e2rdBK2sOMkd0gsfdyVj4nfx5nc9aAxn68NhGNRVl3eS7Rf9z
s/B07ZIECWNIeYjr3e8c7Fl58ft0Xbgw9AXF0+NXo5LTiKWaI0O2c4oEJ55pzeXt2qZu9IZdLj+W
REGuuI9xMSL2+zEH5uT5cjE7u6+x65QoIErL9PjXCp/EBhU2RKGWbyAIYzrtIAACOUMP8Z7rjKNL
l7rMSpaC9vZaZNMaX8bT9wJwTmkDd6bIbJUIvdaKmDj8jNu11MgHQv2/xL9QVuEWIqOoN6IeGQ72
4RoW5bKneknlIsva2XLP1dEkgZfmMDspAv6YfWIPD422NVe8o0jxFhJEc2yX1sNBxLbgjV6Mwaq1
/CWeWSTuLgLpUIAZ694nA1MCZlAUXhbVFQ3G24GB4d9WBYu6yys6D4SLnAKkbDzqR3ubQufasLIn
dyA1IimCL9gQ4sS2CzFDKBEzFquPv79jB8hMIukXfeOwFv6/CMUqGVVICIy65OTODYt5OywyQz7j
KnJt7d6hBF+2SIbj1fIddwIA1E1beiTkeXaheLby8z8zW6gv4uYg5JEqLCKHOvkLuDBYbIw2HIbA
NpDnmez3lN/OxMKAu0/zv/P5/jcMLfKuLAutIstDKxUlo3E266lX3fn5Mz+bJKLVvo1NwRyRIFrz
Q+wcVn8rsxSCBT8nsJHLXFH3+EsYh7W+q/ajVAYrWNUYNXhRWH508C7Pkr3+/jEeF8TgrfmRLR0k
4/k71rjOCa5CbIFnED9Z6J2SM9J0NP1+l2hTPkagafhuNbXy9Hio8O03WSDlpHWvsg5Nn4iuXD62
uGRz2XUpZgoDNtdSfE0yBCMTYMwki1V+m0Kq1OHcPFdYd2SpCmaUndsqTZl4fLtgHYtk/3tlGfgT
7IDUm+FbOd2nBpIclU5isC8xspIMSM8id8HctIUDBStswyAO3GTGB0FKELkx89XhMm455MfqMosN
9E7QO8MwIKc2BAU7fBY+fh2N8NHT8Ll08fPw+vvFtPBD8/0CB9oE0iOaAkBLXPP29SqDAHSO/BZU
oyJMNn6Ydt8EdLp9a2bgw2KoaMmOxoVt8zR34Cv9IZDAjFg23398X2GYuceb01xn8kcpjwo/MBGn
koFIpmu9PNSTHFx3JvEM+lhhVno0mBf7RKk0pivmc4ynpmuXdgaIGJj0CYe2xx/lSQ9TwL7vBaQw
oXkzj/zRTC1EIGNbz0NjAMQguyjI/X5QpxPPCdL/VvnEFT/3eHGPo/IOJisxdwciIDrWG1cpPMyN
Uedc9Z4dRY9NxyUGJcZQbBbGxbawMFCKc4aEcSYSKRbQgFyfJsXaflwoelkuTzy4NV9bDg789FEt
WOLM9e7Terh8QyHCUYVLoWcu0lb+od3luXFICk2ZjWD6Dwho6f7w2lKNNcYZrUFKnYN8e/5vcEQb
sB73rXCy2SsDaYgAsem0unXnGerG0Uh3DarzvTZ0F4Ay0DxghPwgsv3dtQht2hxz3ZhUezQBQ1sX
a+X5uPKnj0+jm+XFNT+7ZlhzAHRAIb4WcSJPmBkq1oM9p1XpF3af7OMFhTQi2GAvMjJi7bbOpkTr
3Ev+Ig61VUThuzEJVaGhXqRWFzfYnGEGs30bduHHVMV0iZSOYFh9GIKYDLEFaEJL6B2tgWPK+3yV
7l/GoqO15YILu/Sf64x+AWU1d51QTknfITI6bviwPhWpUlQMbeTkjxcA2s0D+EFV4vucMU/7j8SH
oo6HQgeJ0m+z7DQI5D0KbXJntp7n29wRF229/hulN02o5DWaiy+vEgkErgViYlnmobd6FU6xXIpD
JKiGiY7kVDS1Pu8NEh2GlLDqBU6dohhNTSnyvKBia3kZQIoyiQ+6RDAWrYap65/STGFeqPKpYDRH
wPJD35aVjQVjqcrOqDMzHbX/6UwWP4qEmEFRMpIuhPnZ0TXXbXp28KC0hjU070l+kVHXE55OLyGb
9sUCI5DZQouMhdt5q5DMfK19y6YXib9RV81yoeybMHJ/Zwz9lrIXJNGkOyYe8Xjon7/25J+tahLH
jpYiKFPupoQsaRis8jpzekIllHDYu2a4GSuglH81Vm3Mi+9Sj2ngOhnoCIRlK7F+fB6HN3JHf9k+
5w0yc+Iqe+plLns5BVdcWtzPkTH0VuCClJyiZs9s/uHnersvq/v0C6CB1no569cGPDOV8vsvhtVY
XPS2qFJ7LWheBYZDO/c254uJ1U5a240pY+L/XDGEcEXUNlyW1S7doOje/bUscWs23MSHxt0WwMM9
TDXKD9Oe117s0xHF2USF/sR3/NKqFmBIhidqUJIiscoFyeqqpgeQ0dZ+cVJ/wEgFqDqcXZuxv6fT
Gl6aaMHCOwOykgWpA4R1qAPaD2sG4IfUtKagsQRzT/FWao3R6vtZ2go7bKa5a+H7w6sgj20kk7Zs
6NkoDFbF7LjC2ei6UKKvEn3n4vt5VTkbrurJBEtu6NbanKDfX8rlloN7qhoTWg4ra68geLpGv4wA
I3EuWKVE5SVf9oma9ObNMBMvhr63l1ZSmqil+ecF7OIgnamqfO/dWKpEpPFsS56tzWVSMjFTeXs5
266WFowTki7AsMlDEJgmrU70z8tJnr/+Tfy+0GRME4T0sVon23wkDnSSn5D6gdJOrWSAMaMEioWz
CFuIr42UfAMGDOVvWqdARDFRpldVVeZk5w7Gs9dNeLP14RKIBh2ucbcpdbEAZuNIdliEA3/i34Om
whM4XsxsAq0HvEiDRZp09jymCM9lMvT8o9VManGsnAyaqA+G4+B0bruBeTTivr19N7XsaGYkN4zK
SQHF+39YhkXNXgt+t1nEtLUXrFY7DDPKBBMPsFyU6WL7W20Rbeii6TRsZxXfVrKKiVzqM2Q55fdM
PTP1X0ia2sZrZv6otcmjcwCEMz63ZRQuHKa3mjNvRGEsy755B1hiowzfByRiBfoiT/UW9R8jKFvz
qJDyBz2omMeSyDVwVZwwJOtAfFS4avHeVbZCNAOKAfP3i6iATnCeaBVHMwJA1ZEoxse53k0MiXjj
5/vdHjuVurH06YGnDx8Hzp95hdbZoqXb4SWhpWMUVdC7JaCVnovTITQEY2ETuW/Z9mMNlIkzCzri
BOHxGKOME1dovoOE2umypkwe3Okoyzq+nuAowAA68jjW5+8dzj1SI51iYyTA9y41DPyyktibuPJm
j7HSGl0pFbN6IJGgfgarYAwWoh2J/Mdf0k+BYfCup5ZZMigy31/82xI10fKmjO5pQz+neiAjMfnM
5n67VZZ5hcBiWSJ45GvPtjKUGn+odJXW1M6+Xc7Kt5lSpKnIGvp8eRuk5mdcp3XYWlDe2s4qcZQY
z/jo3NdcK7i03Q8NV+GeJtapQJ+WTsalLyAetuZKD/XCYMx+tvsRTP02ZgKezQFzs85ysRmK0fO2
eulHHHaUdJZozXm0oBjRWv76htcj1Q2JQ+yJmoQWLK0nHTUcpAcmqV/sj7hawdbdKUcA7aS1ecsz
pVY7+VD0plFBUT2ujauEYB+jDnYjidH2CqAhZ+qr12k68e+ji4oO3c8hXl4J+FyVHjQw/fmrdIUZ
VP5nfpRwxMUGJBND6Sdb/Kz16+6DVG17dAxQsywky014T/UFu/TU8HXkgrSTF+X2NLc2bXKSluSW
YEWUilQ0x5jkx9eG33pAZHad3aB8NOwY4P95lpeVUPaOGVLtKoBFFb5qooGZTC6OSeMCQ4AIw8eA
oNgYanZo73ERBy96yNTX6FyQQa29nMGg2GGRgY4L9bmdgS/yHQdFfbkHj7imTIQK7gbcNbt1bhMG
pBaCUmvIH/Dxe6STGXOeQkqRdju04gh1yBRKBqKG9HiZ/DHf7NYam+wYTI6ZITkATOuJ6Rs42tdv
MJlpGMnJyHqizLUJ64dqqZW9Zz/kaHtJjhy12vnpV6hBYipkyC/3mdiqOtPU16s8KXEvr05dMCOx
2P53n6sLenlRHM4y7+L8E/GZzh3ggCVCvgFNiBpw3pTgL0bQ6Y6Ia98TMrrkLBXmGiKshOu1KoRv
KJeMCZfdWluB/jK8B8nkzB4QRsfh7WlZDpFdPvGMR+rQ+i8y5uu7+LWoNikv9JJiM/RisZzDszpu
PtJ0CtU15NcFJgaeIxL89CivrjURDzSN/9K+B4+R6Gp1RMNfrSaZuMPboFEB9FbUPT/MAxFuLqaA
QX/Ts5UbvzTgGAPBrqqpTEmB2NGcPBxhxje7iUIKakfqcqj1krk3yKQwDNRGkdA/6QV1EHLemZX9
zAKtxQ7ewJOsT4jp3Qk5sOKbG6Z1ack5ABeTWVDUlyPpJIzUCbSCWm/ns2tcxAya4RSUS9j6rdMa
HY65rhgFK3lo0Al2ypsoQDmthfC8EmsP+npOXxRIrQeYMpgHxnicEuKtCMW6oV84BMvuByptnXk1
pjT80vEGiRcieiceSrxT4yHjlbJF8fn4ldKBvBT9W/rj2r2Zim4ciMUL9GyeUn45G3CVRwUv64ip
quaZDpvoayIDWVcl9SRJvKOVyVMME3p3gHhcMwtDxutZ30h1Woq4WQiDtSNeJFdLnvqyVcR8jEjO
jl5Xesb9e5fo3fd7s5DGCstQpEBFf6j3/cJTJNYuGkHXZiBmrT+tLN4SsCjmIoZuY7hD1EYKlOKK
n3OTfUvqfW3zf/ViJ65nmuVAS2fTlVuz/hsvz15vlmuzmMrVhDiQn54DtBlmPVabKq0s+pOJmpiY
ik7eehPlpyc4UGbGnRUb4NqidhLXpeVXBA6Kb0+RpytgRWhQeGwsG/1Kh44u/Bdn2ik6m7soqJyd
FAvuevholMy1YSd6dSCzJnQ8MCO4wkFd78Pkr3cfslemzjwH/25SPmLVx8TUYqMVj2znOWtgh61Z
mGkelPtgiYnIW04BQTIyW/GXHnhKJ3k5xWKM18DDMsxRd9booSr32Lb3vizeTvg7iZhJpGFycuEP
yvqHIdiDwk2dHU01BClNebJ1lWsShHszbwUk1N9qkVIrm6UoTOyK5eJQHQ91XKupDcs/TI9mmg1M
4e8Ek96kus/0+R+yhITpWWCuGs0wF5TN1TqdWzn/IFNcRLwUBJe8QXwzdU3/KOcMoqYMCJW3LgQx
mF+aLHK6QbgnsAz5FBNNT+5ya8pVEFlT3qNIFAmFukwg9qLhdfUvKekvEYxQyuPhAFGId9L1PhTR
iExbU58o2x6rimk22A0CLhhMHH3dw4HtHzicLtcfE4R5VAk3A/DENc6hHJQqSb3FcEoyLXGyiz+4
Nw14OazyMPxw5oTUl50KbqgQXhEEaabXMyMX0yI+h9geslas6VriY0ixjZxo8cEESWQ5HZZP56y2
OTIyRml3gINpnKRclNXKeQh84kn5sPkCgzXknoVTG2Utt81MmTaEKmvnmta8XFQf6TmhJULdvXkN
yNz0BY4QhbdubwDh3i+WnBeAzCu5EKtTIbnB2qgLdeD8O/7J3ugMJNg0XHes8Jc8La4oduigZQaQ
0iHKXmYOlsMbQPVldy5+M4wDVIwO1J1ENegWcZnNsKI0/yqvyrui1Fagndffcqo7aqEJgqrPvJLZ
c6AZI3QvxkWVCHfnvkzGKHwUbOIkBzjHlNomDyYky6wD5zXm5uVhAb098onuRKMGdLxzMeULOWeh
b+VEREECPtn6GpcJtMAt/jq6so5hqXXltltxrBruicOfr7AIvO1pK0LIQdPTq59FcWMyeYQBTDEK
N4aJhaADPi0k/CKWBd+umLpugEJ6dc2/R9gyAV9beyw/AgpD+Fjsz+pL/54v0oFnU1QQBXLl6q71
qyvoJflheX53AOQxnAWAsVmFoPh8ubP8/igUW4ijZjHcnSy6QTch6iHLsy9Oawc4KZKor7TvyfW8
YTF0KYwbTQw6tYKLxUkV+LJp7cQt/AdJbaZW3Cric6bsV8wgO5DAuDDxGPDR0QsDIp+KeBiNIfbB
SVtXlqd7V9ADBboAUN6n1QzuQ3v6lKmf1zBhKBR+ELZGmGcmzIwls81PJ0lA5J2F7S1++qTV7yTL
I0PcHvi7Uvt4td1DPR53sN5Tr00wm/clEi+74ARXgGJ6Sx0B2PnELfLEfC+GLHYhiOm4VOkg74Y3
ImVKqzUxT/ioI8yXTQinuPyq+bH0bRQmZ8xSBgV5UGGm0I5ZIDzxfDA2RTxgxo/NOuYLZtE3fJxn
pxTv3TKrNIGQafnrzb9Ulzr+xOAYn4ByIoyU6jIRPSQil5s3m4I2Z1l4GTmWlKwSHPXFQS7VrKSf
M1ohC71/WwFJqpQPzVAlL3+8PN1m/Xh8joc2QGt79PcnndCpMFErDNzIDPQNuNG9LzTVfqOd35T5
QOW3jDaNpnZ/D5i0ocYvwQAJjs7nD8aq96SUc6Ynda50WebConaoN1msY9ZhKM55qipxWcm/HnDR
QOTRgWGbZQqQUNFN1I16v2eiMGwuvXOHLVnpBtl6dgT9JEVK/iBSfQo8bmRW0GUFBDGQSSTOuZ8E
LP9fEguH60msDHMBDg1R6kf1aEEb68O6mhmZKDyLYIRecz2/erP7RFHOZoQJMoaULlXLsUatrEn/
GhdQhZxO1VLgImkTOM58KUF26K3k1h5bl/klPoxImZMWKBeK7U4CEfUcWlmkgVip1SIDVBfolcF+
9zuLcqQsT5ZzapbHZlB1Fu2Mvjz9YgAlmhf4+jMoQRFTT2uCC4GCbeORrvkL4i70aunuD1obA5kk
DA7T9ecfXsEm5WtjyPkM52+DWvFeIJiG401OBgO7pPD5DteEQVm3YKdinDL1ypFwLgyDIzLV8gT+
A7JD+lSAVHKlNdfUD+oLN69Sivd0KfssXqb4F0hmW1rHq68u9ZAVC8HYFK3n3/N8HuKJ5Qm/4k/7
N2AxsD9ZVm+pAI9hxjI69HtAVVrKmCnliefK3qdkq0oYUbWSOhag4RAFHIjdftHa5zzt1kqrC6Gt
NuXxYQCvcbxOE0noutcxedvRa0q3svRf9CG+qC22cTsdmzeDntvghbd9SSwMaLHZxhMyB3MSJePF
3ZgZlrEI41RZOIn9gKwiPh6U5AuEFgToe1MQerEbJTRvh2BtD8uqnB+iedCp+AY3HaWaBuZiJhI1
BrVF3rWfbVT94RzqzzUZJHBtZhZ2p9MRYdg2nAw+5I+Q9DwilQD4S1XW3M6oUoemnICG8V4/w3r4
BEtQRqp7R+esXNa32cNkkn5Lg8CzlpHyyEfCNyotbdhvDHf4kCrGdGOQ26/d8b/m50OeG9BZXh+i
ssZ3BhMFMtlRw7unZQuVoYcU64JJHbOeoUPOsFpiR6f9JhmurWgMTZRVker7ZgpeZSI0vT6gu2a3
bMyXPjwpFECkN3ju4dtdlugAojX+UVGZIGV4rz+4BhTJVcbYetQ/sIWgHABZX8RXt7pb1LOjZAWY
WihWpyG8vdS1FcJMfHTiZSrsoBWaBdS3XI9qes8uWZWsE/Mv0UIZWIe16iMEpefDEHp0m1AEotQt
kIYQ0WbjXO1lDTTuMK1nGYrcVVGYqcvZe83Te+XKXSWeoxWDgrFGolCdf6/5202I39KtT9xm7vDf
UMS9Wygjh+K/OAt9nOPKLC0+0KHsG7XCr0NDYb+c3c6UyRECzb8yKvHw0vGGajPeKclCOsT9Td3G
X2gxsfnCt6hxxNm1fXsSeUaax7Ntfu30SrBD3qWprhfXarV1HN34SBf/MLKXv/t2iNMS+8bnhwWP
KUfMQcpVrfXRcTt96ZXS3WLK7wffYe3nk2aPkv/RrHE7qT1jJAGBaiiEnxe+V6ophMe2Twf08EIs
0qzqUVGqawnMBaJA++EH3mzqVhxd0JLZtMUyCs7MYCK8eU3nzRpAdA1Y+aVQ9wYBlm8s7Y4AtG90
8OThl+nzkJoQyco5d1TMNxReQOHQrnC46HnxloDjJA0WZIZPvkjUfhJdN/n8/NC9K5JA+/BNzeHW
eKNvWhoHeZ6mGComDg+3HypCVSmuiRnY9RjSpYltZoFoxljTprZCSr1PdM+5n6MUWbLd6Ye+lHIe
P4rBa5iY84OrsX9mrNLkI36ZLFyCMZM2bDfcy538TJaozuskPFqHDP8N+yZvAKGN5TzELDHQxnQu
Eiha+AbdsXA1a8ab9S4zg/QYzHO6H7NLY1FniGxqHLy2y41EvEwgLH1q/dXkN2dbELYqN1PJ144N
bHGERun3QOuku48qouxA24vr9Zyq8Mj28GyD78pO1jrtDDRThJvk9ro0kaPuKibVR/fvBidd2ssD
2VJiruCtDaiNoAYJS9RXLN4rIA2J1Ta8VOJK5KOmLeBp7xnh2x3dAbz1xF0HXmSQWsbxBL3wcUIe
pXRYSm1DiXQoVEAi4vuJ+duy10vEP8iMJjQbmdPTRGmPGqUzzDtdUEedxVMg7EuQn3VXlspvxZeC
FVXsFFHwUcBMVswajQtl4FDzy1rE4xYPtLoZRYGYZb43b269mxGJfaD5XzE4904pDBtZpJARKbqN
+vCA/fsYFd8MmYYEgsDEUZeq0lVdIirXjHXxyfinuMzDDk8vt8/2yGi1nbEpmIREH4ivE3wabRro
ccBQZsba6sBP90lu6Ob3E5nRpdteC91C4J5EZszxJS6CFBuZhqY/z5lRNSXdAcv+wrmqYXsrUNIV
4x+iR+SefAIgqEB7CUO4kMaG13EshoQsijVRYX2tc/+DL+G5pnZqKFxVm5GTqrY50e85Jm0qEHV6
XCxv5iRytlqK2sVCQXM+p2RN6vMjlOFRSvIlunFImx2dQperCoLFqSE8SYnnTiodu2SR5sXMRIky
PdHQ5TzjfS0UVam+6f9388qZi8T96hQggexsUHGg6VFOlpmCFSnGIigVH15p7evUHU7tplWdHd6R
juJVL7G5SE5VFPDk+zF8OB6SX4dOWjTTqTUACoEHCPjmEVPX1rKNmB6BRAL5Tmd888nnmShq1j0F
BzOSJkpWn3FcfCVhCsAZSfXAk50tvv4nGBVfXs3wxLYXWn2JRjHLanwquLQ5CgB0sPx2AkVYp6bv
hZMPgcy7rQOPEmAd8FDWcT3YcEIp0S4QQhmdzRUh8vh7RHWmihco0QwNvgUtag6RM/+Qh/5QrFlM
ChuIFQnqWTc5gX/7FGwQ/HCoO3aGRr23gMdP2UEdnxPzldfCBgNnODMHgFGXuGyNLyedaqSPPK0s
yWBbIEEB9SA+ZP9So4JpLkRbZcix9QGQkemmFC2fJA4A+gFChXE9BqR8YShIt7Km4QpwfB8w3W24
NioUFmt+pWzro5QsbPw2HH1EvAAI3VR2lgL89HydIrqxz31DhBkNL5tiNLC/y/bRJTiz1fJ6ecKm
qcdg6NKbk1VEykWngDQF++ddyhG2UyIIQ/UXzLlTZSxYJVhnsvPAKzQnAq3WmQKqWjAn7/fOaXsu
Xf9JNLaXctCVR3lECSz5vw0WGmh7NCDUKVHXRg0lEP1SjvcXo1z5OR8vJlCTTN1P3L+fEWpZ2pAt
HzjWMVHJJ46Zd/EnbYTxaZqIhlSII6jNzuBZxPF0XR9hY3nz547gmCLyACeb+51sWIfs6vIMRbi0
8q3T0oz8MWYvKSJ7Z1c9alg4UUCWZXED63M6FBb7abrSHezQEGf0N/h/5rZWxeQEGS640rJRHdo5
yT60biltHf47TK2itj/oIhC5wgGc30s8gsZJrV1DvVKgUs1MfC8kQPnYH5baO2ILxVpt9sQkZ5Eu
3gzlXshyVSvyRPeeDC16iWSHaEeU8u3tA779R47BK5QmUravQyf/G1Jtx4cHVPwSq4P3Pb7RhrJK
E3+tOINd8ot1bSaQ0yynuQEIkypW4pcViLdtb49vaw2MqHfQb65ORoYcB3k8idlblFIVMxXxAR08
SKdDbS1fd33RmLz/b5BP/v2G7PoinnW1a7YpYtxWdDoDb6bvsRiok+koFgVsOp9rWjwDTnnNA5Y2
wTb5E+19MtrIXNrN+Pn06HlKHxIENuendHX3P+kPHAWnZx8rUWjJZWQ96g7aemK6j3MhYRZb+kBA
0g7TZk0JeoTuNvGKTdjDpYrX5+W2zQ6UqcfbZ0WavH0ttmzC8745mI6AvFLDY3WwQ4qT6QU19VoT
mjAiBICT7EfvOIu+9kyZV75yRf4yxTKp+76iuLrj/hrv8JmZVqZLVy9+YfBEQ7GmhVGjkItHFpGm
p9KDxRLNXcpWfDjLdJvWs+aokZc/IyoWRuWXUiW587J5bFC4yCGuHogkflXFtu3Fp3ZSt1acV/OV
1yke9HzFjqvFPIhzZd55BFfklN28bB7qxZsfg8qwpN6Qeh0FRFuwa2B8Bq559sfRR9GbSyc4S/x0
haL9fXQCJwZHOxckWq0xlYP9WWk6daVGdetG1/3mcSPtPlvTNy+rCtnIPSELgFSdEitQlwO9izau
1wlGO7akHaL7Oj3vyKSbwvyu/mCplYYveKczISvTN5cjCnPnQ/ceZI987G8wP/RVN3hxRFT/V22G
WdxeoRAYGGgunJZ63mH3bm5CyDI3Kq2xT+JIfRLdJORv05Qbp2+hhu43D0/rxMikcTZt3ZCv27ju
1R3Wy4hBSzpzQ9KpSIEhZA6MO860kgr/8S65pKp8TANAdGRWXZ4D6PlVQ81io5LzfF6KSDEYtuK/
C0A4lMrwd3KKjDzuwI2kegr496JJlmfTIpg6ObGSxPY/qTIeN1hKHuTRiFzlhzLCeZ1t7jjINh4e
Zoc2G0MffRUhwlMQEIGMEJu3joLxf+36lYDA0GTGDb22KBAdW4Gc+cmp3QkT4B4BxylLBef2xhtw
x65v467yPpfVqVmsstDCSuBDt7az8HtXFkvwa8VLckJmgWBpEq09v2Y5MNUXCcfI++pBgCCZIoD1
9FDQ2xeJ7fXut23LtBG2vAUUCwib22XjwEwcF+7oqNEPVFJ3LRiyyYxe7eaZ/dp5vni55q4AmbCn
jA6D2OSGJSiKAJZ4BozIwR2nD/6vKDn/EVQwyCnthqDUOMySkyWXJ6Bsp1qLmN/UkQbfa6L3jSHT
e6x8+zljMP+fFpnr0ayKqItKUZaK2916s0gYV30bJ0PJWEvk5BzPfSV+FpMUNQPlzDJTl15IYD3i
bfhlAPmhpxvO86ebdgs6NFYQGCGntft63MrOecdSsRWwwVH/6Tvt47qcVC0ZlibfyfuZZ4FPQjvG
VfZMDh95Z+rXNaAFYhhIdkgfJ59sXzCnKa4JC7/I/oixTK8vWmdTvpaU6A40HT1E0WAQdcLF3d6s
/1hE8+hvfN+apXATJE5umOvjlF5PZZmEKVN3VsLHXgj9RCUvyBTJ1NECTBa5vMTh4YPG/+np6hRw
kB+lLE0eoAQdzMFShrxKWeRkAGGgyKDMivnGrdbYGthyYQQBCl6thJkSezc9uAuxkupMQ0s0Q0HX
JrzZlemLNi4E0w+40GwXFLsG2Ot3ItERTZIZh8nmxRWOvaLDJCyi8yNAf+LEqbBXDK5B5wh70lug
FkuR614y7rb5kHQKSyfEbu3Jwno/0lLzfBrx2mSzWqzPWAJMR1iGWfDGDReFWUbiwkXtywbvLDM5
zuZpHZ06i/R1MOQNDdhVHuI0ITC2SDvg2CQDhLbbm2Eo8v9pzP776lq1hqocmpoHBIAmgTgK1ZXa
zlv6jw53CNAsCTQXyB49YFuRgI6TeKWet8sGpcTyVNFh9wjz5/hZzvBIBubWBml8zU1DP/AKPjm9
p5cJAC1hqAaQHHD9hvItl0ibZ4MUc3iZqFBe64OvofDxgqyo2Y/qMQoSCoHYRhqZafJvUB1uTM/n
DyDXzqJNXb0vfZq48MXcM1do0TA8XVAGMYZQ7KbgPYgrbI61c7mq6dRPgUqTo1hd7vae+OqIZp2q
v9HyiUR3thEk/nclZkh0LXsA+3oloB9CRZYi4WV/tfjTzoF0Zm17Mo9mlrugiF1Ob4uW9qcgAbPX
+h+YeHiQFGOvgzLBwznOhUw9+UZ7W5xFeL3kk7y5Dcgre8OiPDg7GlV3fboWrm/0I3L5BX0q3MU+
mhm36BX22xUPOFYd5ANZQ30W4IKrxaIJ/blCsWlqOriTEULAA3HhX/jNwInl5FQC8oiub03Pghhh
+rEXCA8yT+/0+zXZi8mzlVzeeYy8p8NPv3Y9WDYHAcVxmz1UF6rHlF7l+I37zu1lGnNvGrsc3IVC
NT16jcElEtUZPtV/AKd07ntzqvOIL8besFsPkVoOvs2LjXPP+02ffMXdG4/y70E/BL7BKUkHmedN
MUOK2Lf6shfZdb1dg/xlmyya7bm0Xc+w1GOBO+7s2Ur8+Rv/g4YR9MUkN0HrKruEAmWI0tzva2U9
Zzz/1RZy8aKUYGrZvFcKrRw8jRrBl+wnWHJvvnTMe9nxZc3tTvsg9wIV/LxIByLhHab+RoVcb40I
FiOOX4rzsYsN4Rk4+7bCnmw0QcVm1PnfwpXFXu/6Cx2M1YKfDWCYEfTkTZpPJWW6EFRB5V2BcOkQ
QIym9lxJHIapoJQxIJNDe97DTcFhpdmgr4rCo8+iXcTV8jQQFbfLS/bO4CzwwEas5pzctaXNMDBZ
/K5gXa7J4BIOtEYb5lHxg/ZNmAEDWootGpJUszla5TCXVnwtZmGpjX3xtSqgSZMwNi24+DsXUZut
G20+UGZtkCVDuv5Ks/vbVFJbGlGouNY1fBUtKAULnogNGVbA14hFjlHb2P05Ito6FdtN5Jue4J3P
KbyZunHZVnEyGeRbK5MCaP/7eJOxFZznaj9VI1LIAGRiVMgyg0JiTkb0/39qT4KTNiZZkMgoQBM5
V3D6+TYAlLMhu9degxlwZKstCTtBHFDHa5g6XsaZOk9h19nLQdg5OXu5zYAjPEAn+LMuJfQKec+Z
XSw0fAEyrbuCp2Lpak7wKtSXOG+rS1LJz8NTNqvZR6UmbuCq/W9HCM16A0OtegUhkY6qh5wH9rDW
oRT+h79u7bBclRE1eT/Q6mYUhf4eATlQE3DJYshKwUmUmlw8a5VXTOmS9GpXwppAmfSqrepBYJtX
o+p/2a/FH1Mu9OhkbSCRR7LJsaLo3wRP1EVKvHD48xd7Z4h6qwYQKhSDDLHZUIlAGYmML4GuUN/a
e97EMn2kNBJXbAj9hJC55Val+sORcJZ3owQJGvHrTOTi62BeN5uAuEwzYpKpKXIJfJY6iGMncmym
rVkA0+iaD8x8iW44tgQAe3y9FptoHMNrCCQT2kc++v1ihfywqROQlnqKDqvQwuUO79+KhFCRFZFl
qPXfXhitWSAOwnat7WDfdas+ptzv0k8h85VH13hWxQ8I9gf3mXIclwPzaNEY4m6vuuvhkKDs7D+Q
xLL66eCFENJsBAeosg9Hq+C1/+uF5dC/ljBUfoDfOeIR4zrTSMa4VD6fkzpFXa27xMiiWMDyNECj
MlgDv+M3UZ1RJPjiiaFHz0wZ7GwRmHmgFVDVIxA++KWWUpiGBGW6CjWN91WrdkW1lDKC98OcTihZ
dYdnTIRDxNsagxXj6Ay6FQ3ApZQHJD1r3f8nvDN0eGoJOtRYvFjon+1STU6qTRFAVicn5vh0p7/Y
kLllE4V8zbVwPe3jUFId/tBnj3jVkFEgeqAhdLHKFBceTgSGxpCU6l+B0JRBo+idsk6w77kRhyt4
2CHfpmi5MnTfBp32e78zb4XH+jraPbbEUSIZ/pb/9Nd33e+s+wtd7UytAPYNiMAJ2CHmBMhl165T
5IwcdDNwdwYaIQpyY7qMim12tgGggcW4OjaW3xTdi77XsSyQuBYoD5L/8RZjb67N/EJeWvltdxDB
sqfv0z7VKEWwSVT245CLEl5lQV27+ESLwfieTTQtRk79boartGpqvwQwJ7BRdOAuXb+MleS5635c
CAKoLOVzHNmnZ24nKX/aTPeg1vXioZw60yPuovsLgbfQ9s89FfL/ND291ZqkM10oUb3efdHt4aGP
r5aYuEdO/qDjJUwx9ouvJ3iuPSLUP3x6vtAOFwvK19CzOR5rCOcVQWLuqRWZ08H4e7TxlimvAnb1
4kN27zcCpy6buv9rV5oLJFrHF1pvVgVmPnvKPlKITzSA1qgVeXc0Qrutwl6H7t5puXNqP3vuWm/W
ihE4a36myxNe5Y8SGzZ9dovZGbauMggyHOb0z4NfnWAr+ercW3mDcucyZEo3PkzNjKP1wQuiyjUS
BMi3uhZVbIXjWKPQsmgOWlYnffAzxw+ofFaKOtPohQD7r+g0d7QexOTG9DAHnGQFSymYuPxuQFul
hQcRfAYvyuW0cc7iE8AANOyC7OSWUjO0awYYEZTmy1nN30Yoa2Hyh/06CII0LaQ53TOg4Qo9TSfy
1f9jCz4wNnTXN/CPPq3221dJ4dMkTemrqJ+/T2j3Y1EvH4D+fKq2obiuwaMK9P9ZoZWZlD/Lt+Jk
1UQykUrvBHCLXC7s1948i91P3Zb7RuvdUmb/wHVL38QXlpx7bd/PL/qxCh+2MZokOUMknm8SmeFD
ENlYgvMLCEjycNGsAD68wpVgPu2dR8W617z7ItelpPnV2ioAmO/BPBb8ECKKBoe/fN23mvccW6mT
p2wu40I5+obcNa2bvUNsS2aK0HDiv1XHyY5CV709wC+ahnTX95g3W3rPDd8W59k6A3JJKMaZ2lvF
hgxst59MCShjayIUcFA2X44jyYDK9vBDClbs3XEBFv+WS1Y/OCmgQKZ8smbZ/BVtyFLrg66xnrV4
13IQlzaxgaqdPsxzPc6HwkTBFfGxnhpxFFmVYAYatvr3FgjM0uEXDCZHQqTJfxxkvB8WE0My58eB
zrqbe/wLOtgSsMr24buVomW1qt1BrsQqAwy5ZoNlP/vEkYx/sWtMTUA+zPVOBhV9Lqzt6xeRmcyO
WvTkqNX/3H9/HHvCw/Ws63E7rF0/CetHQ7xpO0nkkUaOChoKaVoyR4vZ2tnYPr9KORd4id47FkKa
Tkr/YqJzcPl+eY++3xOav4pG8ZYRt5ungOJddod+IDs+mnrYWWMxMP4mVBP3H5tMY7i6Fyk8js11
BGRjYj8scvtfzfilokjJn+INj/K1zGayd/p2xsAnvnMl4NYYoTFEHA9CIKdbGouP2yOeXwFub6Rg
IMC6sk0BLyCSGMUreh5OmAXzoDgkfIGvfEX7kMA/tkZrWWW/WwWXma5N6YmQFU1nbYEWd4KC7LHV
mXCItiPUszdAOhE/ZXX/TEDlitR7HSm+17yl+tNpXgQTAGjA3AvZbFswLQ7b/uhbAT/aSVVjGZcd
8FVWTNg58JisK0PgqTuGfc+MRmPgHC+4XO0udj68pcuoBj6qn5iyDPZL7wuapv8v5rUD0Ui9k/Ya
nMhOkWCOHLzF3ihv12PxuxSxJWtjhkvSNRWoIa0eae2bCRpdCYQ2oWi9Son04gZ+E/5wOrUU4RPv
3dWIHKGwrunVd8WsNMtROHKbRLkYR1IWbXu++RbxA13YSy4pneiqFkpJZiMHZo9ZO/xV6LEeVWwC
haPeFjZfUifsjst6iSPOIXJH5vbGz46E7ce3XPLI6LUjQH4M4fTZhnwD6IPkhp0ksItuJe8PnFDY
9xss0gg1E2kmLZd+kQwl+O14zIweHSjRiW7geL/gZLeHPb/0GuGYlMyePHwZwqH58WFzdK5kp7Nx
hKRUsmSgsZHl5jpbDbgCkKyx9veHjgKW3JfLvf6KFBsfOoQKfFVKz8QIhZRjJPZE1kEBiSwwZaCI
EkBlRkqBHg3WBdxSgmPsQYqR6MUMmbH/gnuGtRTDImciUP66s/Sez0m2qa3wXkfSDlKVS8pKjVk2
u1T5ZpJtv4Awn462VXdcnszQsg2tkfUB/kpPsXclNM7kf02lGG8coh9yeLLns7oVWsDM6+JM58G3
/cNmrOsEc7SA3w2mCgB8nM3H5n7aP23ehb+Au7u/jBnfFhA8ri5gwkf8o8NnAdparubTGJQ3EkNo
hCz5ngKSPe2Vgkg3zQTgVRUZSYECHQnliIql77IQ0e/wNYkvlpTzGDX/xNzSkuAA9bWvYyK6MiQB
Bpdd47wNdnINBJwgJn0ag0Hu1ep8dgBccw8QoEdank9Is/RGHNNJIA1jHi2n2O7i/mji3JQUWz/U
QVQg6l1RC+yVHEtOlKbujc7iEJBBrZ8Pmzfmx8Pg03kqwhvCxR3LBGlmkHurqVsDE1SYanjeSbjv
myYMCcS0cVUdPsU3jog4jq/h70y50srBn4rq1ab3Nd6dmJs9VIpvRHs94ZTCUNCaLQA3ygaAC9Dt
IK8YsDwlzuKMYUsdrUVfyygtZhB71dBuA1+3T2BF21X9cMUj6E8y48RE8gjjiOw/SeFZsj5BW/la
Jf/st2LpLIKfQnTd/jnJiF+IbfuiGy5teyqrzl23a5o5KIgYaooIlhfP3ro0Ol4ivlxpe3H9piHh
/XutmFJBEhW2KV2b0H+923M+kAJPs+e6ePPFVCgu5U1Gbvd47vGv3v4nIWc2TbZtoFOiPcw5S4Ja
/991StCHbMHY3cinqyT1YUL3JQ9cPOqBrDdqIItpUlU709XIYkmHWEwpkJtonV8vUjs6LqMtbV/b
AY61ikIceETt+nkuwhpyW3G+6db3bcmt1feGAozC0pX+wfc+KgHVJNwLTrOxVo82Oj6cxdslWLWD
kkplDcf+6rxRlUpFyYe4PLtf4W37JRxv2j4+/OzMcEvJfNrsVr2VfDM1zPD4IfkeTTDLNW645n2R
zhoZTgdzeI5LyY9qg0TY9Qy2Zy9Z6hqIaOJNERgg+L+vGk4yk6WwB8AoIfrgGBS6lP2e6SECE/aL
s/PxVm3CrDiQu+AZow3vnNxdgXxDv30myNsvt914xgr+KjYy4mB/w0ykwa+5GsifvhKthgOBLTAa
HGrf4jZKxUNZe0WCZy2lyD9/HbHqcI43gw3nKEsnYV7XkLL+T+RTCAiYHFN2SEV9Sz+Tfrbzan1Q
9YewGlZWJEgZLMQQ1P1Do5R/yAvzeLgIbbcvk26AXCjJ3Tv4GIXpigyfVzkcc0GuOMD6FSKZuU3N
h0a4rDQmQRgN5nIBDYgSa1hao0AXt1cjpYnxyyHdHWByT4udXL27xQWTgm6NeL1IO7NQjw0hdzyr
jpbuv23vsNMVH6TQ/qTEYgFDu77VYbkF2C1zWh3MTAwA6jcj1lAyfLkwwwo8tSATXjv9S6ptGqXn
agsws424qpWgMf83IWGP5lOzq1kf0cq+Z0Kqw+m/Q545h7QJZdeB+ox/vSRjGO2zFyJED85cDWVk
sK3YTjdo8xkftH2RAFNlKnBmWRc1GQPl59RRCzhHRlaXzwulvYwvKoii/uTobsgTQSkUEakBDfDB
xpgkViaPlITNR+jCUqJ34uXJH3UohVtMzVWLR+p+QjAH1XaJJzEF0o+YfQtZwPlphLqaW8kNG5mC
D4H4gPmkbvjfoWLn4EpG+PwDM0kDJ3wfjbuDE0R0P1kCUHSOuOt3b3IhNfMobGETha5yZkvTgD2A
YK0fjnqtzeH6Mb0ptS5BFwj1XypQWTeTjgvEoH/rtmKjqNkb6rSi9pqjZQWP9N3qtdXZSfjRbJ1o
S6lHUOq3VVOE0gwYKP+Fe0zRM+1g1fbO86BDLLzAl4aGoKztP27QiemtPOnYkEnHMNJ5r/yS0k3O
kHDQ7IZxtJL/DahIjEZYbtf2fXLjzUdbGD7w4fSjPdfOE0jIjE4Hp3f7+fhE1lSdRKFGss/jqvij
XhtlP6qvIhO8cnyFhq3/WpoSe4DA0599dFZvZCZNrdVT6MKuMdB8McaPj8MEh4gpsWDaDIkt9TYh
1/FUAX6CoVAwEtKsgRmXWUXX5qQhHSf9mi1Kgo1JuO7XyLsKHP/cBInOMnoSP94tiEO6j4lgOtRu
+rMELSypEo1dESWwSo9+o3Eylly48rhQ33U/lp145ii3MBOWgfpTYEUMTnYxA01Hm9bRInmt6LT8
Gwkx4UhwU4KDWDsPFyFsrfrWUA7Kj+uC27c/+qaOO+jvRbcahmAKtPpCTQOAKnRldk1lq8qgbWFc
h+W2lPgygEJZVsz2NovHhWGFLbF4DCS0MMx7eRqBL3eQOrk8Pc/zTzRZNYpMhPXTzXCHBoWEcQIl
hREKV/2P/CkpryagU0I1YUURnr8zX7b0ifyrTEn0JNO5jOJ1IhphY6XKSXFuKFRW/RZxMwJ4dfqu
SL66CEyyYQeXzg8EKN2dmsV09pimUATLznh7MkeEssNJn2R17W9RfwlZoiit6NxRbaX9ZMm6HA3d
6/Lv7AwmvErwx0oaNc87BVSZT7Gw2ktfeeTKcnsihpDUcw8EgK/NaLZrD107N2HBUjEsBVOVp/g2
rs5rh9mmiPZai8shYQWphmQ7vH2Yic/4p35DkY9T/Z63lTsEtD67C8/hwgoBz+9Wh3vjC6dAGfff
KQ0bbTvZ3scCNPoL9RvBFsSsrh0KBZkmQzZhCX753vzqRpjofNg06QuMBX/ikZLFBLlTULFlQ8m3
RGCSgIZkSM9cLWajl06fJ+lG5AddcUL/OLFNZxS9fn2UywqQ/uEUftbhLd70h9+SxOemVD4eq7EP
wyeoAZIlbCcoqEpUmO5pS6H/EwHG2VHLxIk+GWcR8phoCwN7B/GnaUjvI5Pa0t7VidQVZ8YjEuYZ
cwgK6zFHo4ZHVOGuvmFqgeltCmTOyeQuQmaJShirffznY14uU3bThtuqpdsGNeOeTQFDVjs+ttxF
IMyrmaiepNsH5rdNGGymgaUaxipZ1Gi9yvtTpa20xK9C7dcGySFGpW7dFQqnCce8aWtrwblGFnpk
/8XY5mpmc4cl+904dsatoHz8lo+TSkae7ZmNHedolkK7tA46ma7PVCj0ulzhnnXA/dsm7M2Or2sA
+8r8kLp+6OpK7t1O98Tk3WpzL/XHZ9mtNNmmbscwRYR9sIlMZzsr4Hh3IT6jIg3VPnuBUAkQ5TTz
4uBV2KJnVNOFRXlBatr3JILkRoARiwVQJjkKB/TnnM6ViVF+aE8qsJ1xgO8bbxKgjhEmDZAFuS5u
W06qocaBJwgO7ZuEAQXbYiagQsAAKYVovHy6EEg/0mY0RHpjpy3d5009HRRASc5L45yqfLWJ/NZ2
kpHCqWOjhtpoHB2PKS5AwstpxDCqWa4MauNnHuTJVbYzRAZPCeGzXL6Q+OR6sVibmfA27un+twue
o3+GiTd+yRKqkYprXdSa6d83JoB6pXg70Ll4ma0LeTpfs7K7/oQuL7BqBzrjzjjQyjHgjvK9aug+
OWDo9IUrQGi5jcGVnarBDI/wQ7oipmKxvsMp5fu1ZOPAFozhgii8vAZnpx4P8RXPRLelnFW6JQvM
hhPCZH7Sf20i0GfNHgUw7FqhpdLvpzFwv3IAA0Rkqln4E7M4RJcPLFpIBSpw82RBEKn+5VOTh0RJ
p4JyfflT0w8xfzNiM8ItYoe77PlG7RfJL16iZh9HNU1tzMl7K5EKnKwPdMAHtBcUM1SXYkSpBVbn
553KYfx634v8H/kBXjVhFHu7Ou0jbDBr8XuPgF9DRQEfHp/gHXiUwTbK6qSoayRndmsJv5CrWa01
uGAt6hRl8cQBkke3ncWaggp9cOK1SS6AXty5v08a0VOj2WQw1WQBrUuXnrG53TH5uQtfJTHdc18w
uUP2p6TpyE51HX6D8xZPm1/Bvqp3AdwcTMrhH3EPw+M9kqG6RhgeVEW3c1J2xuHuAOFaLhQsyjQ6
UevVMtvLljzAp83el9InAGDvXUatGS5RGqWOX3C555+r7SYrogdefilT9jwYkuM7gqw5J7HTEXci
BZiiswMwEOwsDKBoAUUI6cIkZPT6IWzkVvgaSQX8M/kAG1Re+43L1K++vfGWjU2RrvceDcJtf/tM
MpAdDsH3eZb09YEqIUDkieF9/VINJnLw4L3VN91XZ/JJObJdlpAzQOzXfz8VqvcnlLb64Wa4KN2A
0zb/6yZFbk/XDPb/kxK77drfZUjjxHh9AriST89et/misk/bR3lFtvdw/+0kwZsR4DdGCd21lWo2
gOHSlS9tJBahKIc4uRa6tblt1sHeporX7vwWXFyM6YKMfLjffQJWsZ059I54TM4DDxl+vf6gYJ2/
9zcl9AZQD8Z/0bfYYHm/UPHzmFxJUdcWhObr7SQZjQC+FRpYmXS8GbcMaTRW6WMO6MZ67MvlCxBy
LaCi7sBjg8MKLuRZqPkr0JNR9acTwrhb7CnbU4j8Jdw69xuIoCEi3KW4xtxKQnXuaLtkze3HtvIt
yyvWvqyj8+wmzmn5M4BCZpt8t34goIphl4s6cSK3wNHpFEoq7jdYKEqN+4k6Ol1U5EivwkG0lu3q
Rms028S7uW9DSaJSvQGLxq+5oCCpzUPFiknGuZEVLqIqRBBmUPvUelT0IPCxatLQ0hvNZE9t26y+
vCrl7oPLc/2wzkc3TFrIE42yIZ3YctK825M84Or+PsMZ7tMgXm2Vz8sU93VTU6EJiKTl2/ND43y6
Gzfpun66pdbX08JNNp8UlSMPgECZVMa/dJ9m9Lw31LtDCM27XCxURhXjcfXR49C0U8gm0pTxFHow
iCXNZTeLJfs4JJkyMgVYwB2tqkmLgU3JPT9lb533SKF3lKPuf7QUbrKsPLlXfb/13pmPQedW+xTj
Q1buqdUIt8JZvaJyDdkl1kxQfsbaie3o/3ezqvs4HFKP4CuBVSHkYT8bFzikyV0TvBHqFgQFoH+N
iivEvU4KsT4AsCkXLrFLy75Hk8SQD0PbbKWW/WtaYkNAUioSsxboQCuFNj5qFzr27WtpXxRH37jY
IDWyWA6pO8kcHUHyHmaigbaVjFcIMQ1uT0ZWoQnDUNL2qNLSZweRiMcXtXx8MTE+oGJAysGsLlvW
jfuajUPVJKoVk7RDcbG/1nccn7GV4JVUUxjI3mS/sx95Hc4AUHV98QoUqIhNhO3flnY5UAwNxW86
eJ7G8gbsfW9s9lUqKiuO7bXhNLVAgA89varGJOrau78Xa90B32URz8oLe2x/WEki7Os+OfTmtNYZ
o7c1XyzUs/I3CjbsHAevVPG3suBcEdVJUsHMOqxhSWMVch0cy0+Rv8a+76LVal3THOISgpMqXYMZ
subb3QppotxERlYlGbgvnR4gqwhUV30okD0H+v4Gfbl5akR0Dlhi5uleWE8SUITsBoeDe1J44nOw
s3Hy++jKpLfNlkjcSeW/gCeXthKLAr08HYQUp/LqCxrf1HACSoDAHbfMAq1SoDXtN9aiXzDmVPaO
HBdDNufUQBunlIzMDKGHaLRfLmcu9grOB2DZIBfjY2C3YN7MTmRA/+0euVXk83szH1cL+BMBzNwP
fg/Y1sjW7rB96hDURubKHDuRG5ONtZQrromcSV7UsOvPJptyeVj0bcksurED1Jbu81b49GZngWhs
9vfGr1a8ysvXuTd6TJmZYb7EroYIX5PuAoEzZk5ukiuFvy+6phUQ/CLKjq4hWF24xYXDVTCKp/uo
1IT27sDqEnYnZpFIXJylvkqIKLO4xbE3B/Js6DNUBzi/6xTkdkIkc2F/9+h5JmF/JGjGhYArGuPE
xn1estDmgcxyjQoki7e6taFBhu4FNxyZI+cY1OEI6pKVi0mOpaCef2w7rBlF4RvAiuJP+09hCFsj
CTdEeR0L74NjQWTyI7R8Ht/QMdQaspCq91EePy3NrGqk0VlDm9VeDK/ZHc0eZbYN8ejaS3By93mb
MQU6lt2NTWqAPpcZjXy6FpbxfTTecqQ+v7fkK/ZrpbWGqvGCRGOiPAs3/jfz+lAfdi9RIiiH4zpo
vfGXyhxxUdPFuwbAxwFp2WQPnmqrzUhHvjaQMMjeVZzO/6e32CEfCZ/1SZiOqNSBTmeDJWBgqV7o
ACGio21aMzy5OY/IcKDzVfLPPCjL3HJXZvDWJhoL5ILkOeviezntWtMgUddMwsePxuiX8OYhPVts
c8JOloadbAVpddo4b/hs2clSRVtcWZHoTmBXEg/UEqsD+x/6EYqaTmajiavcsqIaHSGC121n1P19
f5i0zDZIgAGbDZTkb0VtxRHv30qiEVNKzDQR/raXUn9/YxMzOIwZucIIfgLNl/gJt2VDTY3TpqjF
y/HGUM6zTNR16jVW3WTzAtqTnw6cdLq7UAuUquiwKZf0T8QC0r0UxDKAXv7r7eLLv0S6Ifdm4Ksn
KhrWGyjBJ9JylLtztzbsL1P5QJ7REEXgf57pOoizVPn2HbEMXSdEcn7PWovzrG/l+gwv/UDSlDLF
OdQalQieKyon+GPHx1kCWLsxoTdBIfRm1cI1qKjpAewxTM2G52hZK4Ch/z0wD+Ept8+x0PpVtMex
EYBW0vIodrLjlWRR63uG2bwez20U26ngRSVdG45snYmmvbMP+UkefROEFGbZ9ik4XtklPlcyDCz/
pyQwDuVgivuuV/MFNOQkjJzWuoJ5XDsfdzLYKWah6hRplNdX2YY/a78jccXwaIQ7cVa895BwZQNz
NLECZB+zMOgIuDlbDhoii3418JsFT2++Ckx/kihw90/ph5+kTHM1uCAig+okWkMMEbFLyivjlO33
BGHzssjmXpeSLETdT3PRZQTlFpGNRUspX1SnIWYtsPPDuJ/n9Hphezy4rRWQGc61QM879TdS1FcK
dU9Gi+RcaWr8XDJSkbalbxWnF3UyASE0MtGSQkUnaCbI5v/6p/lSFPlLFfscyKmbllslTxUwJ6rm
KdnJzfaUxbr5Y5314ohbabq836m78UVoYXFwyoY9GEMODX8fqPNCumTwy7+Wzmujg1uMkimbwhNQ
UjVWPyaBpmx8A7WlZctqtGXkMJVrSXFsv8Clhe6cNAfO2Z0y4xipbj1bFPwy2NyxA346D7Ddj+Qx
YPNfkqZxWgXFSvjrre64S5DhDch2pSDJZ/GYExa1H6+aoKHt913l9rmD3w8+lyv7zpvUXXh7lXZ9
8y+SZFBrVdl/o427mrU0H2w+ZgJQOIHgD1S2jaM0KOKhgMcmtt/JGhCOL9Fk6pmra/tUppAbvRo6
iYRbobnzS/xDwjVStNSVnAaRxG1nptrbnf/06kfSDmjpc1y0ZOl/itOaTmoNUky1vGZ4yfI07JS8
uMaW1iZ4JeSPF7KSEGYWLP3UcYr3S1vrkhJ0eJiF2xthkvyOPw2BbS7Zuh0bSPNcXYQjNbxqTY5c
Evj/pGvFbLFMP4sgrSjaFYiJoHkT/xIbxSyv88cuslicywi1iNQ4Ri79cfeRgRvUjm2F2XrktBuU
swezZSvt9rYcTNVlLU7pDNhT/W6CobVa+44JRRrWWRtxkqnt0k0OtWCQlE5N5y8dub0j4xtOLjOJ
HUCVdHQOmZcIyVeNZvcWmTnWh6gcwzpK4wr14fLTavUM9YvSgrs4mxjtQPM2AHklOmR7ZkVsAQGD
8qHZu2L0wnFjLjuwVpVTNTczVJDk+VP+ivtSa0oBWy0GUwKDbsNUZOuphgfLFz3reV/IyngxSQ5I
ujJEM3eiesSKiAIFJ0pIimAGfrrW9S+vlkQJsJT1o3Z0nEEpVHByyJE1BblOj0rs4//7lzfOs0uV
4Ly9DLENdsoONXCXVNrZGX0N16HvZTuCvAo1PX3kFjuQbS/8L65PWvZLNJM99uMXPOo3vFMKoCUA
od+vaLFgoUGuvRGzKydMfLKstzHd+llkoiACNl/owqmq3ts5kq61J0Z1Kdz+qTt60p3Q7Yh/YPzl
r5eck6em2nkjmfxYokEO0yxI2IgXCLQpEG0UFbPkFPXzYNx/Gxvd7x1B1QRuEt3XkEloc78qYJhd
GF2qCntyMJrNITB2yN8BVLgnNtr860PEHSs0PDND/PeIrWTJrGwICcqR2T0bpzW7MfESOSFMIPgG
5fA8VOparwbqYAFezyhUTk1LbQalY6Y3Wl5BqnfkgzMV4vl0QAn4MZfClXBzd0MZ0gdiqPuqyqFC
Dz8pBHoxuJS0/PtyJ8Pt2h4SSQ2YmS7NYN9defCW+NN8mr/8bDbphDm3alOHrn49Ls31hnyiuaev
ZMblUO3SaDV8VtFixRie9zE6nPch7mH0l3/FMpeL76gMNKcJNkyhtX8fIAZgNlnk5TROHbbqdJb5
UKIG9qyaIpe2CF5gye57OBqDHomHRe6XI7EK1KA5s7lvwOpDjaojpTAPQlFomepZKKpgjsY38LCL
nYhHBHCw6yB2QjbgZ6vZmb6+AW6BnQbOb5aWIU5Ej/qHaCkjOPmW8SQmJnZc6EtXvIdUCReF3Szb
fDKyAUCOYwftj7qKkJ7sK5MniQIwTBAscH/EecTli6tPO1RwjHbNIe0ZiuxBGPtUpi9QJ49C+nI1
RCFj02JKWJTXwMA1pdobVj7lSVmgjNyNykwFDXNoJmfjmi9lfrl2SHmLOJSh/8VzU8NO0ECmMgX/
CVwIr9gwc7HXdXsyCHqpgof4Hg+D9b+EV56hhNUHWJiXl52LyrJw3KKxY5QavTc+7QhzsBeiQHp2
4XthEXRjELOClAkdiiD0c0tn1yg1HzqA1ZafdywjOqQPR1URdqQYe9w3Scs04musIdRzJjTBktKA
ahVlxSLZj0d27Yl5DhyTn8A9F1NSZx85GuKmL7jAV5k2O0f2oF2o3CxEA/q//JrB0J8BTUlkrALN
tbHdgiRecKr3TT8sI7BOAr8YL5u1VSlPAaN/hTCd8TRSFba+bKKpkB0gE2Lb1685QZ3MzPPt9WFP
BRyAIsc6B/iI/9RnzJDBWgO36GBDbZ0HOCE+DqyqmYlJlHj18PY8Dy4TS8i+M7K41Aer7RdvYFwA
Z1mO1fKHAwvRuMC172PP87llPh/9JFVxuuGBrMD/m4fYckIUG3f5EJpKE/VsD2LSs5a8Pz1oZiQr
7iiLUNcgP30Hp6BdikKSn20JmTVORg6z2F7OHmK6KSgTmvMNVFNq9XM2b/swy8C53JzIvBcl0Ild
fWiUb0CppUww/PgqWV0ir/Z4h9oKtnhBRrC44cd3bhyEyr2SLMdxeX3Ws3HMLWY9cwckLhjiLKur
ZrZ0UTEAg2yyMcefGsHchnzdZRoDPtx4Zz+FHTGg18yVE8KgCiPJASRQcI6ok9GogeUf3RB7VPGN
LLa6YIUTyZw2hxBX32Lv5t2lhfKhT+XX9A3yYP+qhVrszrye/AxyG2f/HPfOX4i3sAuNyKHFvkk6
ThpZ0jdKsS4/JvEtomg5ok+TthWqxi+YMeaGLJ6AiiEAcv5i0uwzz2h2ExBVyhg2HN7zOo2nLCFa
nq2V9n/5RxH7Y25XvKe9vluUs6c1aMLaS1TiBNDyaYPsYW5XFac9QAiYqcyfNZSBz6+xsBIiZ+YA
p3Wm6I7BBdaE3iueBD9S04pvEKlsWc80wYe6Qga2U7TUJQwgBoiKUuD24ARC85ptW+aVQspluxkV
AvmTFyKOa0RnKLFHIV5rWjqMcjD64gDrQyo4gIQwywE/3nvYTjuTf6iq68xDcHnBthCFSMfyXxz3
rUQP8WV+zRNOlhd7bCfLc7v3kxRsOUYtT/7gMalTpLJb8MvidZ6jxYe1nQx6gmdbQZLFGfk/tovt
hhufCuV5/YhRVyA3YOOgAJ8jE29VKR0kW7rRlDozU8+R31tFR1/96sEuhIu7gjDEoQZn6Z9TKiHs
XvLe3CPjcXqJzZ068rUcMSTYeQJikuG+4sfEUGWZs6UV7SbxGCxYX9i0NWyK3sbBlvGf2ngQLBVT
Nt0Xhq4KQ2bcG4iQPQc/9cRX7Ci3WIrKhqTXFSi6GgdaP6tx44WF0IsHtiatzz7MiUH7p8KUNAE1
Yn0uipzku0EK6YeZwV4RkHbQF2T44i9uUpjhRYaSqwxwdRS+jA4QviIXExPypxzYY8WwMwqgwmqe
w3rOTgCO3Ad5194onXRufnZjfStniBPIpuzs5oEsb0QhkCkHptmNzbSqgnTKyWM5sA0GwVDhHun6
DJV7QqtHbTDWfPDQON4YTKiQwra/+X6iJoJIlC24D3lXcLETu9wDYbqId3zV3yAikeFwPBiMKYyO
YaWfIjwGc1AcpyA9iALSeWdv/+e+7moHuysxFIQBnbujeqAlfaG3j11TcZhLUr2WpPwC5rAkuncL
8Xbk3tygxMgsplmql/TR/sIrmOg9C0hMVkJ3EZvYqxXJeCimczIylC8dQs3sUEXxXdL2S14TTCjI
zTQgHe/AVjKZFqKgYdgkGpXOvFIpmAtCpfvZoJP1AfdgTa1KathSM6bvU9/pCYIK8vAuhY9SDsCB
hVy9KRU8J/+5EIJPviWkxyPvKntjR6dtkyeo/5SQgI5OKBIUjxEdPdRvyb5wxPifB7PmCSXcDY8I
wpyRE+VEre+VKh4s5wiA/6mkB9APk64+j2Bd8tIwx+fHWJSdKRbpWSB7d6SI3rSoXgeXmtjEfe06
7gVcTVuNHeM/2FLx24iEsucCTr7P19ggtg2F7aoybLhGScYx7lL1koNyY6Aftqs9x9Np9YV8bd8J
LQVQSv8Yfb9vHQkBJYybOC6LPy8QtHrvrNK1oUikrcfpbmueQqL8FRyiIyDZDCFW3q6p7KSmmi4N
Ksy9kqesRFirIJZECt51uk7wHewMljHduVaTZ62Ks+DI/Qaa6QK01VkgPsMjQXxr0sUKYXvJjUAq
q7FSb0BxDFfqzo+k1frc6Wv3yJ5xwqh6zHIFVC4vFOyng5IlEBNaX45qNXqA6wncuGe5M26sGz+Z
im/lNrrvbpb5pwDRpWvSKgD0z4saDkaeDCQTUUACA5gwyQWXh105BXQeM+Se9v3ETGukU7L79NT3
C6MPGURI9p1pNYfjcU/qiPPJxDwiN/cABzGAsIF/2FYZS7klAxAGFTemODzN8NcjYJ+WST4ZdtWP
N0Nlo92tdND3XlWBcLibLe+YjQi5urLFyDPBaFyqpDlmBXkj96gW++P+noJOSpM6rd18/m1XnTG1
dTHi6kX0dX1l6OEsw2dlFyKIg+Vchk6FK796aIYpHjTTGI5Rq4/eMJsIozJWKZu8p81OGgoBuaen
BtXowP/QN6rxwosnpsb5ucO/U7v2GwPT0SsFtPnVKuizZVJBzEpEJdsoAz/0aIQ/3LQSYfw/DZWq
xx1ZqIinoxGwLvTaglx5ZAWaecS5tow005nKuNsV6WMOhiIxNCqhsBBjUhEDXlqIL2q6g0nwTGEe
25UtyWKgD3SAod0pdRE/mEdHY4XmRSsHI6DsQ+4AB1d9o0GUEIoVrckkLcGbho2gA90dCkGhbjdM
Sc74i5pwhVL9ve0/9BTqc1+l5fV4LWhxQ9zCTj3dT4zxBI9OMFI9OjttreL94j+AvP0ghhfrjyeo
NmynO/ZrZqWLqkj4mUUR67IVsC36HZuCOrvHPb/28FS1tzOgoddCceeTqTN3XUaGvSUfSH3DOT02
weq5OhPdP19i11QVOgkmZnKqoaHqpxHQMgrUIgciA3HRNxJ5gHrWWAd8Es40QkZ5Mu20eMC85qU0
d6k4XrEoEnN0zTnpQlRcVGUgW2e+9F7VhkPgRJM5mpoKCc5imMOA68KCT5La6WRI7I4bUhnBMxsG
NyWc2t+P+5IMIxcEHjRWE6A0KurWdc7WuZXo4qQtGfRnAMtCCjOkiiTGRBIf2h42wJh3RGzk2AbM
ln8R/gygQp4pq4WYrOgmhFMxLJGF9JC8S6kZCz7fKzfZtRsg1upK1JtHDgxMpxvH+FJkJBeozhCV
zow5UF+fmYIuxVlcGNcWZJcxRjnQIXOaQ/IAjn9LnO+hcDUuFRXxv0H5ESf5D7tm+R2ufogQ0oaa
UvsCWZ4NTMXMkIKUqBeuYHGB1xqtb0koU/NMoGn5a7qaqhmHFkNx8ao9pwoe+RpFI49NjIKIYmAB
GDQnrQi9EMuR7G2cQS204CaI0by+N6K0XBDlU1Eo9TUJfGxoVzXQgF8j0/vscpy4dha4LWhIbsIo
ZPL3EZ1HZdMpscnDRBrIOCKzaNAV6yCSQPB+txx/9uxdjGqFm8eg3C2uGv8U9YtrncNziSyWWx8Y
laU6OdiKGE1clozxWzjU418XZ7amgxzkUVGUHLSk6w1l4ctcwdaA14UIOWTOGSS6uNu8A30th2NO
NbazE7bZUwZSe4F5+uMseuTdhLFvSNJNXk0Uc5razp2iWANHv61tUY5zajsU3drnC+NXtO4hm7Al
2UXqhdoGsmhnUW91taL/Y8VY24P64Lm39np+ZupTz7sGmD/k8hR3QpOh8zzwTOMxIG8u4IKVbfOQ
P41EqKzmXcSNXUtQHZNRNS3kMt75vwrYOhhlxlQ03c1ZFUqEYgtXAiQc2fAbBkbzx8Y4sYzC4BYT
M8+BP0xe+ksrWlP5tTE+G10oKyq2QcdRKfPKm9uvGJ3pMVUhttkh/iJnNzC2OODsy7IfN4bpDnH8
B1tSRSqkGE8ajdeYr75FHrcPpMbu+HRH5gF8DjndvRU9p5STfTXuWncOPAft3FW/sTeGHpjDMI0m
1ykMHWckWzhWmT6OTq7ac4c/vy2hXnda2qXt2aLT3Vgs+Ul4cDeRBFhY9G6evh0q94AGZImAhzqh
ZrqckYl5jzFKt8ZYyBhdO/W4KkUGMooJjQXPyeStys6WNDnR8EGO4fk4eoTrf/61tFkK5cA6HiLF
GnWOUIU3c0dGn1rveqy3rZoF8rA+OecFHnweMqHozDAArd6Jo3aui8/Np9/W7AvhIGP6qunR3obg
57oi0aB3M35EjtoFPYZ0Kdnljlsx4VenLj0kwAHT7ULihVpHu+rs1JwM/r0lTWuN+gh8TQvJzXF3
d2W/5RUHdhYYMb3/kT5nz+jg3sF9WWX9xVEfyPa3e08GuDGJMyfL3EEKGkFAoc4aigoF4+qEZkBu
pKfO9AH3vWQTSh0Ue5bIYHlROwRoLwkbKOnUNgWX4kFILarKzp+r4+TmMXGlw9nendqXSLqheSoH
24airn05ZtJc00+LSWgPVRGiuAvS0dgFlmPlsvV3zD++se4K0CJrL0ReRqDoXMICKbJlFSUc2Lu+
2I7Q7mveE31frHETK+mCIDBfzWrOKakfYdbeYkaYGLy6RJFmgLQHqRG/IO/r8MoUqdGTL3MNWC+e
nmewZxrX8k/s9AZx2RWgGAUGXJfkTdIG4fqvCzRJjBjFQaDu7dtBgxXiBoQeZ/IhDdQ8wOjuwxAI
ThGuSd03dNdHx2ydNYzoJflBjX/4eLizl722aLe5ilR9QyOduJKZY/nHSOh8pgP+8XRpYnDI0MTf
cd2jO9jTEE/MFW6Qc/uleAUuwozD0OiKiKWypeqMLlMCHJ9MW/+pQSShi8n/dOduQHU2aOellk0K
H8nEB8PYaZ9ONR1eDObRlM0SOAxokRIVttWNRDuXWFR+iYNya50CB2YGemtuVe1W+ooEHhkZkNgP
2yAoNNAB6lbYO6d6RGXM+tc1UqVQTvFZrEWZFt/f6fJfve6EhY/MchrMSs6yQwg9HUDy6KDgg40q
xIDJyiNEgD0by998X8Yjk00oJ+00HiRpII0q6biIr+WJhZETRJiyWeFPlZS1wrKFmyfmEQK7VMgi
I8XP+pRc1GVzNORPFvFCTkjGjQbYkl6i6Vimg2FxyZ00gHNCTUyOPSx/LKpz1AYU34CZ1sKlN016
m1ZCNtJRGcEl6PCqOfvD7gn3n71NYv3XuwEdhfYD0GEp9oO2JrUCmJGVlKDIPyLWNQTLql/CyAEZ
EkWCCbrJCVtFZVQ1MxAd6WrFnoxTrcQ9csUpRrnkA5Ifh77qxcPlZaqcMksi/jq9mSPRFpZVvyPd
fYHP9TUSG3v3MP02Bkn8lbt2jp0LHsqCZGjljT2x61E++evirF0AMwQl6JFZR4BMhy5gIwz11UHe
Hup7ZlIKDhDMQ7Ib2wyCGJx4e9YvF3IUy/QgE4Gy1FSuy2mmQGc+bGtytUq93iTcPhMuoGKWk2QU
GT2Jh72o+QJ9f86fqPTs7wFYqFs6aIqixL0b4WD0qso2/CR7ZIcKMd8TGqkzO7GGcw8JWi6BRhZh
9DSGocAkyZO1ldTzdfSzRPaOkQEKsa20wrV2lrNaAKwgdoEeCIgMT9VFgD03ushDuvCNm6he8CqG
1BJSz7TKQ/F8KLVfRGdc6tqTbPGQxay4zGW5OnbWszBh1Sjr4LfzAon+PnZNxff7cOyZ2OZyIdYc
JyKUWrLhrv/ZTK93OyJ1SvnoR8nzU82QYJfJuIp+S2aU0wQ5dtfQV2VILstOKjR9jtjvs+zEIWwo
BOAa7WXkwSgYm50L6YIqbvFOD9KpSWGdUOsq9NfMbaQDQrpZpjVDXoR2DVLn9l4zQypeo0emZtZ9
TS2jmGdHJXirjbb3T/ckxH9FumoJBJ4lwvhtXej5QEhCHimnEEikUFbF0NNtAM8MJADqfuEbz9J+
JIlZvumU6s43PdIkFnWLlsHocPVZUn8gbPFtCHY/E1Ptfou/DmVq0WjD8Oz1mCrsIwUBFLQquImm
bj8OrybBNleyTnaHhN48luhxlDmjhTtUcSRRQXnj5s2lwfbs1Iw+cJP3qbTlaem5xWBYZdL8PYxl
8Oesx7JXF63/VdRxCcqACQBdTXrqGCf/t8OBezyxxhQY6C7zB93BHk60v9dcbLgHsMDCljp5l8Wk
OQQyyNil6itfmtRqvKT2tG+HZMgptflfh9uLFthrBDRr1Xf5rAr4W4QR964bRLrzE4i3StE9E1rr
S3fdkrvRjP1AUsXqCgBANekKyHNqKSH9GNJSNCS0OPvAEfkYZmfiHdnNejpT09zMW33yvnoJSWl4
n3J3zAeqgYZSCO29jI5+rvH0QF1j6msLJBiHWij/hJqkLzl5OjDxNLT0cuAC4BLSuhNQ5d47KxaX
dDc52XqnrbU0UdWN/351kr29y8uSnusJ6KtN5eL++/Fhdvc39mfBE0qjFtXiPmPnNnBxazmjycN5
193sW9w+uTxjayCgYMAbSx1b47PRlAdgPcUjnTQQB1h5u4uwMjbpTBIM0hSZpL6ESSxuAIHEGVXi
3S44M97L8XHTYTMeNQnE025qpiDbn2H8+XD1hHA3xxhSbzAURhWziiIjX8p87LhwpbON3lNXnW70
E6G5aTSlTNrZ9PSof4xr2BiD0Bb+nncVWa9wrFUQcsbXPIYn7B14FZ5m3Oq3KXfJ1l9ZGqCyF7FD
YnJO748CTJ28dd7j2kUxLkqdsAOnausi6Rad/61Y7fJ98YZY6DXKzu3tKEuDaU95hE9KK367BsFN
TpONC87AchOrE6XQGQJ6uHE6XJVFKu0aVCA6+TqYVwZ0Qz9iMxPZBsHSPru/VCbqlGZfUuqcq4wp
OvEF+8OqNZKACPrayU9/kyKQIQTrelFHihAqgferBWFlUyRUmGmUxPc1Nu6uJ9eVtScCZY7sZgEe
/5l7baXUaoGkHQgRmXSi6HkUBioZXBb0x8j2TD7zGz/WqPYafvOFx8z9KvnTa/7GK8uDLwK5DHsH
2uYDal3GVZ0AP6Xm/PJ0dJY3aYEmevX2I5ff1VGu88Uk1wZCP57fmCBvFMUwvix+wVQa4ZrNS23D
U9NyfP8IPNoOkt9M3Gfxa7yYQr1ha3jgfhPpcpFs8d7stxjm0zZikgGJhs1Lu7U95HYY0iw5XGXm
kmS4Ar2b+Z31diGrUymw+ncgyN40XyjUweoWan97meMn2mJZ5+8fcLL1NWAegIdxUKJge8SR7IS9
HfzlPpoNivI4kr26KEp9XTKC827Q68lw6i9+jXwVDyZKvbSp1Ep+zmHidKZnyonhvvkqXNRSlMjm
nnfShkovzi++VTLJhWPhSLJQC/T7ROLIf9LZv3yKVqZdIZyYwx0FO4OmUm9uMDfz7nMwHgT41lhc
gcsjtcGZND/okf3tnbbPvg/CDSfzhN59VIW0OTJSKyIzfdiXFV1BGDg3p62JwisOgWhglP5zhY5+
l5jKcp77PpbF8+kFzvVYVybJQM+TSxlL1q0Y/sXq1dc9tGRpEnjNpzQnM+bdyIkeNSBjtj10d88i
nXx01642id7prbabDTyotIXXSJO4BONVr2EXy+JpOK1EZ70N9cvF3MUHp0SE8O2+ar17wZJtpDUB
6kOOh0Hu66nHq3Aj/qQwsbi8Py+JrJuqZy+j9i45fHhbTL1khZW2MktR1Pecp8ONguQ6fhwgbd7Y
4Yr7Sw1d2Ke9TQ2E3uDKn8pUUdqyDwAk/uxs7gxDStyLIYMmRzsLJhzrYe/3VXGtJ86XR4a6zA3n
Pi6LLM33LrchzfFn0+1gKJ/rD3Ghth1iye215aOtRBdHNn/jt9hj+b+5zLH5X4BQlXGAScGd1Hf5
64d1BRwTqTDMFy1ggvST6STXrQh7gXLZa9aN2cxBSZTxtTsMbuy3DfC+rEy9RzntwzMQZ9mlPan0
TfSPiCoOf+B6Wdx66ck25JrRoR21sdtMuF4f/urAeHlbfWOiv7fKeMLDFfxir5DzRlOILyBitLuJ
PjOPmN42uIvLiC/WyGYqpgNWwYgXYAlYqgD9KPJIlMy8rTPknL+rSKw+PeQXXJVbQK1XirMoVasK
y8tElnWINdKrA6zBujDcEuJR8K52/RghMtmIenVPrUJ3zqJZRPlU2AYYUzG5nFA++mOvqAV6e08q
oKziFmr6IEgzxdrYvF5O9v2Y82PIyIcTUtOLKLLv3NfpoOxDUM5JyM1cuSlHFlIFnH5pFMZkub2n
Vgp+Mr6BmA7aZliDfSVFml/D9gYJ1p1xFBZPbCsvP0NvbvWGlY0HH2NwP2FR5gyqmzqsIBorjqtG
Pvki3eVKru1aCPfNvF+XySCrdvDtXNLgi2Q8zosxzSBuRhIVCZqqdReVugA8cwp45BI8pf++PQa/
urjUn2Z0Pi5OY0M+AKh7TqFvEFIXQCiTdF0VajqJmxJq0ZE2onVJoqYRwsuRgts/Qmu2N5wleCKz
iQUqPXPuSpAQC70OF4xGqIyghzGhO7Vn8BKi8fcL0uYY+vt/E2gICXnxrPkiHNLPIgryI5WbdVW+
hcfQr2nVhPc3bv8YQU5nqmX1IEkjjtl26Ygd22OXSqdDgdK8NLPYIIQi2x2teoyJKXlSdjJYoBXV
DRJndPVIRvTfUiHwhED73JF7ySMZkGJ+KAijSfCNTDptuoBt1TDnM51xj+YTvyxWe9EOOB6updq6
M7F07fwMeDijVDfKT+ja1bv9mqpQGhc4LArxo2EY/KlQvDnC146n6BB8fcjjEGutjLFwyOW4NOWM
2m/T7o6pBed1Xaud0qihUS2T8oHQ7SWorkOVcRMzWSYc+ceLMYjCdlfjj6xqUFqnyNazy9zEd2k1
L0yulw/fys9WLme9dVyQQcxhntnBtCYA4NH7wsEmEadyaVG4gF3l8GZlNswR/X3myJW1gLvjASpc
nVbv7ogDJfea5Lds2wcAt9P52QkZtseJ+NkxSVqFx2sHWLfPUeka/ujop0cjbwgmMGmVvhBd8bwI
/GLSbIgEYnkWJxSRnIG2jiB1XUWM/kYH8+Nbckl/4/jpCKzrgnDlfdrHDHpdqZCZedfvGi9IuWYT
/jsZJbCdIaEcxpfp1g2FnmJmwvsSGJoNXpD6B0qRUvm2eW3x5sDaclACNF0jLlDkDVaxL8Ws6pDu
tEmq00RJxZGJxnexG13A09sghJHK7BhPoRD5szdsrUNB3feqH31gG6EZXvm2rxFAWELFZFCsKCok
SNyYOhuaub0dKI/9TYoRBSIPGbyyYFP+NV9c78xNJv3mIdQiAsXIa0lEnPw0uOtziknk4SXjQXhN
L9umDYjrIy7Xtcz/qkKw267KthCIWIT35zvMKcvaQvMiY/a8Dz5JBsDJrt8tjK+fM8V68PTKl9nU
UbTzA/DHYZ5o/7YFrWzVQXGarhlUgrypFhkJ6c9Ci/H39hmR+dAJ+X14AGXuf3HTy2CLIoLfRki7
tCKoUzudr7sgcYzZu8n+aDg+Gbl8s0j998CNwP34KjmacLDrJKoKmS5xZOP5YTXr/X2owjU4AK5N
0fPIcaI7RVYudaJmlS2/z2mBjhwYaVcEu1tTxYHMV5uOGYXOfR4b99xzgjio0bjXLo5XESnZIDrS
RMMlRae8SLEkSTWTodO4r35YV/APIMiRsCYXQV3xmy0EsTl3HhArUFZXVtNX8Aml7lr2lPA6aNml
/50UvFJBySI/UONvibxoycVGgn0rllsBRpOpVcWw/R+2SXM7fBChsXp06vvJHC+9ltKyeG6bq6Eo
DMKf0lwO6f287SenVIqgbV7WtCxsYpbLjxUdUOcGqkuKfZTuSBpujNQe9UqPdOIL44f8PnRR35Da
bfxGl8fcjX4n73hSiToRRaGK8f4+NYKTAlHiMOMvyByyNhabM7PEWmtqAR3avjThqYrYrJ5AYY0d
8fbnjjVoIVxolkO57LWOUXjEwW3zF/g9j7htSO+G0OOoXThCCWThI+8JxL3CD8DTno4WrdrZKEc5
Tq4UqeDZR86Uj8M8rw9N7RgGV2roDOBaiLT98quqqZCRoTd+PxdmE4qh7AjrjDIu5liKLcUpOAAB
4xC/+HUYviWbkQ/OPQHZTzGxtAOTmJGVkP30X6p9megMsS3qTGlQ9Hujt75SfzMT7p3O6dvRBHYx
K7VFhm8OvguE2XmsxI4yAodBFSRetGbU1MYPz70M/eMhX6AjfMrJva+vewKwx1RWJdT9+XIX/vCG
6z3JENQKtjyysyJkT5yX8ZVYrAx0itXsxA8ChXR+MEriQvf0bz4pmdokTY7n7BeZvIZPLiVJsgwg
8lIOpKN7T+p7C3cf+wdGUNRxTPfOb1jzyFlL3PPh5YL74xMqoUbuolzfPq0kE7feXsBSCnNLdzAh
zRLMv81W5gnjUNeNoMOZl7JR+U1JJfrKAKzytcegvMiUbo2ZShOMV8DE6BJgAc4Z6DJDk1ziOnIh
V791I2Iv/mg7ZkGr8vtSv72nfWZJnyP8jZrcYVUuHAVhTtCd0qikJK1k4qr+JtSHtxyjfz3cpUcG
T5KotodtjuRCl9cvQhfs9ObmfX8V4wNuqJg+jUBxjIlb3nDbdIklxpWxd3s6ffj/nXvoa39fuaSm
CAt3QIHtWo9Xh6mikZXtLLxu0uQjY5OssFUpHENfNGQBLo20CVkNP3P2w12i2BoasWOCYNlitrbv
wpNBtW5oJ+y4fF+pGmozwKp5cZZA1kBomDUOFAKaW+hxwlW2pSLYnlgeKWcQPgCLY1PJeDydO27k
9NN16VuVgrJi6C9xnZqjLLgcOd833NmX0qe7G49rZ8eId0TyHwzB2+QQ/GMR22CggeImy0f+1/j+
QEAnBM3ShlxkKKHoXC1az/n3Fyj9AO1uYqZ9N8Mkx5L338AsvpIWNtsJCatIHLuSttrjBFIVFdCK
63IKoJ9J+mhpfn1lsDdR0BN1Kqf2JC/RDA0bvuuBFDZpX+Li4fXEgcUi2IE1GPfRoqTeZdB1+GB6
VSzN/6IL6oQAt8WVV3Oj+rjhDTjBQT5/k0qlhRs9uoP78C+ATHLqGqeO77QdQqEP2wR6EbBi8kWL
wRhYxJ8GO1aa9xZU7krJksuMXYEELZixoMbXERuGMEBOgy5OXzkMVD3zpY3Kgpa+oc2VDQB6vngY
l3sxZAUFg4frXjP6Zgv4hgZst5adPt+rRqVoaexeuGg9hsV9mJAZGlTUJOvgyB7azEXyLOtGkqKL
Ea/a+dICwQPms+k02NH4kAdOyVUba9Zuq6bVpR1zX4FJV3PAuNE7Nq03ZqtbVkWYIFDPBFYMtz5L
tsw7MFwSfp+wLJ6of5UEXfVusx1xmcLk2EA8cF3fry5LsjUURiyICOpQVxc8x7UjNDqLcDB9Q8Fk
f4ncyy0fCO1P6mk6l9NGtAeaqXyox9g/IWhCHOyXKH+15tdufLZc8ECqouE7X/dPUWGcAepeVeOe
vRH2PiB46svCZShF1fhWf5QHEahS6NmcMG2Xw3wkkLMvNMjLAyjfw8Zcl1csOGU1gs0PvHdHBL5m
fWXIj1dvABBG+gniqHcKprwD4fo7TXK2safckV9q8VUPyjzwgKN/v82D4oz7oJ+tR+kmtQofqAu+
HLKvv0GT34jkfkLBCYmS3LqSrnhXOnJ7jCuuAAWIa2idydrUxL3Ozisocz3Zeh2XgbtWpxJNoDwI
3OTFSWRwpMYhxeRch9NKYkqJ/y+lprWU4hPVc7c4OSo46ecDJjSW2KhgQurj9qLdUCKcbeyJlUZy
hJhpDThoBQ7FJbd8MO+o7RTP1hWxgeAg4Y9o6bq8czU1tRKTDcBP+KxuzHHjzD++bJMkKCJM0Bq/
n8qmo59jkc7EKNzDDMHpcXet0n2EZINO8y336p73guwnnR/f1e+TG/puVpTC8qSCko63Pa+b3OdS
LXEEnAKYcNiunsb6ZBjNw3rGzeucif3l0aBDHOtcomDCpe0Wv67xl3tY4rLDCrGIPEP8jQMw4fMH
J8l/1W2K9jmEeS3cYEKdP5kIvRCPahfnyKIqPyuAlsxiinMtudjdOeCS1f5GaecUWoFtt6KZG5/l
913GC9dXg8blsB06yrOv11Ge4gqnPKBN5UlR9MT4kTe3nQrE4BNrM/QBBZ+Xe5qa/3q4nGlsS+sr
siTL5zab9ZopIwaf7ZE+XMUfQcH2vZwOCfL5lfftaQeCCLWxl54Qf874EZoWLkRZsT73ud8VKWFO
8v6+YBJUGsA9JqxX9q7DaREKZdn3syIj4XeMZNh4X/xETHlq2niIQzPtINThcz1ktK8hFv6thPpQ
7TqRJaqZSCexZ1sY7DKoTg19NTzL6ZjNh6ViyJCaw5XEmKyYbSPuUeAcdUVIbYqc2AMwVXLPxsDR
pUAJlkgov0K3J6EbqHhZT5SCJ1d4CjkOpXyxXxH9qJJnRYOozF92Np/7ORSGcXMWH5P+LWQFrxWA
ea/1m2olZDjrQd84+zVYuxGR941MyaGR2AXB2Tgc35yKFdcJ23/IG7Bh/aZjR0I2tmta/On0SL9s
73NopQw3rWI+SuKohp0EnfOeVEG+JmJKJ4osQR2lz3O3tqukyRAaz6iN1UYhwYuqFMXnEcEMW9C9
cRQJTCtLiD8EBckztanqe813qksvcjGH8o29MLq89Ya+yNNCm0QlGluO2VkDsYpOn2S8IXrqtReo
Mp8ANlrymNct9mdSUZcgtgudeBEHor66M3HHmWAHL6mfPPejRHPrvsgla53L8x1kPZr0qFmnuODi
4QlrbOT6hIcDedXjwoN69nzoLUF5YEeP4MeBflF1e5BvXZASHgHRWUZ2UvFJ+LxW55gUo1dO/1+E
0d7PawAbkH7QkzYct4WVKYZFcnl/LpKTqeqpUjhiTJrhbyp/ABfFHwmnzM+LLdyBRmuPe2bWZm/8
zmfNWpwX84UBZ6OonpbenydcxWJC0DGM8i1PCSgYMmO63xG/zLiuRQ3E1Ig+53z74iPUKdOpyvSi
CwzZbmPCxbqNFstf1bNY1JLCEn/UZc46p7CcH4NKadJmuTUQgF+aBS3oSTeX8iojAcA0in5wWNhJ
wB5XvvywJ42KVAGex+vQYpREdLhv8z9wN2fzJfsC1cMBnjDtd52xIE0ByonSQATAOI+w3yJa0uJn
L4fbM567FynXiDICwKIN/zdpnbby7eUG2HelDTkyL6suksE5kKsgmLClwz3JnFOZcRT4i/x9idpN
Ch3fr6waXRb5cED1eQgjo8izsucCQ8GFK85Z6HxZ9u2LqTEyEj/YK3BQ1qf6DGNhA9ywiKaixn3u
Ydjh0YxFq6a8Z95o9u7Nv783zDyQVmOZQTu6fpw0AXMS4r3Z/1TMGfzkxVBQF0DC6Q1dkYZ1Q0PI
xn1Z3YzX/Z1vo4dmR627dWAINQfVB774k6wvpIeWQZSI9jFWcDC2EL9cCX6AVbV3UBypKzkqz3mu
1/SIgZb8EDJ+IlzQGWkUO2Fh5bPLeHgqh2I+J7uI3u7d61V2KzoUIa32M2cZtekw/R/LMYy71dHU
z/WRQXLS/6oQkZ9sPV7r9sfCDDSHJo6ohuKRC9n+8C7GIzuk7NrF06awts7P/P5rZOnJF4FN5Pb+
5dTbY4rNgfzliXBoGUnZ3qwkaEGvuXl1uxr3ICdFV3aW4I556YcgSJdPXf4Z+scKFkDb2Hf0T7Uu
qaZRDDFOyODQjFl42rIvuOB6yQVU8pPT6VN3U4dAsrsLEWgRAG+9bltCFGi86syxXFUGFH2KiTku
P0khAefZigWygk0C1Afp2CZNNetTaC7vX9y8Qp+DvyWFtdsuhdPjhVMJ5Z3PL7IWrttWGkOire8t
yaP4Rk94GsQwjLlX9YksdizmjuAOGYcTghw4Jg9EgIL9M0bZtrbaE4mFgk8lhOKsdKSh0AV3tQgP
8mad9R1CFm5ETwlxPUPh/twxnr3XJXOHSi00U6C2YXLLF5ni/ozB50y+u9yqfbbUVk2YN960G1gg
tYvuwufPyDAovfn0jI5sa8XtaLnPmjKD5MqStTonaRT5fau8JK0BG1MTI5eII5bpVa/1YxTx/ZHf
3iIZ7+zo9xq3HZxqFxg5OtwQs9y6kXarli82NB1aSxoie8oCRtkcw6e4gEGoev5YMRRnSMb5d/SS
pfzAh0/ZkjB2BYvJ/QO81kLsXF9sVvhPzwT2RHiW3flNxIMl1VOu+hc2cq8EJiOJMeA6K1/iH2Xa
Bd5tyKeo/jDtx3x+qjbugphaxLs3MepRVf/hQHiHPnA63OsYVluEmc4InAAPTIReAs1318o+EpbU
KPOKneLlX8v7xybAph96W47cKxcXNAO+kW1zhVEMR3LCTFr6o510iuZSN3DGULBsm+3EwoV5cply
7g8sc5yDnolpCSJR2TR9SYYeoPHNo6Yjrk5A6MbEDHoV6fO3P0MnfeGPPwNCmdSDKbs9pvpQonOc
yV+AeZ0jJzO0n7gP0OTCSwrnBZ2xQAi27o/ozwDOY91EJF+V2EcRA5ynitqprE+qLQZ7d1tzEsWm
2ZXa8SOrSuV3yPXwGrmbK1osXpC4N8Xh/kGwlNAZtWlB1hKJunvuTuzQruwvQaxkdpcXRoDepZTy
bzz7q8+SGdM+0vTEjDAsJjiFHd8SvUAbRlAzfkytEfeF0k+BVMT7aipJt1HIi+GOHxB6T6v+ieht
JbO38OvMzr4qiAw7NTKCpsXB8e2qvfU/dylsKCFomNDvvPz5v11b1Sx++008ywvI10E64S48nzm2
govHwmW05B9BN2EjwOqM+Er7LbJiN6/aRXvvZVTz2TqXfZPepTXJTm0+fNWCYCgCmcm9zUV3ZdRG
IYqRyugjivqQQJhI8VimHuQ7TPqQiZkHHSeeRfpsuOUdKnv3bpiRJppCfdvcJqzenVnH6g9vwgsC
1dMS1XlAG1U3u9tJ6LYhAl0JXXv47/iYa6lCe/SIBdLh7qCoA0I85QWKuaJYYxgG6oN4FRjfaGO6
F7JnItl0qhuXAZbloJLVtRvv/V/afK0Kitw/5ewjtniDz/ghnWkMzf7sr0wV+0r5j4ukbeL8LovS
BOCOfmRc+2ZJTxnQl7ZVvqrbi8XITHWyQTqQgI2L7BoHtvJGi1dKW8kHFFSowyqgyt3dSHCTmkZf
PvhLzdpQ7pE3g/Ntl5He5xuLzPFvleju8Mc2/9zqoe3VaEqLSn7yXSfzZnaX6wk21i8VVddhGONa
3KmdSq4wTq2ZQ45QhZh0COWBgkYl7I4dW6mjPp/mqSwLKbgku0GsK6lKN77ZslSK3U6XbphVC8Kd
smNT59/TE59Zv6NePkiQueP7WbZfkjZRgjaDcp9QVTrpOT80wMLnPoHPn6XzGjzVf2C94LuKaYfw
a/ElyS1HCpDkR+jeuITzl8gNrPqDsEf04/AiM206dSrrr3FdlnlSpP+1IBUsP4Pyrfwij2j8vD71
i0vkNigGfF2TVajoi17TvAhi0uZEA5ZFMHw1RVGFF0+iJrrYU+qULfVMmEHJSLRhDO/S7H0X7Vzc
JefqQe3Anbd1jIf1vk9YJ0gYIty58pjfAOd5sq+lLGzFlHccW7NZY93pwm0isTCDrCcTpHv413KS
L6zOE+e3y7cjHMJYO6NWbsH4VwxiF8SOg+Hwh9l5fDgspcqY0UZn1Jw6hohRfQTSI41ropR6QjGG
bHDDi/IyjAKlB7VywKerM2m7SZ8FVbzval050zIbvNBHZ02lgH35cV//XjURrqpc4vk00mLzdIiD
znrwklfnV44cRNfFsvfEXbSNHk83QeP8ZJs3NH7eFobe0xrOlb3vcDJyl4ES/PB/Kspkw/X72YPt
/PQgaQ2dackE3tvg83wI2HhM3+GXwWl7XQS9dm6elaA2U4n3z0lC47G0y6A79pEtXF00dPNYTJDC
aHIOS9GMpX4YfgMssbl8DMOHPnB58yYdbea4MfwCtHh+rQoJKxUaGm9d8XUeUssx4KA5MtEb75Oy
bqmmWyrPnvrQfBXt372rNxcrrQzLQBidYIyoZGsjDjzqkiNEpnlm5FfDUclSXMTaIonN1wAaGfUd
0TcR63v+u1BDbpF2Z/kB9Jk8bQZv7aLmDiY/5IxzFtVdROoUmpm/cT7n9fkJVbVFq1QI8uXJw6cz
P5FDA1Z8aNIqJq6+zyISe6epi6E6xl2JvfeWPKm1ZfnyXaj66CKKd9Q6qQyXmrdBEzEDLoylX/+5
i4SmeEmgxWTevnYeK4fkPRKrng6JZSXwuPF8M2kqf4rzgIO9w0XaIdjSxA/+WJEMCPUmcIGZAPWw
LL4fPnpzt9pApjX909s0IKKfaD6I8HKWHyRzVgOkb931KfvZEjGB1v+sTCjOKI4VxIe1te4qyB5g
iRl8JDy/Ft4dPr2RLOSlsg5pR93lWtWtGQusW3x8OI3GZyzrdCo0LlUjUpi8/7p3JRdwA5Lfq+Qe
G4fIAeyhNtIWcHIeFeiNDaFigFUOx0O5R1wUPrSvB9tpKICbRGEcOydIpKi4vV823RHRAtKo1yEW
sZN/L5I/ywP+elyKaTGufSlhZNUxpOd/jo8mtv6ZdsbCT2uwHLH8u9yOy/jn7a+ZZuN+PeMNGbQA
CbhCvJgJSGVTASbxXxB/itPyxEzT6jJ2jtThXB+Y22Xa8GXwtynQICMbvug01XFvn5mfQG2HStys
gx9cKLSrhPvZGcZSqyHHL1c1IiT7AAFGy58HIozsShHqw6EogTsuNaQz8H2lThClfG/mdkJfPqJ1
cEFUSEnyMZu8S07Pn05ke9L65A422BDa4HgVM6AiRx35MX7PZhuY+yNk4tWHF/txbpKiq63Q1Oo2
B0X+a2syUXdEE9zjumOJ7oG/PFvCGiKhBx+7KiMRqlfkzv/XSHg4qUeL6R45AQyJlCjxFWh54OCt
csn9bbMh8GdjYgtjP81jFVxS/mdbwA9vIWPlYe60KCWKTpGtp3S4r4acIcFdDMwa3yeXMll1opbC
diguDD38qGIHRRIUgylGd1Y5ypU43zJAOR9t9MH3Ut3uk+BbnSrA4RvkQdQxkoqm6WHgSfLc81lt
Djo9na18uUbqQuyJ6FGreuoOv0JFsmU+3KHm3TJ97UNEx1UXVLBghpW8xFPfKHtpPUN4IHW+znzs
KY2aRvCmdTVQrO6j2VQKbB0yccxcCCgn6Gk7283KqDLH14jTln2AUanHLR2aBMgk8AlzBFVl/YaN
ma4g9YFXQFiL/PCKCPyiRR6HNxNGJFkyWM6YINhrguyyt118mGBxKW20l5kQWVkYdnS7Eypw387y
BGmmLcEF+WKmo7C+s3c0cG6GyR+D0IVItuHJYuqnqXHhAiNW59/+e50zbZUssFYtzAEFwWFdkuS2
/uX7djprIuHk7q3b/fH5F05qHyPl7And829spXTmZg+dGC3JSXCXTPNHn1f4oZgumUGdgPU6Ipwq
V3HR9IXtjq5slz/3zty1bxfKvzq1ci/i7SaTWRVAEZaILZ5HztYy87G6UTOiXwdRXEfxcG5xH1sk
oRBigT0XzuG3UG5OhoLmLltWiRPtx0wvIODPwr6QPjACMl4dhK/Hj20TQLXADO7yLinEaXfFDMCD
wrb+P8tj60NrFughcD9+b1AOLvXzOQDnxypLmVovTflr9RYFivNQZEKWpyPCPU97hteGd/Zx8B2Y
uh1IGXeC64/jnZnoPTLCBoL3XGrJwvwrLQVu7MQNuXCqEPIQglP3jvbGO880vpExfwVjQ6KBy0nf
UZReXcmS8lTXoWqF0IHqr7V9fjJR/1p8riiRMY24qwGC70NhPg1tAWL5DgkBmKUp1FnS0aGjrsHv
WzylKLUxxLrZlnmL9WCjrzWh1A44XBNTZq9sA+0I6ptGmRJoR/z9wZ3Rcp1cD5PAcH37qvCUKzzE
IE/f9EHekSm7vDj6MnIZUW6oNT9T0iODNLp1TdV1td9MfBrAxosK7LNpWosRMJQsk4L0KNaOuh3A
MUofGNA9p4A5Blp6+JMF7rQiJ4WKVlSH0xZAcq/OINlhr1fka81fvIjgJw/7RQhLbuAviX/EHWNm
lB3sk5iQNPShiQiW183sT7IT+/yq520FNm1JL3e0tlxvnICrSEdyv32RtRj6+LQ9YyR68mDv2hCd
dMr9EK5A46C95IFZdNRGSjew+PNhMy2VNJzYwCFvRdYdGM5/BXw3AUN076TL+3Jeh0flrGYecAy0
Uiv8VGnLU/WfoFz4/tR3747YI0fTaXXAA8lO0q8SQ0SDADdQKC897v/QxPpPRWqUFX5BQfyVf3xx
JBNZugZg4nFPFEl+BnzpqvOi0sqHTAWPSpqF/ZVeUEN+V9FPoPNpxpTOEEFE4oNLeHLe86E9QLZv
h/E5dpVk3Z5FqYHTh2WGuwFgc4c1yWI39eD0XvX45P+NZpM3MixwMCcKI0Q12z6gdRYzYcKCjyT2
OmRmn2KKtCewAz3j4Svzs0jMwx6VWcHRV6CgC/t1h45KEuCILUYU3suz+uCkk/l7NZaEnsoY3wDB
mEXQAS3q5KV2RkxerA0ePcXBK0nL6Q51N5aaVYthnwh140qDjZ35HTRWxI4L8uiOljav0aGQzbY5
BxzaWb5JTHIagS8sGzldWrnjdoiHysrNJWg4KsKvXGGEkXEVJi92lXCPGsz9p134raQlJFRO1N38
yCaecwxLByZHq/kv4nIIimutSod3WlhMoLMewPNoy7z3lEnZNjKnj7lRZf4TrtZCgiWgswa2cJmu
OZt8S026/ibs0O55biO2RrmucwXclg/jgk84txHfimFjoDpqFTYP/AhBSF1IwtK1BhUIv4a9lh1Q
4amgYMbqa/h+RDFBuNV/fkw2P8jL8tchJRzpYe0NMtqbxeU98WTOzDVIomYTnpXUZcMNquFRZyxO
DfJ1OejAc8LsVmUTfr/qc/4txJtIAHx1JhPIGVc3HH7B+P5iT8VlEokzghJIZkZU3xu0g6EG0rjx
7tujjmeX/sOfl9bNy6TfoLvw67HSiGdQetYcEAORjVD1tpTC8auhZZYPUzvqNFrpmiRRjIouC4lq
gh3XniHcSwHnyPzihCdjGkgd2ggXISclfTyINagNELWFNuWbuzQM5gnwvfQdXoqQ6zZ8g/+lY1kd
XSzPkHFtQjfLTF5EWmgn8zvCdQvNflcWxVIKNUu9o4Kh0KzAtihB9cuCORrM7YIxKq+U7LHKYM5C
IS7zZgAdNnlZpxemBC6OASum/5ij8kODgN8aOulV0JaMrh897vpP6X4xoCJQw/K/FfSS6+6CZGEm
VJ1LqIs9Pq6UMkJtJmKdFGWG8x2r3Md2/UH5T7rQaontRJovnfELW738iMO6cQwXWw1ry9etb3rB
xWAC04uTTFKcKg7ZHDX2QnpAbENa/zuP428UdZsGATZb71A4kK3wKvzFDE3lPKQYcLOb2XcQ+Ou8
pgkVYhUJoQFqD30nkk5+I5YugwMTFg2G+508j4TEHGhzvGvdL9KeM37uKsLKbnLTgWC/8yF8NxL5
Ahrg7uVy9BO+yVN7DEoh0VtJPD/IW7Py8MWB4DzyewslgxkjulNmudv0HYV4dL28MJfMYnIAhukJ
YSRDm3pr5iffTLu0hpknyLcuSnOy66oQYHmSNVVNUXqLNMEaZ+L9qjHUySHExED4dsn/ANmpsshF
AGiRlaOcBWMF7v+e6JWVpBiGPUP615hUYz38/09ggpLM2Z2VTc14hvpwWtYwsvCI55GsT+pMDOR2
Fg5DXuGvRok/eVl56hQVQy3SiSFwO97pTHFQxvyQOdls2UyRIyjwoWrskfiX2Bab0rSoMQCKlto0
j5W2snFloOC3FRAsDY0QkNsHSbq61CAIGOVN0AjB/imy4lU0jC2cmKYbjqZH6gZMETa/6dohGSOw
saYGkr4ycFlFXQ+6AGKRqmitKFvnZcUmaoTfaiUUKZTMr9kLhyCJme4GAtSiF2x7v3xL+xJBSgV9
1MahpreoIe0rdmohrAvInfJl39TWJcWVvt9qhwSsCyokR19zEiFKxlf8K6v4ySbKTFiP9mq+qtC7
YOre4jQPLZyAYGIPJGqqOHa9I6o564cK44//R+vt+Q5YeKq8hJBMRsC+duK9uvrn91PB6/lp8OcU
RgekYbxHWs5D5kMUr9xsx8xdmhCbgs8qGUvqR9OrKtQ4RrPyzsa/uDx7Vpj0PtDtXCx61MXD18Eg
vphnbEffcIkngW63RABQUedV9TRnumQlbKh5yLipkaNSJCdFmWAqznKlFJVtddGWiXnk0eMPtWAC
cIRaXfncqXStB6MOiI0DLruOxQ/pDok8q4K5MWC+UMMss1EJVa2XnsBesTg3vTBXGVAP+PbPo2Z9
yOaMegUumXiUA4mFDId5DKzF8EIB46lQq6gSinRCWG92WFbOoWbO/A3XAJwf/hbvn42QPp6N2yD8
O2mP9+ClCIuHLIhjjd1hawz1eYcCpEPO4n+9REjVaNnzSQmCrDTNd0CepuF4p0U5u9gj/4B0F+X6
A7MTChXQnKbF9ph33NcffbpBKWllnHzCSdrNmoRpkFL3IUmaYWPhtEtEmsvdbNWtBH5rJt1PzRJ4
z/KuZ9UO4wdaSo5KWSk12iWksXFx/+Nrx2uk6Y0X6+JKDIrCI7LTw9vp+O3IhSaC0gXtcbeBN5gw
fWLOmboc23wNC+KRqBarObaVdKuL8GxpO0+UHwjOegyk7I4YdSj5Y+wUBOk6n22bIfRpcl2UPJYN
oASpjj+ocbRjJe30E1vlZqnCgn1jTy6+9uu/CWQEUZtSIJWykPXHmgZWR0Wwi5xyss5dgbRArtFT
a6Pf2Fm6Vzc1Bl4sM5tU7pUcsW6IYEMUiIvllbDIRd0eqP/nqKkmKwdCtS0zqARVBssEeM0fy48q
LD/nICpVvSMngJmeiMbqH+VMb6OdhShmJo8jw0PIZuQkYgs3OqbiiGNAUZocCiOx2zmL6kOzuV+H
sRjlt9IDiWF55CWu75hrjQWHlPT68iVuYfq73y3LAAPT7XhJwkLtDb85IbnVEx/k8hx9OmQFWSMH
rEPOQSLPJmwgybNdxmorLViP+TFjdzVmaL04zFYnfBQQp82dGXrii+RxLKOfXaIe6kB7rIPEQ8Qw
GPTc/VTJrjEdb77QY1w20+yW3StuEDLbXuCC/gmBdNE7i7+efLJZU12ywO4uQON9/aG7u+YDB5Sa
Q1Cm0ys2fa11S/gXTb8mghFnEFm4llFaxnqmH2pf7Zof/Lli086GecTTtzfKyzI11pBMa/xGSrUP
BjVJO7L/mgNiJ1mVeAPYYBYndamqdBbE1Jlj5ry9oyjYKbYa77a3u85x5Mj7KRBgSGooxIjCrwVo
K5V7G4h5g4T2eejTYYCGWNOsJPsz5kwa6VZGREDG3OuU9NN3XNuyk9QSaI1PNUOJW5cUUURrYUMj
Eou4KiqJPxso3nJpUCw5f1+UG5lOQlchJoSoeGesJ8O9pb6cJ8D/92/XIZf+hqfkvL9YvdOtYpLD
UNxrTkNtQpuoXc+nANdIaTwyuRVpCcJBmSnsa8HgROKAUUNgR2YtlhaEwzq568TSBsJu27euQdtY
Wa+qGtSLG3iDBCbrOAZfl3/9dHYOh6MoZxfyuM35xANvHz0ADhu6u7MvAwbhX263y6tVSZIObuuz
4AUozy2uZlbmdI9yhhgReqOEwOaZ12315eFwRcnaqhKSEMEq3UBTdd9vuvl8pWIJq/Cx+YcWhj5z
HLP+89mVrSp803zpoNAfudxCUKWsZTiczNx8XES+0UJMLhdGbqruzbCqPO7EqSIGIRiPzQHFFf2/
a57nH1aIG+jSQ/RBHmfcYHoTnBlYvNDpTuhHNLJ8l6kaz9+XGOR1IaWYmis+OXeZm7cKdd8kSvRY
2BTuR1wMniWNkg5/aABiJhhdodxZJkgg9nS2g3o/NHxx5tSzkx37j9BSiNxZ8Pp9cmOyJVj76PrH
6tIB1ciIg+yG7+Rtd92JvoxWFpKqK9EhaeXKj87bU8+ENSW5vEuTCxQVjJu6dBhOhFcGTvE5PWh6
Ka7U9kxodUtfL2FJl8kVxjL/hJ/2jIUGTmexYFFXPVYstSeujMI4FVLflF3PQWpYvp4pJWj07EC+
jHBGVWW4kNwxvbGICCXSK4khP5H4ErTtyBG/mpzwMjHK45mOzPe4ZcMnwXRvxQxllqm3kk9pW7bg
t+ZuZhOi4gdJx3te/90ibNuUJPWuvi4yHWenv691fWgvEzzRwnyjdDxJm8+E/Yt5CeKQ1LJJdqpt
p99eLiOECCvLkbdSNmYtyyK9uU05clu7dw9NPQBejouWlfUZITUaTxFjahgaotxfP/zr+UrfTeyX
LxEI6cMV213oV3AIAlrxf1UPElqWRVyrN8K195rj5853woUe3FFL6vRslj1jH8SNOwcCY/78zZpL
H2flg777SZ8WPnAWL0gOHPUJUMumKcmU2bC//DYlAc5FoxM0vFSv8bDYGLAbdH1D2cfyqDLzJT6b
nGAGYODAlrxO3P4gurSaB4SL0RSz5IQQpTAKA/32q/nvV1vNQEJIZOJmcO9jrlaLavqy3BhDdBCa
GdyJgQIjj1DL7vD/QL7jy5ijMH5GRvzdHwE+FoliUy6iVqnkCe9XpMWgvtZokmoeOl7XcFJMD5PH
1kYqDQqEW+ezyCFB3MzfusEV+8TVSOGRx6zfnWYRQ/zCUTXjWCzT9sRIfOJzmATRjY1LCeCs4s7B
15c9RdmLFebgsN2kmwlUmXzLUgi4KTIB2gR/4uoGK+dd/Qnl5WrPDm4EWzouLAHBv1hQeEeusQ1Z
AL19/sZooFsTvRnTl7KPzqHnzLOzMutSvcrJoIQZQlpoKxTnrIlznYEJpdnu/WhaE3RZN5umkuw6
UGLdcPJyXWBCNNCCTXugEGQrN9D0P38nc8J3zmk9p4HCOoxWCfFQkKaccopR9IiAzQZaTlJGUQji
VBG12dS2s5V+fFB2qGJLUmCMvjKibOFJd+6P53t/zIENVe/PU5H9OyoVrJR+SXvlyTTNQLhatEZP
Rr3ncuMgdGlLUkaTNSuCAvY9enKNhIIp1WcCG+fVOrqXaJoPsElf3SgwYYFxYfHIzj4bYYc1sbZx
2f4HhJz4u9HUABwLIyM03HH9+aypqmCSN7K1Kt/axSy48bcKJvzfOFz9xBcdvr2u3ZuzysXxyKJ/
A6MP1v+EBV3DenCsE+tnHf8uv2OvvJt/opLGN6cvtLfXPvbN4eqZBtmbKd8icM+WXn8LweqU8ZHo
4al/N6kQ2HtIzGitoTXqjhyFuk6f0Ic6omY0nJxB8EZQ95zCaRuedTs+dbquvQecg65fAbIUF2Vr
cxfQ5OqV0y7y+cdTpVuWZneAlfOmt8vbhrBGwXSOFSHE6XstRhkq+6F7DE8Kg8d29OWd9uWzWYtf
TM27g7BOO8WTLVbEfsMS9hVQiAYyeOS6MPDChPBufmH1Yt22Ip0G6TNRqVGXJCluBcRsh3cnK+jq
3ADVsfsxg5ykvnAvr4PSFmooRNufka/aPNKJ/Awn2JcHTIJ5CS91dHblXJ68CGIH08fk83uWIsUq
9Eh9TKsNCNjF8f1wpFK8q3PsIzYKl7TDHBxBIakzqtdubP8YqcoEcfOoMmaWUmfWOFVTSHgsK8OA
ghqOltYBF9Pt5SzP0uBj5RFrTvzJ5QnKkioaYG90CqF33cIo1XlJzbmCd0MBvhFH+8AukFUWNrHw
SZ205I78GiM0+yvg05rl6XtgKoQ9ZodHJsDR5jLFtucMEOj0xIvxHMvPrIsEEPki8kdIxs31tKU6
mGFH415G6BLIommTFFlHqbhG3kehfkn+vtefsKISyVhhBkR0nz4lPC4LeNDCEwPaONdbrI/P8vpr
SMhivj2IIpUi4yBvm6/6ZkSgTJFN+hvYtDe9moe4ONSkMBwXVoyoJ/3byPdD+sMZo6zvyuDoxT41
YeoP/tZA0eyIsm0xQ8wSrJYYDPnv7CV1FuKRvLdLxEjPa7u+gbIjjNjALSYYb5vZK0uLAdqISVR6
d4FbDB6lsa11QI+64GoO9ibENlhLIL1LARuk+aARnF35MBUOs/zxNHeD7Jv29nwZgAlxF0vA4R4q
pe60gjOICJoKzKyczyaczGlbO1KuiOTfmjIiXqoD1vCaZgWju0vrHXvvrUxQ0tkgW+zCQua5novR
iLqUKzhMLpffOD15jK3LsCw2659ezJwQOKRPr/QkFfvHHlVtz85G/l0ua/npu8ILRsfoZ0QbRcJc
tVEGIHe3OoUqBEW1MZwMNFsQYezeXg7n0FUb77SG0F6pm/ndo0vK+cLMJ5F2wh7wPyzBiFDCWBGT
9sKxCCDx8XGGXzvqsb5Lbk9ZYP5b7nx4BvmwVnHxO3lNiwiKmNfRLv2V26NsB8zhklBT3ImIs9po
R0Bi+rhaYAI3bSKdw38tr460vsQiBxt/H3wRNvDN0yFmyq+/M3jdGyawKX2I0CRNTXZICPG8KibR
2rlc3bQu5qBbaYPvP1SNAFmj6f33EPczLHAGJn0ug1JlSjyCMz2FNlRf8bTzZEGfi/a+TErExdOG
qfkMo/XWXiT8nzCvxa3Vujlkrehec4LNBGZ5Pyn+4TF12YU2RQBpZ/t2SquGUwj+4L6S4B2w5MPT
3vQMupvgBJLydHQfpIxmeb4H468cI4lcgHMaWKNHHhmMEzZO/MrPUqDpf+uaLyomjvse+o+Tk02y
bgdyAknGTyEzoJtKl6B3MdDPNx3zeUOYQI3SdG9v5k1HPixdr18Nvh68K82Yixho8uvY5NQvRHDY
zQ20R+A0Y5/OVXaK0wRjXlVHTPAVXt37Dfn5P6LKE+QwKmgQ1XAseewW5CAW02HouSS58Sss8Vhj
8TMjIH583mfFQ3nTY1Rq2nktavovmUJpx6nAa6WB/Fw5ulKjZ0j81EsORJLlQtQ8H6tIgLgVaEHg
5er7/BoBZJXw0ULN7zBOEny5eTDbEQwWUXJyASdiF0eIc2yInGoHZgctqZfAU5/8B0eGSa2x8kMF
coVKwF1Gx6T9aahhW7myRyn6sUEpprbXJ0thZ3MSLXL9sbcebfrE09irsWkAcm3Kcklxeh9vffwA
1ARd7W6T3Ntc2jV4JswdKYfA976c9Axhk4V4XX8AQpegiIMm1K1njUHDaCygkaLoK8nSGd9R5JEZ
jtgkWsUavxp+Wrps4IPQgrdo6wmOH/LWVhIeRECU88h+wFvb7SurY1Tyg68OKt/qdOdI9prLnbuV
34y+WESmeC48TD9jvN9qyFXoZPAZyCTSWwjduaU5F41Jjh2MZcAW61GakLqpBUFtckGG5rP6zUEd
T8Nc+bdVqVu16CPtL0YXm3jCL0pMuP/ij7458x3i5+tb4G8xIQi8GCQ3GaUoEA/tUqc/1QO1B6aN
HwtSqZHSs5VDBGgKDH70MiTlIsbi/em3swj9YKX2BtuXmv821jp8EQeHbDYplAS3BP1DgTdZ22m7
v/dastO2dxne1KxxTamhC7QnZ+gl2d0MFjkL/K2xnzC5179CzjV3zTuqPhRe2uJNq9tXb4LtnwZd
J3C7RYZXN1LQ7MZ0Fe7HfL3V3OtmK1uPQ4/V63MG+mFcoMwIfRL/Iw7modyEqg7Bb0zCFjF53qAE
vece4M2WroDUGM71ca/UkpI25j35kfWpLBiNidfP3MOsQu2XcabTMiU9x/4IE2VedjJTn/3yoixz
e6epXBH5MZR11AgsqDyQpkFz28SYnPo1hl5OhPuKHzEl3pxbIKVMnLAKkzLmzS3J7jpkxXDYS4f5
7IrOgjcResxKPwCqXNkYNK/TSvHwQLQ6pOWXt3eiJ7i4BinkGCZXDDf8OHtjSX0AYmtls7udHo05
TqaqbDBVDR0tURzIGIxSrYfMzNvZXzONdhdOPckZEnSa3gNoZAIhYYQ6DAVXqzm9vuYMNCX2Hyyl
/XuRxExox11qFkrabawse4Yw5dNFLOjUYPLV3l45B/IzBQZ2smMfcRGPs4hsdgdPGkD43hdVK6dM
2JSfvNeA8mXnxNZAJjR1CFOL66ZEEP0sStmmaeK5gTA/+hCw6PCEDWXRoDOSrMVLAI7a5iJA6V6b
+LuWTbbfFD56oV48MfapYuzM5bO9Du0N4wgcDc7yCpIionAuIVdZUbf2LhTzhRLQ3Hjl3WCLcshl
H8q4CJGO4MtJFHeqmhaN5RMbZScWXwaYXmwRb6feheYiLzVsmcYtceiiLaYr/Ob+3T1MU1vg+Xd7
+RARwHbHulbpyq6s2j5pOuwtEjuP1F5pTQKEIG0YgFEcnUDs5e8PlqtjQ+0RrdlVe8zMo0JODiAk
DdRdba1smegYIqSRVcLFhnADjCOmH/r4FYW1F9MLwcMkc5QoTq95xXD0Xz5jKRDdj8Br3SWmW53+
UaTpVgse7GmwZdlDiC5t/kWANPWg/XEvKSNZtbzc7SCbnPnmA4pg2R+1tJOuISfupwKZ6P0M5z9O
/T9DgfAAf3u3FP1BI7z1XO8uI8ZC7OJfYU6N6muLwK1J6xeXQskKhCTNEUggs8Bw05cURzBlfFg/
7141SJN0dRBh2WN11m9V0r7IFzkJHcgD59EA6DaB842WxhUGrOaQrKEyY5sqJaN1CBgS7Q70/PC3
DIXJzG2uhI9HmmTsiAOzXp34btQuDpWf5iikAbifcndc+rELT83qjsEpvA68Q7OtorxswxTZSVPi
BCuSgC4GPjZIb7Cs8xy5TDNmW8fG6QecoIb5KBYwOgy75PKbtajFJbdx4Hla8Z49+Gsn4drt5Vqq
fy0d8tNpsiYxBZJiqQckmvAKHwltiiOmjOfL7qOnIsmqd2f9STVGQV/7unEgxLiJk+2QR4z4G3E/
+14iq8pG1JC46Ojorq3tsmxX4xx/wfshCSbDNLTrvFL55TgA0rQk9BMTvGVgF7fWlSajnWqilIzt
Z34WGMBS+n92isbpvNk7C01DldL0ob7QqqCY3DPYQJ8ngKEprBEhKoo7jPgd5SQ++Uq2fOOO4Iyl
vmEnPVOnC3HoPXcn10qOPAVXgtaG1y1dKL7KLW8WZC43srco7RIXnGECMBnKB8yv3cLaEy1p4YvV
DevyfWwzx0PesTWArojfbiOMQAE4ZbwGJyC1DIBAw40yDa1YikRvJ2leXVVmjmX4FUdFvqwWRSRX
74vLo72epavrCxuM76Y/2YX9dfcw4NIfslFjhMwcCStjnpoYOY2wINtpnvXyHIZ4ST/1mMECo1Fg
IvSrqX2VGDbpw2ECMSnop6Wnw+PG5vqQ0D1kZI1xpcfdgzwdmtZTvPKlCgzBoHULeGhDyC6KshXY
/W1lnE69hZsCyViVQo2ERes3PBXhpgXAp8alb5g4dvdLu0+xd+sn293kEiR/8B4/ujjAK051C+6A
cCdAeIdPMS7rEHy7qncS9HclkTuFBI61oUE+3TB9iY0UsuP4FLfzWdgpEBY3f/eZsSHbG+g6bX0C
7LuOtSFNORMn9y03uMg+E6wJ+9KLrIwsu0Q1M3a2epZ10kbIe91+VOEnlvaA0fVnNvWXOhXbHvT9
0q4BnFta03+hZZnAmGLTkRq+7349wfugtSueTj4l41THj8w76D0wkHYvZwK13Ilp93jm/4CPh1Md
DlxqI9fHELlMKHKCyRFes9yu5+OASBTPin8x7o361obDD6Y/iYyXML9IcW/C/mdSlEv24xU3rgWX
Z/mHIv5yOPXt5Sw9zzvE9t2mH+HrdzRoO/7CXFiqDNFyHVChzsmJepTrA0+A573febD3HdHGfUvv
raiK7QT3D8RdI44cW42goP2aQKolvO24svx8Cpi3imAxyaUniIZPvZheZfkYdv/EVSY78HvYZ7ki
UbqyicgR2NR0rKbRCuOgVz5gTEEeq0HD+wbyEOfeLqlGLbXVPDJRQsOPoyHk3so5PlE/edLn1okS
oVCk/RitG6u8OZngIVGlSi7zIMRlbL2HjnPauPTr2u9KJvkhQnulVKvLZCigYJobSJiNDZhEPbUs
Y9N/4jRVVt773U2ufmkiynWjJicYdrf0gu7BY1tOnZlwvbroxMqT6iAvTeQLNWfwgVYrqQ7rOTeb
yovMYFw48xXsYIo0Z8umYmqCXU7CCcDk9Bv5PBG1+GiLq+DqgSU6PWNfv4tNJM3GLpqdU6lu3FdZ
BVJR6yJ5ZjOVNfO8ILoQ+jBcglNaX2kbefIeDkNT38W32WUpkIdJGeaOrSomulMZoQS/jRbwCoER
C1ru8v6Gl+/cWJ/a9VtSeim2IFDbGKZMyoK2FUmwm8kQINs15Zu20gU/+3o/HyWrgRCYYUb/V6S0
4usNeFp8yHffSLBeiTcjejbTKwQXAfOXNNlcF7wI/UW+w7za6sTYijd/VvQKdpY5wZB+diJNoCiL
DG36HX9i1H7hSN37s01cF4UBYjRkwfbar+MMWfHpHpznB8APydfrff9h5cvZcuRdChvuScgw/Wca
VZGkfmB96EBYYcX1J/QcR8bB8o/vR4fK8MoPF3e2AdmMMXR2C52NFclfXRpPdctGHrkKCsYmBt2Y
6MnIZOG7EuqmQpo2PcHFB0bvy1zy5oiMQTJpwkO+uetX6Yzu1K+cwmbpCsvEk/5PYISyxOBY9JcK
injTgFc7BfIC/Y1RqPFzYN1QwZANGJTu5dm3HTKspAC46EI0L2KsyZp6snlC+iQH9jeSvZfObyzl
x2kQwjdpx3zsC+vonZkVAFv+WrgBOmPP9zcvDfGYbNrkeFOWRedULWMONX/Daz5ZpshZbGJD5P9n
FnRkW66F8jQW7dvtbbIlkleBsdhqrkcrci0aiTpi3MnhgUnipQMKu/dvpglgxamqkaU0lz08uNs3
Fk7mc0fAcBwmaK1HfHKjmitckNaRVjFmacLI6jEXX7yAOl6fy1UubNP20vWuOEPFbAj6YitMMKqB
SKTEwbdZdhQvgPz7W3BrXkx7/GDkZzOOTHnHaNQGhLRrKZeLTaYK74pVS8CYwSLa3XiS2tBP1Igj
e2fYzRLuuE2UakrzFQ3I+lZQNjNXkBZjx9tAwAIuQVZGc4lIQbmAV4AqHuaIWb0Bc5xEAQDoI4jT
EC5HTxnJ+1RWZAxIiWEWAVTHSLblFrf7Gvl7lauwvcggQIVI+HKdH3GGPSNeMB5Jk0jZlHLNhBUV
O4iybXlq5P+4eP5k9nZ2GOBzFtMoastI1cRmv3MFwL6l/FUfi3aMMzwzXCyKtji+gn2v3zpZ0qDz
9CBkLHzdkA8yr/sx+DwX9eukM/y1549N7eDSYpsWgcV/LiSmA19r95Pt9Y0EB3xxFjM3FThryOjB
/BCM6iITmYHgrDiHkozeBXB2bef/JwdCBUF6Ow7FLZSqNakmfQPLBKYb18d8tmPi3NirkYA6e6Hh
xi9M/ZjZ5s/04VKhWRqg5Ik0CUreSeQ1BPDyosDXq5BTW9z78rGjUyQREWPjM+Wuy1Fm8WKL0Qoa
cGFGzPUP56/xn8usABRIogtr+F66+ssRzhu6vwojThetmV2P10QecQ/F5uPRwCC5LZRlfRUs+SMl
9bhwxwUDlEzFwZVhGKip+U0kmFXlWc4uqf82W3K6GoChZ9tmW0/B04gez1K/pfowNeq/tJLEIXJ+
7Ct7XgrjgfJIiWSTCFRl4vbVuXBYVsH0UTNJ7+IAGCMx062bboB+ItfsgxDFCpesKf21op6HkJ+4
1/WxXjocIjLX4r9dr8a95+Kb52xlWhE0NfxdK9TcVQY3JOo5Cl60RLhFAiXAu3EVyRqArSvtl7A+
OzomGptHoAb1EMUYJjMGoXzxrF7cjGOuSg9zUTOgz8vGRBU4OU/FPzMqZoH3Z8jBelLBJnvg1UwU
BZNF3dqA17JURuPOqttqPc7gsZ6WoLPA1GhY34pdzmnYwpLnE9oJ+90/OPsplzYaEyL4jMNs1N96
5q0nnu4tNBIG2FinibZJRi+YT3e6GPnVtHHtlcc8benK/Lp0WJFwvN54TlnKxUwh2/vtmQ9w+6iE
qQ3WLq1rdLk+x4BJ9fo96mYHMIqHFVt17tn6vaTBmUCmaZ6o4xi3+lpfYrOI6Tsz9bo75A56TLhy
oUbKYCtlQcAwqvYaD4AeHVlLLGJotfC1bwvgwONEYRS0/yV3urzCECiU69KeXLZGgtiEyFdNwd4I
kysqTOSMQry71autvGcYQoUCBS2L4VAa6Eib7ugRUaLN+AuhTZUy5T4UvqW2l+Rd/z3wWMD0QHX3
6G9nGOPl1DhDFrAT2YRPoR4okKOWR1UcUaVi5vPDKgpacTSP5TILPdXjk9MR6/JywxnBw44XhFJ1
oZjThh1KeQ8YcrxcBGA15cFzJknKgJ8jUe3t4ztXc8E2Bc8JOsM99y2YKENXnKFIoJU25LyXrFiI
gl4ZCS7mmXO1tRUF+FQjfLCxX4KSLYt3Iq+5wkSM59V7pes+bPOojc+e+F08RPQlKVMZBWMV4Ch8
K1A1fZc0aHrCgwj39pk2RTJwFConxthd1LJrvDct77+nopGZ+GyJoCIhs3crJ6+4IwKYZU+GbJqV
2ADHmhHKrImPdTfZ7cHd5MZslVr/WNrI4STNNgFuZ33Z3UUwlhATxKvJkvex48y8M91VJsAY3u0V
GEHAofpzE70dklAPv0LIyRd+x/AFhfjN2gyxDw5vax4w5caSFTmsnPhzGMSyvxLLPp6JptuabsAF
uxbMpYmMvod1/cHmsjS+Pzh+F0YZvyc/BLXU2sDDPpW/Znggq1a2RA7BagJOjMyoCTJctSxUApZg
oD+qP7iXYrKkp3OCh8k4DM9fduy+POM8Lafx42/7t7hiOv4zQo92qKst/EmZrdYiaT1Mmy22ZVUt
YPJBHqt4iCRv1wnh+D+I6peHCJksnAM7YL6gf+4ZdA7kwhd+Ods+srscyv+LHcaTQllRrNMUjkWg
DqE1bEog0X2LVX2n4UQev6h46JPLjcAurF++ezq3ipuePmSLLEFS7g1bJc5Ow+oDeAEgqHU+LuW5
Dus9dGRY8qDogRZhKi/o+es6PsQ5m4Nymzxp3aYowaH6O4k5j4UJs+ohxo5A7pmp2Usk+2LqPKyV
ccOQpZWcNSA2+f9I2rdFCwfoTi2pjqF8yXVrjAuAcmGzc9XPNoLKI8iYnPvdeh5aq5zz+8dzyv0k
FRyi+mz67rm0/2cBM5NAspOh5DMM+1ZygT/EWGMoe2YffyxiC9m66iByTzI0Qx4uvFql8eMcFccz
FKmk84UbWN4jiphtx8JJWrVFqnfwcWFGHOtCUFEXJIuWIzq9H0DfWc4kOo9Ke0+QPKzhNGp4e9BW
xVBL9fYx0FYjkjwtO+Yiu2fRVpXrRhbnzlVIDRUcUTKTNue7wlGIXKhSEac2XVkCb01GsNuRMVAf
ikeeIOwCF7NEWegAoM7mGy24p1/9BKubCBgvwDkZTt/gvp43WJLtckyfEinxfpDdYEzITALrgk5D
iwnkiLM4HXe7gBCrizvNsYuU2YS+UDotu1unZfS41nz6g8RfouzYenwCdnDXoXEmThkFLf1Vku+o
mWtGjv4nn+qBlSg7y1eFn44NQHIhOCq4xFFvPLTc2YNOiAf1VVochr1g6BZqSYpxwnDOlfI8ce90
+V30FJKTW+LHLEalIs8wK4EX3ooymY8jmz7C6W3xnSCom1DUtRUv/8ugsMH3o6NGXdVFiwfguEaM
hJlbc1F1axnnJ8eIWP7S2R24HxVYM/LbE3nTznGCR03cGzvMug9uhzcfypsAYdY4wlqBiF1kAojj
bn0lCaSydPeBZSOaNkj7PFUiVepL+hvco7ItB0++Da0IMOg+P51ao+yu8sLXlx7503E039HdhC9K
sCWJpehXkoWZwW1DXxT/E/HmLdzs3BoLGKhZkaea+7EenVUcugSIpO0d6tZhrGHYYhIzjwYF6WM/
JcYzIItKEn+U0ViY2tXU1lpR29H/slbiJrt9HKfIYvREbXOPsFrV5TEpIvNs0n+NB9pCpGE3v/KO
PneImTosocPaH76G6KL0lNMkSUnra1FL4FVGDKGoWSVO2QLVqr+Ab6lQa/lxQQ3AZtHpk26FnvHB
5uGx5sWHJxqSLxBxpjkplGMpNOeRc2R7wWpRdr3dLdvt8IAP/hAwL5r17p0m0Xu3Y6f+If+n7WNo
Z1fTvzfmWCpb9bv59LvSms0NN1G7t0lUhvDrN/zYW8cbGprROcBCcvlOlBiHRTuFcu5UBB8MePUV
rjCQdFGqvJ2DhZ/8vN26BdNq/pk+8qQ6Lk8yBm/7pYW2qcepVAcqbNO9CrlOC43449Xe3EtU6KWv
yH9q4yQflmvEug3ymqqJiWQhDsQYkWx1kyJEcuyohozN7DUObYJqrhez691Yfm+DwcT/KywmNBfK
ZTWdFnuWXaYOjmFX8QoAMLBoSTTrHUkcP48/my7zi30nusmkvfa9lkvA+JPcXF3qJDJmH/FrtIj/
0ALftiUNNwtY4u5Xc5dySiz/DACGNOowpk46fcTas459tEhB4WuOb5RasJlWg6KVX74xMka8ay97
BEjftrlVht7EVUFnFcGC64c4WVo1xI33HbspQh6ToO0z1dYHJMmKpjCJULrGIQESBkrcTSmydWd0
AWeaN3dZtZemUiBwHijOneT6iDBeJLZoOaq5TFuWkMcMVp75RYLtnerBGWUa4HB0Zovm/Wd6AguX
8MOl2Cs0InqNA8hecW4hc5vsQvkm9/pray+EE4d/1ijZwL0uEcvSz1J0PNRMRLiv0MbgJpW5Yxyc
y4UwPOdlNweRvLNEh/ZEXVciGRLbzNyys0w7HKKmTeEP/m20ZRc2dIJbZ9aeXTK9nG/C+tLQtMNs
cyFBKosZdj4MIZGPSEpa4yNQRrd3oOFebMbbCgS5BLIp3VNEfY9H8CW1yIl/ebqwZMWKHfAk0VIM
/DE56B99Dnun1J1ngbdA/8SxIlPdFre8rnSgjWILURrpcHwJpYCOVBI9tiuaSNaAlK005cAWK2d9
RO/W8Gib+AOj11NrA0Sb9hGjznelRFZUfIxkZbTv6M7+cBkOAE5ohxctiTmjrteYySOm/Ia0WnzW
r7Jb03GzT2rhD7mzxSnQU8eJ6IegYsa6prb+3SHGgtbqjHS3UXuV7k+kaS+ItpakQSh30ZWDygEX
jPQs7K7DOPCSs9O/7pIz6c1Tbhr/hiHJwvZ6ekndIbJED14CgG0v7nx0+8RT/gU53X7JeqPiOokf
A/F8ENxfnkWhSQwlp24IvFdtnFUXpHr4ZTBnP5xZ/pZN5856yPyKdPOrSbg9XYqvCN61VJGkGWin
mWMiClzS2xlBotZWzLltZc7QoOCRpIFqRW0n9e48TOBBcXOpk7TR6y5d3tkpnVvytMF2R+eYFjo7
Z/XlwEt0AX5vgzVGhaXlu9P6szp7/slsteg1SBNHjeVsuRixJ8eJ4v5wtaj0Y+dnJw8bSnOqYJ6c
P6dpTKTSnw5LVWQ//HsR5BHSIEwz8pqct0Vp+g3bzsu17cR9GRIy7PfGOVPVN5GvHyUqBYb6Na4j
WgOrP7oL4MufziRVc8o0vbKNyKYg8TvJ57MpEk5jM+kYY61dK4QFqM7BOAAyqtm7Eyg4eAyHsO4Z
BaEyhHCUs1cEvqUL9z8as4yOv6jzeWgfbO/DcN8vJCtsvfOJXLJIgs2/fIcXsWssKmHzIVCJAe6R
wGCQ/RIdMTbDZytFP8Mcr3XcGTFG2+P+aZ50DI+u3og466jDqoIz0VI2b4Ns2yLaFXTcYTBPAUdP
Xdyb2s/5H066khKROnmZDtQaYEb6Oa/ItyHoOj/jn+cC4O445xrtxXDCJj0uy5FmUvrB/iUw2cV8
UjU9e4tamOS3RtpQuJJlDeyiwVm7drXoHscXMWF/ys8Saz7NimdmeR3MQ2PNkVbddnPHtYJRWPt6
9oaEMMM5cdGoyEohZOHTTAuInH3MCZTXBMGS10lpOEnNmnC13HzwFqY4/yvh5cibVEbZysIY/V48
C1l5SBlS9oJHNPAAvtAKVK8FWt6PtcaqDw1btii4XZznky3+api/nTXSSBaWsYLa/nq6SjW3+cxf
Po0kFcDcUrb5QDUHH3X50G7fuL1bPLGbnq6H4XTQ8p+9uyIRcQ2kZHHrnrnlQRqUNBh29mkqHKzj
wUxPgIebE9yzZ2E+VeXxedVwO1XKKZwmV5529lfl/4QoMyNVE4F1g7P5atpRRg2oLktvv6an/hrE
vlqzKthyXocvM76+mIXeiu58W1rDhj8R3hXRMR2WJchOREadvkLbdPXB0/E4q1B87oGQiuuksCxq
OA2bmPkh1jbdB6wlqoigVFjrtEv4hUGFdqeX6BDLgTzF5Dme96EN69ZBwNXyrecNk8YrvEX5T9Gl
3+T5bmH20mV06aC77rCLFScmABTQoT1EeylYr9hxG5drlsd8I0q1IX/dIVat44fHZz7jIZ7/GCy/
8yo1oMunrN58KX3KTLUr/iamZD26AUHG636MyvnuyPRD6u8j71mmPqszz/hhO5Q8sqVRarfiz1wy
fnERNxnU/AyCZw4kEgwk6hQbVrSzJIVb9bPvLtk6jDdrYJdiHBP2NwGxu72iMXDH+qwiwybk8N+B
6KrYCY2WZ+b4Cx1puP/soZ5tK7f5ySsd9/WvaFLiT/V7skRpgRgaUTxN8bosNPYz1WBpK0cu8e74
pS6vUDMO8LFxpJ1FJa9gA/avv5nYP2jLZ2wHn/0tbUKS/eSOcKOFXMSP6Dr5XbFT0U1Nvlbcnqk2
i0nk1jNJffnFCeU7nbpyzWOTMxWvsL46Rir8uhHjW28kJ5iZqj5l8MUqcHJ3B7SKajdtvApNPV30
Mkje5djJgZoezbcTyNsds4N2lTFaSyKv/i7/wbbCM6LSfdRNoM/kIvMLFB75N0SHhpqCRMFNHGUU
EHwpIlM4pb58HpOU0Doa4kJ2G389HRUHeG4UVUQIii4kz9zQx32oSnPmgoO0WyXqd1+lxc0+yVQ8
ftluLYGhcqTHHqaqFIOLJBcYg6RgiKs9bkUCwIY4CB6he8DHaUnKGLA5joa4oOhthJO2mSJGncLP
1WN3nasFILiMlP6kvS65T7qHwp/W2FqcSQY8qhUtGYdyyuamKY6m1VgbYL2O9VsNCa+rD/v1iwag
NbODGnJMZKhUK4mWL5Ip+Lk4Me4UT5950kwdd8TfVhGxlixtk2hwlwcFBJwx4GBTmNHDqRF4z/R+
jiPdnwOJSmIotrKofUdZc9ALKnpMoyq9uD/1rAJu6T9d+4yCsG3+PDlNi7LIe+OrmVHLnM9hvC7k
74PTQkVOA8UCz7UkD/FCZQDblx46zhQIinvwEl+cxhkPU9wvvNQ7mC7l1Msv1JEwqaS9oHgxZw3+
ETIHJthLupzdriRJqIrqNkJU2MW/rkCcoNmkiGsgw81fX6P8sKw7NPUB2m1YUAOJ+wbEzZmhL7bE
tAhB+Vxg/T5klFKqGYm1mMBK5bliang/kwjIFBNC23ZVMfruGtStg37+XIP6ScJF6/BYQdXLv9+U
5YJX7/KroSDPPdd75Lsqq8Clanqtz1LrcmpLO9EaKwic7KrEHDZuKWRKY4eWTG9ixOzCTVkyEC+I
CPPGavphs1lj47owaCOCPZMYmhUWxHFap7M0eFWweJ/SoORkzGN+FQKwOhgOQovMuAWoSwD/wxas
zRskVlLFi3SjSdXpB56uWAjFghNPE3WZKMacp5emstKvjhIcdS1yOMYTPNOXKpnaWqLDTebxilS2
v946agHgZqqIL+yoF3UJYPvZsZUwvfqcLnX9vZSWVlo5T0ffKGqBqu2ImG2DoqJ/LEUZ4eB/ekfh
s7wRWcTtFcJY2/LwWAQidX4udvFhIVsQivSA4WJeR4j/usNUS5FLOgxav65CxgKIUlglnfZeBCyf
6mJPGcG3KhW22qvN3e+bwcBF5TTDHxf9CSuDxidhtHvvUE1c0CUGCt65Fk0mN6huGJ6HIOQdSX0x
eYpOlmapsJYGa40Bxf+ACQ/nWZNH9mGC1xJb1z6kEDcipVRsvqbz1F19pMfLqvur7dIKyA4D0WU0
oVHvG9gm/2CHlnVlmMnrXwwYp87nzKHLz4lyXMXgqKie0HTipFX7xukQmNepbooZVC8BdHFGdVa+
eYPyOqDMai/kyqIS2qADbrnRWD/hHS+e75tYGgR1lKByNyjkIEd+VDG6DdgXGtLNC3W+/0R6TW/J
bBdqWONMgOXNopCSv6SeAy+KTbBCPAmo7c4PJ3UMtWBm/DVxNRSpiGDJqczuvnsfWi2V5jnpLYPZ
Hm/3BK9EBlkPM3G7u9SEuFJEP27FL76XdS5EobZkGRs7rB7MlBJln7NnbN+JVn8InYE3kCkH3Nco
qyyblyCncTkPm0aHvCw0DN8NxEVwicAhcn2Viuia75IHi1j83cKsM8OSpTEw8v4TYRXzqlYCStvD
qZFKcco8d7vmajVS1q3vHbaKy9N1f1VzdMXYLdWDn6ZoTuArI5jcfYpAobCT3YYQ1+KPuSzbRdyr
jfJldcI+Hc5QAxdSRUrqM828NwfsFeBLIeP/dWSBZBGlbroJ9pwyJF5xrmVKSy+c17cDLQ9FVLSM
+Tfw66yv+wVGgrVGj5OgXu5e8q2W/qt6MrZuBmN+AD4uI+QakWhAH0Ayg2ioi3AiJNFvtunRkC60
2c08uKgKp5IHFkktg9ZMT4yo4pBUdJSTG+KrrFN17Z19pXk2JxCyRITyEdNIyP/+7lrvgUUrXvvO
4gJQHZfpSVbFYH6xOzSwTZ4aSM8LODpiCfZGVCBcUDjt3JI3kEadbxryUQtLb8Hj8LnTxr3sRdrS
pGe3PRj3lmsV8n8LzToCEhZcWkXPgaajl++7LVAfgHAMGvVujIR4cDLxqQjLNSvp2yIl1URh1OjM
nbk1aqylDsfmkTKfea0bLrwDz4CCADpibvi2wAvlTVlKePeWO+ewUiYWjZvjDzcYqZGPBPfwaRBv
0np2Q2/xWdt5RCfIoy95Qqunox49ySKecFwYQaljL98EueLRzJ37tnWxMbszGfrfN0wSsfpRrPBj
Cx3pqmwiOD9TSGJhXQ0O4aMg8G4JVRbP5gosn4u+TUxtelhqn5z9/8OqKDBjKcser6k4Do7BdQ3t
Fb1qFWHF1KsqYFLB9fOjT12qTc80efaQM4rFWe/dFnwYARZlS6/CBTm4TVzHyla6PXJKmH2XvQlP
L/leWx4H48txJ69GdPYj8Qt5xK0g12tpjAwJJ5uvmn8NtUW6AN15UGCKlazf5AZzP04KeLeyPasJ
kgOoum8UjcyucWuF519ZSQ/c80jLs8DhlPmDEYDyRJ0TxgG14DzvveXLVO97mqByIm5M/R6mKgFM
5LzIQy2O4/wyBmVe7pjGqkyzUNzSuCf3sXhxKDTOJ5SstL1YZQ78aW4F3wkZj/9Uy/GA4jl/z3NG
VzGv3uEsrJBvSbRZGm/GFdmYvEzvlzMwx2Q//fqr+ZBFVRHWuz0V1Xfyamxby/1cLOXD52ERuGwN
YsEdjlFP6ANQAC4/H6IK8LwGzUymXV+2at8ApbraTcMhdJZTNuF0m3vFJA/K+xlEvz5u/yHAOhWf
lDkTnSDZ61obzBNlcFQgJdKrKwm0EZMO+6/dh3jAHsQwE6q/Pfrajh4ASgPaCgmuYWM5pF1r/vEQ
eyOym1l2LUZHDRwCPO7WwyQALrUgwXn6SAq6xc8/rsRUzBbvRDuBGglDcSn4n9xxE/NVit2pCufH
1kv3Z0i6RfJlYryAnr/Q5CBvJknIDHSMpyYHKj5Nu1cY1xmTQbv7pQvPENkUqBnIlBxK8ZJA31Wj
3KBIXGp8+ORiAHVfiaVtssly/XRULdWy0nkxd6sMWTJ+tldXevpgC4j3Z+zxjGh8TxafTao4Kjga
YkXegiGBiiu75gIKuX3R6tgQoLjDBcCE2f1os/n9luD267oHftuEAg5cAfx+7ksRqf7EUO40+/uP
OoOl29PgOCRsXAugMLJqJBOpXhxSd3N9S0sWunpsQLVnH99wKGLOT7mi7n9IdYXx7ZbFIiEkPl4O
DsN3pyUgExdvA/YE9Wrde4NH290fNAHAsSMWqG3lbpbU4PwHnjfL89w4tXcVi+vFZSvZKLtRN9Za
n4Ct4DarOwiotp2lHALzAFKVok5FxOiOz90uuYirz//vd5AEIUppmTr5fD33DVFAAKKu82koe3uU
Z2H6MnTCNLX7GwJ3mujkofoTKfgLTIV4ac+n+DwRBxsDoOF6boQzsr+B9rI6XDvZ/IULESImNZY1
1zDLyt1wudqSX8DEa6aQ7kdyPVmWJau0v/doeHRYmp7qQwWUAA8tulosDBk1mN7jzNNxT8WbRkEo
VrcmF6P3axuXvvelHrBkNL0AjYxl3SHqg1sRacekTBSJbOgVLpjerr4zLGPF8RSIHjTzirGtiepa
z/rMoKuqfxeNPRkwsAk60r+dPIh8gKQ6TSvoxiAfN8bqqe2MzYTCaRLf1Sr/ic5jTrKqNMXTwd9o
YcTQ7vFj0l9fzGWTvCB3hlB+3/ivxU03yXki2l69TMRsqULYVPNEI4oRAXVzxpK/KX7wdCfhqnjE
WJaZUVxeva9UYmkyfJChoppoxiFAQx+ihKDvnnyEJBJDQjRh+PPRGXwx02AaVWeT6F4ZLyDw0fOK
Rfid7TbTL7Dzbok+Zb3aLtXegTtTp6aJlMi5CBbMv1T8cSHneFyJePMCydc7+Q4CnSqA7lIbKGhP
KY7DAsdQ+yO39aIYyvg4pXyVPwDhtyU23iPfytTzZygFYZ/1FmO4oyEcTfhCrkGEfrVAlc5thNDd
490yNchGaLGZao/gGv9zoToKKpwokJ6IwmthosBV/Bv8BlgGkPv3I4UsxTRqnBpbZGm5ZNvxCAbw
cSNbaY/6eOjlrRyBsyIca1PyD0VLI7grSvlMjyyW88M3H3VWj28caHe5bx9J2Ssh/SGuf87nHqtm
nSj6RtKqol3KrpFFkUrpBFYMACUK02wx/esG8Vi2nzdxrEl8uV7hbyn1yL9DPPXMyaZ3OwHe5EB5
EXIXX/udN+uOjlKyUKJqFsI5O52qvbiI6xvhydzYVQnM2Q/jUcGzbgJgMkGXJKwzQnwHiE3Bz39r
dSrH7YJiDIDHO1/ZDUcHkoWA2J7p3E6Rz7ki4L/aM055QNCBvQLQV6qHld45iOpjsCZ6uN9Jv3er
BXD2pQZX9GE0/a74GU9xoxBVsHWRFCQlwiIlh4OdYFbiB8GpNtvcpJHRU3sQtcP7SqyPuCdynbcD
ap1zJTKwbf2c7tafiMKbA8ftU3VBoXWhtslzh3TaDYgVoo0XBuenN1BNaoPAYUBWVmo5yMi1/eLV
uYdmdufIrmUsplkmzyUKVd2SGrUMysPAThkQ91c/ZpzQ2jgAdLuMB7eZw3VOqv/5BTxvgxS9moYy
M/9tvNiZumzmNI6Qja1ubhlbd4QkgFGB8nsEmDHIqP0+fnw/pWGODvvVz/jGbflh8IF/DgGQ2s8S
6LpvCZtsQEtq1SL/OyJ6Dsl1uv8MidnIm0JW55BnW1zRxwUsHBeyno3UK3PIh9bd3y0YXgNDsBsc
SRuFtdLeZLazpAkmcYf7157+GKMlMzVYYUJwNeZb2n4HfPwZfd0Qay3RdorpQhN8w9rEl/UuT/Xo
qvA6rBh+uyTKs/8DHpbZ+E4JtCl1Qi77SsUFdzJPR+YeY8x0DiUq1QP9Ee318NhNxWexXqQn2Ch1
oe/lTc9+yXtJjoEQslNE/JEht9hud2ql7TuPmez6GpTYIgQE7u9cdIsE1+EMaF3f1ClS2sijuaFO
G/LZikNaHn3AlNBJec3AANzLbbTsV2i93KhQXM+4e/MUdzJ8mkGR9F+KBtrvPZjxTYDADS6pzndr
CqBwdlWgPTc/aUBZF9oM2uccF1/amuwNMo4WeVN88SsHRjU9ivKCXG25XP2li0flFVJ2Boz948wX
yNQkTLRMRTWh7EaTaCY+BHWhccW87J8fa5YKwkG1zE5qUOYvOm7gXkIj50PqeXKY/3MeHJgifKd1
CLVR1Pl+pW4zhf9eYN8MRr+iHor0ds3XIbFIHHOUgmh2G/2/dyxuKM4z3UUqA9efhwm9FdyXiRUj
RJItFdRd8EQq+6xKst2es/XAPlV+uZ8/UWQbiV2rDGvjAgcRGGCDoc7oqQDrV//pysBXszTm8wOF
nXtgFuVCr4oLB7IbtEHsZXeykDFid7KIVxgT1pyclSMat+dk13RATzpO3f78tC9aopA8Q30D5TQh
JZJi+EmreZXBSKESiTpyjgRMAVV0xpIvSQaDxodCnOJWDnQSqIUQPxreayhTuMiGZfpCtotP1KLN
GVFEElMCIsbWkhEkk3nAlLv3zGkXFNTnOBHFhk9/gETMGSJ3xjMb8W7zoz71LFMp61CYzFha/IuQ
VdRAhmPWSYMLdj2Yiae7ts05vOjlpjn6HkOVHmOGd/26QyQK7P0bdveBgwer6UcPW1qOodtcJBSY
8kPoJC/quYWLCpwJFU87KlKBefirEMtnld65qyw9YmOG20JBN2mDkfUoutRha/Z/z/KVFWN5lXG8
6IYKrSVNQ9jBAV5wz14PHDj/lAHF4SgM6YbwGvCuoA2+makukVEpd6wbuf2Ahkdnzmhqjd/d1u37
jrd3veoVJKf046ofad+CwLq08w1znH5FQG7hd/o+nppAf7ymQYCQJTQbLbzwZF9bV+YwlHlB81pI
u0pPOqx5EVGKJidKe2vLueU7CqMoWz9mCTyzH47WKYufwnhX6e+/9sB+0O4ETXAXZTwRMfHnLT/t
FulEBoXjb6lZNp7P5HM27Z7TkL3I24Ezh2IxrBCjz3cloFhlBnD2aKKvpXJts+ERdkTOAZijcX8C
JKZ5eKxCM93mcwdW620IaoGOIVsL3IZFLxX0V+CYU8qzTyqswPqhV6SU4NiSMdqAsvs7503Yj0MR
8dmTHN8SCLq/YVc1nL9YVRTc5fOQTgBVhgwPCdTmCmbndqJ4FVOrvLaHK+a3ThLywP4RjnnrIdaB
jghSpSOtA8KmNmLfkL6tRUrokJmeEFy7qTIaSMkQerHMa1r1VDUKBYOFG3P3CVAtdh43Bgoqfhpz
xEwz2TSsE06Vpa+f/1Vax6d2ux0b0GStEAPdJ6VnaTtx/IQIquW558DCV+7mFrA6v0oIuK0vyCtV
e2p29RwfgOKfLO1wx0+eBQpjChGDn4yxYsXzc3sGhObiqmPytUhbCjntQe76FWkc2hdMuC4kkQFi
SK7YjyGSZPi8Gnb0KHXlj+Bs7KP3dqGp+QcZaxSkgI7kNZsTNUqJw5ytWOzNcbpqOBbyIQ8P1sU1
fKXhjgeVGAvNpt0zX38/B+HWdPmcyaAsG1OxtgSwQUc6orrHUfQ+65+YLJJiP42cVP9sNpIDv/Ah
iI00e064iSvR2MNwmCOJjKq5bZmIA/3ORaCip4i/LSJjuPYuIY292d1jCVebt7TG3iexoeAJFeEf
Pht/Z3TYvxYiTtDVcaH9vlhnvBToYb5hoH9Wqj3t3+3lssBq2WHKc8Qs+R9CPzbHREGllAuol2sL
/BW/gtI4aR1Y5XdxnAKfa2K4eqKXTHjP2qWTiuxIf8PMW2nh0+NmdOd+6ekRLH7DE9eSb4wa3HTd
Bukvvgw1tLVHwW3wYssstdhGcPoxMjf+G2YIfoC0UECXz6qS2txPhtxOqWFCN8wkdhxDK5WPSkbb
bCrAxU/9Sjvx8lmrZ71XreG/GWecwPo9wGdThJeDfe1OasFsm5LkkjI5m6r+wOqn7ywyjC30AfDu
tORsrSpfxp5HLJ64eb5FY36dfTRnGjSujISTI2oWo9YSmqR3aF6UnLgFrbKM5WcujVhu8oJrrI4c
Ahm1w02PU3LfwlVtYc/OLSgn0pqaj9sRJ/IPdNECMwAC5Cz9Tw5WnM59PTNFiLXGJRxzDF6Jk8Bc
mbIqeQz2zIIbkXKJhpuEm1ajjFiiBwbVdjkR/7mKJzMgyLPBkGqL47wmMmv/y8GOrgxUKIbb5/fw
GMHFSk/lhipOnpwgusG4BvzDUWAgkE2+9axBXOp8LdtL/KSC0PtqWVkx+3f4Uk24tyfDvswfcVOW
qJov64TQIVtM7Pc3DKC/ccwAV8Z38zZeAAZpmfnDwuPmvyLD3Dc6OcBNBdQzUPf+gLqYgddLktHc
fExzLa/E09brMsUIYyXxNDpJoHIAs3joLEFj8tQy7upYb9bH3AfWZi2XRUq6zINYb4la2xwFbp2o
9pIHsBpWLBbpOhtl5Jk89ys7G8d+ht63BXGRe/q8/KEvwoNfAaIcGjg1ihPc/Xq3j3/Z4Nun2so4
NdpzD9vBgC7IlbMqAJWjk5RIpl2B7dJuWS+AeeikEPiUV2ROkdcZjDPN9IvgWCfqg/kLO8+UDa5L
c0XYNhm6K5h8AZ0CjgG30AO5jdHJXCbMdIM1/rEcePi9t04SVpnnR8wO3DaEs/nEFz7nxlT+KW8G
RmYBzfNGT8PospULU/Z++i3CxKeA7aFUqOgdprTl7mYFvIrN8VQq+xj2+us4jtIhczlFoZA7RPJd
uv+GygyQ3P9FVDnsacJ0J3IysKmCu/wtexAIQEHYSk6733NHaOdrMWNllFoNQYWiFrYtPEeQCi2s
5FDeEArhE+6hvXWsec6q7Ev0vPmIfUmWNHIEAmbN5kes66XLQwlDZbDLQw5Gvp8e1obGgMPVlstM
jD4LgwNn0QN1xzP0QH6w84Mdld58ovVNhElybbpN0DMcy2nGiPXIx0zl4zi/QizPraux4Ta7SgBU
hgx6auEKgquH/oZxI5qr1xk43BAyfIuS3XZ1zjz6rr4+AeiiBJujLRBbJv6TwS2uvmn9WYlrSisV
R/TU7MzsS7ahtLnaJbMlTmA976QNntqZUi/yqWlrSRLaKANXt3QpmjjSvG/5oIxTF2ZtQUooZbWG
HkHihxZTtnDBDax2demurtoOp+JiN2U6NmM/wYzZvOlRDODuqhU3Omhpmt04F/TZ4tzrewge6zb4
jMqlqeE/xEpIMzqUQtkxCyrQycCFNmXR3EajRG7yORrKDJr5NnZI2MsHLdziCdcIWbeVYySFrx2i
pnUJdeG930IjI70I75aO1oipb+Nu1oYd7vYqajuKwAs0Ib6yZFWN1N6TiZoPhJcAIkU5N0VDM9QT
1gr12Uq5J1h34mztZ+j2cYBN6OlKsD9rQLJLTlpyGuR1JML4YMhDU6qulp4o65/afaBHCJr4JCiJ
/qp10PToA6n3hA81g/ZR+WKkzOPBRV8d7JnS9mxBY1Zag9e31iKfGIFscQw+cHzQpE/XSK/WBB8s
FAdJWZ4WKQUApJVmNDdC8DRFZFKC2Wy7LfYZpEun8ZZ+gk8zkcuacWHgzlhhY1F1BMEFhWtNnQ5a
SHekwRyAYjLM8g2TNuoqAFGL7Ba1MKfJvcDtQ2y0lbKZyxT8mwrdyFcnJPRDNXdah8PMAjtYnu1/
b1AEu1vjBd46RKNIi1kZq71aUeiiWg+2F6KBQURxf/zmzMT8/aGm7rU8ORRBYyrY1+Xyk1LU1Qq4
PDew+s0V7J3Aj+/q4XR6wOKoYbFNw52n9PpIDvppSp3h+ejiF/9NI1dnZ85W6Y6fz55yT0KuRg+b
s5OpwLzYUtOJhuLV2OO95XpV9dvsqLYccNh1DdGGgRAixHx0P11gN07hW9DueHqWwTlMUoUD742b
oedOAjsJ+16uNgo6+MX7t+M09HZizCAnXGbHmwWTXJKbyDA4RPKm4zDEmJdAGciOLtnTRvvMNV2i
6fc9B1fDNvkW/RpfJHW3HGUsnaCNkMh5GMJyFMVQ8RVBg518/kF13mF0WTFwp3JGQ16D3flXblr6
Mo/npSIaggzHvtruIMDLr+vV5r/zwnk4h7zswU4V7jgONQFTJ4tLdy3Q6N9zDx1idLFpD2GmEFgG
dZx3OD/XZqVr/I2KknUcqBCajqANThBKgTPq5KrqhKATkGeoV3hB6IKZABDSKZnRt/Pjl0fpMG24
xgFPI61dO7uSphoMN1OkcZGLucxrEyoyBMcDKVMpVE+OjIaMO+UTFQCi4JwsrEY2hZFNokQDNsw5
uN9PImFwyJWeZ18Xu3iZzYKbTNmfQ3acT/MeQwcW2tBjKZwVkt85nyx0XTfhmCOKh5pdEN2ict4O
6fX4XmHPIf61qHTDnCV1GrTIt1J4VgA9nuZugmkBI2/a/070Ci7OvRvF1HPLwYI0ZGdG8z5nU7fL
FV+MFTVFIl77s3v7guUQ2Z/edgKujUUn8z8wFOIj9AHAaCpcvPZq6rfEqd5KOlVvkSuDXiclvkFJ
X6BSb2NRDccFcJ4q1+R1NXLxJBVxu2sZaEiH3V7ZBPscPeWBOX+DmR8tmhVEvEU7s2049BaCElSA
+eeVsFjLsqvcoIElkN+0b4t2iEuR1sLXZsveacXqTpzQ90mEab9Ki1OtjbfFfPr93QU2Xbdb+0Ga
L18SRcfsBF+fg45zeZdCrCdAlMPZ0taP5sVKXNjmJ6vrMGxdm8pR6KpRoUzdV1/1Hvfg2mqwVwv1
oA6R5JuJiAqUE19QfYBmqeYv79GFHqqvtruoYCt97BzJ3nLyLdUFNnuRjKyjRVlhbDmA0/aP9U3N
VHo+ygf7y/uKhQlbc7D8QkXukHd/R21pGbUurhN7BXvosnK+KH5sMW71gBBDb0jBFbd7aOFe2tNd
70gq5zr7sYgAwyl7oREASLrXcoSHxXqmoc3jMx6rj4T3MP20lDqkfJ9k/Dqvi1KzY49iZY2X/SfA
pNJ3nLYi2+zk+nslgefMUsVSEuDK7Kylod1CM7pQD1JWup0Er2mDctW1HuxsT3i8rmXgknIdcXdw
wioi1nII2Y2WzNJVFLMY6kbfccAJ92KYIiGJm/4PQzAFKbZHJ/l+NpE5H+ZUzNMpmSgeEd0IxGb/
0mfjl7gs7AkgXKLQpgFUol2v1tQoZQoczQi3WCicbVZx+ZfjShr+s7ekdVWe7gmcnDc75DGmjGiV
xjZ/n6/RsHedrqnrnP+nSBI1DkR/qCqZVopdLih5vxVL67w+YD7N7YNXb98X+ZUu/GY2Z2RLeBbR
Voba6QvC61TaCR7MnYAVND0kTxMNlqHRLb4O7iUrw9aPNGCK0wZlD8ZHqR7srYJo4Zr+IqfmQwxb
qpikNtmpQdUhgejrTBLTzz4rRwyv5P25txZUgXTDr3X0iZpnJ16kDcaKrIVTuGxO/qiUt8Aek2IB
6q2/CgSofbWsUXY4OLrW0+NUEYfRRrDxnWEmX5v51P5DquufEaBnAeLUvAmlyZ+bQGxX7Jr1vl3m
hOQuTlyJk+3W3tI2uHCwc/n+yf+0y6S6xAfwYm9L0RVzhgOTmXK8rou6y/ttoZ9UFTHWFL2fLLhV
bXpvClwj7hDGmRrSz/NBu2e3Oz7H8pAG3KeCLLvu63rRcJhlMZQpTs5Df8WyTQ2ZRfYcIrGUUQUD
ZC6ttclPUECeLc0wZqarmlFmUCGZuJJNR+qQcC0WckbHP9MWwtOv3DnBP5iFU/aB6IG5IO4SAl8n
oPlsYAFmbLB7rmT8poeRKNpz5hFHyOYONCZV0gZzvUO5CXaupbnchBN8b0drfwiPFxDUcBqk1MpF
x2SsjYj8HkoygP1zcI1ysQtR0PdSLxSHWZuJrMR0VIDG421qLOp+X0LHLVqyFnjoREA9L+1L1gBs
2mfhb2OJOaZ69LdrV8gR7P5qKwrr4TYHix3N5tN9vKaWz2AiqZxmBPCswMOlD1Z3dNydrNLN5lwd
2aMco/J8Cbuz4PkZjA5DCIiNW96NTZKQGs0JSc/7s7XVR0t3vNbgB3ODBT6MYXn1bUxCKrwfraFe
UA/7TD3cajn3xVtEdDYoDpwxixAVnkL8VaLR/1V7h6Cqp0hoMLshxS5Vop5WR+MJKUKVG+je9CFn
J4db4gz4lBJNgQ8vh5Icj3AfKBRaFccqjViq5mNZhFgpM8te0QlfHkkVEytsVo2uuwATu5GOWa/l
0f17DgGcWoyiHoMT0lJPadqbp1tdxmX3Il7lVP0mrALL0QF6OSGcc7dbTruA4iwlGnIsr1NV+/ZD
91NjVUzuFkcgFwWvbgIzM6BA/8ZIu3/lWVpgEvHO1cn9Ajx/CUPIsIizT/FsPCRHzL0+RbIJFMgo
cM5u6qVAXof/f8mQKFwsdBiGSk80gY1XkFYcFpkaQLRxbvb6DTHYQaIMoR4mESXUwt3T6kcIzTXA
oAfVVB1UckprfcDQiKSfhCz9A6G14SIV9rkcsEfckbwVhbarF5vZEV4CfX/GfiDxxYaA5CMYPU0S
mY9rr/MTqzMwPAKMKNJDdEK5/EiZMkdnmIb+qct12JvhrcOSjcoSbmuZrRjfJBZOS1hMAe6cgvDz
T8QxzP2I4m7dB1rGjn8q4CGHkwNaU7LxR3YyooTc3Dlrz45RAtIOoXRDd2OhTuMDb9zVJAG3RJsU
zeBUtzvC9vyr6jF3Cg5M+xT5VY84VjZVbFTt6D4KTerKPP4vJaULGRinUDuByDuS6CmIwSGHe3k9
tY+CPfDISteNKktKrtKGBVymOLSfXxqfEO3Kjs2pIBzYFmf8M+jXXdeu3n9h3OjS78vNwxSx/CZ/
dF8vfZrLN6JHStoQGetIm84FjsPW5hAUlr/IX8YFyj8yahMcLnBh5PM/Xsj/S2soWj3JDxz3HJ5z
9WzQ+mJGFmlfXBMM1oh3xcVPzgPQVi+CgKa5F0qcTVHJ0+68UYb8jmjT6fbsDYV6705cDWWYgFgf
Pj8HwhWC54C13X16CpkO5Z2SPzalVPwoYkz92TV8Dx+YI5ZzlGEL03/rjJ6b/9km514c17x3wzTB
5yQf37ep85rS+vFtjv8Varm4Bp+ijoelip/ZWALKkm1CxMX3UnTBXtcAW4ti+NJXrrs6atzlUvkJ
qlVn6MqeVIvckjtYHF8sCW2/qtxEVMN1QHmikXFuBo8OJvYMGnqe4XCuUf+Ws8VTNj9nRpl4F2Rn
tUY38rF0ijiZjBMQUjcmWYOFok7F5ND5mQIcfqw/1YNBakOWIUh/nsrnXuyAkPNutgC92DqFhAY2
41mtuWLpMjT5j8n+jB9Hc+kVoBPZGadNWbKODSq3zk0F97uC9QTSXlh3soXpQjulb2TpC/L+n75S
WxZKPr8kYqdK5CogdNKuA+N75Ywwez9uGVlBdbnGVV0Z8JnEOAVBQWcu+UyqK0k5DVjhNoYW9YCl
DrWgccC378xc94N4yId6eGweDIF64zpZpfLdpeEbcOZW/7ssyaI8ABT3yjdJw3GKQFvCzm/PtGMm
Pl8p8L2xELShzL8GFZQdJ+uiQyAU+uucfoVNRpoOiAuHF0synm/0YcaaUMeAi5fSe/3qESG9Ptl+
liv7HwWgCeheX2Ci1qt+L9DHtCxFgsCSwRA7u7HUWoEJsN2ixuX87IadfF5jlnp19QSYrXkNhlw7
MBWQi8/LKo6IjnuzLukPkvifKPYs4dGahVimJy+7AAJ2O6R3L4dPEJVO1xzG4csA1EH0c3vTB+Sz
hE1LHIpnevPbNv0m1sQ8sfG7Rx89GPRI9v7qij5OB7iK1XS/fcab81snnZhY7l0SwFpTk3R8eCGC
Maz2HbPgN/2VA5uAuVeKW6A99/MgFKXc2DRyHC967PuJWr0kO9AJHL/yLUox/svzT+RBBp6rgeEr
7DgHlHCM7SeIr7EAjWaicvtaFpnZluW9bNHeEzlhM1lQXc03rnNMuf+wmZerxd/5UbD4TG5YGWdh
hGgS0r40Mm2nwSUzTommN/1dCbZ+6Xmdq3M+jEkn/nZ+Oyy86N93EXXT6q6UVTLN73E1/O21I6j1
YheDASKz+oZA9wUiDQlXT5E3eThevBMG31NS8cun/HfRbG50VNycFAcKvndhb7fPHn+jqBloHBcm
L8s2Lo4JlJ9dYiA/0TdRK3pYJGZ18VNw32i5VZdo0gm5eBfhLrszPUbhw5TXid+X/7WhVqGfRbBw
nUsLk8zy+uQjPdS5vNelZJAgXGX7UwMYKYeJPQlEl0c2iUjxzUh7Xhlcjl/oeAuWat20UsQJ68mC
TezRtgP8ZBL3RyEG4p9KqZWd0s4/+0Mkx5Ox1Jljn2QW6bHX3wjRodBZGuwpsxNftjihjwbo3zJG
6RVBpBgtwD58qfshO1jyasj/AjnmmCuksphG5AzkYsrLZhBz4vSxObVtS4JHlMrxWeKKL1lCB7LT
gnNfql9n155wWnbCVqBjfkTpv4JB7k3miGKBUsra72tNQZEstK6U4ND6GVINFzDjvv/o6UxHX8eJ
W2k/Upbxz1gufYNBVfl8nLXoFFMEUo1/PFB7Av2u0G7c6XNDZjiBU+AjVSK1COHRD2cgh3xqfmvG
VhBh+AWrzYL/lE3xxIMSpgOMnuoVeK10myttBk/I+2pCqb/7AqH/vLZLkkyZjZQ9MTgVcAVmO9kx
NKb1iu/PxF/OgihNVgLONNHFTgCJx0Yuln2UDQo2INdY6kKOHdwtdIYNiU9y6IQBjj3O7tFPxO5c
sxUv6OOv6xtyYFEGVq++BZ3cyTEqUL06jylMkzBQpqTET+vOEgMHbhyfUyDfk2BBuqtN7ipmY0zz
4B+o6jux+oQtYoOM1duAOAXVgSqJqDysNa9iGwZ1cIa9YMorx7/GkSIZhR/q2zO6wF7JpjHmY4NW
NOKfRdWqUInJk9xgRxf39dkZACtRelAuA1i42XPj1oCnAVkEIJUFQY1z+jrGaOtWm0w8IygbJjo+
2KURidW+1Xo2NBuARtJ2Qkm2GlMOnMq1Q72Amkp9fyYHYn1N1zb7MUfd2+l67tCz8hzVUJW+mtqM
s1ojsL4hvWo7al1so7JlYLFflzKIZPrC3d4gzpR1zecg+1yL7QTVC6cPJ1KIgyELgdMi+Rl9l+2D
5hahOg+YfS4j5BBIgncnIUwvMUEuWHH3mqV9jfRPx8VoL0Y3y2UkkMGsQnwbklA8P5d19M1cG8QF
Vcf7vHASoNmgmbfxO2YJdt+e26s8cIk+yJxcVvUMDd14W0XTFGyy9k0JP9/BaIOdBme283NaoZ11
JmGJN57wKf1NW92xssJqSXN1JfQ1DcTRRIyFiXEXzDA6lFYM6m4t05xi3QUkp+RiY09EQ5joxqhR
TeIL6IpK7AY3gpR51PYEUc8OEw75ZfR/zKz4TB9zvDQF7OHRv0IhvH7hk5fnLKRQCruC2kto1IEc
rTSs724AXw/5jx6O2TGFvtrAGu/kVFB2WyQQl8PKBlmSPG5dswFBaBKrrJ0D7T6FlKkIdxQGl1yU
IPbygvaesRS3dEfcablaZiL3y55nnEnglP+rJGOrjfvbgPqtoZoDvflY4Lt7c1WsI3qmPS0MUnoQ
8y79xVUeWY9bfL1gwYslzcvi5X9G871xUPIC2upQkM+gMi0m8PjWIFNMUaH8mPDXTRYed9FjDAbH
jJNjKsIs+LZw0dqJNFY25cG6goVoZJU/GQfPmyvshAFdJy7peygVVjomjCLJ8WJikqb8vd2/t5oH
mijxnj+nL0e/T19+mfKeqfuIDF0e0i5t4jb7nfw9Zg7j960iF+M0M3343G/VQKt12FqA7/u+O3eh
pQVrXVDhFU+uNCEZ7grU60bHJo6/XHBAS//I3NW4EmXf6uuqDKIl4sGKU24V0GylB+c2A6Icc+vR
wxwvkVXvNFs25N2NJrP0jXy3UyZqDuVAfg/j2DXteiSI+VmPJM/VTMcHHpZy6jkvo6xo8TXJ4IHi
nTYOWuU64h4Fw7J15gG97Ai33/yuszJwEWTWYd2cYTsSbsDITs0Eh0h65sCjxzVkbr3tvNQ1RB33
Wf5vETMY0b2p9yHkeCbDYV3Kv/9Hm6GyeZb/BAx74PayeOg4F7z1TbK8LUGZTchX1RIFpgsLoekN
9O6ioyy4zGYIcS363CbjidTPjTxpbKejuk1ZQhvSFLh/JZS3W5NTk3he5o0/PZjl+YjsVP0N2Vtw
nPVAFb3zFJnlB0haRWT7uOfQY3yYVhjxh+ofdTSKDZJNpQ6GS5St0mEn1kmvQwiRQBy2Yn0ugeKN
kKzgmtsDKa+wroaawXJEJHFQ6EHeMF+leW/kHVZjJ00GGz/yDSsvbJ4Uk+uArn/x42HgJmS/d5UC
4jmnDqf7Sr/B9ZH4Xy8B5LDznJWD4Fs2q8dTlsTgV2UtMC5RwmE830BEIlqmKid1Nlxp+9R9yi9x
cu1SBbM0pxvErk2Jw8sLN/Uf5P7OsvlxG3iTXNLHon89x2lJClhbphAi95jzovbXZ7tfPfW/lEzZ
wfcD2iAY7Q4NMvnHaIZP49ukyC86KPqhbIfa90+jop9JUDiSIsF/Por00eBNkeHy1ES4CJKGOzvS
+k7RQKa73AHSWNdtZliCAh4/tjctSLQEZKTCeCxsegSCDL9QGrULLH5QSv1lQElO1s5etq2nkGm2
5DcCMHIbRd9RPdYlDxQx0J38AsxWDhLli7PXVfkJ/YrW6PpIjSE4IaPUGqqsb9e2vwXTFUtcUkl5
mVtc3WiMNy7cBLoZfE6ArkkeAahCf9uI/oBbb3If/wfLncioD+dUvZVWtZUlwbnYMH7nCJsnIxmu
egNc6xr/OE0sbWHwkY7HQneOlQPjEm3Ukte41Qh0Uka//JYqK69FTbKLYISCM4NoEz4ThwEiYBt3
W03qWbMNJzib5CYJTrWjDBN18MrPN8DqmreGA5GbmfnS7XPo9tWU1J57pUoFEJE0pgzbF1Z47AgT
lu4HhO/0DDkuObZ+NGr9w6HapWCma8KWvRO9findKY8XRzCICMEBp9o2qXMYjXQH3E9FznVU3/8/
kgI+13a+KL12KtMY8HRw8W18vesusDdFMUjK5kNi/QxszHgz6qKznONszdQ0gO0Mm4FoMfV5wdWX
k88ZKFb+yYE/xC3jwFp6gdfzskqrUb10eCWvIYiC6nhYjirtTU5IyiEdmaE/+mnufbpFiAemnZ0C
s2kpXIDUMCL+TZyQk6dgU2ezzlohvDmIjBJzokFjD9eO+egMr7z0TxPC5g1bm9Ar26yUkmqQOhXx
ntyPfhNjs1Ejfnh+yVG5pT3EjPgjl2w+QYHBGQli+FcODCIgI/yRgYwY4cBhbZgmhdiyGLWf9cLx
/bHOHoPUiaece1eUu2X6dLs5aUV9lIK6MiL1JZ1i5agp8RyhmeqHGtvM16b/zLRsl6FUwhbTvj3/
U8lTY8sbIgTMkUGy6etPgndQw4rSgfSrYNX1+Zj8ItvWRU+Ko3lrEy0IixLHhoEHY2aV/d9lGUpg
totYLYjiC6vaoKzlcL1Ek7/4/u4dMFxE5sRhCmmFNanyCdVC/Qt6yqcB5eTSGtlKaPWGIJ207tCJ
uAbnMRnFCrf3C5PUkyxMHgdr6ljomNNpiyF6w+JIcuDZZE2Bcg8dkW2YYrSF3zT+YoXjRn0S7uqY
WYef5pTNGOy77EFWu1QA9HrTxfOSd/veICDx7t1a4Ui9vPwhGYRwytu0GAlBtnyhfGYMQqfyoT4r
puXOJz/cDwvXJGXe/5N2sxC4rVHCyj8UJnqzwWs5jsDGp0QhyCNaEQHIxLDGNGPazMqpV94+O+mP
s+4+OUFScmo+SJb0VLHDEixwO7AX3SDUIlNAGJj7ec34dIVzB/vYXscMAvVuwNyjYnDv3Zm8Zftq
kvuknCKSqKVVv5ByeAUsTXerkeIWyPBR+HybhhMUW9CTa976hNJe8QBrZYI1/2Relpvz2CfS/O2a
z7i07QhoIsE7jLBmyOQuzCK9jk3KkfPdrBnXGYY3ko9WC+WuixDePhQ4vBVmHq/JcfcN5lvQezdn
Y8g2YwdiKcj4Z0M1S+zz5mJjKUmqBjM9rHghMnY2NkRSjctRLZ9qBZ13g7HlD4gRB5NUqGRN7dyl
O1m3Mm4d/As1f4i2Q1lTSOBVV55E8LR7OG2bQ4R3ZPGJPbIqSEmt6Bl19ombxEMvMxZ94rzjSHlx
Bbi28DvyUTaI60CVAHAhW8v6BuE6VPXWF7dtg1HDwkB3InNagau7npAQQb866eGoyrI6nlIGEp2x
2IpfUPUwIwvGEigh95rgMoo48he1alcwzWkmLHLA0Gjp1P9Q3tWWTIUiLvwI5+yEVE1YRjU4VEgX
CjsXeY3DC83hC1cU0bSbseCb2XUR1e66kzx2VHrx5Snw/suHQeV96+mkiuLfSeiFh5eEAgvPvRPJ
2vFa1Vk0AEbhncOZAqgW7I/TXrfD5qkqEmxUobstG+Nr8Kmf5MM/aSNCBIEkqQDlXqZUcHcvxsyB
NmCmdWtHSy4K5w4Xle5d/nr/kNizhY7ChWxc0GXs3kTiBwkEF+zjj+cwQOsHxgIAjFi4Rhb53c53
M2i+1QgYnTmdDlC0jGtHaaNXt5wrmw/H/F9GescQhInz5C+TkVJ+aKqR/wVx6UHi7hXzVSMj8ivV
wBSOAp8jP/ahPkUFCMKGgDUDirXV9dqH8acnhPAKckCyKZjdh2676B77TiyridEVuWXqltQrXcpp
Q9iaYMRtNQU1RpSiCvG3f34mjWkr8InCj878lw9to1VT2dRq2IkxLKabrF9Fhrey3J3Ku2dTABeu
eYuIAzwS7XeeKEUCyOEHO0UpCwlIAKoIxvt8kYuZupxeyFqR9U7hdEB/ZDGB2ji38iekRmXWGoBt
wque21LpNBLTNeWblsqNZkzGMw+StPhrYKznJIZEMWDE5/EW8Zei6kgTfkeAVCHZAKau2axAW9ET
H+AdeMxps0EsuXpxSih6fPM9b0IjL8QRdX6pFRPA86tHaScVuNnS429JZ5V2DIwP4D+35hOVTbdT
qzzpVoPAA7plL3GCreYTPon3MQbYn/in4XjmmwEo0850WgvGimtqsB2uPbW75WsTTVZ8PSakKUlg
uorgTIbZOkthsdVpAxF5LrvEdJBvkesHHSeTN6OWZsBnvdyJYoW+6h0Efsmq6sXTKp2KNG5McUCj
zjf6QWK2ia5lBq2f+Poht2MWBwAgsQIT50rrYXT6t9YWWf7BePtW2kwbf6apfkrv1iNLh7PLgiHu
2fkD6rb8f+G3A/cArqZv9Dsa/xqZAIAFQQlOJBDgllxjezJcsI5qgo8ssN4y4KS65DgbrRlyOJpJ
J3QtvW3XgOPpyEnwmSABfiM20fG9EyCRa3Lsk0VaKnGuy+mAB1l2+jnI9TI599t+nD5aZ7FhaAEX
YtyM45HWAP1WM+FO9au7hSxmNqSssGRn5uGc4w9cATGylfNVsmVdXPk+l0X3KNfyxB67e8Ljbfec
WhsfYJcHGHHSwvcjbGlLee2WD6bvspcJi9HvebCFoiF+rgGQskCNFMg1n9aT8HV1wMJebTdrsuaR
2x/MNJkg/QvyZuQhUFZ40DFgTW650yr5IBqUbio4Einy6c+VFd4sdFEA87EZInm0pHqDDKwQ8p+4
4y7Rft6ocjbFAT+g18tK0PeC7QnWCz9UUTyynGHeMr9MNNwqCI04YEmeqm+JrCxx4p88Y49qe//v
/AmrKP9OlnhmI36e8AvBIh6fV/Rg/m2PCL7T7EXPtDFuDLquY5nKWYpzpubtg+auzhBm9O3JAPH3
yQ8pAd5q4kDTgh8euH01QN7ZiLhLFJPX9LgAgxBfYopSRmueb4g7JP0xfPn+7R5rhHANhcuMH+CP
e+Vh2MNFkyBgVHyl551Mp4KrEnZsKvYe2Ns4XKxmrFtXxxRwh7bhBhTq0dCEQ/RPmxRq/bhWCHLa
7oOoTy0Etcg7wpZoOhBQqD1j0xfA7mhGOH+T/y9zMPxuB0KZ1a5UBCKYu4S/IGVxDGJTAPx7C3sB
ZGabgTMTB8R1vKrMCqGRL8IoFZ+N9bNrVGRGrjmDx0nbyUo8plsvKatn1akRg5EA48grQ4PO+gIH
A9pXlzXPDVe6kWCAcs8vajkPpo7tWUrEFiC2WMtaTMLWdoJvEW3S+tiThAzQ/F6iWiVMmnOcTim8
ZkJ9y/297MQ62QnT3y4ncZN34u5UrsRw+Ud4mgK2PHF1KIDyoMgR/rmLbHFMir7B18FMmpNTYPi8
sNNIYOt5toxXEpDK4cbaWLCcLcQMhmrgiRoTcqzZOQKnTieblTpAXSP/Y7EBv9uGQVeUh8SWV2fx
2OewtoaTMkl8E18A5YRHBxKUy/uqkGCNsK5YaGyMjBKrYEr9dIVdgX7jvLrsmt7Emd0TjGVw8mGe
BA7HybhFkEHOBCGoxP3BGBlwB/j/qa4WO7eJv731/4IPM656E2Uvu0wHOJ5SSKmFUTH9r3XAM7eZ
N40mcl4sGBmU2A2dYJu3t8es6BxCZa6IgQvSRBKVjS5I9HNfFZbBMzO+dUJCipGacI3Lp9QuD659
eQI6Ujd8ZHrFAGjIYra469nmNg9uL9EmkO/KIZPATjSTebQ0YM2mYexrCmx48Ql9mP4q5z84WEtT
avsTlm6EmPBmUxn2cAJmN3KPsav/PZCYU02tzOFyT6pDQAXSyPiuH6qA/sWgx/zgY6ej7HSONJ7f
6SkYaDO4GlYhEXoUnUDtcGy0ImjXbDECbMTy83n8v0b2hGDCSXcnALJiibcTtCfKR1yIsmI1CAeu
MGMZxvPqvi6UsEsxs2kLLLP9eQO+3TiYMhk0yeCfRWd3tyQaTlP1lainxoTvIe8G+grLd+VUWveG
8ZHyFCWvEoBnOpXn1GikodufA85VI3EwwTYM+sb7KydyiUDazvCmhjtjuDSgbgUcC9/A1KDmlA2d
lFxzYtKH0KK9ty41fWzKdtD8eULnME6wShY/uqw06fd6mfgVQ04nkNsYLGpgJu4AiNshnBrfkhdf
dw9WNRvIuRNW1e6ym/JZ1FX3/44Vb63/GE9AsjqAPDu9arWjspUIlaqqLZfX5vBSqkhXdw1QT6/B
HdCRA5HPvElaom7Ck7n8uzFbF3l6leC0/w7I06xvndMDHcrP0lAqjHleNUtIf+ZRxJqrqIgTr/ia
2r0to4zdOUf6GkYL2+aRNTGdz7eze34PvyLKIvRh+QWha03QDxNhWcLqlfU9SuXVA1jpijeC4MdK
W6VpZmJ0Hpp41+T3/iG6o1pKn3d8gqEEf4NM7NuMYgGpKn/6e1vCFpVnnH/P7qZh4Y26WBmQiNFE
I8AIWLxNynWhWVL3zfIGaz+0Iw148BI5YfyfJL5xmYvhUIV5KPRxpxvkwhc2/l3/PlE/PfDmP2Lm
3cgiihdtz+RuMgFaRRhTEtRyV1VzfP/vsRUEJAC4RF+1tBhp/HRn68aU14v3IjjWZHxbuCk7ybgV
GAm7GCCGCSVehjBHvyRcIWZQjzYIcu6POHdJuSt9+GwPQK1K/lqz7epiWUWzul6xwz8NMCgUY7av
5cwnWphGVvRPvsFEAY9D1RIk2OICkqJnKrJFzmvz5py1ubNAjXVqS/jl3X8nx+ynaSvIRbGNGoIT
wZ25JshKdEcB/wQw8HNNTsv06sH2uf/t7GTDIOB6I1jgTQNUNGV6imqMiRZXdUujpkOvjVNmRsvn
xY0hMtMldX3cpZlJYveUTJ1n5hm0HSWSBxF9ShJa3mqOkSzfs3XoxnpRHPjAQb7Zhd3+MxetPqZL
/MWzwh3Lj/tUXFgHUpekgCpXaqkrG6C2x8tFkygHmqYiUTyhrVT/tCoA5193pAU2M0X2VabgbseW
Mg0uhCwOhZExXip9fA6E+4g1XbUR+93UtUKOTAIecPRESrBWue0XgGsXHIDloIB0CC6Ob2f0BiV4
vJBssPN/Plrb4WP8HTGYEAwDVffPxVK/RdbTaYzMEusP1MOBvISo6sMFW2KW304HDpWfXnIzf2GK
fojTOXG54VDpC7M1rSD4Cq6m+ERzzBx5HsUe07SYJrppWsqzHnT+auzM+fN6cqk4tANKhHun4EWC
6j8dkdViiz/vYZd9MywYA3c1vfKs7eufAmbL71Ul8+t3n/B8iNQmKyyn3y12KgxEfIIpGCMs/Z8L
QK6eYJbcXZKydKpYHD82/do1lXdL8Uwb2DWgAQrp7wIZBM3lRdZMLDMJMaIeFQj6wJXm9VMTUi4Y
Qo8+ISKaz9w+6p1F7U9nrGkl22nt8NXmlH0lfO2G5WmkSPOyLSs3LQQbzQDEOem8NYckupXnhVvp
Rz73vncqZazWJjYSnkoqYTT3/+5jeQU3v/AsydYpZ7y3X5g7R9finZ+esY1Q16fEUOmL9kWVPfJN
fJLcJXa9qo4BQ206ySZI6tOdG5NufBnFM1gQHOhnvFfbOwRg39Iw/8x6QaEOLp8Gnti+xaMdyFwP
II5zJXVMnwDfQajRiVpySTkFEZ25zIm5/frg/2S/XzXyJttR8y6bN3ExcBbQfHabrS62i00XRXQu
e6qv4170I2j64h4mb5AuNk9MPQenroRSvCid3KbLCMLM9OhXCaN+moBSM5kRxXdfKfO+FJOXybnS
97eLshDAnWf7Q6ZJx4DC8lbrD1uPYfBbwpw9axKKx0s//ItbOZNSvYUvzfhNuwI9SxKKz9SDn5i/
/FYv1BFWUYLLJPBx3N7UudGoOgyb7Gb/PDqm9H/iZgMGmHpj2SDqjOMXgsvhHg6h2f6MEcrcAir/
nXauuW+yJgVHPx7ZrRHbsgwsvI5API7cbCv5Z0ToWD2CtTlLCbVU9HMpS0cVRxp31okoRXPmm96B
X92YI9CnvykdphUtD5kPfN9iCqmHg1+pE0NZvOFIzy7PBndr9FeAvfyXLXPRFDUgpjfg13Ey5UHY
ZeLXBOlgwtlwb5lQsEDX1Yag5JY8wHzOVsnwX228mDiMUASvrhp6EWFws1aNh4K/enk4C168J4mS
1iomnuDMgeLHeza4Fyh4MZ75Txjx0R7AnqPHRII4AGkmQRbtuKqWCVdruSQFZiOj3QSBEtQdlbOk
3e5mCThhlyxdVN2gRJSCRAC3H+fWunoHJEEBbG/KgeOrsQtdSZidXT+/CcV97nN7wWMbg5eZ4L+o
Fq9HoKpIcrVX7D7oTCDLqeaSi+4EtcYjxoRpecTb+udWmsv80PPS5x94jx83jeTN4zP9398A9eR4
uPpc1Kdrvec8ND6u97duIjo7g49oBpsBvee1qCxz3BNMFIUUpPWBAeOrcxZyIliAdbp6OFM8W7/9
NfgWIqchJ4szAWdOFNN2E74OToSxOo8uMOTm4/bG1ekPNlNwGdVVah7tdozMfH3MWIG2OM7Qq7PY
o/FLp+zAGtjSui2aKjNEYg57hqlc9uNUX5IUlJI/8XcV1M5l+AJylQt36tDXeDFzxsHMMVDO8+S8
fzSVRWgiMcQt6DZV9gJcdLZWh8pZih0USls4YtOI5nX8S0WX33S0NAvgw0J6B5TGDdcbIipVHIvp
2PLnqfvE1ruwcFa1dt2YiWl5uzIqSK+xnIMdsQrEVKu/uFBuGdryef/48qUvDVCjHb0w2AhGyHKt
mXSp1CBRUb87/waQhcA/GFYELDWCdsUnyBkVLcVi1/V+XYCAOmU5bXEG7lkePYsoZRf299RKrJ12
wlTf51jbJF7dNhpprL+BsfDfom8Q20iZZ9QCiAwPyRXtipJlWLuli4FVCTpLdwx/9kcjATXEZSO2
UeB5OJaGgjFKDKS/0OXqJ6WNdR8TC6VzFm8baCfmk9QiNmlDZW7KxPFxIPHF8JrNHYQS8yN00r3W
BHXpfAWqw00fCHvFIiJRb6vMvINv83TrA3KnTIe3PGGPmtvvP1SQeRUqbeVBf2/Tog60g2/MVJBU
JXLGGUeBeKA8CYhutmygFLW3V+FwYO4jb7I60ZykcY15X4rjoLZTrzKPIKBW8/V56AFsObZk6RqX
3m1iYVkS7yJT0UHt6o1oya97q+G5DzL3w79W9MG+3BIDOsnJhIP9y5X2BQc38RBIJvA5dEXq+fWW
xI0JSrNLtykKx5SewLoCjWLYeDVl0JK6MXUc0b1p1BwoNmEOnqra+HltOw2t3uGAuAqQ8XhY/ASh
fdA7riuq82a/pr6sdfRfS8y7psMFjmD3eg3zpt095GKSvUkAhIz1YcXg/ycJmiV+7rPJqVp7l00Z
UF8ARDBStHX1lxGfCeoGaYoedaZgRvyb6dwiTJt5bI+p85WrlNJvLGFGyUz2G1H4Qpuuc8mWBs2s
016ekwFEviFx/eYCjDnx21qHDyjRWqjICMCpz8CQ2K3iZjpRn611D1hFzqNe0h1S0Sct/XIwgqM6
kUlAxQXXAUNRz7ZOPmWJbZDxVx5AZ+Z6CEiuD8Y1iRp5lbPUmIq5O4JC1jTizaGqk6wVOGGl8xo3
KMzJ75PDqGbD/GlY/emX0+ra2gT2t+2On3Ec+ZQr6DjLDnsaIH8ZkCpvYKZP7MGJn9sgq338Jths
MuZdm7XOCdZEYzGRTK5tA2+/aF6g73Hm/5jA/uxfWapar8v1DyyiI4UBtNIDKyLn3DFqy2Gfk0UV
w362sZk0snQPI8fxb9Qxj3SZriH0rFvgq+H3DNZSthsk5FYH2C6QVYldiUqZ2qo8fuS3XgJOcZQC
OQ9SsNAkmt3lQAbwY0nyi2R3r/ys3xd4DJJH8Wp5BUditDTfZ40bTh6GipM/S31xT7kZ9YGrTB4c
nfaMCu4ykLeS55ZmWDW9sz3AjFDSJelVl979StUb5+3WK9zEGmoy7xnfH9oQOHhgIsDdN/jmbYSW
Q9d+ahYg1ZGZBi87c3RAjo6k6MayxjelZW+zOuVG0q9f+PYlr0RygiV+rnywOURojZPfKRS0Kkk9
dTdzk7/WcpxLOGew8F1pr5FPEVIrl3wJvtgM36xQafqjZCs5LWgSc8bOIMlpxmeyvzwc4RQzU80f
oz+ukitfjIKXYpxTr7IRKlLiC1nf3iGgUXQ+MduZEeu27pIPniWVKYXfQtSY90TgrzkdCVSfkMv7
AVCcBwdGMa1KQzzjhP+kmk4/qCb33a8/qMS/yoK7Ku/34oIXy91m9bx8JnyQw/MfIEj8Vta/Qflt
d6bN1aW5qEg8H7tvi4bUj8IxUAYUqHJ6nL/4bm6k/jpOtltONhU4Ny4xg/KA2G275NJz5lx33tfL
m93lzFqbwGhBDXPHLLp6+941lmfn2UyNT0yMgkaA0DlbksNPM+ga/b5k1pJWDUnq8BhQu6A26W68
gvrMWmt/o2/HD8Gls1C9nab3+vdSFn5sYx6dQu0zEaGFAUaqJEumdBEqSY9J3mt3JFVUvNJ9Lm4J
xeIiSbRZzxxcmFN8jgogJzkMgZLKHhbIYmExGVsH2KnQf/uYr3WFhvn+ATB+ApujjMShJysaVkRl
h++RQ5gPI/NWVIyoMu2v+taJUjmuR8xFL5fKG1P93/HwW+L9tJcHpegF9zbRij42wKh1HXiyMVRY
6mH33J/mABuXuL090jv3Su5IU6X3kpJigO776fU2QSIcgy7+n9qRY4K7okvmjFl1KoiWjBQKkr3v
VhqXXxJxkH5INj0ZjlLG9u4piCtGZAeRftYbxVm3LRrv/Ayll2MzpCqilt84DuRguOk1AGJBz5Ql
Dca61wEs3FOEyiayRkIdhCkk8afJQP30iZ+xPJGpdfC5AyL+baoTM19WM0bqEdqNzFNdezk1pNsu
5P2QTdoUQ0qenXpsDs/+EcOWS2bnICyyxIW6dzC0dW3j7obX76Sr9QMptHu8L0NIBRZ1OJNlBlPj
uttT09krYuE1ETyASvjR112GML08shIWw1xKfoT2waIjcWupiOnefiDxZCnmuYIEMq/zi7nB2PLZ
s/fTPReklcyGH+2mHCiHVU14ZRL+JNy/M4siMA+QW1F3D8iB0B2Kd/EbQBqYJTforCR6aVGcunRZ
890/tT8713BGC1tbBscgYtC3w7+VzzcYaaPt9VKF4XZ4QfWgvsXnrKGQ6rwpuXl3w4EX6SIRLH9w
4CC9VmlwaD0BvS3tZ71eDnntU+IZbc/WebPOobIEWf/2t8XnNn9jWixzrNZPpvKhhinl9tth0s4f
YRUsld20iNtYQ+fSnElXeZOsJeyyUvVoHhMKJ4EqbmZLbPsKJ02B5vZLjtQO8eK0nWx0Lc2aGz3p
PzFC8wFJav48iZSLh7tvfcJV+gFOk0E8xcNiVTUfDqdGoVCK8YqgU99Ry68+IXauAGy0QyEj33RL
Z5k6vpRwN9oZ4eUHCAJfKLdn262e1vwniR5Ulw3TkpGLv5jAzFaec6xUHZ5vMbkTvdnyzRDgljeG
bBB8luWZ83nLKaCo6R3fMrMv4LGTGlqpyQnEYKGq1lQtJAPltOBA0l2OeDXNpORTMYjN8ZrNtVDc
CdYP3bC2g1PiMUHcRS2rhPiIyHoHdjZAS7fAxL/4sjhqsFe+pjlXhHkK3G0ZgnJbrWgeYJOcwE4X
80I6GY/Qrg2IkxRBFurxgInFksxc2zLenNPoOzgNNWCkfsfA7Au2ApmkkbVyqhaX1SunMpkL0iqS
STC+AiaB5m3qjPlTAzZpnz66sTjGjO1h4e9valxNFl/oLxmwVEZMO/Ycy5a96DevaAnuYyUmCxMC
5CN8EXDR350CVa4RB2Z2TWbgbq0w2xaEhNp461oYzpLQUy0ttKodfd8T3IVzOjWxoKhB43iMY+PJ
lV1rkjFIifaMdXURyJTRpk/Nk+0Vl2fCjvH6EEpxuTFjEKOq+YQ/LJ1QEveMQQeMyDULB6qx76En
+PTgUESBt+9qyiJ90U38SwAmW/S3oXvAzRxn89EATjQp18RF0xGFhL949Khz6I/sKOYsQUdxAFpD
6k9NH0wVET3zDyjUkRnOaSYmvrvuAlY7OYj4H0SPZnLi6Aped4rg1B+wbhyBDSNoOpcQEZ53jP0H
MgRDsAJZ27LoPTnvz06wSG+vtuEnLJWJVu7bN95xmg2Xrui31ifFTpoFOqYWoqUVJTxRwxhO1hoG
lBCKDtFLvoECKBy93CnsyXa90PVEy99o8dvB57WINlA36nToMuN9gnlwguyyEvK5HasNWIuIC1HF
QWDSHGEBRkkX51K7E3XAeMPoRiYJuzhrqwUBMdam/z4mU0F2eiwW0dYsuLbpVLMUKeYJZMNra6oA
yAxYvoUFF/0AHvSR3a/mGIODWinUJZRgCStA9pyP+3JxG1X9Fj42DQG1iAaLMII4usK0z42gjBdo
9FD08fIwHrDD1vGRNIYmiZaclqSPHAeHJ52qWk2atAHSBlYbU6Edau1pVdHihFwmjbXtqPk7sjvq
Dhcp9b4Kirrezwh4+M2CYTj3StC5c3y3ylOe0mvicWLBEZDcVqfMfxhpfV8bOxP6606zDxAMsvEG
khAnLwe+NnLiYnb9g43K5lE+pImzRvXeotATr2O5Y4k77zL5+O0xU/Dx7INpfuzZfnZP0qvkyg3H
TgQFut2Kg2H8cl0kjy4TtFam3zYgeQFOHQMJiVq3eQ/iWYJJPmjCMjtde4G+WRfA2tdNoaBO0VKi
I8CrtwD7pyMu64aVwKg8uJiSmKeP0PrQIMsnzDYmOSFJQs1CdHGThn1P/6zFhTgOgpMLl7F4YPZH
na8WRyWe/h/ZNzJufIc+KXr51Oz43QBYRvb6gD5oHf7AlEOJ+2xmIpAyEELfl2J2dwLUgKNEGW+4
N5S16tdhFqLfdU9oYBq5DyL1vIkg00lpBCNs2rjKRKEpJT0RKiGdi28/fP9QHt2mCdX60ZZrEtaN
dMOoJstxZkaUqZ/1iUVZQuXtJibPrvVEIxs+kWZTK6cFGNZ2r/idf2hkfBLgLGGwYwGslX1Gt/EZ
DZiNICIqGiWXXOKVrxyFh/icxeFPgb3pjoEyboK7DgykyTnWM1b+a8Wfuh0IpKlnzbiI9D0JhYPU
R0Kaksys8S0z3NBf8zQ/FsBOfpsGXApAXDSKR3siszbniAJuWGWYGyl5A4bjXKWLFaVkX9PiaFUc
vT7PnQaAjcisAei4NaJuTeXyNvHe3k2b7dO13fS+B0eqdouI3mdhBhr5UZdgj4oucnKSK5yDvrh+
Vy3b22SuYbH1TQOtTcjtrpDiQsZSoHqmwBH10QIRfIEKBd9ErivAJRRdE1vj8AUlsLJXdL/XZ+NB
1c9cZQ3TOlY+ChvbKTXaIQN6ZsWmYYGjbCwsAzu5fA4Z3JNr+1M04dWHPcfbCGcW0Onxu86UsJoO
J4d/LJqJ2TXJWUp1KvEY8JPK5juaxEfgAekSyPHqvBsvn0+eQ7z6sP6FVZe2rzJIflItCQNEfJvr
1lRgVL7jOE96HuL5wq9zJgteEICNVwQEoNOQzdZljcWVlnPPpWMgBqSlXBZKfnHatUSKB1Gn476s
kdnDRJajENIRz3gnfNwHQUZQxA4k0I4TaSGTHYstU3ZdK3n+bJWlWwwUFwb1zhJnM3YvKJfp/+1b
rf2M/ZR6pLVmZhGzBdbFKpPV/1WFcML+Xk3l5nnwAJiSdaZtfmfPvnEpoMOTv5X8szHJJSEoVx05
6wZHjTKF2mebGazdj7/qvoeW7H3OxSQBDQqWixdLzf9wpEwRroxY0N1zXIrSrWQQWdEBgHsxgcsY
4h7VITiBQRQORhhYTdOkLy4xLnaDu/26HPv9OTlWIt86Zz5I2O3SDheNLcvYuvpg+E/brNspXBwo
r3jH2Q7yEk6jefxu1Muu/vl5cWEXv/XZ+Wc2l8t15IisqhzWCIYi8ILnGksxxormxLqGnB1JEzsq
eCP5/A7fIfmm+jxBGM2MC3Zjlbi0xcXKktLABYQbv+WBXRg+WBDM3Fb9uODHl6ILc09o38uM/hVH
fHPwhdjukISHkxcHNO4erdVrZS6jfod8ANvamDbStJfuZEc/atSJvzaSDpLaJUH3NtNl7ramy5h1
7h58wclYTe11VGTUtjedSykZgKnTfa4hqKfcig455SSXyYrgnDZzCNPzsnJeNJH6S6GqCXdMxjz3
+Jr7i48cds9srth9k1PpP8tAu6Zm/3tUrJcCz0a62/9z2kEwLdWQr+A79p7OZfUVT9JMW7TA4Tge
UTWxPnuMP+uu3ozQ0GYWhL3kxVZYhQbX7YVLAedgigmx5+tBfJkjPs2evI3cFx4mizHHrQvAO0y6
YmGCt84rNgHpnBOnfcdCSfP3a800ABn49ixHx+YrgOrAKcOVhL4TCU6AHJg0gpKjUP7b2xR33ivN
WmBfG4zcOkpTU/sda8IqMBc5d/+4T91q7P/1f94DqHVT94SAt45wEGa4ySRF+8BMvAj2V51nf1oK
nmBeu0VLNZQp1g4sHqd/bagqz6Q7NQB0jb9JcXFn9R7AAf0OZ/EUCwZL5YAIMHLr7RkwNxlVtt8k
9c31wVAHLlvste/WneKKrhaW5bs4toDLulZsQPOKeM4wbwxyIFTucbOaoNPHcx0rg4a4NqmVeHRJ
FX0RCwrcKuD7xPhpH61hhFhgBDqPUWU6hVauSUS/HazCOJZcH4IBIFNDlA911Dcer4rTx7Af9Pjh
+HQ1owZOW2KMwIELgwJNZOGfxrXhqFO2kVc81QmaDAcwrqQhDuiQ+/bqlzWSY2RGVenb4xqOTi1+
aFzuIexQvJi6cKPa6o70D0tEQCSN3MOOR/CYaRSK0JA09KKR+6CtJcQGbelo6FBo797uhQElhN4Z
ycpKmWPUkdNpF8xnG7ux/INHe79k5QRF+8TDlAedo00DavdzyDwYxLqIRVTcMPYirH8eu6cmV4HX
R4C6XPsyBNU81XseggPesu5wEIKXMib2lGpBnMD4oktqIyOctAzARfslp0lRI3qobA8fP+BdNGbS
gx/UGO06NwLXco65gU94Mo4oE/OJ7qggh7oR+ee7AeBryEl6MzKWXi2bfG0i3RdQuXLTYs5Fd6YN
imJ6wfeo0nn8D/LuAbURl+XDc+AkxabGr6bQCnMhjIl50qK5Zix+0mpB9/OjZUU8hUcde6dd88Zd
hHulVD0ZHX9KGgRuFl6IRo0zrxnyzzds0i8KN7aa4q4Vs3tKyw+0bh/csYz161y2WPip7yfEyykA
1hS4y+BYFb6rjRyeen4NutX8xqHVF+0QO0gDq43zRniBynscb2Nwb5cuG+tT3bvbFMh8VBLoJ5pJ
zfLytxLXWluNp2XeVSxtkIUgCBPwHWZrOmMRuAvNH6+LIbdcrN10EWc2xUXs1FKyqW3Cm6yPfHUW
jxMzA2cSfJdEXEoW160zJWKulnH1SCa82a9A2EMiVSkJruep/VkWytAcai8FBvhgLPIFhrSaWtTm
3KrkWMbjdUyTI4Hvcms2Hr4NYHGPXGEFZGULsVmavjpjFBLKoOKg1nvlmH709fvjkfh0GBpYDBiw
5ZaiVBUrD2+okFSiZ06F8QlkQZWGeuAZgD5qvuGtvoSToH4Coz1sIBgGDQeENI4njnwnh7K2cgaN
OikOh3eyuR6ZdtBTnJISuGT6B1a3onD8Ahs9KUMYW1oLr4gL4trUeJ0NXzZTrjz/d/OWwjJ2p6bJ
r6mb8/6OSKcVp4yVWCJKmaZWlmaceP7YtJJ01SgJFvoLog/TuaWlvCFpiEmutn7VlvhWlII6IEkK
K2tOkUDEIdr0yHN6wbQvhU00G+Edba5eUnHh3GtLAbZfXgk9LqWwxWpvscQRyR+gReTvNsmmDngO
CB9z0EnVEdrwL2R4bqRrF5UdqusHfvcMH+KwT4NrJt55InfGARJErxLselFCe8zfqBxzAdXmdSj/
+wamTKMX1oVJ1o6aROr+lJWLogu9wX1CDJXrSsV0CTHIK55iLs3JtgPfEkIR9yAUkrhHt5u5h6Pm
1igOQmOXH61lMbM6fPQjGz8GjSdsHEF/oFCRRSUM1Dy+yucFfWhwZe+u1a6p7q1ZaqKY9O8dVu7p
zdkuB0prwArMVQlK5wuKX7Y8hopNZUr9s11FdHqhTdirqgQyAoSyNPamDl+26OOMSU+IHeMq5NNl
t2qrFDy28C4Fn4e3pVJCHfTc9kYdM0DZ3a5Fw0BTtFNmwkCsrw3T7pWtZKqprbAPNqIhP7mkdcrV
H+k0ggm5YYwNWcIhWPdDoGAP5oKMNwNjAMZ/MhAHHfZvA3j3gLrIKMN6gv+x9j1vjdnma7AByRpd
CMZe+ncK+V6Rn76RLjPPo57TuXocV8t7NeCDkeLHla/16iAVTKM8S5+DVVXMJfqKjkiGByil80/r
906fJqu7CCgh6Sq/0RQjFCT4SYAejtRcUMtbyVEnAPR6Cfa/VVNdUncq/YlbEtPCbLbOVEBL9GkV
wUQweQfqGLrm4fXRZxV1V2Bap9mkVlIo0fxYK6iqT+zO460CT0yQYf9QaPGk4vMe3MuLJfehARhP
RZOicDSjxXAT7Fnc8AqZ8UU0PeOx6xT6v0+00330tPVgv/0MTZunJKVpd5A15bjyCFKN2pOGCFr5
L6LtFFSd9vKkOZhE2JrUPDzpBsRfi29lHtrbjMvonGDpDhtdEVdsJo/fK1pzMuavwCTriLiTr8J0
aa9EaFTmHqrWIXhX4FdIlEoUv1MCgfCzLpLsI1aVU4F4yh5dsE6Kuf9SEFS81/SsyW1tEbihVPdi
KI81l/GO5A4q6PSW5djmSUhbn3HlNFuyi+6F/xsGetLv9hz+4oqo2idnNG0FdGlPlx4wwlLpvzKP
OB6Nu7RNPlHJ61E7+wzLTA1QFfEawVVBMJL8U+hci7Fzszr/Ky/BWUIHUOLJHAfx+zVPvHwH0r/3
k4JrO3XxFsuf9ypanJWtrD/9G2RjgZKFIrIYjE4AwN0/GkprKe9ffg6ojypdIyCaoWPFpEeq4WBl
6XLkBMmr1FoVfZM8SOdGcUaTs9vWQ5PI12H+h24rbV/o+QQ4u8rQi9yrWOCFIjaxGf108aQcSY8Y
zOdHcGNA70UrhkQmWl9bRyOBTF/2cy70DeuygbLxabHEaJcBtBbYkNGtAYqp/SlzjIq32GEDt1i2
GK5UB2X7MhZK0JijuNfK9ZHXyIGOCUJxTdX5+S5ve5GQXveCv85VSp8OcOLOn0a4kulcCxMuvJOA
oJnFB2XhfECr8cBsQeDxi8XPPNKVsG1ROsMYW1NipEqv+VsoNDLlQRkpzcsIyPsil8zDOvOHQpeb
MO3bwtY5KaAsgTd/j+wKp/MmplLl4rPLzHdeF1PAyfR+RbonWTwbUlrRGmZKKpoPkmupuuvMpR9z
aQeV2kYkWaMeMVgz8RW17+3stArDKFa65iZKFWNgXClCGi0/YuBlnD5l1qqp8kDk2SqVjgC3WYG3
0iKNxwc+m/w8BfiInc8u9vN2r7pNPIftwep/OdtgdFEqxXXXjS31mNl8pG5IQvdFFPDmf2gy9+1r
CvRrUC579Kh7713YI+5CRfjx7FI7eqQi06av7reYg0MkMZ/WJwMhFWWHa2ZjAVg27c8fj51P8hhn
mfBlxfY5J2gZNpex1+TbNk7fS/G5LIHj2NxfV2sGQrT1+lgm7CEaBNyrB9vI8ZVNz0p8Eck7y/7Y
HBMi1rRN+lsbECTktjLswl81LJIRLfD7ozelPTELzt+FxbqoOZ5+MKU3o35byH4T1GQxmQCCgpwo
i/eRKxKNVcLp6UH0LenKREeE7AtlOoFfERGAI529pRvbEEZJzJIJ5JTK2T8VLFq6l+Eycz9QW4Ox
k9wW/r++JMchIdykhjk/x0YSxQvWwXBvA8DEU94kgl1WbdPq1AT/bBAKeufPW39tGrSc93nCUDhD
U6Nmw7vFAJJzoD7wZmLUAO4mnLckviRa0recYAsZ1DKTbmvbQon/dKclN4ZT4nldM0uUNXZ7xIm8
8Tm9bopux7lkdDabu2dkP6LZhE4D5TIKz/go+MKtcAuZrS3B8ACP88FBBcRLlm0rK+fFT+w6VRph
InrXz0X6LouIGOm/R7cAmudcGeYjyW8e7h3kwPwEAITwrWUvdHfS/Ui/Gv2gYL95xwBY2aojNcMZ
pTnJVqXWJyZvlzOt4cIFKr/lRQvBL7CRiJkqHA7qymobph0UcR0rfz0VLJhtYFR/X+E8UHN8nT9v
jkPY6r9L1fHkhnqHQ2WPuPqNDytm/2/MRlpzpiTHb0u18aHfNUDik3r9riu/pbUVwLeUd4sQTNNC
xfOL7q2ptvpgLcqrH3ER/TZa58GgtO/zQlysOojKhaEOrNjSfGkl0b7FhsuWIuhWBWJToLADjSb7
YPfaD7o4Uy6cUVtHYCcGwuSgPRMUPiIbE+UXvOZ77uxFcZq/tHfgTu98WVBNGesLk3WNBtMDepww
RcGxx1Z7yntcjpw201BYIucaD807GtoF3GUMKPIc1koa/UAxQj/6r25hFJ6s8q+sDSqAwtrhNKro
ZMSkvaQIxfkrwNGGb3l1qaLWVP50ReYP74JmYNU70U7dDqS32ow9dF7qx23GDs6QFXQBVzE8Dl84
HE7URHPey/ogrQDB1Z8tc7UxVC2C0DOrhyJFrspHLvFoCh5p2/6FSMozsVBT22e0C3GoNybD1q1M
MumtAZFlMY5Zy2y8J1UzuVjnOSR7fVN9qhX/1rML4AwpT2bAnNLT4TMPZrZllh5OV51vBAb0SAjd
szYODiJOIQjEmVI766+iAV7uKF5CWrftKo3gOFunlQxtEq1anVYmjrK6lGQYqjkPIlrC6o6bZBVP
sB6tyLAsjf8uySY4BqvKKVI4Z4P4bnS+utmtibVAmrdjZMmK0qWNUAJl/Wuql8ZhX2zqyMfF2sEY
/qtzQYsizaZKjRAcUEjJA9GHFCh+TdUidzSicgB5XV7mzLSvI7IH3Pe38cxH7Io1gFZyjYKJVoVX
TwLHh/KLiqUli6ALsiM9w3Dge+T397leYXTf2Dlcm04+Y16XGgDsOPnQ37lVIxbaGeKL4XZ23Bp8
Uzpmt6WAQ6LIl/14pHImZB8wSWqKeRUkzNkMXgwrhYLWGxagDS4nPxBW3e2Q/xTlkweBPI57vtEA
cCx4bLmyKZuhjNgAWE2pIoVtNDAcIrnA1hRajGxi2btHFTp3flD7GaMaHqjlmSNR9B7btDTW/U6z
Lr0SWIKNRpub5+M6aeEMJ8LkMDWH5wHlq3sdqvcHC0euLxYVCo3h/PkoQY5lh6TEO7bBN89fbFK6
+2NRjbC27lKgyqVvl8FW9cL7mn6WsH1X03COYWWasFMcDks1q3Y2CDdEWOZm0ADI0tJf6M8yjNqV
HqM4xZRJTTIrUk+Tjyd4FCz+lo2JggmlFf9vbGe/cVSJexfq4sV1w8rfMD+X80dqKb7jjjNrgSb6
0R0pouAYsAi74ZUtYMMaf24uUZLeoaj1fQY8VkmXmsqU4xWZ0QUF8ytFfhXFfTg3ExcOKlCSD5ov
FjozmXBPi2cAZJIS1KnvQ0MS/sN2jXE0eSTj/emCJk1X/eJ9KHBDlz1eqPXFsuBSZcMr3R0tiHl3
qncqSbo9GDb6U3E2qmr7SlruP4cGcGRgNd6GrTYphaaEtUBR247WZDB63eA77M4ysodcZQvRt+mO
NFwsCszlGD1T2Fgy6KBEjk1BPhf0rh6XGI+YCEgQi67oz97V4tRDTC0gztWfLcr4T3PBN4Me20mF
gkS/ojyGz5cEfm5sDDWniyPRjSr7xvMJuutRXRBqSpjUqscmtkXMeYUFVAaVwu7Ae6+y1qs2uLkn
bimVbJq2dyUIQfylf6wfTYs0zgXow+ClbhuDYCwG+fhnJIGS0BHJ5Q5bZ+JTiJIRH0kI5CvQoIlq
rkz7KaJcDz4PYAEs2YKXYbvEh6BYKEFFaZwMxPSL+t5oyNjk4ulQ2h18tCyw5N5WSlhOVv2hzGJv
rtxp6DzhSwEFhov83W4SOk4aLqeuvnayTal/4B6FjtY3jg8tPphXZR5GtflOFpdvgdpv0wwGHGrM
N+c0yCqipTb5awbCGoZGVetv0ZWVYAx42YutJVBVpJieHo7R9ErLq89F/lPvCW/YvyFtL5JsqdST
Bl67+UKZK/liTa10xGJDhYhiv8K1DQ23JLvfCnxNx60fYrvuDuybMeDcjFDPu7uoUlc9qdiwIY2j
xWOYxGubCayaplXkdpGaMWRXQpi2TNXn+Vj6plu7mqv+7Uf8zvlIoDAuBijgZ2T/X6DlxRozar8X
lmVn6KGeNH0HtxB5nQl6m5xbruryrcxjkFfetzTNyROMQNbHIp9eCwqCNoN6SB5O39uH/a7m2WjA
NLkNiP2YcZjhDEi2T11mToS+FeFSO3gyv/xBIGUzXUlq+95/ZloT9RPyrXxz0MigTjhljxKCTmaD
KIb8LpRmCgvQ8BdI1yV/IItpSN7d5R40li7Oox9PBm1WFgOvYVGWQlMDPRP6XkoW4ocDZgTxppfV
DCD4ajAL43OCEkAQ+qialvhRqJpYzHo6kpJOTTzuN4a7mSzO6dErfzK2Br1+604YC3b/BcQ0BZkD
EyDaKp+wTXU44YjwWIv9ULCDXgvc5fySxmzHvwaCFgbuQ7seJfV+a0SkdHHJIvs2WhINZem1bwIZ
lMocXdC/oxaaUDTpzfevVRRNuTrSNzb8fSTfywEWAOED9OoQSN63/m45rdoeTELYJtTxCyIIPRMB
lpWsOkX5M8JO0qXjYk2frbTAgLYDO+lb5vArZ1lIFo13hsSwvXs2dZLZ8vNd2u6YpYWz6qIYBYf8
H9aSFe3FaOkVGxeNQDDWpL5X73h4Fq/CA0Zny5bm0upJYAO9HkclfcBglxTXKbh5TP6Ng9KhWi6p
kk+WLLbErPGd0RLAKep2V+ecDWEdg+uVvjpWCVO6hAznZuJnZIVLiUA0TacsL/wkJgbrs8heheIm
0YkNdFvbCTCAu8RgmQ3/SA2Ic08ayWfeFRN1it+jNvu50h8GCvddmMq/xxsKWQCWtT2IF9HqYDzO
7UodsMRUnTk6M/wzYcYO0Y5NpC2dREabUJzx5XdGhYsW2GON7H6LBuVC6d/2YufdGrnE/vf9J41d
w6Q96rsYtRK01tgGTrJzBhI1BkMFrZ++LnzOThOXR5cI5RxinoQcSTlJ/2jJrEXXMyQpGL2TlNLF
xrhWyBAyAfKzP9vOmxmNrPWjz0tmaK40SCxO+GlWj4xhMFn62CD4F93z+z9fZE/lBKhn0y+5YsXG
nnxsK2sgOUR18Jxu2TMz84EvAQqDZvPIRHvrhx3/IpSkVe31pjoLSJ4oY5gVYGMf85nU2bMN/pr3
+Hi2TZBiuMcgVEZJM4lZgI/kDRfDDAwSQpOHjQMsqIYoEL98SzVsZSY6KhBDA/uTqd8assIr3Bku
8CT972yr/YFrex+WAYHATx+tI5nylxk7GkFh7eWRKvWn0MFDDpovR6aCapGT3AtipkuoNVyZAPKi
Yxp7Hzsh47JmlUUPN/xaNthefYnDOYdt9IRAQomaMt40izu6C7u5pw/sYteS2kQr2fOfc3Vuf3Ii
0e0XGqpjnKRKKBTfEk1tVmeA0VhDLb78WoP9LwKJrPm5cGINv+E1BsWZupvERgMi9JxndJWbKxcn
Z+eUl6lPRwtJzW2e0jxjkf6040PBGTWBm6uefEekj5UOy7qJ/HLTGZ+3BVCmcPzHDle7dBf1U3PQ
a28Jj4PzSDUgS6eEuelyWpWv8yPpKBxHnFLquspcRSvt6TxWW36Je0QpknDm5VK0zJNYlH2a5Ske
PkjLLHc0qd3ZsnhoFoGlhYhRaUanThOEHdgpesMo9TB+g1/dZLyja8L0GaxART/fR0WtY8ec3xcQ
AjC7JkgukJJzqS/YrtkRrG9vwc30q6Uui96JRiL8aDYAw0gAvRH3ik8pvAx0rFQJy+6oEAWS7w0/
nze9uYXEayImGkfTeQF0zBQ30o7wTRu0RnSq2oTqDxhqIYdu6ubo8W3VU1aa3MvpZSZtXJg3DfWE
1fmeBdqQ9N/YMswOXWkScO7vKa2MlVd91MQgvFsWC51q6TSf4BOCIvEfshnYkUQe0tnmZ26mAK2f
/X4/LA0jC680PES4zvX/8waxOffS/rNl1WRGhQtfPdsCR4EuxxIeWllh5oA3sXPVI6XGthljcCwx
9Iurg+wFPpNBb4uKXn97U/arXFqBa+uTvHQIKhtwgeV/pkyZcuxzVogwGNXWGIG/vJFsExPtiGiL
PKmGTl9KpzSI4p999TAHZ3TTfXgCfvOJEY+HEDtM7wJc88Yt3zH24W+Kxvd4pMg1a1hK305nzaq+
OK32wYQJ3PpcEUThi6L9jvvURXvBn3uzJUWOndsyvH9K15J4RB4jviPki6ncgCLNOlhdR4AYRVFu
sj/RbHvTT2gGEuVgcwniyrLyVg1c2w6VYReY9KX+2x/2ObzMfbaMcI0hlWV8UjzaCmD3Rmiqd3E4
U7Ic9hEaxZ322skDjJWU3p/GVHDqMCek1NNN1p5TLPfTtvOn3bxUIlt5wOV8VMP5sl54oXrxMJfR
eiXeqMK7AYQA9kYpVxKH5F6yVESoGFVQrI2HGAAPOiaSEf0lLo2eADjVcaAInc+xUMTiVHsNo1ZR
r9bTYamPI/cXUqTShfaFcfGjPg/TORPIdcnIynHOGqpwlzpOT5N1/TzbT5BIZb6bsQaJOsxBbnVc
L5wYlxaeG43MRzuXN38uzY8ZOdmQ5HlSDt7o7JGdzUrZzzK2C9SegI7NFHSV6/V3ZegE/TQJxcPu
nYj3UvGqN9uWoVq5b6E0wWsCQcVHMkWxtSuYc4LWIKFgnrS9MT1vW2K/N+MFhLpt+T2mGKPHurAB
4jfC/tbi7llbEOgdsUa6Skpgfo6O/jLAPX65nWsy2G9bcBY1QAxWqhFZiaTWvFAcW57X+Y5JKJRp
oYR1ikaZ6+z28kPMcmFAsiixeHsbr9dxGD0ztNGSJNM940+8rsFS3PcwKeMHLT3a6mXdvZH7IkFS
/Ii33QhCCEI0hVqlyeZs54JmHK08zjfRAw7niEiB+hR5Tm3C29PIHxGsCqw+fpFlvEJNIg/HDdXX
yV9bXhAUCZXAvC1kwQLHxiMXKINTBnqYH8xfL+7XAmu7FbM3p8NV5+5y9oVxSMXFnB54LYDGFlOo
RNNO2hzaRn9O9uZwThfhDI51UvGr1aOFro/E9VeLJrugYtFFNv7WT6JT+9jkVsMGR58VWRua50s3
ZbpB+uHWb32M7qbnDws05R03RifwQiseVL5fF0AkQCrmo2YwoH/469R9+RdD15PEGbbYXe0ZUsXs
C7n3zx3KHAM2EPehQBGPS6phVkfXCz7APiZxnvqHpaBzhYnZxqt0KNluh1sTxjhWHDNkOMm7aT8g
0JvFQF2qaLHS5WpMNw0UIrJlpSg4oMTiikLc2X4VIqGssILhDuI+UL6u6fwE6Vrbs2wg1ynPKqBq
xoDyQ0FVNI2Mp8Sp77LRRPaQbmHLVeKptKQvpJHx6U5h0i1LcFVhMLXb6A4a+eJkSYvOpv4caqxR
O9am84lBDPzBx5JX0uEboORkkKpYZWJj+4IS0WydzVN5dtCQrOJpshaRDWMuuy+XvIocT555pVXH
hmTY9jny/G/vSBCsFBoOyTq3sj/KTUx/tOg6f3NUcCAIvp8kjF58b2PkcRPpqr9Zz+OT6VJTY31k
X0PBBaY5BnzAq/ODmOqbhWNGwZYhfR8DXtKVEGN0z11yr72kGhpTXgl7TnUcjaSr4TpQ0VUF9RFY
hkPIHPig7JKaINXa7GwmmofweIP6qo1dFnB/G+bDyS5d+/4zHVyeguJH9jYDtu+VH5tu+2AWGfzr
pU8lO2i9SS/ScDTpZpxKGX4vPY1DbeTUO3nxKkgOuQSVV2JjvHrSeucPbD7ONpltiL00gKM/lbAW
L9L1VuOGIwBZGDWwyw4clEh+p7gH6Ze/ym9muk0F6/wBVRxwvx/lyoLSIXzcqHI3IBejEO3tOFa3
rdnzynnRBxGaWw8UBNod490tLh2XxXbPvawEyE6EHio950pn5gblN8b3e/fUTPNZwLYlYnFjjrdS
N8IEbYVkOUjO1C/ooTqCUjb6Qo6gwi8xSfpDGDohGpAvwSS26Yun8w1x1G7YoeGJm3F+s3Lges7l
ACDVfHnMu/l42EkODXvOfNm90PYbfexGc2FIwiNuLlQQUiFDAU3olwhwVUBv9+A7pXnzkHS0RJ1F
yozOFz+mVd7ATFb08WN6ph2jdhjS06aQcMJg6vK1V7Uh1+ne1LTJbioHXzSUgtT5viaLn1nDRoJa
dSxozvFEn4zxsAzNqQlrzkC8Gjazda3bwWb3zz5oqYh87paUorrxSBZtGj1fH2kQKgQfQgQomVIl
i3oW3UnwH6dTNGrlSxRuv7TyHz20XhdMGl2JeASXthjVQK90TrMJglG07j1MgK41FN7MZ3GVD7FC
h6Uo3WKjrYJ/VrCxma/vSI2GA+Fjkqibs3Zd5FNmMPLvrugdBtg8YHfmZzwpLzD7a48n7mtwOEqH
OqTrJLEwUdXEnAEYfQqNUSgrH3Va+L1SmMtPEnn/FGI6tQ3cKcMmvkEDGH6f0sxZIngv8Qw70ebk
H9ebxBzbXPfkpw/o2PkF/6pGw4ECMkIxDX2RxPBV7k+u1cZQjnnyYms+7bGB3WP4/ekCxkssfTor
0bEgVxUQNThIJZYfs9Q86wg2BMrtC3IIhL3pkdeW0dj2c3BvMZuE9IX/FKX4ozTALJ4UAEbwkaRT
QNKNtG/yAZOdUEqQIYLe4lBdDFT8mONynfGylfDD0Ha/ZrEWOT47FeXXNzfPghCoU2eQCVcafwmJ
h3MP/cRSrCZw6Ol2P6eChuxwr1bLL3GV+bpes806OgH6Osd/MEaCW/jP8HZa6XWBX5cL8Ej8BGNU
k4JKxXoF7tC6nPq5VfXzmpttHsa2pBcrIa82+/QGWHceitWAcOl0zg7JPZqQxFXlw6/F2QGGkcVo
TvtR0TCJ+6iT/Jez3x6CrI++W5mP//FeQGkRAUrvMd9FpmaQ0MdAeFE0YMNN8w2JlfDe2y0BsK/3
yAYavC+g2EO2UYdWh8abz4pEHcEvy9Wyj2zJTcxxDpZ1/ao9NrvqAZcLDT+Ucga2d8VHd2I07p0x
eN7v34JjQiN601NtsFVu4Yi3dY2mKOpHwabAH/Ws5NQhcKvJ3BQQ0qB0lyIhVcRb6nV16ZP8Ch2V
hDwUVo8Soep0Rq5/n+6cNDXP85j1JPUNbuIkYly77HV2sq1Z8baWwnbMIW5MzqItsvRuhrpt+JKE
6S0zwMCJWmgdsyLDn6EYWa1hARYyk2IUxlYpn0Sv/D7BpzqM74rd+mfiU2/5+B+LCiJqe7MHv1Vf
Hu7G5YVUqPqESkQ1583ikhnD30DGjJQXh/lw1BlQHWKfKirDRKKrQcR4rjE6AolmyNtCVuHqjtZ5
7+yqM36mh+lJxDcazXtMWlOiDYzfLrd3jf2QYS5Yo0aBfSnPSyKWeVf6zaoyM4uTVnPaq0XJAWcx
nC9iSwJ8kQdIeevxz7HDST3VAe+tRu/sjIJgFcXdPfK5kMFYLUWODbky+s+Xhs5Pdpin51t7rF9I
5pyjXlzCHJm8U3o22q39FdVb5G80beT9YoFdRiyNTqmpstbYgt+5irxz1jBd8p86C/5+0B2TgqNk
qzHfOgUxTveNi+SVnx/VRLHfdxT5zd26dFl8sZHoA/aNBaXrvEaUJYE0DkhARU/Xzl4czne+7jrB
oKHSzYCORu6B66gk5F4gBLrWRJKcH3PdXULOHHVADvv9bTheDMiUXW9fE5w54O30iAGZMb/8hl//
FuXVhgBiSdacZDr5l4h73DrvghrS/8c/CO8Gb2Z8i2SaLQUHR3Z/KHXuLUKpa8U//fguTzbEkmL7
LD4Pdn8xC+Q+BuPmouBG2Z/wQNzlQTnWgYG44YnMcNSkzuiLa+JhnyZ6PQn6CeEe4FQJiYxE2nPG
cZ5hwSHO3rKrTgPgSbUIdCXxAbtpSB3O55s6xfPOnkHgwuRtIYlArEfjavKEcR3OhUBFsuGosOzT
jgXGUv5J9/X3ZAVqES4l1wQXeR98fx/qFNH9IdBjwFFWz+WEdNAzZ/hf3DsgENQJb+yiJQmtHS/m
Cjq6jQG1dmhp3WSlZgakAVixjO1vmmPMP9nOBbU0rx0AwQoFZ/1ajNaGKqx1kU1X8lrLSr4n9Fuu
UEklF7ilwiKr11+gt4zHTAisbY7DXaZU+AZetbMeeCJNlCwgiQAzdnqa5YvylZJeGCTAk1OI3PJ8
6y/iU+Zr9JwV4tbuSA7DuqVwtmmuQQdU7r71Whaeh+XygYkR6wC1+yThdfrG6BYK08BYBQ2MeSy3
jSgwEUM2ShkIAPwhbeMs3C1H6FrgXL3zotgiijzneRwtPGUCeM3nbu525KWYrej1AnzzO5CTJFoM
VMnpVoa+Vq3yLo80CeBH+cWCnZe/JHXSNnRoyhVHXx1oVHAkUfi+bNhjmVFNAQRM6OK33Z3XHqfj
+IhCAjU4fj61w94/cvbUsehYwdZQWlxEOZOd4iEijAeulN0dcoB6W8aIYMlDG24GWkP1oOZYdKse
Gb/V/QiCq1tDo6hKcgth0nsDbRtGJ/C/nU2XG4ACsIM6tM8V/M8BOQmVHlN6X6OO3/e9KGsaTTvN
YStUfeuS9DX16s1lZMmVmhVUyteRt/5HNrpCrLbcPyur8Ol8iHbplO3oDPBu/+OIlioTMzlO0YU7
AZk76t2FK2nKe2b/Ag7vMVpBjdMekGr07FXsaThtqGZvQzhpi/zzawuBwYXa850a4VH2LLOy5yMc
eveWLEtuX2h2bEFdltTjkew5VTKbOEANM5pIcW79Q9Gjk7KuOlQy4zV5JJf70PAo5KJSjNspjHyu
lP7i9LaqqVZNckztmyjgBtSUdv2dph2V84/s+jvZa9mB3nO05zz+Ea/Y09hqgqhlLUTErvQeItXl
HdKND/4+3GGIyO3gzDATa0lfY/uibv4pOAJibnqKA3l0xwEpliO89bT6ub8VnpEoN5rc7LCFWFop
Ze/uUvbB9uc4mD9FeQg1xHHeTZsuif2AKhiCxqn7NUT0iTGxXtnvRSFOjjTmdcGnZQa6nOeLkj15
xcgwXOdr45s3jHp2rtvFWx8u4p3PFEyhW3J3yTKCA1quSrvvzhSvW4TVTRMnHuFhbO/NyhXV/5+v
5nj9TP5YJ8NV2bGA3+zap2LL0BIXhd3wgJfqA4cOr+J9WU+zFzlWe/thyDYfRMm3XY7BLo5BeoKp
q1120A0EGLrfrsdxd4L2scaGKtNjKVGgiF3/8nSfxHdg41FBHwpzb/MwLpXSdWA7yl9s/1C3ycbV
WfmkP0dFWdwa3JUi3bgIXfwDMjSXIXndOW4rbp0YhrN5xDfbEKXM+HN7stIqjh9ulXYcRXPSFdYb
1aGHlTN3Z2J0uPzIupCkIHNS08GcJcKumWJHLDTvYvDKpic8L03Mtg4iKyexIaedZfkfHXNgN2Wg
4FM8lns2uP2NTv9gzUPWk+ubM+bPZnhrAqNHz9c0rxdKl11GF/f+Cm7N2+KL/8GFQ1tOOcKe7VWR
eIkC6HmYqjO68Ndw6O2ifregPPzlYYm5Xomg7POXn2VSEDuN1MrV8cD89xNtvrhqsehqSXJhopD2
GESRk0VZXtE0R7kU32WhjklGsCM7VqCX0NM4kEIQXWecQiflGJ/7TP6p5r73I/lqfY2Fp0+zqNU6
IOYqdGDwEkKNN3UKn5WTzQ503SpnA08W7Ii3wQH1ASmO015J+LZ8l7maqoCazTKz1PRoGpSXd3ZV
1risFbYWMeqkAhfLz/S8OUlRRYrsTSgXic/qovwCmBmteKddvb+ZG2rFjYl6X0b+/sVgATVNR5pQ
rDXfWU4D7vR7hPvQNn8JNHF7pP1PeSM2DP325fJK9UOTgT+LCxgp5M7JsbkeYcB6usjYYJJhae3n
hBBSRjiMov3xWltOIMClLNqr/GqtntaT8mHp57fZYCu4D7o2CGyMbTCq/OuZYo3CefBik96T74d4
ihtnBcuTnhDhVo8eawORqrO9bGTmVKgQJ/nsdNmpFBHHmD6L2+jckIGijJp+hwhJ2lU7O5y4wzvC
mUSrBvh68nTs0kSuYHsTjtI6kNM7EAezMAJ0qYyamJO6CQ2Hc3IVtLMGIW6Z5t61qVqcAuQLh6/e
EyAdgyL0mD6X10KazPsRUaNP43wZHXWi8t5LGM3NsBsH912TgzzSPyfO00umLiOl0ATqG281CPEJ
cikorD+F8ms1/VRNVh25iIDYmGpt96eOEIVtCKTFlBHwKcQCKT7Ywt8jWvmQQ5TSC0Bhno71nySs
qXexjFKXoInM6l+AgcGeC15phvRT4rl4Po1Y1qtFehdHDPm93fPUcOYXP8gnNf5oaMnDIVmMwuWD
/OJvMitoaDufg5sBQFpK+y+LDrebZLJb31wCXy+U++jynC/PZYPFRmv6T8Oly4Sq4H79NMJDYRli
930Sg5uaM9psfRN+0rvR0DP2tciTMS6wl66TStG/nDG5SH/CWTT6hUudW82lXXwmNmKRt4ddVwXF
iM2Die2M+ta9NIIDffWe55i1u9rzwD6Hzj+gLhDQVmngoGhKL1cDFNNqDwOgFTWk0bA2/QGO7zOK
wkMPENCnE2G1jLfeTNBlCfERcikBZLeFE38xEz3+g8srcngrdydU2q7NF6kgATueIRrQIO7k1uVo
wqwgujm5yU1CY6XpAurpDo+OS7OnGQ5s6nRiys27KG2tkWU0oLsbGkD5y2bKUDXgAbe9dmd+L1l1
eo9BvGrRgn02mMa2Qn4/cQSahd15+jC8hlZhsaJ8Rh1ZDhyNYt+J4BOv0CELrLdROYCJUtuCi6z1
AFJXvEbg+3hvfeDF3Dcsh2DWEb2GzIms4qYhqRiR/9YDkkWVwkKsHtq8HCX9MdZBxN2Xa5bgsWRO
J1qJlxvmo+uabEFLyDXx6xlYaJ6kctxmDwS4D1teb27pyb5h8wt0pRhFynlI6nVeHxeDC+dphn3Q
oarSmpJ5jHFBpQ6uLGTzVrSq3vFLvE0X0gom1cta86YVXGGA+nflhaKcA0WfWhCgCfljE+otl/3B
CQh1Q2QsWOMD0jIBAWd21X6Q4m2N9KrK3O1PAk07OeIy7UjdlAyKR+ryEzYG9CaMy/y15WT04v6/
L5LmNYLQbRgxMwQbhLUA8YWiePt2Y4Bip7fEDAXLGOo1X2zFRsuhSF1RIBw0puY5cznTlLrkoHIY
BZVR6PGyU7dmddupqtLqmNAXTH2120PkvHgTe5gEcDGNrtSbGm3evT0TLOa8VxmNV602xncLpXEE
nnIQrcBOHlNj2JOGJmlu5aa3fwCEr/zl4pDBMPnf1dlD5V7W/qFrUtoF5+Rot04+fXExYynBDTkX
3OeHNhatrq8bC+aa5/sM+ntQlLJSNw+5tYZ94S5CsJfQhkUwaDl9aoz+Ol/wtJvHYYUu5yUNh9Mz
q1oOOYfgpbbXdThH6O9KuJZyp/i/hOAGuG/4fTccmRz0o3JVvP+vsmXh6HwjnxmM/tZWKWNrtFO3
6hvssWXeK9/FFy77QpGYVbucGle2miKG9VmBxAa4Peku9MGSCJMhxYEzbn7dNrPhfUeDzhWC3wj4
tjpMlJ1gXyu5wjjnyUbI/Wfc5UzTARRdodaUPR/rdcIO7uvdCWi0TEMYfvFnBzMNUBXB/Cu2eWmh
448cxnDV7S920+yUpEkkBN+j9/axQFq7mAtvViBb/tPz48Tw0fx2ecgEsVlG3iNvgWy9rZ45WoeC
nOLkaK2vHvzv3HfhvH8XSFfc4t028whQcWyQd3Pjv6vRJ1rc0uzwQWKZP1W2RQHYZApru2AYbuqX
lHdgy9FkCowVbKVSutIjZ/T+A2PeUS/ltBoT/h5mveiprcs7S8N7LQODf/SiZ6sxG0Ojl7+qLVOi
iMIYCJ+chfYm9iOlDenpIbX2pZAfV41nfqCo7C+4zQpRaEiMTF0oFWerfOe3HJJ75fTZDbMO1uL+
96tJJDzsIhVlRL1g9wz7POQKPDtcKUtcDjJMJpTbGNlh3X8L0tNXfVt/V/C/imP43nY3nCWOMzNV
rz7IJxW9V//Qgt/OeCOreBUsySohmHyz24sbaUPeRtEZj0P5Gt+ppvm4p3U34S42oF3g7Y+Una6S
qeh5ZcZxK5FIdWDBKXyqVZX3g3NCV06q+VKE+/ZFBLU+J1tej0BoYYgaApdiuu4oPq/ejDBMtZXc
8XzHkATSjOESJ5zu4HGLzGNWYNQxfihaWIm2wOr22SQWoPcFaKf97zMgdaDTgQ6Y7+xu7S+XddAV
WP2ncN3gAt39jiSsvr2QJgjVhvzZwG3FaBO1DLCEOcvOM5T7PfULFxWJhGygVC0RVMmYVfXr8NF9
OPHOjdwSYMTYrYM0wYRTbaKpvQco5mKHyqdSE69tNFiQGNhlPxa4lRNGk0Eap4nDwsV/K6KXOWI8
P5st0v9bmky/5RzL4V9gcHwhs9bBPXFYfxh5ifWMwgt8RTtY4JXogDdxDRdGUCpM3acGe+kPwmFa
tZzEVSOsStFiTWWWBWxYzwr2u+w+AB/offPhGJ7W2pDIrBWggMTROx1JpVYK3Y3AYBOEJ4g5na2O
HIyhPCuPCtW0GXMV8H6LWRbVxNZRK5PrW8lyG/SLMAPuMilssoshDBD2mHXajI13vPp2moTXrHLI
Q0LWPUczFMLsf9baW4xSGKuL3B6VYNYXY48XHr+rJfNfJ8JJ5b1JnBWkzOUR8hwwZkWgUaj0UdSK
a08haUSY1MrXqRa17CiqvvWMVrxsL3So8uUyokgFkbq/Yquh2wzw+xr/jkx+wXr7VJnXlGfSMd0d
ejvHHI7i9Bo7d53gtPLH+fp/62v0qQT3TEk7OmaJk9GI/j5AhF2fSb2ATDuXWKd160YU0P61poHI
3wjTkfOeS2aRIcngZ98kV0BoTS4WLYjCsGNAkAuN3xVjsT7u+wgbndAQxt+yL59G4Sr8asuJH4Vf
rEDl41NEI4o/U1Bp8s1qyOsmfTL7pINTefbCt1s56ZDMBjkbL3YoBGsDlyw4GS31jdEXNwJXhRJ9
QttuRkJ3N0m5wbNoM5CFuFk9xcU3/SlxFXiUrdadE1Aszvxi1iiHJb9ohGDKsrLNTNevspY2exRW
XSW3qGOZOp2Wecc+JXZ2MvBvaC/RPdYONROdw5lMnetbO5W13MFcy68so5EI7zODswsQSMl4/e/c
NG25v/eF3WW+dlkHofXWwWXSPtFCpDY6qn8spSfjtC1EpSrv/bY0doPxeBdWik7MnrPdp10gYJxR
KS+0y0RG/yfwMZpL1rTW2HPa0CrFk9WFp3KmyGaQ1bvTtEoYlkEQEtYFfSJpgRGJryKyXUcXhGci
9Fd/YTZNtwSxdxa3yoGdwD9AzalqMp72yOd8rAxYfncfTATwPYJxzbpN0TcUKwNRROegnq1QJZdf
Iv9tjUZcL5+pfBOXAhskzjm/3lz+Eq39IYhCC7gVNGTAwPhIdpEe0VQdd6Xq69D8t2S5iug5KgVM
rAviqx5bKQ+GRMjxgf92OlXfhAfVMiDOxPWZaA/sXDrasroUAfiSO+bzBfKdrV/Gk3NH1xah9Dwa
OUs8pO6HFwgaF8Rx323dtUk4aYkC4LYHz8xpr5+ycX0Q5bACktyLH+q2RI1RW+y8WBZiQ4ULZ3Nf
bo5u7eNYQmAd/UHrtLPMpVNd3uTlXptAFzM26bEwqdCtC0lhuVSgFdmpAZI60jdedSzJlDSBG99C
ht/z/dHQIdVIc3pDaunHV4am0JWJyeFVdZm3/1mfYGL5pHZp9QrwGgYPU1jy0fqZJgJyImc4ELew
vpCZhaKanjUxnYky2cLPbZuDtTCNFGI7m3JTuGwUnE0VBeLs41TleiX4TtYNomMadiRch3HLupz/
mrJ7OPay/+JM3dBYkRX0TLiMyuLoqiTU66T+Tteh7/jIFXkoQq/4Jtrj/Gfo8Rr2AmcdmWMzr4BI
p6Ed4l6az22L1sUYxjSlSBwCdcD7rjKMtviumxl49XYU6KIa9kzWGXrx8w9pWWTTD6gSwBVLqgNA
wwsg7+Yx+9XwiYwH7Ncyg0XHS7uFh4f8WsOfam86lgEMdbVlUb7N0XMOsEBHSgsA1vOYqo8Tkp5x
yXL66LxBYSSaUWMXdtNhyehcYAWZpYFdDZtLPc8sWxvLw9vKtgzDU2j7WBRSRX5PDFpjMwKoJwqe
YT8Jn/Lq07UqbScD1McB7BflfqZG3o5QU3CG7IA0DzqX1PnMARhUu35z5eKPrcYxGy6KB6W4i5GP
FEf5/fOKvIDERStd5Aekfc6dY3BugV/VPE+DFXaDXMsDCNJrfBTF8nab/rXDx24E1Ul+rCWLS3g4
VMyaPB9t749LG5pRzVu69ebFrsIulp05wZvmDsFYk3uotBdyk4kMa8c/oskk+/OXDi4ig/0j7GwM
+15tfxaomRrVVIVmAI2BdI6xQnPw41bc1/d8BpQoVkVW2abvZYGzagA7o6OKTQ92JSCOiS7B21+o
Y3EpbApFhkoJ69EoFr5U6NRRhB/GmsG/ePbOtCFU2audF5BTBoh/DAKZciAH5RCRbYHLH2B7Roex
E1jlkjfDN7C889bnhFwDxGpra4tYxzhGPUwiQz/erwwj3hlyTgyM3SGQL842RHsgsTAka1JtOi6F
B1ED3KS4/o9uXfs5ALI6mAklcd7bsatIQx0Pw7yq/q2y55uicJI6iPFLhcLUZP1R37R8S8TBCMvt
15DW1K4ETbiiiCk+uGNEAkxjZQXsEczXdMWNJ9P30df5u0vvPPKsHKpExVYc/pVnefVfmqGwaLvk
oCFof8EeqUQvt+3uz1fTpOklYAXj0rBI7h8daCZnLD/keS6l6DAQEW4pJbgqpeW3ex0u9AKyCPHi
SJhfJ7Qb8iD4pebtOV6Q5EPlRtJWni9Xk/Szyuq4yHnZwfWUO4EeynvOPD4M78R4zZCw7gApeUkK
1dNNRcQiVCPGCq8ejelm1EV7FQybVhOHBsJq2OXaG0YXxk0fm6qsiVK0gUJrQ97mdVPcT3yK79AA
M58E1ESUt8Xsbj60L05rKC99nGxJhBKGl7VL86ntgwCi78OF7GF6GHQ+SSxCuoC7MA5+P/bfcd2t
7VvOVDJnrEhlY5cEWf50ptHlrdufuyPbZJ3FR//WpR3sJ0pym720W+SF8kk4/JFKPjX+K1JnjB6w
r+X4JJujcEhb97rS86hPLNyjqp6d/QctNE3xuEXZcRiTVE/Ym+1eA+5O6czmeN6GNJmn2pjWzpXi
PZlc4cPv5pSW7VgorKg8iGRUquPbOnbDydfE2er9vEJqqHzcFJRWo8FK1fKj0n3z8XXeQHw5PMHi
UezSUZXPlyeVSKde2Bvg5KR/ycT5B+Q39puKEl0WLaQiB4Rurqk7fIPtDzVOoqcGF6xbLPM/NvgO
lkESW3o4JZNe3D3psgPF6LmEK+271jKFaKbbNI7ePVYOo45LbRL0rNPuRWuiIc/FcuA3lpJ0mi8H
gz4Jm9k5aKDQkP2d/TXIl/QTrYw/Q01zWb/aPxWV/6K8FgtfpU0ZIsZb5hP0Hj2WvXx732/stU+A
V+nQnzaM85mFm6NRwsNM+x18TLP83AHSEQmYoHpTsMOcHsgNr2llzxz371ksFXigLt2yIBGN8qEO
jRQI8vfWrvHLnEnQV3NnfvNbLgvVh19LtJ7g+7+7zODihgnAl3bsBe9Vjuqa/9f/tzrGjzGfHgn1
D/u/4XlUaOXEqFLV+JJ/8H8Tur1zqdwbmC/ytx/d3jrGkfNf5bvRjL1aVVYxjsnmt3kqBNUEF/Jn
VtYSC32owA5fwyvFqznW/CAzrgqaFX98LhWJ9FSgICXaGRLHd5ZweAdFkLYc4MtWONqzMi5V10Gz
KQ2Qdj8bVFGyhrDpypcF9R+ze6fIkyDp7BAzu+gP60eHkcWo5+3FChZWx3a8s5jHisVihy8kRPdN
ydTUbPWWs/uGrWTlVVkLW7CydB9cOf4xPeyPq3D2SVysNLL4uhAErMeP34Dl5DXrT52yROyz+Eso
Zu/D9VE2ThXn6Xt8d7NSbhVxUkYaoU14GbNTiXx1ghuewDJSULrHVhGxMkQBm9xzBLo28IrzJsqA
8VpM9i/53gLP5PIERPq08LgLX2EpVm7QtnTnTibovbltSxPCbl18sv5/jSVIZ5ApiHgjFZnhe1yb
kFuov7to3OQ1chiHo9DVkbMv5gOrAEPbe2zMK+mQy9cXsbcVQVSi0FVd96BLo5jJ8ykXcA1nVvjk
ccilRMI6oBNrGTgyed+/mqZStCvhUVGUB8fxkHqOCWn/EwOuY+0qCLminzrU339FTJfKGyx2HCVE
aHi7jxaAM1YcQIp3NK8Qgtt9lW2fHqWEEsw4XNr6fAP6f5m158SUdCOdKZ58/SS+fr8EZSjS+Dpi
hHhSeOInGK2jyQ5wM8/UZO7iBtjrKadn9sF4XEuo+678HXivdemt6mMumGrTOLWc63hGv6WGgXIh
ZK4CVxOfIc2tX/5U9ys3REoUtnr2S9EzCRcKhUFrgvl75xEHTZ+PnRNU7dNoBnz322iKXb2e667K
dQ13dKQcFzb3sKFr8Vow+fVEDwUBHMjqB84LOeGNyClymiTpoeP7Bmhl+XL0rFdJChvjOeptGP1N
/5BfdhJUVQE1laDVCAXat9th+lahsazpcaL2uT3q0eBHNakicgXbHDnLQSJ2Jqs246uvsv2NfiRS
/v45QP1izC7i1bhd/zDf/KrvyC81gwjarUn5JdnPacBYUf8y5v/5xSdKupexFCRJFs39pZSHyEeH
JumeQTMI/sYGAyxKlHnO8+/zDM6H76fBuu+s+xeiOTlCnVsRgeRgx3WuXd3IX970fL0wlGqLiIP5
T91dii5kMexdz+wh8YqIFcUsZVt0MCEvp942D/Ydq22CDBQz6pd48HNuMBmWBFrp7JSaE4kbV7hX
B0Elherq/gJlYENOQQrbrhpDNfJzEUwIo6Psu31gC7X/W1bI5qNQJSBil4lqBIER9wzVhMZ+sh7k
6D1+QXIiwM6704ADw1RzZlsFnq22kLxmuIxKvQppYC0qQm43kmK18jhYWh6CPRlIrz6lX2TpBcGn
lDKSdV9uhkh9vMwrR1PlHwlJq6aZVNZE+P6ui6gMRWWxyh0/YpS818xl4uus86n64qcQfR5YjjXn
f60YsXM+cL5fiBFxgavzraQbV7AWk9Oo/BxcJXQsxe3DYL1bC/hmCYwKQie/P2dKlAM3pQ233Cjp
fULPg8nmOKmZLuoMC95Nq6ZsRxDRyxdQT6qT1alsXUehvYIKbmNUu2DZukIaCWOR5qE/upbow67t
qMDzG13+8UkcsHorwM4qByaAdiFMi++lKmjr8YWs2bvgiNdjONzkgHPfnMZ3rCDL5lHB90MVH8lm
WngvVl0gccRu2NIdlee7V/Fj6DapYoCDsgovT1mM71t9IFM3Fht0PXRVzfg6q/u3frfTsByQ9Jun
jztZyT7VZc6/Q4ZpACdO/n+hoj05QCe4coxbasTF+PjneFTWLF6u8XkwmR0yBkr6FBq1C3yLK2Px
rD8mWt8jSxiCU+cWT0I9cgaJhcth19k3c6YIMDhy9GMTPrR/HIA/Wua4Sl92fb0907GtRQzwNUhs
oa7Wqfh2SMzKA8wVpr7ZnF7aJk3yDq74PLqWErAzAtsN28rkJlK0LtEX4RwtvrDqIxGTuWtV4DWN
n1UguoBFVFf1EkX1lYfhG4SKnPyI35vu05NasRC0dn9cu2fddRcmdq+1k1cq+synII7c6fJdXmMK
i0Lw4mdo6GqTlGXyjd2gumqmF1NMXZTG4sVbyxoIKgSjtvGYk5gIDFV4q7swl1nuswsPWXVA+nNv
3BpXQVOLexS1FX7wfY05vfK3E9UUrOmrXC5DcFUaOy4FxBmF7Sb02+ibPCSd8vrcKGXGnn1uXTtV
sg667ARKIBC8paibY4tyKAj/uPn9U2IGjdbVJNagoeQsh/uULkx9EIUYTWalBhmoprjPRcxo2gdd
9Eh7HHCSaDslllvtJTAzUULRMBB++3NstRv3aKdTlL3ZO5oGYvWj8i9xDOX3X9SKGY3yP6oLGBKu
P40Nu2cY9kjhame6nVkZ0FFECJt07mn7gMaznbXUQmEcaSLVpK1nzSmI/aHlXT0MTV7i/jBqu9TD
6sYEHT2phR6mRNh77b0ZTwmVouuY4iJYT9tm0qjTqzDtgwUNyKgMKXk+13fQQu6C0mGtnQFqm1x1
NGFPt7MBJ2yww87gSVJygdZIWW/EGV4eVnmNbRuf2PPZBhXmAUou8YNkz450rT5YzQInC42Bjo5x
o0bjFauQkcb+Q0OxsOWoo0mjMbwgBJgCOjBXNMfiRMkDgKO1NAWEeM/3wBWwRBb3lY+zD4voORui
A8dOZJltn7rBr812W0ZHOSIqXlTpkUAfMly65kp/ikfJUJVzKw27amFxW7Tg6s1K/20P7YEH+w+p
dncIOgUe7d5864Ze5CvutxaqARavmLhnGHCA7S4Ii9l05O1I1Y7i8u0drUWEWQiWSYTugT1vuZ56
ifMrXYLYyZR8nykSOJEHsGO3ITSsRTwVK6wFxp38S3/BggYkeI9FrCIC8HOPx5DlN2B0Qu0NoI9B
mENnxTPulyNYTFvpWjD5s2Ro5X3YjDGfUD669DuCxD0ORS3OC3prxzsu4tb+AEOiOekBTcDawhXM
HrgsHocOGCiynK4ZkfdxDp4UMjmxZk4gVfsnOkWQGBUb3VfJXJHqcwTWrfoohVnIQfIQNPRTNI/t
dEOGHAiv7XbaRu1Q9qJAABmxRCOL0kP+wyToXU8Rv7U7LiNWwvsmaN8nDgIuI76VXc1Gpdbq/zwB
PLXWC2TeFTGzP9SiqCPK4j+TCV8RM9j6z7IPwATmre1retiybVJDrOcPBBFD3UwA4HrDRUSN0XZB
jIbJknMAo+mzCUr6ne/ngm4ZKqEwsdWKoqvyH1yJwBLNbfrZulViPB7bXaDvYbb8dAFl8FcBTwNJ
Wd5yAZrBTAFXjL3LIlIfdomJHPqYV8+KEjoReMwJg81NiqyhhizA5XmJ7El7K5TB/5QFLUGeanzo
m1iHZbTR9lcqfvRYIWI5/IbdF6NTRxnm3sBKVAngpYXoZJpQm7/J2cCsVHfqUMJ/LjA42iEokVuY
K7ZmpJ3a4npJ5ByIJMLg+YOt2xeg0xUonOe782S5zm2KVjWS5pEferNawXOs6l2ub14ie+ClejGh
fE9QyhNSCrCRZKtJHHjAGl2clTRv96ShzB1jtj3vppfpN+i7qgKxMgWUQr7CAAdoKR2V85rduNda
C1ImirSqQemLaKNtLEc4sRq/X6QV3thh9nesnpedDZ934tNVXVDbPCRNO0qgLNSoCIMXlaNVB9HE
egt9Ywlc3MaV5O7bbtBZ9cvleJhGFXWS3yooimp0W1AgYwosY+tHjcfddEM4EEGu4sVJL2jr0mH1
/lau7Q7DKsn+LJuIZ2XzE8t5xQj5D8+2y2XR2CRvxkE0mta49N8QO6Jcii4+up0cz7/p0ntbFzSw
aMQNl8bEHhYhnUq7kOTDKDbfg+kDNTPT64AGByh9Vt3BFEqUX6JUEVgp/lEkmjfTG2LLVMfERTFo
fqJunXLTFsvlaAIM4qAVKY0TAsv4oBDuPbFtpVTi0N/1i6YxOTc9Zd9cSWNyV83AZhYMorFCFKyL
5d/NJBcoq+R/c7HIwWXffuKbuR4cAXqkGI3llrPyrl5Lrf3i6g+WRDDf2vOevhxvOLLU3yWzN8Ze
wPtLLzu7JJoUtQa46pRoMW73S+tKuR/ivWa37bj2QbMbovCiAMIdFbLpm1PrQUgRnGRfOxozUQkD
1sahQLwh/EAUUsHgdwetPhyH6Pt7hcXkzowDCW7+Yxy134inWThzLmaFXp0PUp28BxcSHHIzvf/s
EEmh4zQFbpgB+pzyPSvJgtRPiPx1KMJ09IlcvjVx/v95SenGVI/AiyomRNAE2SoiasQgufCYceH1
8Yl5vG5ZNjbmriEwux+pUeSr2GKxkxlVg4rMLfIGohM6zzEUoMdjJjjgu9M53VhJ9cS3dxu0SRXL
y1/xTDmHTkWo3BmEb54EdirbLovS9+BIV5aIFXwN/cqm66xLeoqTddrjmG72EIi3zsEiOeEsjLQ2
jCmsKw5nzUqCUPeo6OC7eZQO9vf8GfoiuVHSy8wZNsDNHweWZCAlUKJzQ4Sw2vUf0/Y8Cd5dhz8a
agqsnZWEyvzP1iiX0+ex/9PWXYtTQpFoIi+nriSO7gkeptTK+oXDTez3dugwdO4aRWFihyFQ9xfq
PCMuXf6rmfipvkKvmxd6xbuB8zaoWV+vHxQ65wFEolvrPmSeEcdbpzi9TpIryCe2sx+7ATQGk1kq
HbkviqRZsDIZwO/uHawHBmlsDmWXGEmxJ6wpAnRgNpOzjb8cGJtZ6fFP6XbwQNee7gW89VV+89tD
S+SBPcpu2vmSnsGbTs4ZZbKHkVsdE4vxBynCqrdI8YzbdZ3bQUSJGU/GMmBgxaCTKFkF5+4ssZ00
foyDysHFKNgbiLAEDQDgYOvlIHaGXQjV3uRLyqW30GQWA3UR5+uA/Hl1Pmxe5CwxEAev8phzG4d4
Fh+3919seYSus14OnT7lXDGU0toxLm5UPRKetd9fGU+Hs8GFyOe8C1EMfgo2HUwJawZs5tYV1pDw
2AXljFVSFbZFXd+Uj9qICzqXsJ+iGGuBBVaeVDiwUIGQLzKZuq9KkbCGoNsQ2KYlowslO9xNISlg
o7HTeqY/adae2SKNlL2RUrV7dM9jzkz/kj1kgWzSS5YBbxO/eJlXR2s40ueJOopchmXqebMd8Kgm
oGYPixevvRbdM2rVPqMjwlezD0AF5TAaoZrqnyz2HN2PhnFNV81xRRn7FhhN6oLcWqxppg1fujQw
FS5ylptq364z83xJpPB7Na/l3ch64hGRcbIAbm4IYQxNYI8jKA+cMLL0pln9yAmIDRc0a8UQ2ASi
SoAF2Q30daAkKcEwuVuaQk4tcghHvXOMvBOytOr2r1wCVoI+lEew0S9cHMRZdWORTk7GEdZR1v5l
V14+suhM+EL48sbHVzDPOwXxTUwjUoiMpvNchnF45wy/Q0+xCVe9cJgnANVxFBVVmKa3f+giTrjV
hK0v4wgJdKZRcwEPwGGp0YHdn1VM3NciaEQixxRRZRkrFVzQ5BY84WWc6XM62GuJpzdmK7bKyziQ
Cf64ErSKY1tBr5Ra1chA4JAnDm16HR5FKiELU8J2BphH4rWliHlnujl8c+KM86/Kh8MtaZdZxWH9
Cah8Qo1kff0bCtnoHv1qwIuwi5uqWQv7ykv7yndNPCb3IozfjvJvag0ffthKmLxmPXksqzK5DyKj
3R+TfnFLiQeWbyHK8qIrPDZrGi37vszzlb6JXaKhNHCZgcWkDjOOkKnIIDdKJlD90oIXSZSF1DTN
N+YszdpigePopuuImHmLCTbU9ElXm3YMnjz6iWXUCYly4HjAOhieOZUz/kkqi45hVBNixKVp2Ov+
ynnLxO9t3udLVrSzyZIkUucIdWhKViqOxthW/mIwHG3E1zXAb/IiBvdttqtGUQhtLRNDVz1yNWyF
qJxewjphp0pW1IgCty+JbElZrbaOqAws+5pq50jOFCypg4VvO/AFr8XwwWuvk33yNCdh5OL1A2+F
Pvm+lDAtva/T1HQo0oE1OkEKInp2zT58/8vgCyvv9TnoO6fulRb5mJEezIGDXxUEX6eHFxtYQL8N
La2PbazZyJzTYRLEemhvGZK7XZDX2TwECZx0pS0/TCWyhIdQ3uMnejyZEM0Xv9rfA3IdYbn7E9Qw
naygd5b3ra+HUfNNEovicujjW+4ULr7AomIfXSXh0imt23g/2p0oOwg7a4/iN1iozzY8kXtuVX7O
oP8js3vYNyDma7LLpZJEMnwLShz34jot1U3x37LZeBTNapDD++k021we4YFjYzzeu+j1ktiNvQoz
2CitL9Vt6ZuPPcued4jItChs1LUNhy6Wf/0mT3oL9n+OBuBVIjh2jxYtb3xTTpnmtiey4RqyVLAj
843WgncJkTTDfeUnLbKvjV+9mMULXCfcgR2Yvle69A3MUHtsx4D11fsKKrXWV3px3+086Sn5WRNF
H8EikuUvaI5pCLlgGkNb2uJuGUcAVz63wvb/3JM3bGbkwvj+EP43AkfX9o8YZeBYV+zg4mpcDpdV
7hFYXHj4nqRBIg9vCIZx+CpAdDw4nWi++koIWymbl1wgRJV0Vzd+cP+MKm3uEGCJI13pHZebrjRD
Fj02t4gkbeTh/lFHMxORcqvupltbuglLsC7cGjPn9wODRNYULa7sKiU6nwz+tSUh7L34HE9csMk8
58uoVuxjWxuQC5jmDuGDII4vyIZPhOmvArpIkwGLsYFErSdmKqRkmSkQHqDe8nHgaNPMj+LSNg3t
SpvUrY4oBOae15l27aX7HE8krq4ETykAFmbDoet7NZPbE+RbikLIOVPz2jcC4w8rqT1wYfXM7O96
M4aWuE4vOcuBl1y2rPZXB7RJu5DDoPSsDrp9F6g/pCJkYf4y1p8sFhD8lWlAPZIuaUy1PuJapWSW
yhAcOptVGHvmVysg1Y8puj/brWA3PRzk9Xo1+99NdIDOmyoK0gLPgnCL1APQANTuaqx4RnB4CRSw
4h0K8CvKRERL3z40BGMG3NcHASXs7I5++rDAYZPB5BIaEBpznMcFJbKDEv6C6Bbkl0Cf8zHrSMwL
PBhuCx0+0oUU+BR3SOL8pIz/7lFJ8jwCNKe7pjvOgEqFo6udClMF/jjpxWHLsFiBOZFwnigqt5tD
RuCCiuT81o9MfdIL1+NuQmRIn9lZYNnkJh+rC9IyF4NkFCvU9AcT9LbmWJB2aYot9HfcY4Ks+i8L
+lM2RPgH4PlT84FH5krTaIPCPvkYTemgWna8ug0MHXNA+bON9czKIMt5el4RxoWg1/9JCQCGNBkG
Hv9q2HgY9/V55dVT9F28Ko+vOEi3v89dvBoKvX+kEwbSxHOcGqp1w1zX4/6cHPtp/lq5HoWCkCLZ
nDIHXNEP6ZHD1bJx++jcK+o1w3+DAnnzKJGLXzRMXyRPOGZ6iH0M5r18/jUjVkE6tCvqaiTtD+xG
+a9YUiwERL3AFfXzkmgWw4kcFUfqwX6/yUUZtit3znHF+GL6ht1K380YDsXX3t73/B60uc4TbErK
eiOJxfo9szHJQAlXIDLLj+8BZDDQ8ozg8oLrt4Gapi8umupOl+LvQIcrDaSnF+kVtWWpXSxqzSAz
vB0a88HhgWZTBmbLoSAcaYl07naDgaSCUUgpajA2Ps1IVqZu0h1qraPpiU4awc5wys63P/QeE/h4
GwPFZ5oVL9eHUbXqcTeqUc7Zk/1G1aKc+a3t28Ojf9cVJVGARhZHr2kOuzqMutDJw0+xO0QrMj+8
bQAHTn5eoPyKOO0OGftJ29IoENPI8bcmOY/xmuUB4uafLL1vV60f8i5MLvMFmM1ZihmIX9lR0cC0
4d2vU/vmQahIjkBKiHIHzkXmRF1EUgT+LtRCWv3hUQclQJc9k7bHecR0HWbcHUNEzny3vsySB6Cb
7Df9iQI1H5GZJvRZHwS8APgQ4SLRXXSNBBvP+kLmBxxsA2nREFGkk96/GAucEjXambA8GJQcSO7z
R6/ttaZC6c+ZFnNNRbNssKNOLrzi4IFQxqsbYwStcIUUVr4zsH0RP0eyH60DzJIaIHynsp91jJaQ
248GdREMC+pRXuCvGGWwP8llAXFqRkdQXfFhDaLSaVYd0PM+mqVAIyH/LRRkP9eoHti0XnhQT0th
pExRTVupNWqaijXpLLAp9gYcWD/vyDKFZCAD7LnTaFLNj2Bmg9+eknW9MQxGBZxgrS8pT9qtF3MP
GUmR+K8A+ql2GrwxsUbYLfln2kgE7bPZjC3obczyvLHOuLKk6Htb/gusPFYjRwJh46PUo56QIBXB
h9xcgOEbW4jdIYFfe62VQj2uj8RZLxr/YHa6buVUYF2zbhsTazrdU1u/75X3t7brMSu7DxwUBs4f
kcGVWzlj+vRTzK1lvL6FfMggT1oqbcn3o0Qeu5JD1H0PNZMrgntQgbM6KESdaw7G9YZoapsZKQvt
Tnp0FwC9Tau7R3CnA7W2GdG9JSV69Hl6q2gGb3Z3kFOSfz9guL5r2+jrc6Jibj0/8Wnwi4ZdKlL3
9B/Jgp3D0InctX0I2wviC7I0wVDBmzBuRAQVwqoHmpy8JnV0JjU2OgQBOiSzJEn+Z7XmiHlm0z80
vyxmp9oKvMAa2UXdJVmbeIHU8rlsi3TsMAejXtOKUHertgImsoO3+NGIT3H74RDfPD1BILvvXwj8
dT7220ixtXIkjVGkOXogPYy8jucEnxW6+8+ozxiE0DqlqIb8uSIBRRbFKS2AytHIR+BEvY3vXh3z
q0eSKRv8NAOvCpkKwP79F0CKiAD/+oSJgojIzc5nCnFDGqowO0wO2AhONHFcgL395r+U2OttNozU
rmykEhSnzjee/XYcYdJI60OWA6GJVBU+7uWmQ1bfDqlckLebd2ej0wBcsSLz2f/2jhEk+2iMMHYk
2dQ92ItV9vLuAc7B7zyRieBCUAaqUHRwYxwf/L78ScQTZOXnSpPEmJ+qno2MRNA7iJ4Chw4SDtIW
f+EdtSMM8QjDgOJSMsLb4fyvhCFqQ324fQ7wsUh9P3Zff1420OB+eEqnJX+u0E53mqK6td3J+pos
DLbNHSYcEbKeguiYdJ+UfjKygrS6QKABCRLQT+8UOSvsYAnnlozEgMxmMk8cGmIKAmGO5o7qtoK/
rs1+LLsFR7sFtYDeqegLbhdlu+RuYfS2aa4IZvNMA+foQw25BFJY/CcweM3fgjpOqE4MKFUsHcwo
dwQHep2AVf1uWGGMStZNcnqWAXhkms7kGElGQNpsRzOhd80srshP9HMxp9zp+I3ZG1wn8hbeiv/+
8B4sLtkfd3fExLAJuxCyVbhyPtVUDoE0Km6fDuonodmDJyxPJOf3NXMdIX87ujEFDL2tHGcs/uIz
CoUBcPgdrXbduzI7ENXDwRwgChKXMmvMsT0Url/WPi9UUP1udXzUPJUYxVKED4zD8pd8MZOjBvoa
Mi2i00hUOoXxULfCWYk0VVG/J4gtFvfqekE1LkT6gdF0q2y8RBFFD9uMgQl2/98Plg+gIOAZvLwu
d9n/IGdxntEEwNgoBd1NCK624j1VmKN6Pe/rMAkuGnAPO1t+uFL/Ibm2ztHCf7NFz3LXv3Sf9ATG
4PIEpAFwODvvlxdqqgrGxBBOGmPOI3vhaaRTfjYuqOuKO10Ilqpmt1sw5Xt6jQpSjSBsXe3SAU/4
0/zagjqRx4Q9pv373rqxXCJ8NOHYmP09jARPASmYwx/VxUwOvC0rbRkkF0Xo7LhTyAW2+c5rnvuQ
yzvnlMe1RG4dFUKH0dqFR1cUh/S8DNYpyn/HlWdpjSHCsIIWRi2BL4s7rYFcZ7OQ4jzSSUERyRwa
2kguJWRp3EZuYYdgeDj1RCLefvvaCOfncftVBZtbWRXTP+hM8klQSM6AmJ6yeAnUqIsCi7OVJtQG
o/OyEFjcFffz6vGqcmqTboXoqnl7wgdCgmp8TIBSmVeJ7G35Kdo3hTQdIhusLVJqLE6q4IxJDzbQ
ghKQI7HY41s6lOnwIxS33QYbFFTxqJGJWdKmXF9b/ltDwFUXgWi/5zI/MlgtlwfdAbY8xmFQRp5u
CVuq5A5p1eQXBMIedDH6LOkNUSvWmxRixQ5sjLExmu7/WLoDnXnDB4u4a4TNgzAbPj1mN76eOjNf
og4CfOsXvU65KXsNU7QFSPhD6/T6QgvkIB8FamMKAKri9oocpjRut5j5WxmecZbiw2zwy10TGXER
Xz2aDqjObfjLczd+n0moz/3U2URc+Adk20pJJrpwn48AlnRRdncYuXuWk98VjawJsfa/9yGpD6VB
qKdhg5rrx8FMRcoC0hU2TAXnuRoSrFDeF+ESPhNsmjErycoPT6+1EHkt1MqU+x6B+9CGBl/JUfxz
q48d4i1WJ2h7baO1b85ggnEQ0SThWziEG2RMFB66c6cgCxGFZVZK/4b85RhKn5ddUij3ao8DC6oh
9s5W8wOLNjQ2M9WCBh0vGfgEm4k0D2aMhKRJlUO5sPBzoau789rKiqGvWTKsz8qsrpgmdNbpP8JE
BYnXAQBEgqCraueA+YRA5WRVM9lKa1i0jNa9fLzSjrKkU5PIGMFTPMUCaDpIe2+5TGVZO9eCk407
erlPXmKg3ou4yRig0zFLvjGsFbCuSFmrkje3pHcXtIEOwrxvwJv67QKHaz3NdXow5a+LXjQceKwa
PiLq9rGhMpPRPNsl+JNmgDSH7mrHcar2GiwIgfwVjNBOhSlu+sf626dQ8tEOt66CQt15FQ1tqyzB
Qdd8pdim+ksdh1AjDBP6N6/NaGc5bxHaa2ExK8iupAOBfKQYGKMUWoz1SaeWGxOh7WVT+hEPGBs3
4qVHiFVuVC2c/9+Br5AmSeloZYbPyODue80cAukJ0gM2rNHwRFKZPD7U8qtc5Q+dmTf+OCF3EX92
jqigGczSjDnUuR4a39kz9f+ldYvJUVOumUvs8uuhh+FM6zGrW+onymgtoQ1SaAgWqwNtn1X++lg/
LN8RK2JJ+OKTUGq+5EbEyq/F+nuXq35gIWZQp0KwlF0q5Rbvz4sQM9Fi+8FULv11oQ4GZP9fdARE
HAgFId5eV2P3A4Zn0LkxJ9nJbKsWjqHggLwL7eV7d7Ymqe+j1s29WgLi6xvk6xNxKHUG1UA/uKKr
az2B1tsVUy/RS9UbLmqvFLDCDk5SKEoMmpcTeDnHIuCdgS1ndfFH9eZbEa+sXP/coHVOqQHz/dwa
rUe/QQP6x642mZ22PkwGlXcGIzRcfYgta6dM0xMC441bTZDd0lanLKtrPWYfLuJEuiNpBfqGpf/m
2tFraC01xBNsDW+OybZqCqmzMD3jrapDaKhMNTvHvk9yff1BqXHNwv3JgOzfnseDdeHR0GHo5fr7
oY4PDFQvd/N9Svh49yK61mRLu381njpGnvoRqpEcYgE93KuAwSTHIeN2IxVkzKIQZbtCzXi8DrEu
orW+CqWYd9cckT+gVziE1EubbL9lAkw99Io5+iVn0w2ZFZ9hOCBQVHpPbqk+bx4Bf3j9jc9rYvXh
Zl/Uh3nh/ffWQir9JhRTvk9IUxJhDGnZ1splYqvQwVWiwt03TQXQ010DrFZrV3JYxTTn2pHmCRO6
rbSWGxLO16AhoWQ3n8Ye3wNpUBwE95Lc+SwFonxASHoBOCcJaRoX95qK+8elwB/cKJc/Gv0uA0Bh
kVbCGcVI3CtgQZFA4nOyvCp/dItsQtRPUXkokaLK5fbdtU42S4jk7quMpc13vZLmbLpduXUcYqWd
RfXds9M50LEcYZWC6/IQ5EXqy5uQJU03de/lZM9vvyNSHTORscXjJdM0SZny83apK+qZdfGeWRC0
ulRcmiAkHT7+SQMFsQJue76RH7iffihx3bEt6KDQ+IQJuvXZGrA57HXdSyzQW+kl5X+HUWFyAQ9f
Y3OUwJkRbcgjUj3uMQq8ufbMrJmSQoNkmeDjPLvshKetSNNqte4D1gEy1uSY4Vww+hxgNF3XsA07
mFvsL7QkgxRxs3f79/D8f9XmfDXDL4zjMUksT8tadYOYOXoH4vHjmLLml1YShngWnINfGvwMx8ro
oxz7tgxcPB1Pt1yMOeaFAfEm76194sT0bWzbHEaz9v3qM7kRQ+E3vAfW3U5889+I9+fGvqKl7pC1
tv0JciWBQc/4yrGOAsqwhNbU/fBo6Puky5ZzTVxckJLCVNRQp6O5INtqbfVQcAxuBsqXGdK6Nz6V
XHn4Wn5sZUG8PTD6l9CbjdlBX4KpS9NwSM+8NdoW+GB+FRWndQwKKWXbX7jmGSVQcyoWvYXEEAQf
2k2Uz5jqTvWgtfCL6kgJlSL4NeOnAvrutTK2O2D/NLObHtx4VZgLiI5xEEV9CuxfExTAQd1mFozl
7Q9RzzHAOAPed/2EVcMb7eOB4blDOOAyF45BnBdJ72tUx5tzrmbnNs8DKWoOoavZikk7F80K+b7i
G5xKslsBG/8aJP+P4cEsSiLsSQsptl0HLJxmGDwP3s9eYejNtqHn5GPptpIzSx8DRdQUeM2fMxO9
O+GBvEi+Z6hc/X9pX+CuQ10kqktofprckMo+gPhII4CdWgGsEOCI5Os/9vHeJL8FHSPzpAmf8MEH
kd/5cUWApMQcyfHqfoZL4H9lyQsZh9E65N+VwHjy/ZcVAvT3IHpVEoRxACH7OJkbPdZ3Xd9Fwqkx
bt0UEyeE88tsBK0DaTZTmlSePezGRa1VqaufUgivEObuvzE5xRQCRftAYSukdXFgHLcnlEPpXWhE
3D6lx/MJ+KcJQjwHeDdouXHQ1l3UOgeEqh9hE5QyD0TM0Z5gCTNxsazosUgqFJTmE+NccksTau5d
D523GtjwCJ8vkHmfrEdH2nqa0XAm7Fdeid5ffmxFgUaFGiM4DDGoJTpIxrwglTk+AoKmN39/uToE
BdoMAEPIoK4zqQYnkcqygi6+DHD+ycp5X1A6sFUGvH0AV1hWngacP/eeZOQZ8dVUB2aec4xhQsno
Qz52uQH+bUESp+KSixeUyLxYd+Go2RiNnniK2966aVFzblqHKrrVTC7IWYnyVoByqCZ+VCeSQZYu
0XLqrLI/MsAK6MekZwLejdjk5/Pz8bH31lCtFU3fFO5TtUvKETlfNHAtjF5ZMLvilkx/4/Fwvu6i
yWl2Sm95a7eSR2tRnsL2hYj3T1ErqvKteBQmwWwg3PQFHlq+fCc8QOh110J1JTpMUKWE7jfbCGC7
4Idv/2jvy4+DjkWiRfWTvMaX7JgJ+6HCXzldydx39IxY6immlgfUYRGmcMcP0JSeABm2saBWB8ua
dCmUogmx/Xuj2CD+kUB2IYpWolP/E7Wldxed8bPZ4iAzKcVUzTjHdTUFQuxof17WovsJ6K+PFPwv
ovFGYh5wgF8LSZvO3RFsROiOz51KPsK8Kz2Cqw5Yc+sjUGpjig2cv7xGRhYzQKBnHzrOxBB3VWRg
s3AD+ceciMiRhxl7ELuMvaJ9JDcSyRnqyOpEkegLkDkDkE76uTRJyLvwgN99hhx6QBzUXmPUO7jA
qRYzRcIaPTxe6FhG6p72iwYL+4mYHOJMF0+bnQNK0OMZrwo8JHnOJJaEtUNJ+8nSGXc+F9ETOnEc
py5GM7R68ijs8VoULgJAbmsyGAovmsM7NuaX3WJkbeQfeXabgfEQMgI64DyK8HpJFCFJgJExYvy+
X4JQYN9+JhEfVvU0NtHeSoMxNt+7GWn5D6Zo6mNntWnsjAlYXwJrHlVZzei2P78dmTROpfYs1XI6
Y+D4dscGN2ytsEEENxhzojw41jIerDdclqaXHTtUK9HDtGGJSreaMkwnGDUozeVTS2PBNCyqn7IT
0J5ES/GsawgXIXLfF9XHcds59da2IPrFSv3IuA0vkGvAEEhJN7ffqM7NNqfRw7szpYuA/idsoB93
uDLGjz9jttNFtvr1IWhP9vhqFV0zpJGQO6dDxlCUYM/5cEFDmm24F8ArZO0433TieCEvnf/aZpKa
kMhP9O9YDsKNcbiwDEgPSIK0XxrXmkQw/CzInW+azAHyAHZTBIp4dpYJnPOWiLj5jd+eYKnt9QQi
M+MkjJqyc1gQMn2oeVyzUK72LGePhtGgV6PGYRbe8DxuvtoWI2waskq2Vfk8O01GFHk3E6OlE2Za
cWiAALUXqdAt08tccfzMPmnJkj116V+rlmIlwmm3D8ibifPJ2JzIVTcUP8/zLrFYy2BaA1NA7NoA
2DAQkDu4wrmWccKHFqdO3Lny/b2LKAFXhve5vtwa1ANupxTnE4r9V5x9Tec9T9OXBS6sKNhbvKAy
tASs198pjYqUhZrFxsR4NVVScVU9w63udjPAWR2inMJ7Filh9T9I2jrGeC1rKKGyI4d7WCPFMHHu
MC7IvIfe6Rnabx0kuPIffAICyUY8dYScBwSXLW8WzH0Krz8T1Bp6Ajvw8/I7R561uRejiKKqtALa
bzwh03nwg78ew6GkS6wKxV4zfqMWBCb8gowEwkb2pfwbsmnw+C3ipp9tCTxtv52ZNHXQc29Wr9Z4
yfXeyB6QWwLE8FiWcQgKJKqhV7Qw+ai4m99sSr/2jil3vPEIBtFltpeXcR1hgqRi+/SbXIYpeXsD
hjEE5WPwhsq7801RtIdxAdhoEEz4G317LrwbrVIxq1lv8Hsm08ipZIeFb1GtpTAx6M5FA2pFC5nz
j+Tuig9AKayPQodngjJLbLxMjxvB1be1e1iVA50Dn4SChN9BHu3bF8/wj65GLlyCalCMgwuk8D0I
q4yGCPeidfh6C8IKFFhdy31NsFUqEYoH2AieoBQc5EBF3gx4b4uz0VV+taJ+DuEecrlx0+0ACIgv
SJs0gBvUbzdP2LRrJnIdmhAwklZ8BtWsZkd3x46xANC5fC5GuJ+Pi/THYmz2iSEF8USa3L8tg94e
d2n9AA5/pwXrpqxNf+5FYD6eeSv1jbftQ95/vK+ahL5wW9NOjsmVnpgaMFVMuPiaWhIQIDpcwJ1i
pQyGaZZAfSon+cjuHDPmdFrQueHCYTziiYxHvpADmZ9UJOF+zpCtwXhs1/SZbdvo4vs5ZzpWpTBe
KtJ0Px9Jv2hhHnh7iBQuEYvADUqTvyYsX9GLUHAkz4Gjup3jcFwj+af9zUf9MegPqklZrw6M911P
7iBKhTRk0U68XYfqvWLjyHxDrcDGdIPieIMkqHl3fo5t6xHMY5rXfKdwA4CN2nsJHwJSZvMV/V3a
D7tXc8v2Yj1EwvFaVDpAqRFCTCw+IGy3zyq8WqAhenUcpaCOo5BGULJkEiZzkOx5Zr2Jim7F6Ioi
hfkzJOdTwLh4EtxMRU3vokLB04t9R+N8/MayVHZqDgXEB35Az9/wJXD1rQONMd4tzI1FSEQBBMEf
gu1p9lQElkHQaJJd1tGMCn+sedy6HXJOaRm5B6kl0PDuHiJx0XcneY9glSeFkU7auJ4gBZyI7+N2
6PNIcenTbGMPyzj/NNROUfa4osXs2H/8NuatpN1TL6JgnRMkfIjX3ZjfKlPsAPm/qWwjvD5Y2kht
N3nA7QMV5aNjvN0iyk5P2c0IgW8fuc7KZCWBEcwofz38U+7kVZlqTeW0v7TYwW50n6Sj12zHjKWP
s4Dk/XS5EPYYD6C15OPejvuVqIQ9ChnvbukheFdxv1kv9YVpZohEA/nherRQthr26ZBfkowX7bmB
5Qdut8+XTWmqOyLqNRIQNI5WrFH8qCnflg6OtTnSInLqi5oPSSGJ7WxTvApAWMacQ8La3lIJJ5MM
GyDjMhh71GWemRYBr2wppCi271TpFwvI/bF/e0/WXMoDhW+WquuQXjyZthIlRB//M9ukEkQYQHkH
aKbltlII7mAU8kUYARCrsBSKUyo4+y1Q3kM9fuCze6u+jtmN5IDqhqcpOMVdRPSOARFcZH1wXEa2
QEl//zFFzcTdO3GoFnYs0EBwGxREqoncyhCCjvtub6m4qFIuHo4ESAderLuA3drMSuYeSIOa9t6n
M+bha2Pk/LAgyZZ2saCv1vZi4s4p+JuRdDdfKIzdjI1o1obqd3gFojzjep7138Gb9n7zjQ0dJFwb
MT/HUxqHkkRIgkEEdrJnzdggtqIMuHc7l1PSBiVjJCQ7FKfe6UOreh75rUb0soB41IK2ObV7RR0G
SDPrgX+20aS20faT1kAO0N/xPwUqY5UF8l/BSyRShBE54Shwag+j3UYTsISjK5xO+rtgXqt4Al51
kwOTUbH9VE/xPIoHCn3GNO9MdByjlxVKmyXIhH9bJ+BcTU4M1dTp2dDiQAi+hrIc1xW4P25LIXbg
XuvOmcryzQK+YRdI/hcOOEti5ba6UEqo4U1+Br/W7tnyZuOh4TBHNr4Nu2oIJFKiELHXPy5AIsXV
9kelF1IGCRX/cLAyptaOsD08+v6Wim3NgUbLV12s0MABdSwrZC8SSWe1ztY2i9pI9eYGASXkaX7x
F4ZJBWJCun68UVErJ/olR7WHZNQ3WUytle/3FSoOA2XRnYLTeyetaWpq+Q8trN4TXfB+6HxiRBUR
KAeUSZf3QLMfCHYCHMVFHUba69UxoJhIMe9QatrVvGyKgW41xnETC04QjoHXvs28pvCp8YTyC5rE
55nQ+TDPIAoZ0t/7wjiJpT+ptk0X9QUJORDUw3Rfp/bpchcy0TTaPMw0xvTeJT+dT30sJYK2Da3d
ekBtgElH2dbn1jL7ADrYHLXICVoa2HQ6tg3PQYAhshao7kXk7xDZcd5N94mEvEcXmmd9yUSidwS6
5NZRpUdBrWZ+rb564qrxy0+KTtlcZ00yQoH6g0u9kanPfC7yxH0L32Ca/wCL9xpbG0C5cK7t1SqQ
SljVoN8ZU8wi+Mmfoy6A9/ZutnRDaMHWe7beFeuxPLkZmxmyAFztq2SQpnXWjlegedg/CPW30sUA
OsSmPJQebqx1qu3k9bUGAUrGBkJ8B33Qf5V+ymg+CFXirBs2/hE+rFk+F5kTGyrZFpsm0yGF3HCK
97wSibVJvq9jzNz/8J3gUxx1FNKYRz+RqQYAPrF3AKmvFy/zuDpii+k9LNlRhvg8VCGb8aCMYkhf
5XyNgGpTTfyW1v5XzdYbHkcY8FjaUGlPa/ODgUuf/dmMbauY9F1quKuCB0UaHKE0bheN4K7QjRe2
ZuXIRxvHnAnCe4fZmE1nhsPle31zMYF5q3BPgjtX4D/Kmi2iujoHMpP6NqaGGxIAAVV2vWAADwyq
Vgai4JkBTYu2cGsmCkAlCatF1TMLQEh2MT3Qanemlom5ivuYDk/s82jtHqzqwTeWTmXAiCMyW3mz
eCMQyOHT/YxQFschaOPe6R6w2rTO2UcExuT0NS5FGBpDg9JJfTgke0ff3wEt5tFpnXOG2fhkXHrx
YDMDXkR5MbaEnENO+vlqDUs7bxxSPiLU4kAUBaZD4prcFtUQz4AHmHdfjCMEbDftRmZNo4ygWPyd
qienvXPx62YOWxLvqZg2YV5Z3s5SsRFXRZu6qGX3HQHaV5zxwwxiFqwZ34Mx4hkDD2/JpCC1xRiX
OVoApVGgwtNuMpQWH84GWtC37ulRhhibmqx1gmRroX1v5RJkoKbXTajaVuzjBOyjkWu4NA2MJzQs
yaWlezUtu8a6+OV9JHFi6bw8LEaIrC6coiSmo6QjWPc3zvXfPOthZC3ZUdLv3RYQpcKfFEyOHNfJ
JB2/ZVaXS30Tpt8I8ZbIaWqpK6lzgs4G9cMbj1JQjuvInt0FlskU48t1Cu4PHg54rT1D2DVhn9rL
qWO2LNVTa5Z2bPqVlFqIPpf/wcCM6TeoDYoBG40nrmUwUHzG6VjrxskK+acejnTfr+A1dxslMIh/
ml4FmTFEVfiC/volS5gE6fm4dHzzIqK9vOcn8r5hBO6J4D6wVqOo4i7tLV4qizVKDYz5mpbHhSVJ
L5pwkP0L3ECVqhgOkhPpYDHdZ3m36kScCwYWtaf7um4/dlNKv/JM6QxUxLWkwpdTV0FAkhVW0I6r
U1baIPxAvdjSxGN8S2d2EosJqomgUJPfnGpXi6kJXSagwCNIn7FXVsYahQWnxCTCB1ZOCEabBtKO
Ro4VIu9DEt3UOrVeNgbfcpMFzr54Y7uUeEFM1Qk8EX8XXm21+Q0Exg3O7D71dJ+FMlX5m+g+akBk
yiyywWOhGibaB0kGzXAwIymLuFPpg2ihzgmtyPj/M4Z/MMVNQjXtPY68/j+kPmQB8qnWlFF624sl
rkxSz2QedslZI+3kkqW6O4eXZj1cbjHLCmCrmxMGnVXk+v2bwE3PPv8Ga4aUOA4cTVDDoBFGketH
uXpqas3XlRrCdFY26Iv6k9Hqh7yRMS9mjbBBco+Dk3/b3vsIEHOyAgKskIYLSlDBAV9RWPZYz9Y2
EkHj+kXhrdfTYFm6i/WRebaRQNAZ+VZOLS+UNI7SXv2Y1Ht9lBej2oFyooTFWBW2X2rm9xiJ9wKg
fnbxVtAWNgLn6ebgLmvDl/iuaLUC7GA5Q8rfV7TErY0593r2AEWT3fskjQDmi1CbK1XzJf5JzeuV
RoRKwqwEUs8ZwhEjXUOk7t5hM5dJ7eXOjM7PPk/k441tEiLEpavse64PCeyQkaal3eE2CvhZZcf8
RqnGwYo7CKgKttZJ6wCUQ/GgCSVFLjfjTUtIj4py//66+Hux/0/jcLh4olE4bvT1YKgW2Nt0B9fX
H4ssvYXXcdu3a+KwvQSNMlMnPWsS40RKMOGtqjd0UacLrNH/+lBPNALjxGD4DvseUdJ7JSKdzZ5u
fkW1SbK81sNoXRNNeSiXzWDthMeW5nOUtNNI1qkzHuF3G+fGQ6gHMbzz9lIuCU+ouHzBJVkGNEq7
VPXyC4LOm5OxtxtfLYhYqSwKFMJwdnMUBD0WHXXq3Qz9J2DdDxzGlAvdo0mK3TIEQzqW5XIFz71m
b74o9pmDsd3PBrMLLOb3WHGVag/JpSwFVlzFfbebZ0ytyDRUo+ez0JKlqyQwbEZDAEASzLS9f+Ul
GXQDrHFKX/i3ib5HozNmj7MYOiXNELDEZH5yKCvXwnVyAxfbkcA9oPi35L4shznP511Q0B3IOx4k
8Ch6wdF1ZdEdwum4+GSjfIhwpmjvWetNDfVRGBCAeTWjd6xZUeWD0lr54J7OTD1oeQrWCln099Em
TNbYMG5/b9UUwvthNoHgAbROJ83SnK3fcQsZLlK/K7tLGcu4D4U+4U8kNDXAbUQINpvnh9A2DmB5
nTsNAHyWUt7T3aeXJ1oAK/l4NtBbmHIRZJJYM1jgf6ZAgvzmH/QlkCTEik2B1x69N/+9uxsFD/D0
9nU8BPYifM3d8OaNdQ3Q/gEbC53VLTcJFfyiAWe7tSZvRpT1Jd40JBu4X9cvYbCVataBXYFV1QDQ
0w99DeHaLx8ZV5gOUjgxrXsYAtrLQt7I4AJpVknecK8EJ4TU0TYNrkaJFXNScaC1SRvpNkEQa1Oy
hJVvPG0b9KVUZYrZ2HIMODEge4Ly+Lq/i5T0izX8I/OZe+mjdfD3ROHvVxgln0RGDWRiwOaoGyED
ZY3PoB5gpw730YrrL4jX7V+JzSNXmnnI8A6TJWkwbefwTbR7DSa4oDP8i2mnzQqiDrQ/tw/Zt6Un
bN0nqQJJV9SuVd4cbXsjF8KZb2v224oZW7rxuWPjbDWkJuZo9ZCvlqAGGhScXEfNmXl66N0R3yOV
tvTltVs8jRkX8ncfSBMtNOJVRHzvrIEdEvJP/s+NNZhI3t95pqROuxh639NOmHaxjllyrMwUrJZw
mt2ULgo1OfoIjSVIBiUscEGy0oKiqWxGmG6kNVogJcex9eY0Rv0HiC8djUWkwVciuOQw0vuTzq+u
WA+9aW2P7Zzfxf7XpN8EXCpBOj7XosVEzIAPe7vZYyhZMapn95hGBptX5gI8Or3B5jt0G0rgvTpv
V7Yvo/uR0eLGJsDqf+Y+AQ6uFmvV/wOmpzMdq+iq+QTPH4iKhPbwN3g0ffls6j8cT9vaAASpscN6
OPsPAxPgNPJD3SaXz8KSC3mgD3QvDELhSxTF1Dt80jnCMN63IaPTEPU9SMlhcBe2ttE27opm6c97
vC0fCHf2rDqvKx+xuxcqj3Z5gHGfbf762QRRX7fFBV4H0DsMc6ooaPkg9UyCNEVnGws88vmry/NE
LR/pSaCsrpANTjiUbFcGDCtBfHRw7L15JIDFG/ElXJJl2G8iJ9bBAFNQPx9QSsLk4Ve/v4SGSdlt
zmcNUiGbXGC5Ujj7DR2KLRwSxfG+2D2d0s1whiOOPdVNoFArbPZd84yk/GwAY3HJDPVkcnxtoeFh
mF+kuSUUH2YShc8hdLF1ZChLaSkwAheTBEJwT7av5FFSffG9TFJX/BZTDERBmfqlHg3/JBs1NnOj
tcinBn9mtrcTOU2+I4FyGgc8XHPSFNpEt89JTLtNtlDWb6Q7twxswuy2e/Ghg7J5Yh+mvnm94y2A
ugYDWybBtnBrdqPL59rs3C/mQ0wt68NI8i//3AAh8JyT3/CicZ7FyFxFO1+xgT6A6GghGn005Ete
8JQqCAnUSyAaQNsk55bIp30FDsNl0r69u5K2/BmC/sYNAeOyMvqW9YQ+cRsTwuiPtavk4SAaXWKm
XGBx1lhXiGJhLpeE3eltDV2XFbwi8lFR30cMCCy2IPcv7pJICXGYFdRq0BFdZF/V8lexAfaFiV5t
ugVxZ3TJQHLDUCO9PEkGVEoENCipK1I5ZIEBXQJT6iNDiP8apOOYIUNTCmtkPZQLAx7KtQOVsjv/
Uhrey0za/fRNFtXO1pQOGliJUrRFG3vPcZZYqf+FNb/sEvZUMu/0/9C4QTX1uHBcv74zfzFXO0Vf
xLY+fpAvpB2sfOPtqSVaZZ3dDgQ0CSqFD89ev309fMMSWUxXmw2hFWm36jpLNpZfGgat2XVcq7+k
u07k0d/fye2Y7bxPGsJ1H3FZbc+z7H4xW0Gcioc+R4UcCNzFgPoyvFWk7Q01i3pHbgO3dAev1PyF
dtbNDItMp2Py76DteIMy24ZKl6jSP+2zTtf+4EqT5Ggif7BmEz4C3wvcLXzahBZ6n/FR26xmur4C
40mKa6QD8PONlHbLolBo6DBScX6UI45jU+LDB5qyKx+TUMtEuBe9kqbneznGlnb6o38e0l0dV4tf
uZZ10wBcKoBfq/7ZoOHB3vXoMxIJoryw1ZE5+ntRfF9FUKs0Z4Bw2ulLiBw4v7F+cZLz3yBI9bJn
ndKC5uTdbepJaTeOi5yVHKvgwgqSkNgtx9vC8v+ZLI4ut1vUTr1c+DDInh1+thCZaeevUnwPssNo
rx4hrMekzsO8nlsNEtMKj0kIKv07XBBbacBcQFvHD++fLs0/F/IbS3rUSxVfmEFaPdXQLFJsb/y9
P5SEDJM0FB8EVQnFqCYy7rEopnq+EoKS+gmM5EFs2w7+TAufr6ww9fH6Ng4f/NjboHuTcxIT/ptg
ARFoy/AHTsO2HkSTzQSZC2aPixDQsayR1DSQDnv6+HUVV/B6LJsv1gqa9y/mg6nq65vlDeu1SP7b
Mw4x5LJWrq5S3LgVQfOtJVGZXpJPa/5Aa+NU9Nh2Kf5sIRbWe6A2QB9IqvME1w5Ax5EAeRfMX8Yo
3tO9ED4ZxWzrHMJ2TdGpOYls7/xI8lwPJtr2cq9xgpglykQ6i9xDulX+lklpeYapPHIqXJJmExpA
urVLCVGknJPHvh6lCBET/iV7gQ82UyUHfJa+N6guBT46Ghgn+F9AZBNBi32F4HBdYOZr+0Uoci1h
SByTvatyO6+/UWNAzqTe5lSNBCmDxr6iC16+++Xg9NeTnP8zAr9Tnpe43ILogZxpRpBRsMSSbNof
3uoYWa7KTG6h3yAG3Zkv2Sva95vs4aUn82vNpcNvNjzjzt/+9RWmHVrbOSuf283BSYRg57TlUXVl
JiV72UvT8MPNOgm3WhGf733VaSefSxWF7UOPrV//YZek+GvXwcHD2qO5TnUjwFFPiG014/7fT2Ms
aIo6D2nlRfat+vMOppjb+iAKUfZbIw7rraOLtBS1E9p5bYY++oyXv3L9qYcplnfbuWB1ur58xRbS
rmLPHbAgMzK2WkugruWEmmnU2LyONHdrQPUSnitVXb7iTZHRmZpLktyLUt4pFZvPNd+vg6gAuG7e
TaxkfJOHKUDvG6aQfsltM1Tr+AucWrkeDLPMpcTjHUmzy6YLEm3T23l4Hhf+TcLSHcUva1+mLU69
U3af4gPN8CBz5jBm3x7BSiTGI3dVJhlRyES6GoedpXogacAh2XBjmF6cTEckRto48fBLSETqRdr7
EWgPewVDJZPiCJ9kUergu8EQdXlpJfhRrOyWWyEeS2UjZO8VhUJ2Qa4hZjDUdXPeymJU6kGGdLcd
HttvshCqRUAu9uxDoiOl9xNvwHk+7FBH7nXDinRgjUB8IJP3PPwJdHmjLSimhPpnW9HPWIadDNPK
gcLLG29ruLrEG6JAd2+IlhIHbvwyldAIPtKVV13LiLdA/ODw7c6yOBYhiKkME6P8WVG0TFLufn2k
tYEz5YgVgtSF91/VgY9HiBytgVQG0qqsD04sX2iYa2HrxhvmoGQGvmq4qz/iaAtsQSsVJkmIj1UW
z6QN0rOosnvxGMwdiDNRcgLhCnFyjVLASL5zHp2cVvucM0r+o4u+lLw5O6EOpXKnTpQV6gUfpTLW
aSRmCWI+UcjdvPQvkxlAnYuvXK1BM078MvXBqyWhdc99j2Y3oEl3+J8A0I0VApuZlc7frUs3CXSr
1c/adhS/ToZKVM4asQ96wl83UXa082n7DeQ+uG/5PvLlrJjeY4+aDhJqrE5yVxWnbpZUxJxtEHtA
KrY5Pc0+M1ay91L9jj456iNFGN/KkAlqiOLnFL0aKmt2P03CE6mDfJev0WbyYlmvJbtlelDAvSOj
zToe2jBm+7k84v3kSnbsZp/DCjcc0c4M6ZlClsR0EpQDwblMssaabLcrnXZainHKoDEIEKeC1oTJ
xS3IrshLZvKALQBf+agXCIudm/PEN/hCnQoL1pPI1IPUx/D7shgqA5PYgS1YkuMezMKqBhl0op5X
uW6W7BZeQSSm9lotT297VlChM5rIa1WpRyOcdc1Xnit9j/EMc+oAq3v17e8ZPXWuB6fFU+DeEMAD
TrO4OC6pIoJsWyaohFcX+ETwpPk2LNh9iKohYAzD3/yQtTLdBRv9ELBm53zZAn/PPuep1QewNRsU
uI1J+Ft/NSzOHRrywSpE6evoiwzxb2WXXVyutXqj1rtXLmZ1O88BswtIkYhLhOuYWCI4PrG2r/ip
zvoZ0MJUw9HoQjouzkjDezaK+SnZt5URjzuFHXI+0UwEGloAY1JsVTtROLDWCtsNa6yKXz6kAm6E
34qJWszyjh3DkczLioYKn+ZeIR89b/oTgBdfLncMfktQHDQBtgm5kRTuqxkwiQUrViUbQlU0CiFw
ompY1QEoAMioFlRkxGdhPBLa7PJzTnQkgmwQ20h5nxTEdXg+MWrHB5idD+Fux66dlwcOuxKMH6tr
mw6OkudSjrILjlBC4BTegTyvecP0VHmTGk0svHpyocXsrWk2g0ljjcMcXvL2oTtpZFvzeMw5PlkJ
YkKebSfC+duuVXEzBugiH0b61aaOdiSbWUKOUJu4m8qIddvmReKQRyK6pcSX9gw/wOD2/NlEJPJl
6XahsxmFKAbi9ywzIEZl2ntRY4EQag5Ekyy6eVVvy4czUnwC7HjubZ0xab8yaQW3/ViO0GMKzBlm
8JwxzQOlxxRpgLtj21wLWgN0V/aeDt/roQXMRuoOByK1fTVAk1xv1gsaR9gjM34W4eo8Ixz/uVIq
17MwcLnco2O3fzfq5btTvIZiFbwOF2IX70hyzt6ja2Yu4LZwdw9eyBSfv8ZLQabyiFMwXTTr+rsL
khgDZC+swv9HZ/M1DGcZpoavYNHmLbpXz+5lRfFm9nnNMcYSJHz/5/ovWJxeADRTIoJ6JyUrUaqc
kEn7DKuEpJPhmC0vi/UPKlP2g9DwHNvvN8H0Dk9OBAeZdKiuMUszC81ZitJzQytUQAOM6gj33bRe
j/r+9MixiS+gDahlAVp7rvAVR42SUaizmnpEdO0tYCKhFUj7Y5MyklmXFx/kYWVXDiMCXVkY/Z9c
fHIc7rrutr1l4Ahuc5epxx2nQHd7X1oaq2PSUcA1QPJZ//VHecsUmSLXcsjfzP04k0WCv1SnDtHA
S+RIbdFX85m0cS2aPipnFhoBJJ6SAUWJnFYTbyzK+2DcJQHU2ceVkXEkSuwI+JcyQuQlINI3Z5mw
G4qPIVyH9cl9o4qAN1ujCaFVUJi9cFQ4N/y4RRG00+yZOyKd+TpKYDgmSkxOEqFCwEZykjog2CUZ
PosVBiXOjR3kUzsgRLGyPrTs+ILK4yAHWUjGcz9kr/hmJ4umM4FWHfrDH4cCaoXGi61m0kh2565h
QdR623t5soUlsBUmbhg8uPeeE2ainWJw7Nv1XAz4MPPcGT3BpJ2gyDbCtMysCbDBCNJ1J8ZE6mcX
0bdNFHQ+bXbXFZw0SJSMGz3lw96mepbnCY1iyxvlzdP0P3+yEVVvScJSmOdR3cuRwvojyjrOkNTJ
y1x6suS4c8TKpsjS8pgp+vekPW4t6DSBhgnOs05AE6vdc7iw4QY9a09Uyy8JBeBqUEkZlf/NRqoB
0JFtYTw4Zn7/SurHvTPGAuL2ztsB1aFJzj6APYpgDafIAbtiUbr9X9/TsTaWi0LuYDlZQgfq5xvU
lkzox6FdPc6wLfcnREn2Vw60saIN537iZiQ2h6BcWxuF/CPb/QHshmERjw54LdYcTRLREGOXSB/R
xqzwue7c026S8Ttl7DGpf93qUrfwL76x6C9p65VG9DMNxCUjxhaLxRMH9OGvPGLmibmZgLop1EZX
16xCO7shUzukMpGK17/aM8TaOjMdYG7MRYEq88W0kwEI88NlZT7JaSi5snvayFT+Vr0VThYSBhdM
zTak8A8KB9OsQt5gf+sI0Rc3h10NIRKm1wzA4TaqaF3DqYeijZG9KVjuWlG8ZeP2bWJbtTqKRvrN
bzWACyJUB2W9PxDTFrY8c4CL+JAKkAze2g+kiCt1+mK+cBaSqQAaDai1qXYf4TM/n9HNwiPY7Fta
RGUMGqQdQOSjbtICbrV3kRb1HaG/yg8cg7E4ORKDYICfxFtbj4yJVZWvCZ6BEV+hZ+HXhmjVWjUf
9RK0Hc76bKBSdynTCXL0aok4pMbHBwQxNWBYyzoCAHwI6nmRXwwj5d9CbE7/NHwtlpByxhq/pXIC
LbupDAZWtwfI7nq3/h54MeW8y+McmPGQpWY/8NLQqBgnXHEBl8W9LjtXv+ub62bAG30OpgnfgNL1
0fb9JBU+ouISD0Q49JhWmX3A3pLwPRFn9LZtu+sHW902KVB0of3hMWgPXHqFpOxaVzLdIBUDEL1B
h0/YVPHDQdB+ZqA6tYyKp8f4Tb6nTDZvfwC2X4Ua6NxzjsL/fVMiPkykBfnT5wh/+qksrVTTCjda
Aprc4YaIYgZL3DOqGgH/As/Fl8VkPQbhi3qhkRWp2Q8CbWif0QXREpYZVr6r3k+Celrfs1BMGjkg
O1l2uBUhsqjbLxei7yQzUSHyPHIVtmmSyelVduebUok9z7toRa3ZaV5MKmfUSlKDQBGrfMAM5Hf8
E/4JS8Hl0GqWo6rIs5FB3C9n1Ekl/EOnz3al9Otm7UutQEhRdgYqp5UFV6oFRYs4uuYLeLnvloUd
bpHX9EXk/WUhLuA36kU76K2pSyOp8ZyL8hhIiypixKYXzAcn8hSQu4J5Dq2Rbg3ZsNXL3mYno1HS
cvof2IdiFsDrE6RvY2W7XNm4wUW27CmwTRZS1NhNb8Q5LA+Ega5L6ArPqqSZJL/XfPJlzEZXdYyx
/TmOWau4X48DDbz6c1MmVFCk0A9FGKs96EFZ9CVglpC478YAZNXQmtpW1z0SJXjhDwzJZvdIvVmL
x7hnXxTgJcwgj4Nf5V4Wg6jBqHakHeK8sxiX6gT11OodODBmglZbm8k7L4gBvuGdvxNUQfK0xbev
6hno/Ws/PPKQdZhJ6jjqdSBRYrV27A4Gz3BX6v8m2I0TYl6gv4xigAJKDay6IXTaBdDvxIdy0cCb
4W3LXwz0ToOCO+vTiPsQqK8BnFwfw1z2yDahh1b1dK6rPUk+OUfWOdGZ67fjblGKj6Ku1NxH1wpl
6JHvkiWt9O2Z1MGOoK+O9N+/OFUrmL3C+tFX4FUbGG20/4fP8jpcZmKlBPt/+PGp/N9ApImG2RMc
AU9Ms0aroi3AC34XuZH3P/57PgxYQS972huqbLUfXXCuwLADmAAm3oTLJDFWPYoW8j40nh1E58cC
r1E+kq8MHoeoW6ywF1JOn0L5pStfahYOF6qCfsMwbTq7Wozab5jRRbl57Tg/CXcWJG+ZU/q7TgLp
zjIXmrjCiMixTCpci/M9ou23qDzrjnx0cqf63b/OYNqkMLi30WkRK+t0C3TZmlmqsTkMZsqv9vkW
F8L2VxbKUvePcmYuxoqUYqTj7+scnfRQjCJsajQqoxB/oqf51NprCtb5iz0aEi2AeXeFARvrYtzI
BSpv5/Nq25Ga9wRXBcrnSIVeRXHV9DTYmeUNDAeRUlmaPRhYrK5vmo2ZAEUA36v0iJiF6yEPI7wZ
P4kEtGLv10Pw+6W5H6Jyzse0ascxSkFTn53kmpKvE6gANqd3WK5re9l5CLi4PvyWnCSuYW6BFWNA
ehc1L8LcB0KXRmXWhPurYofy0PqTQSajq8TZccx5heTyI+Rh1yU6fwpT4v63TWFr1LjwEAn5aiBD
Eo0405LCOHXcaIACbw2JtbaZiHdcEDFaWESc8+a4/Sm0YQjRg941OCBmErtue1qosUbri6pS3UfW
3aA9y25ftxJmndNX2dEKtRkSxtXrqg4sMdSAQw+Z69mz/kOG+kO15hOtf/js68oBfwByL9jCV85H
f3ZEuL10WL5zAVdcKDK27FVK+OsrhqGh4pwintfkSy03q1gWcktG2ob2ZNGCEWmRU4gocQsLMI2C
kqySAWUXgJpCL/YpVoLbE966eSEo1TrbnV7wTk8cEtH9MpgM/wFceZMONNvWEKLBr33O1IEM7uYH
fQ3CmNMobmktGyJ09rrwLW4a8UJ1EyyS+fPowSfgMWPfBfPOaQW9nDn/Ct39rHxSWMsI1C5+g0j9
X0eIMXCidChvu74xc5adcIijZbhAt7/f2zhXbJk33wm9mM2xgPnSRVwjiebX/+t3Pb6MB00s/8ZS
5fVUMhcgnur3037exBOxLhYOtm0n4I+vuWyh3UY9j8P2hNO/MwecrVzXVjyszWGnL6Qc7aM54E/y
6Ib6r61rMkrLNuQj84z++AXiUM1RvSaQgHts0CtVeeIxA0u8Yh+5Hry2PLGRvlWSPUqBLgv+L8B3
bGD0jMXYarxoU+jg5aZkIyybffE1W7laPQKduHt8AzqRDdMhim9l7hY3O1a1DFc7NS3WjpK7EY0S
4jCWsAgsaOyVD6pSzfi+ImpTpNJMvMTpBBNF4c6AqT0Px/N1WOMBr4drJln4uOCZppq/LVmZ/OKp
oBmbY1cZuelvWp2304t9+2b7tNdYvwcfK8CQyevyuZjOavi/tfTeSzIC9wmhA0dk6YZoimtpX/4b
soivXrE4GbW99NR1eLSyIcMBrPlPo2RswBTDpSwBtZjM9kwefS+La3XrZ33bf3WCMpRUm0Rjvrm3
kimh1NiR2N/7iURQeooUNVub3Tf1QGB+LC3FBVTuWla4RPa25HNtzQvnZklXiR3HLP+m6LlS34aA
ZoBPLj3cXDbQYyFMA71EFIxGYMYcz3cXx/nBEt9+iYUOxokclDmD8hgRFpnpfYYVBUgqQjj66RLA
2Z37TK8BKEsN1lOdcrSv8ujpCinEWTlT9SLO52UwHwGKeme2fIzxaq1bCYV2mfP5781US4vBlZo5
6OklNNL+ioOY00OPXOFNOnznD4uq9UtwIr9klx9RqIqJPkFBf5wCI7BDr9Qw/A7ipEb4zEA3yZVe
GA52CHii8sHMsNAvTEa/7wlFU1GzdVtkgSg6FHlIhtdNd+V85kNf0WUrqdgr7BtMWjAdBiVD9k7I
QQIz+vgIfw5xO1QS6oQgahIDljPGzTl3Q3tObK7d+b8oc9umfZFzQbFFeHzd0+5JShnyEvIY9fZw
lyvgbiILf1HgszPCfkLzr9nkfskp6Dc0s50LY1CnFrY4c5VA+hl3IdEHByqJ91zs+rF9LC487Gvw
WIIMTtoipUdrVnFxOrxXrgqd4mA5tjX/hZBQiBZV5ySjHyiReUAH+XI0k9/sBPMymxL5Q2gXFP8m
Ixf13FtGFsUKWfQWkM+aJW5Al30KG0anbiTTaI1Iux08+Vqt50Ua5c498gn3W8zxgBhjnUHO0e6v
dF0H01FkQcAT+m4SgQNaBkPKYbkf7Ua4NvrSaawW9d5h6ck86dFgCMWSIfm94MmsrbfFWoBbDdk3
TKv7BQuNpCFUfU1zk79mSyIyygEUJVYE2Drobj9NLpvv5pB3Cs9losCz9iCLqHyiHMh4ghfxyI/4
CCzJbOJeWG9utMZl9e07/aiuns+/s3iWLRkN07ZPVNbTcDv/rvdWUPrOQwmqEV3CLV6sz55D/xCf
lALUgpXQXU7VRxfJ7PCF8dM/7muJ+eX4m+PHNDuK1/92lsXZHUoVie7XIzkwy5DWlm14NdU0E+F+
2ebA3tIkAtKfqKnFuRk1UAvNHO/1p6T8Z3ChDtJ44Vc5HHc+vXp5NyuIZMPUrY6XD1TEgfKHrCj5
TYp1YpXalXXlvmoJHm2LxCVGBUyTqEVkIy7PBu12+qaUo/6RwuCG9RbQMFMj5efRluQdFuP+bjMi
0ndiPEWmtzChGOyiW0/dLQiJi5WiQK+3ZTqOrPYAJ2qpaoCiGTGIw6XQUTLyhP1QTNoZYZ5jiua0
HD7pMkq1xTK5mSpOhE6SPvrhJeavmuIB636y+w7bnXT4XWvJzjxCkrw8EN39beHPfz1Zc4S9aQMr
5fP/5F2YRly25axg1P3nzs4BGwqoXXoMr8/lXicfbpS8RrNfYB0oKru3HwKL+Vu+c0fs2jD2pzRi
fTA/3axBACT2YcnByPpAoaDab7Db66BCbDxFBOJTeMTJyoxPWU3g1IF1IR7rzgXpxEYvMf8s4Q16
IfMq1KKdWxqpqwRRP+zYWzI8Wpu12iL9pYOskG4c35vOFsls12E8XlCA39lYa6nyyTRhZ+A4NsAj
aE9UkJa2J1KJaxSIyYgtwEEf0neFKtJmn/D1gQAp32lRbSxLHXIp4SV/2uKdpzN1HCkASZkQk886
acflYgbPw1q3R0IrPHZCi6o17oOurswpvAPhtGRtslq1G6PjOcOE/t7vrusGQrXEZszXYUeCepdN
ZMtKLWqQGcgGhAOrBA0xqcr5npUY3dYrrVh//BY9SCqdQ+lZaN9j2mnvGBIMPiXsP8NsoKaK8YB3
kPxs/xyVL8g2swLWrDAi3tSes9QNNMJg8YoTqUDBPyUlY5FMk/1CcOrJd9M67KyuewIjrUpaavQK
SGklh1zgRZgltbIonTd1wg/YkXlNl9LObcOy5rSJiu3tCTfWSiw6DXlHW/jj/NEImGuEX1xNfBtX
tfdyw2Tf/gm8jSeXX7j4pkI4woqXZ9qTSCjorG94KiFl8H3SbNmuEgRV8EFQCRUZuCMbthomoIxz
UQgMjt8kdc+NM+huuLu7a9JTttN0tG3OdHJf1jpSPno6nva53AlHJxpww70aAChYCHdYpkJFhqZn
pK9r4JzgnGGBMuqTOCGtkbT8Q8ykO5Z942Ff7bAGIn3RXrkG9htw2r9mseubxY6bG13dqIFdMzpM
33zHt4iVNiPD0hw9GqWsRuhafSSe3BuLhuC2sNYLo1eBKw+humX4P64GjG/JJYqAXxKDihUwdfzr
wzhhovcKcAafqWeyfV2LYaE8eWZOhWfT4bKK5y87MvJnksirK7sRiH2xY5KmT9lZJi/giSRc1B22
uLhzrBgtN2MHgCZBJYC01kjAOBYgBRquS43cT+DePkn1Youn0EcyibU97e19xfwe0bN4rpOq1AMV
7dMFoFKo4mi8njQyTHW1iw9PRw1ogTsiTh0np8XdjHEyShr3lJLGLn3HqFIaIKcJIeACvGB17oEP
gfQiq65SJ2QfOAaxrH9RkX70nPacT3APjSJcaQzoCY4ZCDG8g29cLlAUy1TsqWhftl/H0GW9Xvqo
DCYb17kbF7KamPMzLJ3KYjTFd6EBnwTex/2UoqFVyU16JJyaKhvSZnUds0wvZbmtLWrehm/dpIbW
UdxnxvlYMyWVrs9GUqJlD8pow4odS5oYA+OxW0Q+moiU/v88R+pOL7Kl5yE9MybdbHtOJl7BXgsz
A6FchtO2PtDTZNVfiuGlOzB+yDIJTM73Wc05n+otYefDGk3nfGFOOK4MVg8xJ+deTRwWmWTSUVeK
YQZeo+8ljtfuQ5HurQElivnJV8tmFsIuMlxH6IvfatP0ZJQllN8au0/hPQ51RT3mHWaeyDf3l6Ue
vHVru/tHDNgRJJkEOWRswG4jpY9EsHnyfDLOd52LsJWB9ZrED/9pRD+WasqWBOLJmqWj2feavZHC
QHKBL2nPcTfQSuVGRbn+JliT5KOUKvXDRwyOmnFA3EO2aKnepYCldxFsFAHeZ2ZT+FlEKhlucX+O
m1eYQpbMswN6bX9jrO/NUaoXSC6E/jaTlff3YtkYam+SBplZRWG/5VZpQTMLouNrCZFeJqffyniG
smSrR1Yuuouz20i4jIV74RCVbhPXT5z3e1lIREKW+cnol8Pq8BkLs2TkQucFj5pi3niRM7ZmIcK9
a2cGUFxoeWhcyH26LmizED1Q7Ycb+Z5nbDlX3uXBBMXFAKu3IXaInIkCEcJpznXPG4GSkDykn6sE
lZj1hVNJLCBAW3JuXDgOE3dQh6a5wFcvCtiki8RFGyQb1oS0r3tYiyucYvjQA5IvL3XfEO74R6Mb
3QvHF6TUzIx2VwIGO/Ls1nKTGXIAL5iW9GgHVI9n11we00bB4noBi7lfgu+cZBECVN58cdJTVoWV
6/zQJ7HM85Isn4Z+ZS5EZ+5KHGCyMRkbnXgy/RYwVQAOo+5pLVejrNbYpdxsqHA6pDGIutKia4Wj
edBMJPalezfmQq1MtUoVh/bhWFFn9VZZ8hDXFlMVxXZWs7mJhOlnPtWSmghHJVq8P3gEUAqmx0yT
WwQaXu8tNwK3WfBmexU9SW94qKrRZjSTXx1qPgrpXuyY1sUU7BzbKpim/AxaS2afWp6p1Q/ry7Mc
QPvm1aEAxC3qe/l/1SHDq+BxNBURQJu0S2VYMvAQZG2CsMwWdELFh46VsNc2QgmjMZkqQet9/KIL
b5MncQdOg8xtH7aYSXjy6rbOcVWc04v7dcQtHqitrglawfnJyJOuGCMtcY83FWAVIdBomOPb2WjA
WEWT6m9B323imQ+7m+OHfJkcp13Jh2swkhz5MsjFCg3s4vbS3EJB8LALYqGJwIRSmCA91ADOnrni
jTdCEjFAvljIkJrtPUHVTOJ9ouBSh4tynxIksCiBKaJ28hK8H1PtmpFkVM6dDBVSUMm9Beg+66PW
FrqBlEHJ6YUNJA7gebreYF3II2CrYEi+Rff4WMfP2dcbEjqNGaOyNHqSu2nfU/KkqUqjQvuA2Ap4
vqbvEpm+Ealm0YLihDsfx5/6o63PdBs6E/8hTZi+J/TVfgwHE00Y1zSqqu9xWLCe25EI2cQAGwHM
eJC3HjqZpirET3NjCW41uj12Tn2mmhMXkKx/dCCwCju5csx5X3PNG1EzEcSVS+hhLjznVLAwsGj5
rWiahctA9jBgTnuSOYXKHtiOevOd7nyhjr1fIg6XeA/w8NtaXWeckTDEIVH9ifYcUDsurpDmca0p
Uu0OqO1CmpZ7ZQM3MtKaHTwP1Pc1E9LlWFMPRcMRRSsf94BlNn4r8NJl9FeLH3yscKzUz+m7PpF0
+XQeK+3KIMYtgpf62sltRVx9IL9glwV9xrQBUyz0YA04A7PfCJh48CBNRlaLMLEC8VCqYi6ddWAH
V8yCxI49bquILwWItdvW4Q9qOcc+z6C+/IpwC5PH5enVzyn4X4wCcWCupmBpcn05nVRxqLeJNzwo
VdXvIS32BFsyVAHxCXgihIPh0uXvYI6NI8LlgI13H3yA2cG/RT2Ix8qqAPYOc3U8pCttm0ewH64y
ZUVGl6uFiAJj9tK3OkgqS/quKG2OF1gGAJeWX8ooHB7awoDz+Uzf/SrKbtp7zcJACyBJWNhbstVo
iZLDzHwPMpEzQCM7YK0BZu4QxNmdBAGVC0ybYKsd2EnNIvp2aiO3dcTNYwMrJxFcxGq9P+CUiL26
7GMlBU1saZZn0+xNOmAxWa/4HRccAFjJAeaUdOKWz+1CBXlgERotZLnZTrbZnFOFlY/Q9YJiNPTa
wNK7g4HpnPRVaJZfHRchVZbV5zwjM4aKZryqcuS7JeQMCJhvD+qJRkgneooeO7t45vUhbf0lpNOY
SoXmn2loDD8NcUgorkQ5cToCGus8gsgEfHBHl8dGC9zD819ZlLtlSqgWcjIVKzzhZkyaTGb7WZ7x
Vrc7t8eXoLQCwRvbnXB6pjbqsKlpF1ADLX3KX+oVKSV5X8NczaPc6em0bkzONCRULohU4SaGPe/4
EG8UCl4CsPowtOmhZhPE6KYAWlHWnwr3ZLHFpoQ7pCuIGunkqzqwXiHRRCdLcjXigqqfPiBmW92P
3v4/RoBy/acH0BVYUpiuCSIO5cUHX+3MEvl6dr55WWuCCe/mkvOV8tq6vO/A0I6m3iVtFr7L9uu+
AuiRzAE0OrK2/vA+OOFzm1tHyr66GrX0AIdSAMVfGcXaklHqXcAmVRfWEQHd0mCai8AJ7XkDrAKX
wKPISWnkTtRztMqWlF4HJS2DopLFcv10S98IvI81Yn+zHVDbjJCQl9Y8uwa2qKeO1MzH4gEuvhkA
uI509x2FV+pqvZDCBVSS6A8bGASsJ9eMccZBB+cyck9mJHH+7+kw1ImwzYHAaOtfY2cfFwsVyNK9
ttJVdLiBDqUUD0F/LDrWFRxtY57lyfEGhut2oJH9lGQCeYN3O/0AcVj/qOaKtIkwTXfD7jglWL8F
MY8rcaNegieBD5OtSNDhlLgAsz+wKEp4fCvAP0ueVBWLEqQRzVtv49Ayie7K3Vkec7TGw196tUB7
ZVDcWZqd31de2K2DQwrqGftvmvizhVjrOsPt8F80NkCNK7lZrU5Zs/QJ66t5tx0QvNszDlTA6Ty5
K2AFPca6tyyKNqcSBMKnCe5H+HS2y46fU6gqGjCqyjbNZqC4ToH5S3KqTcHPZOisBxPkjgNZs+TO
J/Vo6a90vw7wvhnYszJcvwFoTqdgUKYcOQdfyznQTsXbqM5cGTk8WE32N/IRp+2SVcLl34Ie3qMR
u9DWz/wP/4aMbXacvYPQ0vaH4MJQ+3miO7wQSfGzol/A6p7uy/duP3yVCWfWWeF2hhzd1gmLpiS9
8qg8bNyPmEA6Cww6Wxm6rvCpjE0lX28H2CynFqOIsdrZLCNWLGalFmDz4UF1PdcahVOdpz9NvevY
walPtYyKpvw0N+nOO1VoJdR2RFPubvL1HkextmudPZmHAMYmQFN73OhhUqUQMlysVqZr51ikEeAS
0uOXVi00McQ1O1FubCOwEHgRQvOYDfRHLIZmZRY9ysWDmxMnFuqeRb2picMHBga3NBnVgXRPIpIs
TMmqS/pjtZ7QxUtwu0td0T+wfxwbOkUtlbAKYFjxWTjPaG2PgGtZS1qwybsaQeQ4AC7a4+h3pVaJ
T1RJJXemO03Z0OqV1rRgGt6+OjtIDqpaYK0EKdTU2xTI9gP5yvjYW43jX49qnrdCLd7f9WQJcMBF
IztqY12lP3ww06SoSI1QiNG5g5lU/5+Kh7InEVpjD71MJA+RaFc06+wCWH5W5yOnJLHoaLJrWwdm
nStaN9DDbaYUkmKKZin0SHnlUd7vSRVkEXvhO35/aa7DSNqJolbhgo8mzCZAuxwTDDSKEZqR+0Dc
ovhwVSRrD8Tn8nDVDcg3V76Y4+R9s4f0tZoi/V9owHL6c1uB6dVblW1sSnoikHpr/A1VBXj97tHA
YEPEuZCjTiJlBE+asXCIZPz1TfWzBP48+FVSE2+9wBNzhGySdyToOgjd4PXu1RWUIcdQ2qx0aE8s
opOm6eLyR+15jumeEPAbQuQksyZ6IqQLeeMMhfX9gEHnW1BqrA03tsnZfkOAUnxTVYaWe4nK6pGb
rQIGSMWM4zh/oj00J7OCBLVzVGuPk3aCYw7nmS72Ygcxo3dYewlyv+t3r2QkfjBrTVi6YYpjngG6
M1gf7Bf79XlHbH98NXCuVy2yNc+SGbad6I0jUUrs89JyVJOYcA6SHXkLrgRlI3duXOuFMMHVm+Tj
+DDnUEww+ZBaX+m1BGPowgfUnj+1XMAQfJzPa4tq7hLbUE/AUvtCl4OlbZXc6rlKefXksUWeRlBj
6XvQNGcyaJAYzUMJKdmgMeMVNGmlJmDYA+x9uQ8cwZph8txHU9afYiYZSDidadraqCpJ6Hhl/W/r
TB9qSAAakzyFZ5EhWnt06Ovqeddy9Ludi9VZNI80bisWRBfrbxz1ubTxAdoXgKztRhC+l9sQjx0r
mv8uQMitQyaLzfYnRk+PuYTEfOZY6CUboB3NtJKyo4w/EiBO5P2Gf6JCit7d1vKPscpCtdS9m4+h
0xCzx0uyOhyytx6FrvMqZ41hUTxaWV2wEiM1GVTQobTf+CWIUi3N3GA1tz5EYGyUJV5B+97JhY40
kfb+5IGGfV0PpFuGTBrP2cQHruNOFQaM+EcArWIPL+BT25Tta/CYVXIcvfoBdXsUqs3/eT8SnHtZ
pQanxXzq+t1NYM1tkR9mWeb/tknYaynew6PZhUl9vVmPTwob7LpwPRyOKh/GUIkKfM0rq4duxFoT
Jk6JHZQdbrKfup4wIwXfatPAibo+wBo/+68RsCMwaxdF87EfcDExFYmOK3q6dTmb9Y6eUYZbEdGI
zwq4nGRPauhZ3tYclsfe6Y4EhJfifP4fq6DEdCml5HJoYs0VU0UQnXbdKmbr7sLkokt3QCsXdMdt
V8jEsSYlM1SBibIarg1klAMI4/OTiuqSMzvJ+jrvhbT6pJSQITQyAorI8I6xn0vM641DBcPz7y2J
Ae5l7i5YvX/jUCkUjnPGS/Wrr6A1FbIE0S/uvGL5DSalqU+3QlCA7Y/jASplF4igx2esTcCPLuoK
PrkbYTupNVEoBdn6AewlxWTfCTC+9eM2J/mnYaCePOqpOSJuPxFj8ur/1L5B7NHABjl3bH4z/qn3
pQW+yQBxebrABChMr8ZFMXcF/HbexMwKKBSdPsKwLy9jXKtznaAuPvzciJjfCykRY9oOB+s+SGv3
x6aXStj/eIIDNz/BmlrbqfCJa63tcTBlu9vC2aw8LN7BwI8I8R+Nl5JnIAb0nhPXYgHMVl/vqP77
wzORekf9PuDACyQWdpRTvBGM0gevamHNseEPA85MGC79FDIW39lWl9Wkc7pCsWRl6rmmkQfITTmm
EdlwC/9tYTzGPuX3lPofcJCdDp9nENkCc5wj4U/vBjFiVJaRXnoOcHWhbwiz8U6gz3fskOxoQ44a
UKCMBZ7C9z2hXZQD2M3HPhZ8JEfWJh26uwDgBrn/SjRaJXh5Li+RaSyaMTnL7ne7inoqDF6wLKeO
a4fIgQIMFHyYUeo3PFjPC7SKjkXGtj2eZ8Qex5suOcjBoYPNFRTVfFSrv60pUG845Oi42yu+3XVD
Xf1M6zsh/lq088FP5OoPlH1+gbZb8wz/CSHc80CQAShvmgYFcFUB4zZF1TVDkTnkMegAWhZeI838
aJCmFakQn2Y4WdRP6iqBsLnHnfPtUHg1aERwerkpPxNKlf6WiQUmaKHZ46xp3riDLhFeuU7QWFb/
Bhv9FkINubFZ94UCQisg770F1zNfl5Zo+9uFBnks3zCg5C+ZfaBlVk7VJHyQZD7IU770OOyi1PpK
IZcp7tb87xRHtqkwqTYJJXCWgOAmDc8dukeMJ0MHAeM0jn6877vrP7qGa4i076yJif7vDgvg7itv
T7fXzmkJzaWnnybjnk4niAoSUK5U3QvKtSsghoL7Jrt/2y3UNDjfo5/DdDCOepbLl9YSNwXAEdkG
w1BlN5Vkr4Yh9NmrAckknIGQy6NUotZlA01JnD+V70FoM/ptLGOs7yJQfcoTcS+NmtBRuon9Tvsm
vPqqu681M+XGKIWpHguw1cC/VhsdzsDGvfWrIziy02alPFEhLbyakmhQR8Tez7UGI9IE4yJdfD36
a4pAc+nZb17wEtTPN6Ddw+3bm9b2Nd7TQM1p3V+oKzQ/A/DQ620jRUZ2Sr9ZZxvFntg9TXeyPbYT
6dd6638S2wrwQEtJq7q4WQUCLSWuqtG1yi6X00DViINLKWTpOFEynWcqFTWuNDK3T8AvrrK5iZZ/
vZcH8FMLmHcFN3eDJubAJqNKW1NIFWGPS0+tUQ/x1gl5D1wlxCeHkM2ge+alLN8X2oHHaN8nXgKa
zCqj+jB0YFExdvF5Mu6qSskfV+df1jpaTTMtOilPb+NuEgwInBnBQZX9oyE79GCqFtIVvJFdTi0C
th7qpX7e4ZxhJ/D7EjzYL4Zuct+ZHkI/NR/0aI5ivwhoPdV9kRZzQsM3BJWElR9+QYg7aVJyNPQ7
D/CJl4YLK8s7fKQF+9UlT46iFxTymZgZiPqFGFTNqcX0teCwT2ieDe2E8AeTwDX6Jp6k7grfeKpC
xceaBXkJZZ1VO1x/CWY+fb+BzxTCsgF1LMD3OptgbtL8oenM5r4yS6+xSuWTmtB/TtS7MDELQG8t
rD+qkKZtDjRKNO8V2hKGlGKTd13iNKLk5hL4+2pRkk3ENDxvVkGpLevL+LQNBVqD0rBMONH/5l1A
Dzgqi5jkmJYkqGn1/eNGqApsb33CbkYxms/5/ATjD+9ZAzUz8cT5F7xgjGryuJwV9C/laILXZHes
2rBVpAIGPHI6CGLSY04cJ6sNVmkambyhT9WR0N7EvfYhywHc0yXYJwQ6D1sOajr2YGW1Ri1pnT2E
s4MwwnQocgxNXl3xV3L/NEmrreUTW1MWpZgamGzTohZ6voXvdngvr5ZbyIr7terh6NZBs1KMVOei
k4Et8ArPWEtNnyLXr1T7fqgABh2ch/C+fbFGB0NamsRYPkiQ/Hs14RCupRP/X4833oRqUCBm569R
gt4QazhY3Ecz1uy4YeJgDhcJueznSaK3atifDhJvaOlD7JgjzhXUbYCIG9eTPg8vdbGn/oXRzZB+
jJV7fOGs/UfYbM5YR3LNtVwRfUP8AklBdrK5Fq23+GeAdiKIIvy+hhXH+ZaQD2mFrEzKs46ErUUT
mszxIga+j1hqbVUTTtZ9zxfwqpVKssKPkCxuALsJDvRkPDJyz1iAiT38GpZPrU9w97jwFF0ifSaa
KGK4TphnaDIcFKBQKRP88WgOsPoady9B2ooUhZpTT/selivPRp3xfPblSVSienPy/4aQFzVINXu0
tbjAjhwgyoo/UcTwc04envJV5e271lY0stQBVMeYHJdtNkJ83FfVpJcomhUrnjk0F1FoPcQq5InA
lGM9r53fH/DiEF8A2Xlopt0O/vbCHld4qD3HR1KdAX2CBguqAqMcckt/OubH45bYygl7znZcPavi
M8esqSyL2GpCpAQtzOs06XVkwyFu/un/5mZHVTZ6TauR9ykQHX/nFUgHlmID0UmxM63/K9YQWfAR
ivdNbQMkOGGI1pXdfYkQRlk8FBkJ38TkIjf/6HH7Rr3IMtr+JPpP0062mSqs1acAyXhIbL6lfWzm
+EjFFHlwmFQKdT2YnGgb2PCZOZXYzCf8UiL0R6t4wmzqTcSfUMGfuX0ssOfVNq6aoZgj+JS2imx2
zGFr5VbFQJEDs9RiNLkrn2LrWAfPG9pG+A2mqlsslTy07dXqO3mRfidQDIwwUCqhM7Xo3f0A0vC3
D4gYy6sfJ2LvzH8pGfctJsw+PPUyn9/1xJLQffr/OaFrzBaZ/jpPO1CmGMItdpXfLQB8/pPWy3tA
j0UTC9E7p2OszV2mhm/e2KJJtFTJWVV+R7Ser7rVGndOgzCgaw9y9ZCbCvPjC1LwJ7cJjY9kc3/H
IyfjvmJlFvnik/seqbcJxlccvTIlX9grTzxxtL2tz1u2ope04dTpYTTk6u1znKKNnBxHqnr+TeA+
rDJD+Yy21nNGZzHXQ9MtA2WQKBop4BCYwWBJJKpkT9Z1rCwKM/AyRSYBvYg7Qpu7s0Z6szQg8w5K
88PlBxBnij/CeYp9r9fzg2wY9P8nQLttKQThkdHpC22Vh5QRapY+e/GFmyJbTLUxims03tB5MbAj
Mhzc6mTMdH0ISQAGXkNTY/H+psb+SFkW4jV0AwF8ZI5mqjWFVDzqU9Cbz/oHyGXJ2lNmXv463aQq
/LNwEYwat74VHqwLregA5T6i+cPu+P9vqLoVrohZ4aaD6VmhXpADQ0AY50auQY4y+vITRE3u3+e7
CtlQ4T1amqAomWhN1im1aghECOA/+QzH6rjiEK6FAzI9dYqmjYEOTc69eHcQvBzyQfW19+vH/L16
M8b4BOyztc6JBmY/zB/wEl3pmp8pmBu5WU8GoybgXpzOtmdhYTZV3smUgaB8N+XqTO1WpNzosYnp
dFe+3AuyMG+4xKIfGRKV5Ut4qkU1/2OzkumQJVU6JW2TvX3wt/+EkOwutPbpNchZNFOAg9zpMnR3
G5/Cr+rRWs2mltXtz0oG+u2TmrtVbx9YDOWNCo0QeoSsz7jxIgPuv+ckjcaWCBpuYN5aZ2lTqWgP
onrjN2QczXdwazXZlhzaKqs4BeS1WchRQQjUYsUbcNqwSBunLP1rgXZPn1MnJ7MukgEVntLH83uu
qaR4wRZpgNe1vxfedZQE/w+p/4YkbfNiSRSoyJleo4Q3PerIkjXceMBrFwrWySkZubvsu7UjOEsb
ZllYoSg7fvlkhQs9Z7Zv+Bh/+BUeTOyUo3RewyKL0knyzMEbJrCyMFyDr4/ib8CBfeU+3Evvz4Yw
CP7TeXnwlMi7ePY1+YY5g8X39JsM6Yf0lW9/0i9cEKjr5JvY3MtlL9LukZViOTwmCSGJ1DZVlprr
AGsrv7Dl4UwfWuZeG8JGYF2szMFchZUNJ6OBSgbFT7DU/dOZBKy38Pxjr2HeK0zNYdRJeUMyIv6B
77+VxboPipldTBcDFN9+R/bhX9inGNeM84s7yN1PNMTOpVlzzAykkMwCLgUQsFEWDfzpZ3uQbUTY
UdAXCXyTioXSIEYEhoZ5Thkh5khA7BNoqGgr5Tzw5E45Unr6VWnVo9/0ggF6vuhfTJc5v8U9Mdu1
vro/7q9UEqMcbloNImGHbWCeqO16lsatrP855jA8pT6pnWXykVzQTFUv89JOCseu13dSXY9hDDNO
RV+RSvhNICFuID7+4oLyU7AmQ0CaULpGy0xLurR/z5l3l1NI1xhPhHyfGuyzydprKuJnX6BTj4RN
i0UDWJkmY56Y8CUU8M7xGUEtw5SmHpZhpsd3eixfsnzkE6MAvVeOMQ7Z/F09AIPOlBevKO42qspc
xx7I4caUgDJMeF2KG6zscDW0anI9JdTb27tSMRu/fKu8SBvfsiY0pde1XtjvUJ4qA075B1K8xC/s
HJwtZLTP3vpeS8YPImnU4inz6dYq5/0d0TZcl0hImE5rdfXPf/s+m9By0siSU3YHdzRtzB1A9Jkj
XSXwzlVrWT2C+47VMinETrvhrReRANGzDhSN6ri4OWxLDoKtHw3UDEeuJYzw+ZFDtjJtoyuLhFN9
KMFTV5Abg+TwdldJl+xg722cbWDVlutU/SM1X1AAM1kwqSPnadTk3Dr0io859UQRLD1NpL8YISAi
6vCfCacFM/hdRUHDCC6qLLsfAvQWsg6OwRRhXb6mjcL+KDgz2/Wg/sOk9uyJnwAb+S5j2hJOfvGQ
lbH4zsZT6ZYXu9BQfnls9XdwbHZugrLxHDThEyE8vH3VwmEjJJCEbjtdfhPxvhAdtmWBgty9Umpz
qtTcRR14Qej4CiV4EnKtLGFFJ7TxJOZBeHugpEORwytrej+umSvIHO3Qb939Hs0d+oZsPMI8+3fT
NovbJI3iwIL3eOuCiP0VgZs7fSAKoW1PD6ZgVOFPF0ip8WK+svpX9iXPXQs9eTHP7W1oRFyJigaq
WgeaVeo6tDEZIIgxAs3X1gn9aochwOul3A45nQrIYT/Zz9wJaqSBrgOYkVgVr1nR9NzvQPfV8KG1
+ho+vLXWh7UOWLrLRwrNYvpP5a1NlgWoXREmKxWtEmRtmg5JxwvsoOGcS0yeiDCKndKkfbxGF9k4
p7GoTTYz89tkjEi9Kox+Ab+6qkr70Fa7bcWXDA4PfXWfSgsMpczf5RZ1ROl0XvmCCgoKSQzKrlxL
jH49md9gBDMTBHQSbh2D8yUdiMcoplcChKbBwnUdKuFufWrG3QinHWfDBGk1q7PdYQ4FYGI7f3Pz
4dLuEv+gN+vUemHoAK4Mu8oru6y8OQ9YreZYAXMKvtRF0D703XDnahKkhk46g3yzk2W05nlHOOEf
b1MhWzTLBNhvjGeOp130xJcbQmUTq6IcgmJ22DUB0n4BQkU/sVH8yA1c/aZ4DkQCUg5ySINb4UJs
/dcs+88fJ2W2J28Ahwx0tSc1iLo2qw8ZjiNK2YvsFNkJKoAtgUTOM5jwwzL23j6qCU6GlXZR9Req
BZnymfUZf15OLrcj61lCGVORaKHY8ygz6wkvXuI7w1m9xsn63d+yYFabr0Z5nqIKDT89oXv2Jj6g
Yo1wx9iB5MMefpazRA15cCMx0wFEwoD2RQPBphRFFLZii5M/v+13cEnFmprS9yMZaZIEYhXXPVjd
+6cZvFi8VH9u7PRiVgL+M3HbS2QQqDMZC/6xHnNWdkPJRMFU0c14uzSz2ykZg+tWU/WUXO0humo3
EgmOXR1TuGMpeJ7A0P1xl1+A1jPLV+xf5V2SM+POof2WFSPiuYKfvHNROWeQPjjE3vEZysgBfYOY
9q7lGcWOoGVw9rs0nyOcJXFOVUVyqJrJCzXdJitMn6JIRN05B3or4HtcGLHnogFNVqFUl0n2qynD
012YqFLNy9gHZ1fA7VM02rEBLdDuug9SMq6HBvju4uyQnJU8jWXPRhcp63LD38/ypSwFt8gYjJ19
lX/Dxs/cNQ8oxydmoTrwGhyEc0XzRNSGlJcHa9OJPswGV+ca8ihmnUkGG0ufdYKFjBo0yMoYDOxH
rFM1F8nySZXx+i+J76CfjFSXB77prgAspehJnEaUMqumNpru+BOih97mQIe3HBJhohIyev2GQudq
PO3ugBzJMGubUFJ/S1OIC3okJL0qSIn4VGk4IuRL9rXqFOndmj3/TxmQ9V8yLx8Tc2CC92E26B9x
bWNP8/+xcQrrUz4cpzpDbLJhgJArd6mL/92lDBhrP+b9IAjCjlaMfrO94izkgzBykClUISnaQ0JJ
IGSpP6bFErp7ekw3LyUBTUbj6fbZXgwxlW/oDTRQt4vWOcG+KHQW29QU0xvNir+PdQN4Jp0eGMhV
lbh2VGd3276sNegUm+tDhrDXbbFYKq9bwcni1BOWdANJasZ0wvbOCw/R+RyAV3BYWZNGjDfqFna3
nW0ULtkqCfu/CQRr7CCBu0wXOs0WB3xIG6qF+ilBwvFHMAlrIVklZZUGhl81eJFqaz1QzgwJouer
Jl7bOn1ttdI6ftPFvA+WeNT0ppmJZKriPYsAyL4XC4dBoN60/Oq+nPJMOLsvgR+vs2CQuuDNykv4
t8AqDKBAjrMY7ukehvzzgkxj/UXGd+ZswCHr5iNSmULSyh2Qn0Jexff7cEqvrSsCrlNZyIdO9Rxw
NZU7oacyf+YCimEI/v4oBoPKfOo2BwR4t725mtD6mE/aCf/XrFdBj0vHlignxgfEKdXMQjkh433A
rljbnPup6X4Qeom+BjA+3ffO8E1wQk4SdS8yc/hdX8IoelVQxpu+3NFR5WRoS0jGxmhIO/3v18DC
jifu6oWXFjNgmb+JCkM/b8Q8T/d54DEJ/eUIW6x0qGGe/ZpR3WGRWnEh17WgvIs1JJ2W1AtYovA9
QXpnUAAfdDqiDMYFswc4O/CNwxhS34fKFBB83CK6xTS4SZGNAHgm9O5bHxAbB7iMSt+75DEFCUVV
5lWJjGIbfOdFEYGY72sCMZmUL/GRTDYSUJJtgMsDRZYVE+Rmjb5RXQ6Csktqh1NeRg8I4TEM4S2j
NW05H9LAGV8yF41ydVbAWWiTewNQ7AhhWN9n7ebGKg/9sTygeEx8PiqALnz27jJDpgx0D/wwAqcm
LuzUUCoCtNiDBSR26S6zQ9RqFF5+Z2jBbqBOqwaFH0wesxSaNQITVlLiY8Erdk/+C8DPsBe/laN6
VcXk7O7TPc+Mt+rqSWqwoDhKzAlggYUq2CXdz8C43XVLTSAS+3CskBjd9Inb3gya2W2w0XlAcSTr
cT6aVuhHKXu5Q9gf5O+oCyErOZl+KBKsabEWF8uxGpcxb1Zdhu4Ol1vb+O8zlZAJrExU0kU4Q+aI
frGodNQcyAVHbtDBPoCMfa6tr3qkZ1GHjagok05HpoNzNj3l/2pfkFIofMWouU1SLzgmcarWoBUH
wMtNzxbTHQDlXrmwgLRR5QumTKN9gzYF7yXEGgXG4f+pdceiYOYgqJEKfcpMJf8xPAR88kjK+4Gb
Yjeei/OqeC5SGg972iRXT0dtO4VjOmso6bsTFV02jBBc/igzJEx4Q07XYwOZ9TlNqyqBJEeqDPEJ
ey19a7bCCvlVuvndLuqRG6GuatAb++vRZBYCh+Tl5zyFDDo9Qx+JzO074oUt2XFD5lJSq2MEgUOt
6QWO6jktuOxeJgmVk8ED2jll3En+v5UHtDjl7j822JRQdd8G4R+BjFSEwoQgeDHpOTKYcwJZeHoG
yNC0f99gWbFVWkt3PaLVmo97jTUkuFt6IbTudNirlvUXbGTngtnSoZncxk7qWfY8bhV1XPV1flWZ
itNdoHZgNGpbgIy893J+gaFqBTzadpO0TsmpwIWsEQ1NoaITju8s/Kmya70zyXX6YCoxBhCEZPsC
fpl9n0kxO9PncpUgb6yf/cKeDh+C1LuQ0vLg0XXkccmQcbf4DwlGVE8Mlcti+OqXrGqqnH+rgmDW
3BhdR56o8WFxEaLQpOQXSnEtP+8Zx80vsMEYuikL6OGRaGGMCM9zIZH3h4RB5MRKNnAlNL3tHXZ2
ISaUhg9DnXA6iQtwDpkQD0NTouRIA3vhl8tPKIeaBvtwJUsP20yZgUzK2QA7S+pa6W1vYt4miRu3
M2es0iJ7PLPcExpWk9rBIZ3EqWoqSCV5lq2BxOgfcHda4pJE95mALxAy+B6hvLWqe3Yig7zWxc9V
SAA3dFj5u3SXjJ+GoSv3ssuYcfPPh4gYy5RbzvKgOBJeC6435zSKhdtG/hUUFxr6g5OH1fmivpiw
bUoiEYXi6N1Fzk+Lu/FfB6/9goYqrjidHO1GhzGr+D5osMcGhCm/R2U/ji1UoY4FZN0M6umL3lkg
P5CeCvlKUP4BdB6S83WAfiNunO/fms0NzP+67xTfRhWSAp98N1G/w81l+LISugUBKq3YYu108fMF
XwpQTlH4ehweIlfk5NxLnNB/fZlayE07nFsKOOyUCdThvBS22vC+f1k/h4rg1ZVu+oR7QyPdjJkG
w3Fg+vYRnGuU+iYAqBHzPGvtd1K4s+FgvNtLMzfwF8eJOocq/W8FEpY10YVbTsQqmgnH5GeSRZyJ
boahL1vaCB8IE3IETGTRwYbXS7FHUNmdbxST0yYWws2RZW7KzEjXMUsB3hV/4Jo+G6G2gv7xnP/J
4KEuMIPixEZU0pS2/8+j1xqeayPodPIoE1coWh/TgHae9n0IYEW0LJwp8yywsaTAQaRzHk1XxzR5
q9q+4XqHQxr74BOkT81RbHMnZy5FtUZtvudfsFVDtfKYdMzNgtyOQ0WDMogi6+aB0vGp8KB2W1en
bv2SrnK4JMJLK2bYqHn+X9INx8/Tagz/n3F0b3oQ75U2qdzhG/hgJVy0BQ3UNT/zn9+lDZr5M0I/
uJmE/O2pD3k/iJii89MRfxuANzqDfMG8UXZ/JuVqNl53St7BPEiQ57MR9OK9Z5XyAdoDW4cjzNTe
vSVfOB9ydiBWlR/MP+pi03BXUw4YGZIUES9ZBbu/GPplV6WErWWjbI4AJ7Y5W2baBvVUPffPKy8P
CFA4a2gAnLQCUgxyT/o/DiSqFxULBpJwu7BGEiM1gWrkd9TG5YRso/jXGsQS3r/JZUM9p5ASrXve
vsmjw1GIpaIDr5QrVAVHYHqVMlWdsU7DqspehS4HP+MXfDEK8xeLY/6TRYoUcnHXqo8WuBqZLVqb
cFnFofkM2g51Lz9BBBTjxRw3mUVcmFbAaQsGzA+Aqr6hiZDWHXbO55e19XgomVd7xXUtSjD7YsqD
MqxYtL2Uh+8q5V/gaxBmx2ydQL4u5nJDbc+DL1xFQReWiWZwVhDnVdaOnO9VJfmjh3XE5grVVRFf
xewcl/eCbkYnuf1ZxxGJ9QMP7mrgaYQpcZ4YACNXt+w7mjzgNaZ52uoG5iGKFQc1FqcCaO1NryBl
QKmWtcJwHJvi0GAT8gVaZmJ7o4l6k8eE27Pp02qO6DECHOQhE/X5dfiNOTEMxhziywX6ytwDRSq9
pzmBowQoSDpaUxzDoTeTFZf39RWKnpJVgfiCtNyBbk86vuc5cIXhnvcbbBEcGi/Bx5d7chb4iDIz
C7ncLnmOdlyxs3m8K+w4sjiyoFm7u6iq9bc4/QHJCEU0snAp869Bk6E//m763nIPQ/rJ9OjNBcVO
8kaKCvDlRUrINMKF3L2Q+B70xSrPSTkpEsF39WVQLCdl0tx7xqTfqYqhY+RCPAZJ9cyyN5ifTeX8
hzqOrttUqPwTkSkjXy0F0T2u+IMNobElUixWx+TP3YD8Vfkjndtzy4LPXfdCCQzExawGWl8PVW1q
JCFAP7XiaZceyUcYoMSRXjacZ2q65YMhgJKWHHdpHAaEjNkwbD93drX+TZ/pt5DlBAnWHb4a2STB
Gbem6qOnsDJdv6feXStz38tDDLMt9YE83JVcO/k+io5a4g5/AiaDTT4hNkq5zYcCg++WU2YhSY8S
S9VJg2OhTM9Agt6+KOTUJSbtnTys8Vgr51j0iYeF9yr5FZtMRByikZ1Tu4S2Ft5xGI42TsIGBOcq
SqESgENJgSv8ypUMW0kE95vQnEPdA2bSyCguLlbYksDWrof3ra6MDHmykhZpcd4DaIViecgvnvEM
FWbEQDVcMRphJch4SXRP4uhDLMtTojNXOxUa/WQA8q71JMZ+T2k0qBZ4SkHGFuic/azY8lOzJZT2
Ohfk1U8iWBNvWfJ+XHZhM1dT1T8AKuaOJQTzz/GW0LptVzo0nBXOPXIu3/52PqqDR9C1Yd4LAFef
vyE1vNh5dhbT23h2vyxSln1HHjr+EPvOasbafVM4YESo+Vqo3oGFd2uLuIz0620rsggrITHTbxA6
K+wbd4PJSvxnhTqHN4Lk48E4xazCVVIk0M/dWUrqmBjPVv9ocDKwZnGbqjSwj44B1Wc2G9g6n7Yu
85jRDBNRkm1Vzw4Y14QWKMfxAv1rzC98jOgSs8tnGqCvyAEaAQfMYJ3UdErxiKLkDxu+viCXjH1N
3d1Tp86EbIEpfCkm8u45177zxzaTUhPF2qbzjlpQM3gYU34qL+ZVCCJpYKFZ2s/67D3E/gpd/6Qe
PZV1xBFxoc6WVL2G+I3h9LNfPSeSo1cH/IDDij/UOqVJYREQMt25df/TpIL02x/Z63Icn77xP7YZ
ykUyfvUJmlVAbNyr0NXZ52gburVIQx2HgFMf5RM2aez6tjiNxnDNn7kDAusBGFst1qlzM/ZmApq5
fNmlRqRBGC9TWfvr/jKUzfe56R2L0ooiAPdTlTHPOxs+hvdy29w2JJAyDWksCB//Ysi4zKHFLeoh
KdmfWb6rr9qI6bOLOy9q4sa+kP8puecKD4UopT8sgYLrGSZc+Lt0MiYjRkEvms1ALT/BvIknuw9K
oBKFJJGcCKT/Gt0Z/UU25tof75ufuOtQeZPCI50YW5CeDMt2+UIJia1+QTjA4egZMgABWH7QNHTB
CsYPiot3dFCF83gmRpDXVAuxNuVKsrpUAvCcMkkaDOdc+MbgQAxV1NNCjz3sqXA4iy7BZ/LOz9mw
MkrwSFr7jHrTc5AKo542CY4D+X1EznKOoggUw/wDZJ3QeokGyMsTK2jB/+ugWCJg85OcxlMXk3HL
fPEYGbMIMaAGDHUL3mUoWZonEwYrnZJwofZeReAGKcJAQNpQItmKbFdU24EUTJA94qdqfRR9lLry
QPPqiSwURuOc/z3DjdQ6+T8X09ONcT9gNHkqFpJbQvmreOsSmtlHi25mJHDChumMlmAAmzaJWltt
wJvy0fDQo9/9oV3sl5Uhh7yTlscccyjAEApD7mDj800ul1RXD/6qFUuGV+CtMzBVNLvAxnLjeAJ6
OXJBqCPWof1iaQmFNmfWAlqRGH1SdZjS4dZIhxT4KsH5WWCDEp3bGU7akVL3S9LO/z+OAuUuXolA
/mjGDfge+verYfhgSvAm9LkHHj8EJqZIYQWf3PACYV0oNGO8nxagblejrQ6V2rkwE/wcQJuaan8j
dyNJhcqW+wbU+FGK18DkpV0TB9vr3rLu7t0xkmM5V9LLf6wdbseEfcvNe4nas9Df868wE98bxgiS
AcMKyg8w0jizDlnBUGMbuKB6Fkv/PLI75Qft0phCSXTfX0rk0YRu/MFwpb0tYLHjshKa53Oh6gsk
vUoNXnx6UkYsXtNc57FpODa2B3YRSAljToLTOQGOIO8ml2wZOuVLiQkwEzGmKRZMU0tXrU/ykEy7
DdF9bkghXo1yODnIvD9rV4q5O4fi0yffXsQPjWZxfvwIzIr9qfcg8JsxljT9EtlklmjQWqdxrIbe
9/NMehlKdRN2910SlTJS3D1ekD0UPBzRtQcnVgVbMLY8IZBIFSEPMFXaOKiAxtIgaMYQH0rwldoG
K3gyG+v3y6dgWqf49fPVXSFqk4CLl+RMy9+Hr5iqM6wbeuAUdGoMz//ufUnxNxCwPyfa1yfDPUwv
BGqDCp8bSxKNVmN4MxsyCgsCHHCei6fFB6d2zxPpRxv7TOtX2EqxrpDmAd6M7c7CI/HNGYHDqI7G
hbQbQSWmbYy/hXRIi7wTVhlAIgEWyn+6sK+31nT505itTSHyXQRzOOvTbY1UjICTRSZOGumk5dKr
0wBhhzSINHqFVXctHOp1Pw0/kVutjFZdnQg1vcNEBfKQak2faVIUA+xHuDA7zC4BcQ93Y1Yr5Vk3
LgnRYcq9TWEgQoQfHqNGauwIIx6ZwEKgGMGELnbFYigkv7yt4mthu7OYZWZ+yLvAC4+JXOKSiIVG
G4E+1dXex1WQdA3YnKNOBrRdL43+IvKto8d0SPWBGNRj8hJXVFa7zqwlj36II02q9qTtO+zcgUfg
f5px5CCu0z19Dr5d/4wiu3dtPSum+ivxosq8fzz1uiiNjOgCGvwbo9aezmumRGtKsnY9Ji/0BDWd
eVuUPrNETvW5xdKpMlwtEHkFrmdQA6rp2NddPmxVLsLAbqhGseS0HT+6PZoppt0bp9kEvrRj8Tbp
0knpsjZroSCGbmGdZ85u8gitwTd2GI8MydFBozOA22KwB5Tlq+aSnxQw22mKH1Jx2Yxr1axmMS1Y
NdOPSn3yJXQ4lpXWYXWlGGqezTCrLEVSVjzavy7ZYmPVhNCANWxm+LkLZQs2tG3aNL22cJHYw//M
IE84aJUltV+BubRG3PhmGVf1gqa7WXuuQ/a8WOIcmIgAEW9ICqhp1b+MTdhs1TPu0/tcWf3wAM+t
8CUxZNlV/BThnQNYCJsZGA5Jgqnc2ZADud3T6Y+/TAlgGhqycK+6WTkWWZtr9bSr5a+fc1H/609d
mD7pPtVz50sey8orwqeOucWJCALCNdkWdiI9WamDAFgqT/tfSoXMGwfNiFVaHGNg+Ey5Xdauguhk
/n6ViWVoRX0mMspV7WEkj2Hi0yvhOZeveMRAgu0GkircuoHvFU1aUbmpO61RaI5S4Uk0YQOnfh49
Kb3AewrLOCmuwZoHUeg/JGahya4LNa4XDZQxHfL+ujb8FQb9H6binjX1DPrAXsL4IkbNIhVhGtSD
ozwWE6U1p6xYaGFy8cbR6h7PXHoDcrrgg8H2Jfmhj9b5/i2arD9OBdhufhohPB/qn4tBsAhJUhT+
NknNMNR26R51dYIHewoUqDFFeTDwqfED8lK6HFLqkVpUVK8Ns2jiDaauLkmZz/aVvhXKJsxeJk8E
VAGram6rgHDu6xY7sB59rs581AAFkwer8vDa1YiwZC9NqIoI23GISk5jtDU1AaUpnzNrcRfUOFyF
MxnRmP44Ib5ZyvoCiR/mmuMh4bSc9JKZ9IUTIpZWaNBw2SqCIbcTbDVs68zedskKMfmYAnQvMAie
bMeSHvCaF5BhD8EQe3yDkC1mg7Advbol3f+QIinW50qn2Ga0uSZHzqJAQ54JL8kYKi2zsbTHM0d6
jHLE4Tvdyw113jiyNMbAb5OP9rOVz+K3Mh03/Zy1l/jj4kMOdlQ3Wd6h8SlP6WfMh0VmtwwRTZIv
+8NnxAgUcfd8ThRSbAogbPTer0HkhoECOUeOpOJYoigVfwt3KbZpqU/WgKvkX2o2GcBItwjsJO//
LjDjnwU87p9PK+3qgk9caoWeZWRsuNiVqd9dq99dLGi0DheUFmEPcaeXKXqEl8jmjiK0wpnzo1O/
C1TFgHPk0Fl6bEPhs/8Uax1nPC69DYKeGtWLdxDkIjQYCB/Ix4/B7GnfR3NXJ+k7pM6YBzIllG6r
/ZeTkZlHhgcJKeY4EMNGyPZM+PqvJaZoA1JOurSddhk8hkFaLwxAl4C3m53v49QiyaqV4MVEdqmy
IkuflgFy2VZyFWfa/eXOxSwUQ1mMJhJeUi1UZGaRa4TlF74jpJXrs40FDqe2cORMO0Ugd/1h14Jr
jAnTMlLq8gnPgeEEWArWao8w+hrCeoDidlVPZbny5eM42YoXfG6ycFkw3DMH2iiKgY0C3Uj8mini
5jWDiK3ICIyBFZ9ZudFdc7/in9jia6gdiPdJfyh7dMsyqeOLTNRRs1tBb1Nav0+6JeKekVyQzOdR
z+w1GnzvAdvWPH/lguki0q+mUz52BNREpXK0GUch4Y4IbJ0TlQuH0dmURZzZ4fi5AGYWOENAyk00
wDWcymfIix7lG5y9cMnB9hBEFP5uDiMUq55V0+tBfqoOx7Rs6XympfX1XuI6HCPV5cNEoQK7RDWU
IxksJo2G2okvgUYDe/TvRtOjOzwWAY1O5MdeIYEqW+NNwNkf832APRf5Z9FTvgZpp0ZYuI/jwqjr
iEXzM0o0/qzgdla+V9IrdumDk5zZeyjynI2nfLVLwpLCVsbRYXOtUaprWVlr+CTDqr2W7LFXDkz5
BSSE/qPGGGZGDvBZksrUxjKBau0AbdTKgefab/z0oKNK2MXnTCXdhqj2Uza05TQ5CjgodyHr7wfA
LSQOwiF8MrCJHFWgwSfVhMqPspy5pCNtIhuqNqIlXouJB/NuhZPAs5QfmYmnDFyk6DhBCmYV2ltz
26jyZ5Jfd626xjbcdEHuWaNODV4vY5PfEaedFIiWAFe/mZdlZRUksPRgKsNOKADEV/ZQwExbYBQ2
gT/6A3UengLdxzuXQxOGTgK69iKqIOcPP0oNPkp5wW6ezfx4zGMKwYyuRvvOLRwGbjOxW/5gnxDG
GECMMtlqo/5TqFYb8RKZgCs9Qy5eyGiKa69hAUTHdzy+GmXg7lL9HWGIFiDs5wMBt+7bhiMmjRa9
mpycTfZ97n8vT/QOEidCvYarl10/F8JJa/0AM8cGjtIxV5D0QDiJ2sKrU7C9OP2WlQr3Ukc1XQYj
8k6uovsqV6isxDNFnXbdO+RnGQnb5R+LsLN6zjOsabesS450XtJnWbXVPO2wkheo8fwG/6Y7HbPo
VE5ASUCEVcCSlZIMPPKHXnapj2xRFzXaN87ZQZ8XdYwD2s4ySvTmkG+5TpR7CikVhTpy14SSXlRv
YexwUjeD5N1eq5poF8j82w9TU9xkB2Dr+H3OFeJ18v7f0rzrlku0TN+lH0jQeZNlQkPcZr1bGcKG
QG+mXhbr4EsWDvySpef3wsYXo8S8Wzo9Jml2izIU4miJumOclcM6bdyCnmlMddr926/+0Fin5Muy
icJQdJc+jXwFOQ8cwvmHyvn9FAtOTQdtF12JcJy/69xJ28wqwPnu0VdaZzQCg5rZpqLiTa+9EqFQ
Ti6DtdyjexZTYyezws4LK+6A5aIC9+9fMm6nHd5gfG2h8gNON3NeujFdzpwBCnFuw0I05IGfQAtQ
RhFHf4k32wdjH0Mi/baoeaSpiP0pA/5OgpJO0gOHGZNJLs/OFnWLTA+y7eyfCbvwBr+SY2luvKwv
MiTeF3jIAIsUEE8GPgKMjf/Cl+UjaTf7ipZS57yLUZq9UJKTvptwLpIDHTEzqHKzjKDpAAwaPEY/
d2AIqBjlRMoEcY+QXVdquAwdxW8q/W9oRzhn9BicFLk3KSUTUu3yyl45iyODkzsCbOMXOdcH4rbU
5E7+iNu5klZftuzgVJdalvpJtwcRrYnWts4nqvDdYYdjcgJjuK6A6WhZnYOycnZp2RCwRUTt2J44
dg36IFAkE/ThNFMm2mcIhjDtlqF9JE4rjHruUmojJpCKYD654PUVQCHA66hguxu9DBLGa16I6IME
KL+eGJ1YJQibFV7eAu1xN/kxCS2Ck4FPILu3F4KyDIUY5f8rAgbIQkymxpksiMuGnduPZL2o6UDB
ADukuKZlJOfyu5MGwQtw7cLtG75se89v71LU2sIMxkwS2V01iC8tTwA181kmeJ9ZMc0RSTwJ4Q1M
vW0/FOYMB2SMSM4I0UeAXrJGiWbaILROZr/QO+kmxnLv49ivKAw4OrqL3ZVoDfm5lz3hFVFd0igT
kE/LWXGadODDu0+up+PoEaox2IqwZ+7qv/kIv7PXSwXoM5UZd9ElcymWk0usWhysv68XzF/b3zZC
AFB82q2hexHxm5njCQHnx8Vb+v3v5aLau9PhHIHBzTqSeSxcbggkeqhhNtulezNphxKxpota8kCl
jNk53Mogf75OJhrgxNNYbIeqnXuG2ETqRhtf8NZ2nlwGfHvSGhYHSTGwG+K8dtkhFE/RHjtYWb86
SPlWHo3cDEeW/hNtJLdZGSzLA9gjrsnuHbIifrjJrvlWtarTkNT4XZCNHX2wz7G5IyY2Ap9ZPMRA
/XJP1f/6Ohf5wLf57KrJ+kgDjfRY1mDaVpBa4t4JJnQDTVEVDJ/65ctqj7jh/GypIysrQ8+Nyq8M
JInvRVAr6b3xvemEPdBL7NKp6mw1VUIVlEiVML7j7Dqi+sXSZqxgRREsKC0sjxVboiaT9FaN4mBj
UNl5fjIKBKR0YhcA6rb2hH2Ls2SxY486kDEZp97TM9a0z1iChaGkOuxLhZjqlcf2ZAMWbXjDeCFK
hJzuCJOQhXd0wT0yGNfb29MMuBfuYDYFvsBx+D/7ftuhWu7fvfb5NcU/erePJW1SyKmqZV/uVU7y
S3NSru7HToPup7FDjvw0VDxvKrwVmqoUP+E+q+ZZQg6PQR5IdtHoni/zAZHAfzIpqxHxcWlBXZmf
y19MtrCaNOknetXOpLFbaTcH6x+UgxNB0sxpxEQ8Mb5nVBKq0xVYZRBs6POFHPYIkADYxVs2LvaG
7t5a1CbQoAu5oYUU1v+mZ28/1LQroe7VVtIB4uDcUcdRd1fzOrbHurDBneQnqh+i5qvwFKklmM1p
nEteOUEf0SoyG/6wfkZIQwRUficFnrftMV0PYrtN4jDWV76aad7xM9/57lSPfM2hXFdl2JpAfkLX
DJqAjUuFydIAaRReyfTSnaeMp92asR651NDTmH9E8ifHX0pKufhONF/QTLuKllWMk10RafTEj85H
AGuAANfSnJNlWB0bXzENO8X95PShYyvZhHlXb+8Z1dPLJ9AWpBjAAHXF7L5Rwu5ACmmKzX1rkrEg
2dwbdlqjxRQC9myuk9SdktCWfNQ2padRqKds7difdX9eI8RWlBr+RrxeKLvWP6qY3/8J3q6z3Syg
8b6ydnUP8NhzTvxkdtqhIV4QhjXPT78mQm6VLXhrsb+ejmoJmi3ebBO8crTJIebo6m4fMm27kbDY
7mrKnqThgJjgnWZ7T5ky/dgEy8+s1kezoJmx5ISIITwVDLwd83tYXgaqptLWGBMk/0C88zJ5QPxW
z6cLSZLGXW9TviLuLh8zUxcLyqqH/hPy1RWFiLlz5j2Nv4/GKpYDfT/3PBS0nTYHI8/rIA4CUe+k
578rAlb2JgE8G4Hwup4gbVBy903WhfByNBxgj0wu9zIAuwNq6ukVd5TFZkmeTQ3PLijZoOYYWHFh
jdV0YMhZUHBa1z8S5BQ2aPT3JM8gFchgMrPQpbPAnjWWBnm9KRZtU1h0OF2TLlmXrbuXD3UpAWLJ
QgHCQHNH/jBwmFhMHGbX7EHLtsGDmm+GsyWawWs0mqN5ysTE9MN55V9O/fLuObGRxWl+ROZTFCjP
pAPX/7c53i4l6aw5SZiDIKXuG2DtpgivQUYoYZMl146GWc8qhyBNugilYBeuomSgPRZZsuQt8EEo
8TjDWPjQmV7U8b7nh/kD24XjIX+wXbApVydKQ9da0AdtTNUaSneNUVvmDniZs7uiYKoyCQlTQ2cr
v5nsNZCbBkcAJBbxOMW6aFmVew1dQjS6obKOB2HzLKvstIyrr1DhlGwoH5+MTjIrhnLSo1ahC+oS
R3ACI2xu71zEauP+41IL08yCdKOtRrKUOT360PsoDzPEX7eBWmRy9CKLZtyCEEbWhLJrBCjwD25v
YXvEz1XEZoAcKgTb6NSOhwuBV+7s4RalCHuq5eM2ANzLYxhXEJb31jGo8cQOqM3c9hQ983uvpAc9
JvXCxmOTKkEhKxpTlGtH2g+LNcax49g1fj2hGxYAGSVmUSDYFsZNgrzduClAhDJ6cnGfM0URHEjm
QICyq4CmG5Rmsw0YfgN21dThiTsvN6rIUKQHIrdCgZTXWKH+R3sEIvV9YN8D9qAUL3d9wGXEezTY
jPHCtjh/AkfuXGCDKVDQzRO1jzTiOafF2l4xn89hCpaoG6SY4p91u6EheKtL1nQJbbvf6WRwsich
caSH8LQVK80j+y7cgD5I8yeBVMG2yLUTm+okCyCmsfkviJumx+dKYJcGXmr2CPVp5r5PLTwwHSwz
P+/kbzw53BqQPsVO/Ot17Y+h1ZK5S3xxz0Pyl48lhMZXUPmqcQZ8XkoDB/0i+Ja+aTKVPUDUAQd0
yGJLPtspL/JZZuzmbKegdfhjdy5oEvzEyqYtLiZukQYlmqkVZ+2QD8WxVgWirftjd+9eZTZvtfE2
DE+duN9w9tuiNFjLnSdsTBAkG+F2f7RrpeyQMbpRSpdzw0XeCazWiq25eiV/B7kE0j7kTIovJbet
qeyYmznAgIHBDsUou47m+fGK64jBNGehFAEq6u5OrPxjcinydH7cAIVbp6DP9Wvekn7NkJoKJQfc
b42WmvOPbyRiz0CXsiYTusaVauuxNrTJP8aIKu84pRrPCucRFLveGVrTr+GlGmqI6OXqB44GbenN
BsSdmROkI4AXpc5+iAXxhLleawvW4AfI/dXB/ncJ9AXFSoJKHsr6EhQ/2UE2I0G5YtuVc4bdFQGj
txF+g3MyNzbLkp++eKnv1knBDsnoIC64yTHBKV9WszYiZZSuLXqhur1N8y9MlOtRtwTkl5EJRmg7
svsVawGb0+wrvCT+sgeJZIHdJtBQV+rI+d5BR/TT7L81hsh3UNJ5fQ3brAtR+wHGuvcuWtSZoPip
QAzPn0JABpS2kE4RSfvg1nvHU6jxYzEFe/2nH9RoRZLBCA/hJMplEcc1DlPFrdemGmrmmbJfv9yO
gE8L5BsYRBecDNGdGlQRr9eUy0Td+qlH2F7p/dI4oWGWBHpYArl2/Tp/vun1RrwOZ7qbdNw/ICc9
jm/xflfXoqz1qUHXbwXwcYYexyXcgjrmB6MkzsiRVJ9RyXcktVJz3hbMIJLMq3dwKWaj5VQG4JZu
lEVq61HOu+dLy4LFZU5LDYUeKqcwQamwNbhZrJr8lnjgXFkqWOwS+ly5jkZDBHnbgoaIfTvpYCys
+PCq3bGg0ijNtfeLP8u87wKenPzB0IEvCcwVQaGNsPG9fxwLMgUcXu9BDkE8qtlY5NabSfyaaGn8
nxRs2nsHShKj8fhBj7G3gwuDzuQO7rAlL0cg3T0pqfZ7Ifq6nn25xxxYNSSQSqzINyEJqAUtoDV8
Pal0aWjGnRjGUO/fFeZ+mRR/5IEJwUWU6N2sktRJcGA0+/Ktjtt+fF/3b3ztOgOuBium+2/8HCSc
+EBH0mLchhFIGMfpTX7J52Jrx41gGISNNvQAwy3t+i1L/kTkBzEbtWeuL42Yxr5uOv33in6vzTGY
SXgUInXO93EGh4Vmw87M5K/MWl+XnP3cOZbT4dhceIkGv3hOF+hJRc3wF9Cj4x6945awrR43fVfJ
y2DtZzyyHSRve+MqZV83/TIikXjC5YlqAg49g+CGFWP075qlDrwktxtFlzQYT05UBMD6Gz/wmPBi
H7Gx/pl7mWFtOYbASzNf+ymbSRRA9VgjTeS8fvqTWCbdkED2asxeWtM4iPwQSVeDvgGw4CiPR7E6
r5MwUxlv+i3V2VoCqlHbXOxlwwk6aNIiYtA2gctLGCJvUsu7r0YUnuW5F2YZaoJ4PftdYsFWnjZ/
QsZe7hRx214Qfrr+B5ugkbaTSo1AQ0QQPrkVL6UUrC5BveMPVo8yoam2TZ2YN4/KyrKB+GOJdSrR
S4XzXKX3Qjm/LfuP+J6nN8Gnz9pQ646tAs46gnItHEblmsl1AlaJidy9SxNDdAjkm2wID9/gAKaq
sV1uUKOUyOYjFFIQYxJ0CPDHH4evOaeddkoWiAtenkjQZHeAac/yhxOklC9cdGSFJTdDgNfOcg/x
bN6wzmlZUzxtrSIfYjz7N+eIlotnySGV5fpWAwVTv1mpoNLIYSd05w+vdvPo3SZubTtCQslNZJRW
wBXko+bO/ANm8hv0M4qH9CEJkuAT3B5iMu/TNnJKBlEIXb3qrKtpBzEOr2cIkMMqhhfMCKQvoh0c
9sT/8Mhp+2d5qo+3YMX/NNX3w6iuC0g2bpy6kYYnLpuIg5wv2raj7pdXxbOc4OCExkZ+h/93ynQ3
TF8qzTv2aCo0DimuALUWzkj6vmi0Lxpmz5fqp0rLisgGDLUY8VZobny5LvxyZqZ+99MaoMte4TZ+
yR3OjcR0NKnv7GKB2c6TXwvXYn6na0FVV+KrrRwcpIWbw8I3sAssQFzda4fOC0/cHgYqRiZh1FRy
rI82IDLSp+dM0jtFQywfzsvvLQtL4nxrsmm+DFehbXkyV6jSmPNXs1v7WJTc8fhD99IvQZn4sxAK
8WERlQxqQorRg7nqbod+0ytuZn0iwJMWB4x8sZV0LV15NXPyGmIlgdm7cSvyMA+O38qvk4pronpa
p9OAfD13dgGUHPFoq1SxB3k0MuK1N+iOWY9zLBPtor9zndmxTHDa2Li56KSniN3tgL80a+IhD6UU
r6obrdyTetcwb0ZhbOw01N8keBKGOJv7V9X5OnG15L6r1MptOLdMtNU+DXCNhlV7OlSjYkHaHo6p
xhrhNTialikesv0BEbkLElW5zInpmTC/o85d5kJEsQBxm16qQ0oXoo001Pirw2Rwb1RSpXBZOF+x
a5+vYZ4pItOg3iArFKcAbYg/V62B913sIRIajo0c4mxe9Ys4JjSMRgdXiiCXqD/donibc8gYtMNg
ZyWaNzAKiakhLFN2SYj8urrgrM6Y4+WgIxeAZ+OTKWoNJjP8ZklR7pfjgXBWS1eIQEX0QkKgMbGf
3PcTmXjeuyj5OEknQfropJqG9p2mWrVW1F4yoM7NhfTPEohL/AxuDZwsWJuLGHt8AZTOY7wenqJA
s5KIv4lGYTQD6yDXXznQyrNI0uCGY3+pLoTH1tGp4lVkgO86rIjEreUW4tYMydtJxIY1qawmN2Fd
dNyqd0pDmRyJzjgv8Zx4Zjg1PhcqrHztsoYp6miraGVYxeEbCnOsuDDNrD588VBnyR/KExzivojh
9xtgC7rTc9SVGQWcTP/uvCRIDnMPuWwj+0iGWG1KZ6gHqwPYKWHAcEagxkldNlQbVTzu6+qJjWtd
EXxHccnY1nLVkONpvJBRxqXKpPvlB4zqPNvnF1pjeeBlfX23dtVAK20ikIWFepou/JA5FMJhfe6P
OVCuBR/y0tuwPSVkb+j1GOWGq1UVvcKPbRadF5neU+6ArvwStUVDozZk5ZWhejRsTY7h45G/xteX
AYLfgEYY0cGfPFF81/I0KnRuHtmehVeNnABjTZUepK+rf6f5+LnbAfIuaLAl8xPr9Oge2rxD8n8B
bVDfO47pJ9H2p1qGbTDq218fiLVS2+lergKUnLSYqSM/wjcpDGUEifoWxOsuHK9I76GTdyq1upMk
cOsAUAKYVRpjmbRJzN0+EEPic8MjMkIsMYDsD8HnW1JggB1MN2O6h6Z566kelU/+Gg2p3nZh+3d/
K5G4ZmRevwNCVN3BI2MIYKUK6vimtdmI2cQAByVSlvC4W1Yy4pMJdku+cFDmRrPF+7BTGliXBeXC
Npl9tmveYujZ+6scD6L9K36IpGJpp+OpnheHWMJzH1Nz0WRN6S2JheiIhqdbFEyD3gQQG5CLUkLY
YoBqnq2V/VFNiizw2YERYiuCAhsJN0xjyZ+yoPqWogybC2o/dSY0cRb7UHoDG83yyMARFNq7HXjX
qE29oKjLugkLYTDuFGGs9FqhyZNN96kRlPnaEpNc1zTg6yvFq+8FhwDoZ2h0ABHo39OiG/kSbiJU
OypoiG944BnZl62pOneOLlodQM657JexGKKnDhtdffZ7beh9HW6o/u63B79nKLblsuqXzjBfIFp2
os2rUcl/mLutiwog/AJs53THrTFvJv7mfI6IPDmrSaAmnYLKu8kIVR+9QhPwsXMucTpXCHD4O4Jq
Q0IU3givIr8ZwzeumMyHl8bJEK7c215/3xPdllGunyq+DyXcskNM5Kp5bV27TgFxSv8tXlN/furx
gqL308F7OZ5lHe6Qc3hlyLs/miptWnbBL42+XlIfT5pjZ0f8iSvcIfCgVeRTGS2vM8OWYL6RT3rP
HDi+EclcezHQPdsF9dp4gTCJ+dDkWcGwiQbUJ50T/+o7ox6O7IrSvHcTKqHNNCz7qbx1k4v+aBBu
mppoc+G/c7zj+4hdjCIHnyAcDQ4yR943M7o+U+L93Bdho0Li/JuchBMWOMqfrnchxWKVO9KVHmR4
4nQXTgAzAGGqHbkbAN078dq+RmLLcfXdmToTP1uVSExD6IHljww1IDxtBiOVHvsG4CAB0+lynXsp
NhZQfLCDI9T7yUFiVhQk1lFurrgVYJKghyFWWxzz5ezoHM0GwKZRt+oKDPoJbt8hr4qctY2bK9sL
9n0DBUytQZXuvF7xRfo8yoeDhDfesiaX6us+O+HviXX4WBAdEcgtrCnt3+OjsWTo/UEgdg/WmRzh
JC5SI/Gy6IePPWG+mA0N8IUqpJIuLr1NYdTe3edA8P2qEglgHcefDCMUcP8tnMkgFVBTp1lxk/zJ
07YGarnVgbqOVUjAJ+jG+siHqvJPmSo2WkwI60Kcbp8qgIlah+mFcvLTpQ6chPg/fYkqazLaSJU0
/dXOwSLauZPA2THm6+QzhpgXtOQeYyYd5qlUSZmImoIaM+zcKYLXc03P1U8IY183DEc9e0hDkr27
0ncP8g8nfYM678hm4zbxkKZ28eJi2E26apEx4wmvYHPSm5iobaZirvAO06+DYlmWJlG3LiooxFop
hBwqhWWba9ES20i1udUjEL59+FtoC+BdTN1KHCPjuQDl8+zr8PjBMKCpfNCnQKUZiNpS5VRx0rdn
HGpGhB6W7UokooJ3HCqhNDPRe+zBfvOt3vEJBIcQgBWF7vpm36AnY3WyMd+6Wc1nKtipZ6Nt/HmE
+gQLfQf1IuLQxpVP3gGR5poqNupiGCNrqc/1m8Za+WDHVgv0qPrtQF7poUTEXzSGHZRVPINMsBDw
EQVHjhdkpCnHUpXsgRCCAILjIAVGZ++ONmbFwuvyYT9n8Oe854CW9nSuVOqwMm/qsT7s+NC+Z+/v
L8S8fRwC2FRHV8Z+8nz2QyUxfsmDiHktKt0NdKPpICcbiQNwspuYFvmZPyXvBZzOAQ2P2aZzwgOe
rVI5rIAkUq/ZDrQNmqrYtFVaq2DqlVe0S+merTEe49a/KBWdWrlTdtUkRiKukB6NRc4AbyN5fMHB
up1Rl6JGiiGHdpLFW48vQmw9jg5B17a7vucVmtpZ6vm4KsaF1tgJKwYvU7OFbq3u+eVK7Ed4aDHy
E0W/Zoy7CXBmXaXkPiTKs91YRC96nckPDhbH5ttp1uPcr1JsG2HiT/1NejuyjVBsgYNFR7BI1ntM
1WiEBKbEtMJuhNskF9QQLYEl5eFzFMJr9aTL/yfYpW/618zdX/fqLI//W/Tu3pmlV0xuENetGCyc
GTssIfq3Yg5HJtvAb4SfCljZkAiF6QYdsxU0HH8urn1t8AFe3y9eNmi0wK4OSSDgyR3wd9ykAIX+
RolLIEoaGRwbnNOo+wQNMjKJ5gKIUYztbe7QNzjiLI45PPvBCRD9v5G+S6t1ARPS8T4w7wqoNjB0
FUr7RY60GjM4g+GA+IbuOQ/b3LimSP/lsoZmANRors7rPIfku3wlNbdtLAtNSs+DhFCEnw49Jnep
HtkVzsSkIjvCzZjiZy9jHDg+VtixOdFsBoFhABIYh4Y/aQJTs3b46ytQ0w1QKph35qd+wuUG4svQ
uKMkY7v5zTQ0g3TQv1amC79ezFSoLZxYZv01J0tJX3oqqEb6f0ZZQuPgIFH9JbmE4Yaka5BBSK5U
GXf9+CagS5FChhx8epmX10LfIBlSs9usLe+AzsUGLhG3Kn/8xWgogxou/C8Bjho5j7vm4M5DBUWH
xIFRcX6vbpyew7TW8xbg8Yf74xOfKiS+0clcQZOFAM90NB+nC5QRHCzn96dmad6dHS9r596RxiI1
LeA7BRyxSQrF/eFhjNbluRhSMg02kIiDEqYDuhF9GGMWlB7SgiXLYlgIO3w7f50rXKT4FZ8v7whu
z6MsmZUpgpixoS+rrWsszhb5WPICLiZEaoJf8vQDJ+9KrHK4hqHEvSKgGqzaB5T3pNOzlyQ3O1W0
VS19HaX1rGjLV0KZ6fcio8bVUT/+0W2J9iWEAfXDdPrVpfw3Ba/IUnZKZq59J2bSYOI7wCV4XtdE
TIedsDn3DvrpLkIl8x+WjGITbqRM6ulnFp+0Yne+nxc6FjxoAhW3I1D6tG6Fnz2hqFitcE4e8a8+
3hJxRoBDEpMh3n43ROvOctVap2wy6BEcwh1wKbe6hJZWzG6oio1qv4EaCneTl3kFtiiqjZMpEK9N
ZIH/7LvHhfttfKpmPPDFBELncujIMt/DYr3Vol+o9MMHirEc5wKe/3doZ0aBWjhLjIprnplq8aZ4
WIqfjfUoqLldgdESUXPgK+N8yq3B7ulTk/JwXgdA9HCadtdkqrwkkZKsAmx4MkEHdozJWq6bU3Jn
EY+ivofSdn7isxfHq6kAdanUyOfbdZtoeEugZpRLM13tc58EQrb0/Hj3+FLGVD4VuoBrkuMRmIJN
hKIUQJ+b8bWqUuA6SkxziHagSPnFzmgUKe2fkY36SmuT01JK9XIZkLewnuUgn7VrJXMhOASq4Pjc
/7S7Rn/HZ71uQbNiDo88XzUet+yMAxtUEcbAP2JBHdehBEBkrLf/h0SWZqVxxtDsMCjcaht2ge02
FOnhOOx+2rnBo9z/hhzRFhILaAuao3r0IWvMhuCgOaNI/50yROjM9DS0p8H1YMrPuJZ1VAF9x/De
n46gVi9xTi86AcVWJ/mcFma9e+YF/DAAVCNaTgbrZ06a9SZD03+XStiRBVbmgAS2tBqGHPYb3EYr
E80aCQvYAAmRm/NUvQyPky8mSZTBvyqhu6uHZgvQXH/Dl1d2UXGRxGENxcz9OOdjGALJkVCq8T4D
Kz/FFo4pkA90wsADU31FAzy+A9cqI1Y+8jqNnJlU5APXf53JCzP0QpPkD4l5orgh0cMTipHdxJwA
qvupggu6PzW7f2BL78yxKDJMY/iRnVI18TSDED3Pm+HywSENSXXLbFk5jmZyhzED3tb2nFNFcZg2
83zxUBO4R8AqAVoYrK4oCTGVmgq4KLJm/+GmxYt1CnQOrRyH/FtHL4XLCKkyJ5jgZbNWtiL1DmzV
BNOtgvZUtWGot7pxuExyQypXNiA3TbKq/6g25TH63rrXWE9G5yn6MxYuDeqKfomIZZToMNn2YzAw
DonCyMJjRrFhlZQaAUDDmt2N9XHziq0Z73iP4Y9SF0x0GWeX779zhYWRZap1KUkiFNBP+QjVj0uG
YdBGxUZ3AxquK3ZEIzy8ItGMWXmosazONtk9xYK/hmNbLFFFezERhybKB4uBaSdPjmmoVvzmrf/C
GRG9boL+oaRxmOesJjH41ln5wFHoIw7HqKs21f63MZVA8aCbIz4F8HeeD7C/lSdHWkwIX5FJ0DDt
R8UlEkx+fUXhkJqrfmFxA5ei1EmqP/UOQOnDXozCoItph0aBBubTEfxiTin64FLF4B0XFHytbOz0
SGlruzXTDDnYzecPWGAGilhyW4c5GXkhj8CyysSZfhy5YlHjQklGAG383Ttr7KUiQEXPmAlCkEEN
p670oKkrK0SQlMDBroZ31s/hyRY3f2Ue0QNE0aph4MPe1Zx9fQPblN2g914Eokts7VU93V4K7uaO
tLjpMaBkpU7Yvx0I3P4FGy4VY8fD4jYG0WVx72rjE67G2nPr11jtMnlRib21S/Gn3IBjlme/eW3V
W2iXbIWs+8QS/5PB85L/YbvP903dCYKsBJZRf+P6iETNnjJjKraNFXS0CYPF0xTgHKnbVi3xyCRQ
mFOc7M8COMCtWavhY/f+2yiXiw/g/iGyp9Yf7hvFFDsFDzICa7p0O8xHKEm5c4JVNgL4lyjbgrYY
vxJ55evFLlgNB6E9cg3dGUzJBrlpT6uWytY++eQyt2qGsamRSppxwdkStEmC2ru1eGmOhyzOi0Fd
B/yDsGHOtcWl2lX58c/oBWhSiB7HT3rz/e3B8OHpKjtL9kRC/J/zHiazhf71pZHgeqkRvRCIzMUc
IWmklLYsUEkTwzPTGvF6cJvMR5vz4umUKDkwBGQfTuF52iiBpQ5g2jcgpLbckw9F2N/ndfgqIns8
XMjD4gJxR6KUREXwzXXpz0lPsXWRhu8qmPK+sXg4ASqooPWeNPn5NoYKtBHBF8NKn71LFOBqmcy5
fBcNKYQLEtwuJ67zLMUELbY4lwDSA8MShoOiNyh5qKnTQsz0EiRK/XlC2zkCtCIehRzZu+AA1HPE
M+yLalHdgVknVU0D6dPUNuCMWSeLPRzO5vm+IDBytWlM9FT8NJLVFo4zIf1sfWZdM0goXu1eNNqz
Sa6VvW+KuimeZ7UnIuRD78SROof/KeQQ6/kiyJBzRX+WxFF1Tu2Zs5LJj0x+wTM6UlsHovgGN4bV
Fm1iq4CHSc+VJ5vQ0MlrVoRf1eQivVQ/UWHzqbzoOkeGruejbXQfibDiXXvF+fEmorFuiL5Rufhj
JCA4kuAKEaeauvwSf1psdigqWyYzpF57M0ebT7GWScl6fZ/lMBPW+IZwoz/F6F2vp15MtS+BJ8kJ
vzNmZfydF3ZV6Xz2JA5jnR2qZ3i2ZsmnR0RD8qgi5TkpSNazbvBzIx4F6WCtsOfSLgoyzBJkNpbo
kewZfklzqQnHKWYN+VlMVh/H3faTxtB7tqyWl67ZpEWRE0RRF8By9i9o5yKjSMg6OqMGRFOOGfUG
r2VCKslPl4JQKXkANY9ht3/wsyObA3pmwK2ouVx6vR9wjggJzHHmJw+EV+ixoS+BkxQWIwJlBeuk
hCPCGx3prBrtJ87UiVfrCe7K2KK32THuKEfKqeIfvnggOnlYcli35XJHeSVkim4rfIOIzgZ5spMo
Ms22xFIdrVwG218dyZ/g9VP9K60DMTCWLrCdtPkwfJvDLlS0lPxLQE0W16JboCnO3CtPX6UThXPX
GDF68/26keAiFR2c9xtePQWw+4HFs6xu3cufZaHyNCjOhNyHkcoq6wInl8RBZY4Y7OXej0qOGAwr
58gI4Raoh4F2L1rct6EtYqIuzMK90nrjiWaTVl7nOp4u9m6ywXdKs69MNhh8EX6SEAz1AYEcEW58
BOMTn+ILc40q74tjWaCrPAUBdiQWEjw2WVtT2eMKsQXK5u73zis+g5NM1w2qe8AbuaU80w4aD01B
MIHbhaA675jB3unh3KpJiePVQp24N4Fz3ZFQ9MVRlHsvDWI4AvAFpuTJY9mWdOCV1mD1uyyRSB47
Ubjl1tTQkYKnBza1U3L0WyZqM/3sh5N3SsJ+GwfM/XbUVkO1N+bDDWs7NOGp4A57XPZUiMQMxA1t
7a7ZMK0yRiNVfbpg7sV0BOxPZoSrnj18j/DqF37yQozHk0dLhHidKTBxt0cl4syCVP3h2kJIwFy4
OZy+IBmlsZh0Ow2kxRYC5TxxyLU9KP2q/kDxPzi8Y0ek3p5N2/3Od0geMAiZ7UXTIbguw+mkiNnW
p+Dt6ASLsjuAJrp5X+7AR+tNkiOoqgVaIZ+nyUE+MhSeEot0CuigNzvkvcEqr7LPvAaRfzK/5J5k
FVf3rujO83wS0bF+iAHxUc6HZf2UKTU2z3Rs0WKThynEQk3BzAGikPAntAmpUerDEQ82uQ1VA0WJ
h11zlsxtnx+cezqe8SkqvWDl7MbusoFbV21odDberFk8M4TXJPklRCQOL53JACD9kRQrFMw3vdco
WjW1fzllBrJOvmS72mbMOu/5WZiHDIbrbcvQC2UfhbGk8WeNoxpPYPP2OyksadDBORxZB53NauPt
PQuDmMeVwIF2CiNx8ivgCZwh42dIjd1w9shrgoF2Fw+vPPHgZUZfoCIM1b4ac3sCFfSUGOmr9CvY
3W/Fx3Rfq64+MjE43yYUg86LFyWTNRDjD2ZRgMp2wn5PM4I5hUW9X5T0vy1EXSLTR5uNCrxhazYI
MvXJUCFRaciY14ur6+IlASFF3tYuHftC5u0Mx4lzS2uWiRqeJdh/Tqob3RbZex26pVeAv4CUYnvC
LmK34BCfNKoUMvhUImElqFajE+5FxRlzfhSxheoQJvLCDQz4JGSvd0Z2QW5BWL4gxpBV1kSNtqem
+A8p2nWX4kAAQceqZfwknh6MYUDL+zZZnE0BgSc/LSam7/ofeHRUgZA7Zt6vvhtYVhG+dyKEZtBL
0ussPxFZOXw+n2pSwt32/zsJ0v7w7layeGw+f+Ao9NM+JEfjyalDr9xKywAFHa5SYU8urmkBZVY5
9xvvvhC+aiIwaEVl82QME5OCaJ3jVWRH+1nbJUqXsa5fc1KdqEAc+qJcJJ9jx3E/y8cNY11xY+ul
C6F6n4ZWLlE1acACJxg6Xk0lf2A7Ca619sHxsNesoPjCjIvlNhbSGsP5hhOqChMoX70y/QQa1dd/
SGM3zki4pmL4ACrgksiMbArOFpKIwr3+ou/QOiE5kwih3afcg6tNxJ61glJKiF0jFZAhOQr5zLXs
i+CNrBgGwvvY4DLJEZbLl8b/kYqDpMUTNl+HQ5uBdig0uwQQFqe3NoSaIKw81jofOP8I7ShPweu4
Blx3m4/OLaWX/mMKxANsUNLknlq9ppc8c0/0+jzT16+GZASO92XrBetEc2zmci+2hB+X7zUSKNKo
p2cB3pp+x7FMVvZTSKBt9VCvnZakWYrG5UR/lPTfUqq+pMiw3alPPyYnxOuv82CGHiR5ZGkoMIJ6
0WZvrnh+WAjaGRkYj9Wv1pMg0x9/DqA0Wzu5pcbaTbz0CEGdfhuvAzgWCvQLmkwlMRRT9YacdJib
UqDnNnTkeptSEX4ikwsSJw5zljQAxe3z9Bn4Hqc9QY8OwQNK0mBR+Wu1kouRxxKIA272Tnhon/OB
RpwJRGUyMHisB0L67ObyuJbBrI+F39nnYRepFmdLZMsRgnrLB01ULGCrklDz/ADjJ48sTAHQOPk8
KG0LQFjdfgNvPIB9kpg07DmPt7mgmeKcHTElVLp8DHqKsJb6dSUDwEDtCyLDWy21E6fP/fyr9rXK
ZJH/CFUulci2mKJjbeL2bRyxDa58p2pP1TXcgxscnQQOq3FT4H7gvf8tvwYA/egsy6XwOtoNkMs1
Z1PNPwU1G0R0lsnRkePlLqOWLf/Xvt0MXsU1Pg/AuOKygJanDY0YGpJABGLbw1gjTYgZATELxf+O
Ncjx2/rFlranXIRIYM5KqRDoEKi3K2skBlIkJxpRLOFbZU6V0leUTBSaZIIVTt8Hl9ApWk1mzaYG
zRFKx5f+zYET4hOwaSePuMWYwP6ElRUM3U1QEWMHutiN0nELo9SoPSjKUl+vHyzUpJsGYMVC4n0U
s1kBaWwmmHU1HNpXfii9MhtrUKsdfW90ZChAn5OrlnHtTNCwt23RbrdN7wszd5UTEuVLRhPSvCs/
y3fZC2WbHFGP9EyYwSW+v/jm8eVeY6woWtRCFeihrZMSUZE2LsWI4iF/c8AW03gc0/7xijufKgnE
kTUArdeC1IZN8Xrqxj8zTHF0WpPI9jaYfai60P4HJdQSMWK1x6YwSv+tGDLJCcLcdrRLiEE6A4uu
77b+4ctnLiqsCWt+aCK4CGzJ+syXRuuv916xwmBdvYVt8RW6keL4HEPakC0QzuA3YXxuAROI0JpL
rndwuS0KGWk4r7kTY7BBf9CEIQjzr5WSx+AEfQfEYFahALH1niPRkZB6E4U5yCVtU1VnBqcIN1mg
uj714yPSJlz5ZK5GYEfMQ4HvwWIoeeF52Uc24TQ1Xetq9CdJGjtddq1mG9hY6UiIdSy5OO4PtMpD
cqmV6BnfVSg5x4BFdkTHev1aSgJ1D8CYc17ciuFgdDLXiDQQ9AUZXol9vfPSw28+5sdAJiCFI3U9
F4ag/28PPiqnno7S8cbI9X/MxKkpLFQpiL/vhAjNW9ZjzRYLpEcSuIdgfryJT9qkLe+tVyjwaIOW
6Rys1CqQFHMRIklIkULjTMEFPBpce2dnmDbl+k5iQgyuvyGLay3jmnHuzhDtGw06eALmM7qU8Psy
44g4gI8vxcRyK//5vbbclMUpbd6m8LKFj0QsbU0/SXW2XIYvDF0Dt44f2VhQzXy5zdlKMpsBkQ8V
LfBUX83EGdswescUpt99lrTD7eIm5gu257yiEqDEEI8faXYW5c3WkpgjqzPVQ91A07ORhYi/9EvF
50d6KlAxIB9R5XXLVGDv/v1IM/enTpSeEhSSDMXRKbM6wT0Zo4GAnQNX3hgi52/dDJTc7UpWw3Xj
jynyADh50J8GJByrG4FTYnd8uQ7BUl39dEIHMETzXeSfD1EskVRY3FGvlEINFZox68PsRMERdYmb
c2lJLSRKYnHQSjmdjhGnlPgwJ2EkKLCyErSKlv205Fkb7ggQuXNPhKrMDZd5pbe34Qkgkm206OMh
uAjprICMkLmff6h/kOeUPvKfNv1ycafu/OUDeIjuSGRalYvW/vJ6up0bZa5uDwRtwanGYe0ObBww
kn92ZwT75lkbOsMPlSmSrXv5FJeTwQt+de020le78FRIp7ZvR4kHoF/zHkdiVZgBigDmB6FMUxB0
sR2SKSjnAkO+bXg16db1d/j3PYM9iPBOmsSjxKXP7WzGoTsqSJgs8+dZhz+05bNexSLZrtVinR9v
QtwV/9RfCBtUc9TD13hCIJ2X+5zJGljx5TdFN21MeG6CyJgRt3LmM0Qm9vjxKCem6lwE3P41dKZW
J1WKRHgDgFhaHQSb2NhdwJoYp9N2E974w7lLjA1WxEwyaL9hUqTeGr3ui9j62fiNN6BMwO8dVzyK
GIMHAKC2RKHXPk7FR3+X1PAExwqepuvCKCF5/EFPMMshIzrSRtLWCB2za9VcgrXUp9OvXXLOp3nY
QMD95GAjKyR4/9d2vHiLDhyfdLmUCgYXbP5QxXAlKAxq3ndjblie1rMG1Bd2z+pwq1Pk6VDylgeB
CcK76yaTjctonHBMGfGtbQwdealTuod555eECbcj1g4qZHp6yK8Vnz/5mufBvvMuvuxpOJUObU4q
74pgW3bYiycwb2xBZrHfN9cqCZrzAOMXgS0ROrkgx6cDtuHvn/2GIbX0jjDbQ1MKmp66eOXomJHK
a3kJmof3ZvzYbD0TeK2om/ipdrJwhseZx6bcKNdavi7zbbdbcL4Nk8M2SGrOVrW+May1yAEuEIpr
zPr8MtLtDIjnarH10EU/+RuDD5FVYsTLUUHGRjTzcL68MW04XUcmR2CRcXwE5kYOPJAsWGETZCaH
m4PfWR3Du0bidhvH8Ustne90lVJVZxz0e+2PgbIpoUvE6CnLB2iCADvo1xhQ6JGwhj6UcC1oYawX
uDsJBQkQ0An7hIvsawNtTCpUWA0BN0LWmadBF5MjKeeL9HhHQKUhOOaP4c7Uh8XZmcQ0Wp+hkNkr
4SzllOj4YCP8U24nmuWVhmkjdqzL49PJvakoOK7WzIixDDVvFz6tdq3YkvOqI6GmdHvxsoOl9uEX
AnTTiZY/4C4G31RLf+UaxZgmibDJfMvY5pBICJeHF6TbHkqoHvMJzgJzcL9uzoKBzIHjmgW4R2Cb
yRKZccWaWVlVUcxZdKy+6vp/FmKesF5xlNBQO7A5fP4ssFIVxVDNLNBx4qNowJyLILbulwnLXIqo
77ePn0+G5n2x26Gs6sTq5OzT/ZDAh6N9ii6RpLteIbOJUy4KhTD6qId7+wQmnUZVN8KBdqvNoPz+
8VOy2hwlW1c1yHY/aRICFF1Rmc0dE92u2ufL/TQrimwv8oCNAQ6BONTEW9wV8LaCfJclheWxroXk
s9Kcxyyrp5yu0UQkbC6zxjrvzr67EKI1ACVoQPnCwnokKp+FdwObjrhkdSDasGbtUptStTVzCLoP
TxBcMCna+jWFxlfJxhip6L7e+q8yKDglMlVJ4nsjk1uCkENjvPejR2Nh46XNPGoBFlXhtc4MZsRw
9aVn4tpxJwmZ5NNoE7hjGvIhKPWajqBtMgPUnoDuSlsAuS/uh0ZQ9AqEQiQIqDoSUKKQHa9NsIDf
nd6LGWB3wv8la35RPhYifNvQ796SlTnl933h8dfBrA/ZdHLRB4fE7/xymozDxwXHT7luVH8FysWV
1REUpdDuwBQSnATk+UPGl3OzfHSnruqnM1iCUuGOyBYA2FM54HGR/tQmUDA1Gxmnx6VtITGj8NO8
4umnQXdbndbWBJwTSdItv0mu0YzFo1lXF4ROW0J0Aetq1+uzmalGYSkgmVrzMvaJCyFjOERKrYzI
yFIicQw/UFg1Xi5rjoGpZjWnnYvTqDGbHXjxAdjgnzXgDQQJZJMdBxJHjCymYdVOvMGz7HpUiagO
THWSmrMRT+6y2iMmRkVbzjPKdBlvV1OZKFWnwwkiKgP1jETPREPddl+XgCzEyqN93onLrkwWxe1D
lECJ42aMMLiBW1uvGvZImcUbjvOIztUdcORncYvSnbEmmNV5PtSifeUHpV9MCfeCU5aeJV4Z6Ri1
V6Mmj+SXz2/++sRny36ITPT5ID2KX0ux7FewkVS09V8+Dc3qw5HREOmuQYH3/6Qr6rGw+FDPun/E
irrYE2xYsz/Qc7zYKbiQqTAQOyL2GBX+TBpBAGYiJS6fyI0DqtYnOEWNXK4kQC9RBRV5TZuP3lXZ
9f2hLR5e4tckRj2zNn2Z71YfI8G43n9q6uXmuARMP/nH2WPb/nXjldB2uZ9tIImvQl/w4EVG2n/L
/vYU+28/Xk4sCyLeuGiZZ3enw5ezbupRG/ovV6jbbikcKS/JcI/9/be3xe+G/g1nVFFHQJGM5IIt
s4jmDHbt9/XqthpFFMHazhDshlKdFGpRmQVrGZFpuaYaczcy0bwGQByd4/Yzb0P0RV1DToTw+Wtz
nnWF0z8bN3TmjIgbsGe/q7Dgwi6/0E2qzr0tlhz6z03k5lqr1yIZNwy8MnwaNy1YOHmfpPd4lRqj
RisSgFGCDf8fiFSozqM3rdD2YPxlpQQ62qrs9BMNPi8wmQM68qngnppu2lwHDL4YyKbAd3gZVLfI
IxSROerC/m5xAjUkhmi7MVW1WGDiI3dasCw6pIN6DfhatJBv7oEHwncnx5NsuefpfAdnXvfkQo+C
VDlf29MUMYiX2Jmj35Vx4PFEWkOMgD+omtQuQcorMuWTiDxdyrBidVtur7hpIZ1wOCAR9hXztPMV
cnTQpmKyltTwKecJJvvTOn/FLDVrkMQWprPQB4DWbyFjiNaDAopJ41BSXE5dxcY/aFKZrsl8FDTk
hLaEeJN+QbDSmBPB62Z8wq1fpaMfD1qcogpockTfenVxQrYvnfKeV6BwlXyjW9fAOkRNeooAJy9a
sLLNUT8AF8qpSQLKV1cRDXHMhHO+x2gGef5Yirau+Q52tt3nS3S1UwcWVf33Lym1jTLmDP/+/EtG
KXtMda0CQVVYLHsOH5J38l3dAdivEuyLm66n0IhB3icVZggRtgZd+OslkNwZDSAQTYHAgsPy1IP9
B3rgDacodfSvsK92xrk+1OxbmyzkpACohLP8I0JHEEuedIUP/vy4BW3/1FMlTN710bM6o5CjHhnq
HBYw2ZRH7lSmvFGYQHai401IUzgvS+gX5r75Vn/xOjmzF6Q9L2zFwZ0ed4r53ykQrQ4JbDhuJ6ui
uinstpkCvOnLqLDh61oOxTC8XEWKYOSaNQXxZ07QzarbGTX9y48YXqX230AINDCpqRIZIzTpx/MY
W1E9OmDWkFZuLAJ7xs5ZD8QIwABVMeC6vIi95kDjgBaNk2vPHOSslwrBpHyZZ1HHYTXDXeZKJiAz
cN5GgTz3MDCusaRyH6xZAZ7fVxcTFpsc82x4ZBWuuXeDWPbC5uI3eGaBXEJ3lcWw9lnY234ib7K9
VVx0VJ9d1CW85JVUkwitjS883FnFQeMzr4wLdOEZe2mO/GhW9LlFYIAM8+ks7Q2iDYRKOSdxSAaA
Mzetx/QZX0I6+UNb6bk2T+R4fXM9kJPnz99BBoNyBzFgEFu67i5TkXEZtnxXO+geqB4puKkEpMAD
PVQmJItx84uZBw7qZJHARW65OxPKmKqovQDFMi05Khh3S3pALS9o1gzTawfrNt2LreM+cUXPzdlZ
TImMhPqFwxif9uLM28/0uEEnSnZfTeOCVQp4xikXEUxwPgmutifkxseqndX1vgZQCJPYYseDEVPo
3Spkus7A6e/5Wscksf59kWNuc/1Kz/QtfhtUii59N7QuRCoNULG717jYPUA3eiEskma/hJ5nTbTl
9dOcxY3J1aAhZHcdDxa2J0roGwB8qYw1JpKC9nl5GeCd46zIHiBRLZ3ZKMB1kY00nhxvjX81QOqu
8EQV842xnJpgOnrc6HLjtOE2ah72Pf6ErEXVgTj8kJBczTIah7PgxHnaVkqV7sz7Q08NNKyxHPFC
/Moq8YBj+IDE6iUryFzYKOk1TvmtmmP6lYgx3k/NvVjnQII2AJ+SkedIMIP05ylqo+vU5OW5dj9d
JLhsiWH6L3JlubTgaCzQKdTo1UZHpuYRacTehvLwHGkoFYi+uR8NPE3jpLR75PXSfsOg0/NYUmwW
FA1tmQEaA6g9rgP9a4f1UVkwLUE0Uv5/v5dnZwDu9gzCOmr2o2zSY4IYyovTTjxgyBcw3pmelKLr
Y16MVuLhk43OiSIJ4qz+/8m2rzTYFcOf5kv4/U0Pk8CJirfIdXr7jzX/jLrQoABDMiMQ9MhCrhjM
Q+KuF8vowahqTrQs5Dlm+e7l9743fdc3qLgCgMPLV6puGxJrWqC6bOqZ+cSL0/NOeRvEJqfHTWUV
Oc4FJXxZWQh1vbZwrzDwCjGOv2ygIm2Ixd6LFW0UenuX418jkHD5DC/0DZ6m+ne8UTzwzn7VM3p0
S0LfHJiy+v7nBXe31z8TelSTTT1DIKvfJTBh2w5OgZdJlRT1aMLkFgLTP5I9TWzZMzL7z17qxOie
x+F+RfMd81wZroPWVKccb4bBWz83hK9R5T7BwGtCsbh9I0dP8VDIKn54w72xLBG8QVEqPXVRELel
BYD+n5BwwlkK0Xr6Ziwp29b9KvDw8LSUAKltWcxnBKL475boxA/zi1pIHuCS6OLHK3GzcS5jMFXb
sGV9IllS69IA2EqdAq12cUXlCTCxYq4P9N3p3ZD1vHDBUFkqUG2guZ5as09HfXWkdNn7v0lyz9kN
EYk4nHmIFBctU0Cpvm0sisHpSEcXK2l3CdOJ22DiNf5jbje5CYlaRFhNDLRyEp1k+0vAo5FHR+tR
dPYIoK6A/Cqhewcf4ynTkK6R5Ir8QvUPoHY8tGFDeDqLkB50byp4FHDT/+KdO/hgBiTJZrKV25I1
gWNqpvl30nXp+NXUpJS0ug6gMTfitf2sq9nyr6sTGy9uHOIvITelgkZsUr4hIXW/71AqMx42u7Oo
em6jgB1aMsfMjAKSY6do0QCle7Z84yhF/gnl1xl4oOmAEmT9sWg5vpNr6OxP0sVhyuRyRKwZczUP
aV0pMXu42QwVuhonyPqN72cqOtJ51mxtVrjtK6xvj1kxgvbtC89RO05a1n2ZtGgqTsR2zCx/Zuql
4JLzsIq0l6x1nLhepMpiui7JCtOElZIy6fE2WlyXD7RNaPb+hZfU131B4L7VYyuq/LUhzE2T9wfu
yEiVRf4aPsmhriqQ55fpsfpSw5cE6qjtQ3R7jUDIlhi3kF3jvv65zHTbwLUobrBrATxiz/dAWNeV
27rBc03+341NXwgJAnrqpPtGtFQLmnlfQoQhErtoSQPWdUuh5iY5NVfcr3QYkD/7uI5PELsao6qO
6hzuruP2TtPbzrViScmp+AUsFsWUBs317M0RKG4S5opwyvGjvM83VIcb0xDj8AS+aZlC8IJexmhp
1EHnmCSSfirO79JvZgroyZhmMxi2eHvnzLlexv/E3XMa5KYsEChmOGxwxEKo/5NLsHrf5m8a2a9/
bc8gwARR3vbAbiV4zpcsc3fsuWzB8pEW4sQSbbBWiNTgnD+Df3ml6ttzVwPHaPI0EQpzlSrmAiPj
BSVu31KZj8Zli95ybOm7n7U5ErrjxRwhzExk1h79pLMoDfIqwH4AjnAi0pAJJi1ju6vlctCKVwnU
RsEcVeF7uEAaOqJ+a1/yzEc+3z0zeXWAyOQjDwojfbRT/cHbDpB5P6r3q4MpIhaiFpEH57uKpOfB
uoUnFNds2qbeNDazj0Mnjjl/Pf7i22ZdkUgnnpnqsdHPPqZCkUj6lgn6w8jQEfcq9z2Mm88Shys4
SGR95Bj7wc/QR6IQOkoKoCRL2fGKSCo6mdv/FWlyVqsIIvYvVg5/AWRKX+EXvnswbx+855Lhk56O
BO2qyqts1xTpgh02XDB45b3/pdPaqJH+4580qNjtxZinx7PmbrDJ2W7pZOB6bH5fOiGoJDaGkHsg
MYi7BX4kPaUdQ2zUysSERWq78U8avdHtZVUuZZCaLEomHsXBrgPKE211FU8jXUBuSg2ELd0Rhc+W
jMmp6BHS1c1D2zCxbShG4Qv1NQDDLDsBIzwoMxlsKQgwYCx6W944aWZRTyK8t0I3roYwmLWfam/M
F/QW9q0h5+zqkEOvGqigRNWf47S75q+USbPGUECoRFjuvO8fljnwqkgLKNopg0peG5WOFjY0GEYb
FT9NKD69PtWv4q0lZBEEMSQbo5hAGoxEfU3f9wbQmSbnPqhnSEveP84h76LA44WQHSJPdvN8lHaQ
EKWg0oBLdRlohsPeLmn1GLalBAZR/xHaIrEPj2foM1lVtwzN8Xe3wbHWn15aCThHeeR8HOylOvHU
7TbBlsqVzPmiwiR+CcOzFPqXVUBRPp39gfJgeFaPPc5ga/g/GVqXETvv36dlOt9edTCEinzz9ALE
TZwU+fzhG/LMky0YRSFT07ssLkUdWtGAkkS4qI+Rm/AxVRK6WzQcNFnLGuWXX4g6ifU7OCRs7Hb5
B5q8ehLOLyYfCL60pZ800ghmBVM4BdsxBk+tiYOT7G+89DQ0bYIPHCzuVc8hxWwhhKaMweO2ZjqR
9S3oTTY/3sFv/1IRc8nCvQzyu95/r0gltjLTTpCMUfsQzCozNX0JDT+nXZQNxI6F1/aLT1qyOKyH
mVHaEIExlUrZShqBOCtI/bO+pKc/wtcT2XGf1/lvH4Yhi+wcA4Fglxou3FhJeo3/YmC5DAJ5Oz5m
GVatxPXcSyEpgWp2X1E7IhmBe0n4PtgnY04UkgwJvWG9yeHPmMjtWtKvWhWtzz7e49x2G9whEOAU
hSurl2kqG5EP+v3QDS6nmeCPQRQAWU+6NX6rFKf55qwYwREvkIo0BguAIsfIc2prVsjWELsjKo6F
4Q0lz/cJ57zn+iuszR9YkSaid+IDts0X6tvcs/j5cSaBJA8Nn5wAReKcaDTcsNx6DEyTV25cembY
t5r1lUw6FuLLTvfEBLIC1HQlxskoJVVsL0oHSe8E+VdwIDtumEcu2NYtAM6pJNh8Y+5cTVbeUIWf
XZiABezBRfRMDi9TZkWCCcHe8k4UueK/qAHwrpT5VDm24aFRW6lsRFfHcM28vy4Ct0rN4Pt9/L0P
Lc7kxdM6dF909tLyk/oBC5YfJmnI4p7QrNDpLOpS9/U4t/AOikhwxgtuPWINr3srWHj4lz01uHco
eggNcpUen9bugY805iOQ5GRDk/iT5Aem448g9Z8VYR4/VrWI4/K50vJM/85P2rigcMziO0QflKvf
XZzEInFcMhTRqcUGel4ldiBxAg57Myw9JW7BVvztcLS28VVkk6bKAcjuOz4P7MSh9pmQWJELveaG
C+gLLiPzyxHGqSw4NxEpMegWS/up0tE0uhwgsBgUXuM00148D/OovjmBurKmJ58kIXtWbSgT2a/N
w9SLmF4mitY52yOPi/XVlxcxYbgml5ZgEjBUYEgCNe5P21IIawoJHlQzuiMNYgKJqx3H7jXT4rBj
TGvbx+ycHn9VFN+d4lvpZOLBCbu+8rCdmUswKbLm1QIw4vm/fEP/UNKJf4fGSMx1mpdnUMhvTsm1
VKSRtEwPPMgQY+ZfBsAaOWJBHQoM+wHzH7GoloHY5zwqn1157Aa2d0q9sRFeXwqLAXDCKrD60r0M
xB0/gsRYNjIQwNfE3C6c7erOb6xiKGgJSIn8/R9nEqM6Dn1yoUu/6MjPXQXOaNSUUYwGKrilLME7
dfYYddvBwElQALeHexwhZRLCCWMYirLNZGedVDn4CydhT22i0o6kL/iWtEhvKVV41+dCZqjzHkw3
BUpodc/zZRR6h2Pg9/gO5seM3/dUa1NTCLTNCokmGtpad2YU6hTW8bDkNgbaXkRgDjGLQVD/mvQK
80D5rqiRCVKzZDzNMtnWlnez+OR4GeQLkW26n13TX1PIV3ECV4o0OX0ukBzNT3hADy5Z8DJNzIP7
dFaz6Cqpj0+Xeqnag7Vqu/w29pG5ryhWELgkyuxe2lHXJYi3J8yOVu+BiGoPopK+CvkNScv3GhDQ
nQnI7WkY1KmS84PuIt67O4xuSHslgx/nRJ3IXFzH8pHMMA5jNC8TUrWQZJueP+U8c0D8tsHeZ8ou
SBUUj+IjVoQAwMLU/stoP6P5j+UR6ChaMf02NcEwx3Aus4IrKotY29Kq884gl68QYgbD+QV6oAxK
i2s001L6AKRFKjtnw2w6tqMFOaKo4HWleTvuNCvkC1TqT7FZwigRXbI9UBNhS87/tf6TWurggk3g
VI+LM1sKNr67ehwuey5NGeqlfOOm4TRwa21qyLR9xPATavY/VtAT9W+HbV2bCFchFgmnvxVMep39
fpApBHeo0Brw6gnYYC3JL+3fWEPPusP8Qy2k1Ci7jGbVB8A6s8INjqwG2W2aGpH0IfWmqsVxRqJB
Uvc7L/nlusPWHCWaymhRvgY0c5oP61jiVMtnr76Y7FlnAr6R+Y/MJvp7YBPA+6QURNunavG9MFQV
FqmSWU3/CaND1Zq2OVjuityroyepUDMcI58JtJWe+MKTUXdIO2KNkiinjftMAbDivRz2DrCqwbYv
1IaWCrJliwFBHetZa3M78zghxlw9SFTynnOniQ74aInjJvu1sHNArNVQx8i0BOI2c1VmwG7VZFAX
5fDCdgmVyAf3a4XJSUpYqZpe3l7ceM89jNjBmfmSr+ChoPce9zXApL65VvGi4hElkgKCX4YixFR+
FeGfBUVt9mL5myKrvU6PXQpAonA3OPMqmb7kSjNrCBAXLtJUSoJMVosganH9TE52TF+gcfFTavLt
LojBwxz0Ub3DuvBs2F9DDAnm5ulfWEcJzaHRpRs1HG/vIt7iceC1MbG0AXgcRWYKuNp82j/jYWVz
GXv6118w8Y0e8hiZi0mQ+STG4EQ2b5+OeuZ2Wu2OcDl8dhKMhWp8uohAGU1DS10rhT35RG6tNUau
XT4brsXAbrsxmHsZCmi1S10+ykiFKvRJNL0GoqFJFPRgwTSrJHANXP4LxrEyB1Vjf2jmG4sEQTJe
+r0SoIgwNzlrcHjKjcuzxCiH3Q4mWqX0QVGgnpggLRXYH5mhE0kIcBn/TxtRfnWJrsTZtZRXui/a
zWV7/r42RopSRZni+SgP1Djt8bfhyYMLi10HdXEmkP239xbF1FzUEXGndOCQpHmlYTOxp46aK9Hm
eGmhQtGhGJl3lUqPCtx0Fy3ZlLugObHOgzFVRm3GsImg2AsgNh17PzF5CZnLbXl3P/2jdXRPnDqp
0mrJ9JryCe+n+18xNFTP2yI/sFZ0xymFrkEFtR4MscY/pry5HUOyXWpkVIOTCk1HA/r+/6fdRv++
ly+Uqa5uunfcUIxoqqFMRlEL5tnRrOzMmS/QWAZ3SX8LcsluQlZmlSERyVzzXo2BMRffd2XBzoeJ
XPvglEPlnBmZ0qCAi3X1aWZCFmql/3Z14b9s0Aq1otQqqsZu7tj35KiIfzQawHjCYitRO8dncUG4
TDFs8wUm4X/ruQOYOpGYXwbkFTUEltIZdeXEF+siZUpkLYkyM5p435JvKtQBr7uXGZMVOUWIRZ7t
a+7E2WG/vWe3s9XKGqiYLIBEXSe/28pOLXmNuFqp3AyhiLEJtm67z5jiG5mNRJ2R66G6ux5ht2kR
8fEMDB5PRmsluYFm5btRd1c7V6gvMDxThcQ0PvDKd23XpL8Tv1FtATo6LT//aqE3zjWFMkaVkBBP
oVs/VViZiQ/H8+LeKEwKLr/28z9DQINhzaFAqKeaPYfUoXwXkptW2Ys7mH2nTsvCHtm60hr4cn+4
AT8bImxduakQ3NvodRezyyRAv45KKJhxIV4lTxeLsE3MLVLLyqh76LagZ1nhVYJmXiuNOfzy1dmE
PxCJc7V81hS3/7O6xqnqcszqeAdZC6c/ZAcWYH8OAoe/XE2AYhpmKnDZmpIiw4TqHkabeUI2ik/4
bd8U925xXUuV3Xpz552eEaF7Ek/VbWXeAx/SbbLuj+P+424YtGYPYXtsvoYE6BOaT88GfbyA2NTk
34NLhJ3HPULyze4noCVCiYlcJF5aTFqiq6phUtHgCiFtrHCDxbmPdFrH/yh1vJVgjSP/lkE97I9R
tRzPvqCSvKmpzL5WnO/zAbxI7jyhE//9cNX+NGxRwQnOIBUU0CV5BAr7Eluf+QZC+kkwQKANgXku
fPMyAEurRI1tT+qXlYFjinWQIDROOQ8EsWSCk9TSRbw2DXg2tsI1EzOed95HMDkdCPtRbX/VNXAo
p2y3KOYIVI3s7SMyXG9er01v+7dZa70RfDec59y3M6HhPgPQOeLCXIBFTzUEaKEbB5uiqhbIC6ia
Q+hsX/YBAMEEFiTEWm7evhmhkBgaDUhn555veyUVw6iCP+xX/gpYx5Ktm8P16R34iP46p/RPYGoh
rdxPg51fepTdEyGdiXIwB51UI3r3G8A0rV8+0zyi00TINhD8PFq4lHY09BObwNPvl+OjGhu9B7mt
BRwGctm8hiQ5KW1bXQSRNKVwVxM5y6ePoCaTxdUU9XoIZS8QaQpLs5dPr2s0ACUfNeAZkNmRUB+2
Q0Ja0mJsunKHJRfNIDMn9ZojHyeRVq6zgDVILIPAEKjcUW/T/KvObSyfGmhfywJfRtBhp2sYpYq4
b931CntfzMK4oC04xBUP6ZvvKssCBUvbar5FeovlElkEpRFqbAPIC5HKOjL2UaFMqrYDgu3A1VZK
gGAO44mr6GgSRW3PivibLfhXMYilWO2C7t4T4ZCP6rGLPqu6CmX07WnnvOQrkV6Ua/FKNy0m6zPr
+pPrNQ7pe/NVOwc9/WqouBKeOmoUJ+916Htju7/HDv1L+lHN2T71eNrNX+gg3aQr6XntAJMx0CPn
wOfJgpbepL5ENFvkrabHKZvuRrW7Go9b/e8vHFsD6WiNoBWAs2vEWNLLHe2qIbDj01JOuCffy4Ri
U5a2RFtdxWxivJ4orzfxwP1WL0WjsjK3Lb3qGRrcxn+9IHgchrK+T6v1kGHHlmJ2FdNo5ye3rZcj
LAZHEbqLSyFoKbf3myZVS+6Dx9op48Ey0l2OPsMGhFHTBsFDAQiQcOXB1YfKzUVenrTNnEXI+L4V
5As1Od6ENrv4wwkhm5jtfYgoazfPyU0HamNw3RPo8pzw7l2xEN4VARy9iJ9FzWS0hVUeHzxdXnXc
f2V4OO1v12PP87N0Y5iFdyFFJizW8vlmootXQReR+1i+cZlI7j+XRPmYW17W+1FLkU6XvrRtyHPz
mo48We/8TiFO54In4Axyhxfpb3LfphfoMF3rGUdM5FFdgxhKHPw9fATdYqPiV491A3R85Frtcohr
5nkyBUC1uqmykdX73Oybx3FIpmD3pWNz/8DgWrMQ5AaZPNHZcJl+cuwi8Paq55ZwkK1PIOX4un8P
FOp4xxghzntOENeKN5ghFABNq/vRjJLor3YaU/L9TPlMY41teqY5o43B5yByTEoN/PWj8fUxOvCD
Q5+qKemZLqTf+fD0lQiF/+Ys+8luMt0H3aU8wHVo+Ki+m2zubV1did7739buKaWkr2ZuuUpueZJu
x5+/IrLlAFi3KQ1QskhEPT941r7T23hk24YtI7KKwSU0XlVic+mdc8aCia0vh0NjMpxsNaxb+0RN
VO2uXOnQUeS48N016pjmLlLTL0GD8600zIheGom6yg45bO6mce/qiv/5zx7Z0tm4HdoeJmvdqfNh
ih07pwAb5Mpe+zjWBhi1rpsp75KyXOh51JAxCLQvnUL2hMn7TGmRpuQw2BvX0+tpollx7R4S4P8m
w3LEv9a8BBUNuzmkphEW+tDX8RNweV5/HEiHVS1ZE5qa3fFwQqdvmxOXELOYZuN9FS559XPv9smG
fBuJmIFF7+AvGsWVKbAS0U9EoQHEmfookIfpzPtL+wtp7iUTMnLtaZfNcks/3y9hCAe3HWZulPgd
BhBbMu1ftGzb+nDt4eZEG/noOWART6GGJDEkTxlCGCqD01kIh0ZcIwZW8EcHePOAJqu31Kx0BNZK
kfDkeBE6t4qSSc45BiErzUMUbkfGqMs70h/9bXHaR1vMxgDtMf9xfqJzVw+Xsx73cfqlW/TFDDRG
ozVwOvi9JGpFY19HRGLzuKK6x2TD6q3RAE7Qufg8KGqCQYRIgbUF98ONTk5+BiLMc6k3w88rFO+0
9GPzhIJoeRdCjbNViZXRyPgHnNItMzc2KrK7K+KMhDgUL31gzbFAIFHdyNENrOZ7ckz+lSgObE7k
kSU+ypfzzJRfXwQVkzcet3SCquPydkUoRmiuqD3VCrADwd3rUCDHMNiXOEd8WekhWvh0H/PTm/po
szSYAQXGKJyUN/qQ6Aqke/pNSo2UEmMDxpmMIJdNmtyweJfIfWYCUnywhLsdIVq9pvjX+xnpBLQl
Gc8RveZJt1TTZ8rR1Gy1s20p+fiGhs+zA76if8m8AsJloYYmYu5Ak7zBP6vYNU8/ZhJb3/J0bx1Z
jvqGlVBOrCOOhlMiPyNVef9vglb2ZfCMaKZR/bFLVfl83onlx8DzTzetR1+ENlmsOVuPUjkTCi4U
JvCT+1uOT0Hy8hq3QyldvTwlWFx5zbAakE/1v3BVoXR99OyjBXgDd7KhBkxfd1wTWgumYa3M1E4z
ZJqhHWtx8tEb4KYJFPkESI/MoFn10voU8RfzobMdfekbb2LspFo1E+t0zgoVieo9Raq8x3ijnX66
ruXUqCugsGxTI4WSouK1needXbNZTBj9oPXUFAnM1JehWWcSA4xgfw6ssmYBtfr6wDQttfPObFTD
Hj93u9VCW+Id1b7i2OvfCWgk3GxCu0/1gkhtGyhRBjvB/E2MnpRnFEo4nhYkuO1tId9TiYEeeppO
k5eBlH5beB1Jf+gNGQ1oSBUL+CiXnaGH8frxyfbZiIaiklP71rgNVmcs4mZamBnSfsnaOpEIBWfq
L1fKAKchsU1P7ATSH5xUHw9ZfpzmV/n2Fcd2qTeQd5J6Av2Mf8ehJNqJ/dTiw7z7kjZFS6ps3e0x
ZLI49xrG2OvXnQXaz1J88fhdcKNIJD5UA4Rv86QHB4q2D6zZIfn33tkq1IX19L96kjagB9xwxtqZ
JC4Pzbhgn+5nvd1ydyS/bikdTzPnKf+4e+S7Hg+qmdyHcrhnvE9w22yjbcxjbd3otLr7THyYHe9I
EOOXiDTanO2X/AZkLkii+o2dvG6ngzmJeWJoyTWvnEpUyvenDs99Z8SgcnQJdF50zzIYuCazn/NC
09s4gkwgwxQuA5StVofP7zoGq1EZdqhQbu3ywUh+KFLbKJGvHkaXLpuN8CVRJ+7piWUhH2/HZvLL
CmJIEBr1bOj2/Tt2UA61S58tNCIShNl19VDbxHzOhw6bOq+GmbsWsvYzOKcq8a9VnITrcm72bORs
p5cG7Q2bXjSFkNgv5DXxIzkdyPeUVnMPMomufpJgpbQHEzuLtx7d+iDtbogaRcisjeFNCqetWWeS
kuf409xIE71AjReMXFAZTGqHpqfssxQbb+SpEP5C3hlJiheSLItYIncPFdZu4BtfbL7zkRJMtvIe
Apcdw1yPSl6F3ZI3FQUcB7WvbvqfbKSwe8BTuMvET6j0ANUdHF3QD6h7VD5UDegBLmz25De+LFs0
UrbxyhZ7lo/le8e+zaU+dLW/FwdX3ZFncVHD3gqvKB0psd3RmlSCSUJ0wd8g1Qvh/4eBs3mi0NB5
YXGoG+eb1hi6AcXN1Y/Etel6/oaj460mD0lwfZhgVUA8RfAL2a/vkUGFzkDIEL+zkFHlQQfqJoU8
AXm7byevbo0tz8EaB3HYTaLt5FwBG/gh5ZdJJkJj+3pVIx62tNBHe3wSZGImPXTUF04/vaplcDU4
LsN37CCSCA2Vw7u98trWIa1zlc4QdLYkOH/htpqD/+aoYvopdosqpNRL00QlGICgM/mE9n9/Tmu2
FuuBDevJczjWLnEj9gs2XbQJ4HS64siqf7VOK5XfQXk5YmRBHXhDHsV2L+T4Ya2TRJAQheRgX9OR
w9YVrrBjmZRDRImr3yXMe/eOc8UY3mG8BnrfKpWCQBcOvE1aDfmpe7iVhLZkelsdFodG/CB3Sngp
ORD28q2aGzGUCfuLNSqB+OohqZXygjZt8gY057Ennpllrvz4gBoz2AWsqFv+XEzgWLKBS7ltb74K
sJykb9PTFNHOVv3Yb8eRqHTWO810P677aiN0HtX7Hyt0Mer/2L4AW49Lbbf7FW5AwchPYx+omKsC
98OzdxW4ajk7dEdmllUjeJFCU+0psFJlIBkzbZSm9f34bs6wvkzGiD6bCLeSDVNjs0EJyZqFGJjq
mTSs+2DOW1tT4FmILHart4ouHbvZkiP6MHQMp7/VecUKKXHA+YEBLtyU7LMhZkr5mD6SLjcJ9p4R
N+fRivtS0r9PeZkomQn9LLoIhxKhSyBctaxVbX/10OBtYCwtNkVDrRLO8VNPaE2/yfNgwVcm6yH0
WF6/zG2iA7oYbBv6aVhMuqzCY+UK93j935VHjHwDBMwPThc8TtSublSpXHedxfX011xQzNSGFsEO
GYEyax6nptmenh7fDXYdQVARUPK5mKvn7NNz7+zjrRmUWq+Z2qe59oQ/pH5vkRBO3pwEUU9YYR7r
C0tKLesXbk1ZhGqpqcacqZtIWQ9egmfKDA3m3lDVK/dKQGW+fc5oGzS3KeNHF6vp/2HaCwRsvNoV
M5G3+DPdImUfrWM6UidNE7YErhlcLGVJ3p/QtPd01tsllEUILt44sCSnZ1F/MCxeGKrGjYz60I/0
ij5BNre9sW7Mfs34vqCdsRP0eaxW6EjUCO7ii5Uumq00gFw6FyzS/a84kdFpGF56Na3Hasv2FPeZ
JQ/BqjD1gdIB8e4ZNd63kouQl6PDUPdlTqFzXxIxTCsf7Sms9uujunHzf04MdeS4FrGfkPiM4ozx
OwxlQxmz7tQyRd12ObjQqVhpOjiBCBYm+d5+QSYYPtN8mZGQ2SFSaS4VXWRGSlYv3z2IF0eGeEcO
wx85ytkGGCQBWMtyf8aHVYxJ6uDTeXYvoeH7f8eXn1V5p5VfTyiZjBCH0yPgqs2IYPUpwahwxMUq
EsT1333tO6JUVrRKd54DkwieLxTqvepKs+bsho3/W/kWTBPKT0I7j5KVqVMPqANjXth+eO8x4M/E
9hf3B0cvgdybZUVm1hTymKyiCs/BOOJDfc1u9hgOc3msBfS33PfJxMvBwNEsCWBIyD0FgAYDB7Rw
Rbzf8mXI5Zf9/sqimO7920ylpAdyFOm538J5xK54+i5VB9c7PV4bFPZL4tPiKpxHwFuEOC6c4vcV
b5NZ5vUxYGJs6xsl6o0raeLaDdbxkZiZCCng2+Z/BhAIbJ8HR4Xk3U4SxBKXnscCI1b8xHjCChtx
3JuESysr10joYqA++dQrnWjG3SP9Tr78r59XP6GWEENgWZRRMYrXfkBRz4chXaTrrYUnOZ2gdi8+
3X2GrzOFHWudFIc1KwZihH/pUDhvinfVE8h98b0Hd3k/YxRVqu2XfB1uKsN99AuQ9szQkvq4ksgj
T1PiFytWpnVEc3L8X3wmW1ma9P1r5n2p2w+IMIo6eu9g+GJ6ble5itW3mGRLdLFQiFvpJI4eCnbo
lC74mez7+14IzkL/vcL/SHKpkEWHD9HeJFd5AuDqdt5O3zt0pmkr234jZlogcQWWL8p9vTbFC1Lc
yeWBwxBB2UkxD+caElWtCHkhy6hMwJdf71f8oLqtxvzgjDkLJRTeZqzoRgpYU9+v9HHCjqQDHj1E
hlJwyH5mth3MNwLa2iH/c2N852z3WTKyeCAlmuF5Es51F32RDoht69aLnP1wQvrqSH2tdxQdgIoQ
Clvn4d90P6NNVZdxYqtU3sR+lpdWVOvkd8cHDKWixASSL6VxF2vkXPLZfKoTcLHeWW3pavepB6nQ
TDP6S1ejVLrLOjdTg/ON5OzjSIR87p69/f+VZzHaqJ0k+ta3tk19GcRrWPTFliMRtaWCBDAD9wcN
8cKfADSMEODa/fNRDp/61+Os0U8TCpNQk+NqZ3XTNPQBUzof5Rv0rdF6KdSXwlWaVUGK0HQAGf+j
WXJxmYx4WU6aAcjQKTP5seUoNb1WHfncO5UXaV/SVBfa9ndfI4KtCVFUeZ3Gx7qF98rCc5vjmDXP
JGenygK2uMy8g2utbJzjV0N11Wb8s9rIAE6j0Zbe9wC0v1p6oG1U6oNjXKkGKTUFm10wIn2nBxuI
BT+4zGW+0W0LUFP5hImr8qDIzSnCsTFxp5xzqt4M0XYfznvUneDLmSVXduDgXhomUkbudPRTTQfH
7Hgw0DBAaipdL71upATDniAHLZaa16J7deAeo/SsbfZtfnBRGqJEoQFY/dAT88JOZnE5rZrMcTDD
EDGKUuZEn3hTPkrHWMrKSVBH9hm1vACg8+WK3BvzE7v6X8ZJLi2WXT+8yVixVtQiBOfPa0+Jl6FF
0wF/Wujbjdtcz2bUYQZCOQ0WzngHpDW8FmbojpIGquHqmubn3PAWVmrjPlD+pjzg/lP+3L/Bj4bD
+VOGDoRv9G22o3haTonuklryF80CHHjzVrxbFYiP9PY2DcscIZhMFQ63cySr5rrYNBN1X8nM+ytn
lRS34UxogIP+WVFXJ9ONT+X9bU0FeM0TIy6T+gra+PbvYo+VXioxMJ8CmFpXXthcf3+Ul6Sj2izV
EE7Eq5HFfNewdX9eVL4vRsWvdoe/T/r+YSbzN6Tl+ETNDu0SINRZXKjxhqJPfFsZYn1yC1rHIZCt
HAsqxrICTZhePXm9g68ldgeaTI8LDK+JPx/YtCyWee0UEzbqscapnZPy8iumPP7RGslV7b80PqID
MaDqB9shmygkMXlUADA6xkEOCqyma7lzigwxzJFgdImQWR99UtxawE7mwr/bOD/gA7Ix4TQ0fR85
KHMiyXWcKd8is6WSCy2ZaDGGmMc9yMFOwW1DuQ8XviDGQVNIeQCGZsT5sLvDKKjjkJ6BFvXnEqZA
/ha3u0pvZbbDt8zBAzZCvpzDFRskwovzBIXyQqPkxU4xd238zSns8VNwOmTMYbUCGjnoTEDUdf+u
E07rqZG9cZhEpNAzMFUPTollzJCavXI5/CgKI2fQUuO7iBjxwwSiOQ/fxgfgG+hDmu6djbafxd9V
0L+QL52lv3nVeC6ppixxkQW6vPzrmdxXdVGbO3nPnmmim2JtQTNRH7vEPe2aJ0AjbUIz+uZCOdPt
gNN0MNMxf7d27Ay7fRzoKFW2JO7w6RKp3Tp/FOTc9b4TFvvb/AcnJMAIZRYGMCLjv8kzfLb49idc
PaAi+x6IQGLBwe3Op1XWIHCWtQAOMbV3VxjO8QkMX2xSBxvB30xqnu2TzkI40ntTzyYoukI9jwR4
Nmjp+3aCJXeAnz8xogKaeYhynTLH9hzrAxwVSCGIFgZjpLBxL2m+hZ5jnynwoB6AVnnVxF7ziVDm
q9G9o4b3Ej60lbC6JQiqKpziwpjHkClPIfUsGVx6LCioZezNXBXWjiVahDZUei6cuRZ7sQUGnzxv
VLAzplHKIoD1F4gEq5y2c7FVfEqHo70SbsAVgmzuYYxCEFYGcXD5qAoCftTejr2uPi/FZ9sZI675
M1Y2SzTAhoCwouVIxTHxdy5odCV0vgYXeL5MpSb6XL0f64RFmIettLzHxW0n7eP/PIGEps5TcMLx
UJdEfvMKsLIHapmSNC2WkiInuy6oXlzoVwLhY8MPd4SEJq6tPK536FCoucXLLY/J4QbSBTEvf0f7
9UhkwxACL8QLdSVK8wOZHFIGUOvjAgzG7fjxdZyAsb1JT9nQH6xSqY0LouDAQfx4PnrEyp4u71Wv
H+dP7VTgyX3nWBBR6/btNP9y861Um/tC2pG3aF1YXdcchy1K6CzV+NMfpnLtc+yYlsw35VNqbTW8
IcS1ioUNgJMy+IqeW751iwBDzdmjaamO0pebzPfdUqfWgAxGP+1yGrV1epq8N0g2bkrSb/TiWby0
sl/6XWrEEnhaOsW893ZNVSkUDe3Hiz31dpJuuYj9yRNlhYul2MQvmzW9HBhl//vzXPNhrELK4F3c
hFQGDhai09SmqwtuAY/YktJqJg6YqW0ubFRGuLsiNbABg/J3DDLXq5d4wYAjQvTG5AYdBLdzNZaF
ILAgm2FkOrm78UY/iPxEIozNRTRMKjEIsktXPH3YTnLsW5qrUE+0vSpYJl70NJSey8yo5u/az+XC
gwdwhpImhADqJ1KUu9I5GMqxYe30LHSYx5rrgVlsn83yWNvRTlSucyrqFEtKybPHa7AVPZWYDNLg
k56MPuOG2WXx7nsQ0yUSjT3Vg8iK4JE9hxA1+cw23TdN8LfNC9hiJ97DrC6a+QTT657Va30dEdlu
GS/wBlvCD2p5xvtAQEQmI2L0w2ijZRj78HD+vtNohS0iuRpZTv5HwDrd6MxnjU0G6o4lxpwwSTK+
Kw/Oh+IA8qYcJ0e8jFXRDe2QKN7iGKE5bxR0k3OIgYq7Cut1Wmr7JM6ilsn5VCYHtlVavR9QcRfg
n/s3GwZZSKPe+n63MyVo+imC/dtoM/WvchaY4oBn5u4vYtKWMkV5psxOJOn6kowhip+aDDhi+Zle
XHtypY7073VuEDTH8U6SxoFR+eryftvMEKSKoMo9WgqBxHn8GcAmKvyeXppIU7Y6FyVjsdvMJ2hf
ylIRsH2tchDuClOOcZfl28wbcihdPX1spNwF4p60KTenbl0ucPVg4xiTaPi7pWkheVi9p9nMiQd2
v1Ul9vYbOWe5EkcJV0fQPaqDlp7qSlKOk/76pmLxdFcmuMMDDV7o9kOZUY59jvQ2Ztvltny8u8Sh
hAlXo7wRZdayeA1i+6zvUBw28JpE3QjuffmRHRbUn9czxrEwNYK486iUyfNRkmmOr86XV4RNmdVo
ERiGr4SF1EfbcDd5uxzt6RzaXD2F0UPCqa2rN0P3Yko4vATYnz27rp+qp5tauf56xQNv5EXbmSZM
D6oPLzPXCWbjnDzgtnbPvtOKMb6pcbQlkPrwDC8nKqb9DLY/q+n80bJaDwS9Pp/tQ48v9iaPlOJv
tBQIjoN4WPNxcPX+Z8BUaLCdeLpk+8kL0ANEw3KuNywnYdiDMLgbg8aqh4Ma2DLNaRw9tIn8161G
9r+N1qM6uyHtwuZ0UZeK3yX7rFdvHLJo3Rk41pNlqRPoN7Oi62oyYtmI00MnKTnSXEeVUOCFuEf4
h/Xb3PKWLvuczOLyFHr2A1JJlGKa7DpkiV6at49vdMODZgTrDYv3i/wLlTtUQdTKCV5GhmTFVQG8
ZUL7+Xi/fs6iJFH3NVgwMRTzOfBJBh1aw1w+wRg8ceHvy/Ic5n2xTnS9+AGSHdz2zSPb8Pgbss/j
hE9tJDoADwj1KZHjVKDbYBlSohzIA/OuqYZZzn78Oq+1ycYN4Ht4d5A3cPKB+TKPy8r49Z5PxoAS
g/CQhHvc7Aqq0ZIwJZEyKMsP+IdTXgC2Z0vob8kDfxBY9r5bkDxxRYjj2/HZ86fEYbXq1G+cAbbo
UqhjKfEHKdJuvF8Pu9V39bq5fq3cEynEhiZcHNpVoNZeKj4rRBQwu2DSNTSt101EsWN7VkzYbFk3
ohQuZ0TeyBoyJJZUFo6vNda4nYDZVlq5wjVmmE2rzBxXjmfswUAJyaIyqh0rTH1yADZ5SZZHC2Qf
NMOWNQq0Xy/To6j8UAAS7Xm8CBT69SEe1a/uTlAHGfcay3miE11K9snw/aOL+6DpMmttA7MT6ojt
T9uivqjJnYW4I5ApN6TDWj2bG3t5Ox0+88I9uGb4snyasyhSMh/W1HE1u+6yw/EggVWuxMW93XDt
DxB4Wr1t0ZYiKrR1syh2YdaPPadKCo4Rhsn0wmofi626Vk9FPCL4/sCeSrhSirRHe/Ivgq/ZIGvx
OK1yk5ON3VZNGY3lezvXs/x32GAmRhqYRhyojP1wly+vTtuPxfEeyuK9mTrt4SPKAi28OqF88VDk
XsANJKPp36BZm45SCGbebBlFhoUrpHoA2uOz1t9RCGxJW+8djo80k2XfJNxbU6BSUTkKmliJXjGM
lraHR0S8mAxgvD/5dQl1JCLDoQV719uXNfMZhIJZpSVyWLxbEggWta0MBq6Vyx+bdretl1FPRfzu
CkDs2+KMZkFhrcmX7KXqZXEaYcciR5uUeHdRtcMdHfP90Fbfvf4l9Zx8wOZ7tetEfcnCDh2tvdng
M6WlKj5hQSOgLdyWQYmrUSMacJyjDWL2a9AwURiVReu7m0mpjqHPln01ceron90m1j5n4G9bhoy1
I1/TtP/UzpGlPzRxH0rLgmu7YbrN3fLTnP3IhcXhOt7g+Q7MOVAYU0O2tmcFN+kUM/51I/l5hPLf
HMEPWd5uDDxtRjr/Y6f0pH96KbxC0nRUqK7lM1RY3D/gpGM90q5rxMNqqa8iu/FiYUng+3wWczub
R1ynDQ2/HZsHcUvmUDbf5peMRcCSmHxrE327jSXWHgD2qrDPfK4GZGZDJLaXQXlHBgInBFxSi+Nv
D9vPTqWM6JkFslfYYt6/yrX7jeOjnVPG4QYPoTOL9QLeNXKzJQfOD0SO+3an/CAumCsXFHdfSBSL
gmfiNoGM2nt1YsoUftjkMaIF5ZnMPxxF44jNKWweJfVJTA8NRMeA5MSsbw8l1rBKyp/gSvvmmB9f
QYKMJK+kiPBjQH51Eqn3e2j63lJU5SQFWeLEm8CfVsf/zM6IQoajce8+mlqDhiGyLFIF1AfIAZ/S
ow90Augi3sn2K/Kpyb3UU/c2RTtc0LSvKkyp0viEDnZTYZEmjTbMXTrOydaH5TJ07DOZEDikABID
oEeE8Mk613O21nM62xzSdfzQV19n8ej9gCD+EBAApYcBKUsttMdMd6+b9dU7VewwNWuUko5JMy78
ZUQd3cY4v9g7+ikZZgZQMLstw/h/pMAbMuw2nQmU2aucZxXQifrV0PGJs24MLBnqcZtrG0ocfxQh
6GPfP4PQh1JWlg2DsX1GpNo17IHJL9dkVW720EuE5SL9fMx5AX9aGBabsXbnTFpcxP6I10KGHA8U
sI14+W4+XPA1ioZYAGtnI09QHGEJx+h0MONth7kzs6LCBAYPIcB1pLqMQ8i8UX1si25IVWaufX4f
FwaaHwL7qmVWPIOo5mdKcEr0U2+Le5zf88u+NijcTPILpCYOohUl4R2NepWnZ4QlIbQIqxm2swCb
0AQDk/g9++iTHE88kNnJlzKpHhirkxOeSOK8BddtQ+wpyj2aT7WyIGDRK9YmqBFnQA4HP6lm45Hi
5llcLhKd1mOye99iyobDWDO5rZoqccDWhIBiWISclwORWcpAXozr8xefNN1R8+PuOtzWtwcY8nRx
eZYui+L2yhyy+r8fUO6vdjO9rPkIl6hqKq5sFQ+dIJcengC7ey/bfTBxSzc0S0YsqgJAWAZ1Y4MU
xcud5fJzmdyZQuZqeMdj2PR0Yb2FZxuQuIBCt9+0JCDroOHR2HO8IuHkEqEuGF6b7Pa4rJbGEvSf
H1akdM5ncOwYrMhpYiwbrut+agLq41xDZgub8+ir4i0hTdgQXGVHpZq8vGvqrmrYKUOSBfQrM59j
FjGT9HWw2ez7vq1jy1BnN7dy0VOLfSTbyFNmCuxK3meCQRPR7yu/OxAkSoQORNZC+nKridtqbM+9
8KQQ+mD8aWOX+yIvNePSMQegzWkGBIQ23rwKL9uLrbindJBQiuC7jJ30XFHB2+rvaoP+9qXHlgO+
iL3xVFPALsvPXJgbSYkeyIHcPG/qrcSR3fqmv3/Kve4I0tedzvfNhib5+EOTYiGfYWLsWw70vms6
pPvCPzszbPgvMQpohS0Rb44AzNUqladRCdhteJ3Ay9YWqbzKARtKp8h3mucdr6cBAPeiGfKf9UZt
gWlmnI6V5tiC5sVSJk/xVlCFX/X6p/R7czLOmbO0U5LaqxCxVoAn2OaBoTKU/Fvn9hLl2c2loQYi
beaW/1nZTUTdNpb8+N7rc1zZG+WWO7+dsKGGvWjA/xqKeoljJSLsz7F3PLZcBmo6usxpvR/TKf2d
1XW4iQd0BqXj9qWO3/n735adt9KqeRCPOYH7BF12hX7B9P/Wa8EVmBI4mTbKrMGv15U98+d03SeW
KaVAY7fubFSNskEt+cV9buIJc2tENjkzzG6ORFNqbL024Nv7ytcE4YzL8ozRj5mX2Ku7cSRocMre
JPBnMP17M+fctEyl4ocrvpF6P0NPFxp24cZhx64haozcI8ByEdxoJsrPkAvkHlWiM8bMydt0tHwV
Wo2Q/sRWN+/CJkxwOe+LzqdAw3/yDtISo6dGWAy/NfdHeBY/OFHp/IBO6CBy3Y+OxEjLFM7YSHdt
M86x+fV/Uz49yAOT4CvL7LeUgMtANz0VlT3CCbIy2b2QaHo1DP5kSp44d+r5hdZHG9+rR3QIYwbW
yiCScNCeucpYoqtsveyx4h3Htwf4jg0zShyZY6egPGg87PViuoxZ8yuMl8FIk6x48EIHcq+EQ24a
YtQ1plg5J9xK/ZFek9a1+eVX8b5JWZktTuOilf5i+u6d7+fjqL2VKSAyhpNot39xFsjLGAwNbUAv
x12EXPR5jv9UNtF6AOzLXQeydaG2ybv/XjQIImtXoMIJOXh+zcJLCytCn8fHkHntDn/FIAA/VRXA
0oyTVMaTeZDhAYIdc9WzcuuKXcssTXTuXYWA4swP1IDwrZSTj1O2HqBXzCf9GXSbNE9xIkF3UKyl
oXzeo7W02BYXxPd8tPiAL8MP1eGaTq6yJ7HsUUQ/Kv9EI/V0X5eK8Wu5nbiy2Cum4mjoWZi3yHnp
f+TRkM8hiezQOxpeUax8gS2l5MsXMxctCFWs+FQ/LzC6h59lXWC/4JKmrw4f3peb+HFvb2FSBarG
I2YTYyyypz+B8me1YWo3vnhanUd/HKx6atxkMgpBgRrD0NCh5AUgstV4H0skTUFHC6Crx0AWsrhD
9KkACmKEufe/Ks+JVO85ETeGygQFakeddmrRHrAmmr90hVkvke5xlzQuVn7DJxXszseAwfUb7Rlc
7wwLBMg6E7w+sysog/YV1o+25VSMFmks3DvslA1t06EvfDIh8zSY+b0aKjxc6kFSoTjXGDzUYvfQ
vFgp5CABOdvomFDcqA9gkUdqB/I5jbDqmVMcXXTF36RGqVFRgiuoICqySrz2XuuO9hXPbseoi4sF
76pPWj43looGlizJz3DCtko+Abg83vHzqkzKgBYZFTzyRPb82i0u4y0YMuvS5+qziTu8k3olBQFX
iz5FX/yoR0qW8UioT/NYa0VcsqV7N8qOkitb+eZn3s++s+zXo8KIuTJj2WYveWjvdQ0BM/F5yS5K
FCVjIF+efQjQ3jx8ON3GTMBMxGVCAQ+ShgUNqaKrKE1/kmqnGO1IBr0ttelxNA3gwJU9RFA1kwVB
RRgtG3EapQupEZX0TSHAVpdw0Y05cS/EGxZjtiJmZ5ZjABFrkEde43CfaJ87xd/YbYgGwTfm9f/d
7HI7NAf/DvBqxTe2ewLFKwtcRP5yWZU4CbFAYVGIrgmsJ5U5YRZZHAYL4zFWfY40+pWcS7kUbhSG
L3x2Xp7hMfaG1ouLpiGXz0ApFaIMJ8U0Adrs7VJJwJ+jgzi61GIUEx/nzNrWg181IJ/uylVNx/VU
HaDgAVCMYfag60YPqrg0C3zwSM9xivosp6UwZQF7dxobI9gfcI8DXe/nyvgD6M+bR2HMJ3xO/Slo
6vi/xmLGT7OZSU2I4HnlAnfrwSnsFW4Plpn12B8Qndd9OpSnwTtK2132K2iaPuau7tKvqo34qstc
E2a/mkpGF8+hcH7xy4s5Qw7a4mqxUapP8VI/KjLXXUMA48Ko1uTLtmZB9YSZ+biXSaKErzQlE5Ja
bQPMLxsaGxgUrnpaR9JjOBU1L19imST4q5Dfro55mnDCHyUk/pAeutROIlNBt1L2wZ+peajqZ6V2
EuNLTKgeW3jV3fHvKUn5gLDgNrjA3KtjHAFw8nOhOTCUB2v5dRfF/G//fl00SUAzOo1TqtqU/lCN
sKaXSCxVCS9A3GuFnw4sHeBGAoGm48KkZbNwpQaV/gP+t/9LVczZuZ2SVjT7yW9rcKh5oRXab9Vs
WZryOtr4i/buvH6RHmKBT7Z+kFm+ldSdA80CELqVwVvygx5ypG4DyL/I3qqSxru7XP8hweWhf+VF
OmmAsoGs0TDlvR+1qAMDFbtojz47TcYPVTBY3X2wXDkRTJI9OkXSq/QqvdBsaUCBpkBGu9eVMttD
5yIc96zujCs5SToPobhpnCTJjj9zbecC33Xh7Mebj176u1TJS5io9RF5fdOivTV17l/vE4OxzvPQ
cxUbtNygm+JPqWoBwfxltXm2JPtDEmsbEeAe8SefrXRiCxyjApPgCOkslJWx7KHM6f61dU5AOfCY
yMfIm22f4JRZOnOnxDLoOvkZUvFz2OAEkJCzkMN9FHTUDN10SVoyrmQloNmn1Jut2zZsPJf3eK1j
KpvrjTtW6QvKPkXKxHjxfMvV2P1Y1aq616Jx7wKISRwJVD5/le0FAMO7CofPXwWj6O28hBfWzFwh
4FfNV0cjzXT1j3SX8jQiv9E8/7o3KC2eTgfffstTKFRkI0Ooi5thdYHTt3nUu42AS5NAOm+bs+QA
nwvZm5G0HrFSBD51NtK4qZ/RwsX2Pkij5XfFfH0o/mQCPCq8ZPlmIBpf9OS1EleHCPge/MrfYqIJ
37QY9xxa0jMxzrixj3844/Xv386FkQX+3b8hUgBz7K3ezE/nz4ryTSk74kNDJCOtfRaH0mcum+/e
ejxCrtUbr6ikJpIe1flpvo5PwpnmFPGVJ8EEyZ02xeVGp0GzviGF6kOn5b13M2nIbcSo3UQw8q33
rTIzzehYtvBzorZ8w9zXWzf5jhRLxvY/IclB9Ie2bx4K4f2QWJaCvvaIZM4zEDDKuptPdvqeMsdb
u5oJhUy+FTmIU0cLACYuJ2Jbqhw/w8Ad73cB5a5CekT4OtXf504Evzkukr/2ChuIjB2bQZK54ACn
RdXuFGOUJLr+SeuCheMTGpABZDqBORd5W2wJqrP2da/OGq4LOc6w+dptezHXjXxWjugvaPeBNo32
WXl8zohMD9gjZDOAKX3N6kh4KibqF3YCU1Tal5I+IBQaDrJaoPEJriWAu0HkFttItJbx6PqXU4jP
IGEeYhhyWO/Hy++jm+rogt2b1e8kABkcS6+z4kLPbMLjH2hJhNr551LpxDoJJ2BmbSOliksCCWwd
1Aw5ufdVJYCXy5SZM3EUbEZqXsgZIsEcVtM9s1Jc8j61/7o5SPd8A4SJxkm0pibApukHGaYxHAko
Xro1PeBY0YLLL0OhvtFuN2Wt5kL4S+Zrt9wND80QDIRQCMvoanogyPSoAPRfEuIla4eFDT3vnTKG
ab+ZSFIQfZ1ZEjLshlzzvwcMLw+OWLlQ+EqhK8y51JomW4ETfPwJZyr/5Z/xxCbDvHTAAaP+ngCC
sOwysrbDNOHLo0pJorUImYZwAhp5cDSktuEKyloq0FDEhSJZmey+BAb9hwnVlNkHz1XCNhev8jt9
7Kw14PeMMbVDXly7Tl5W6A6wenrLuSrHb7u95bDkzn5rB+MZ/sprq4S48QnhguYKOiGjJXCM42Mt
YjXSoUn1dsbIoqu8EnFz/fWQc4qiz8FFRH4iX5kq7Ox4EQhRFR/e8vfCejBjJz/Mg2zhATKcePbi
vuhwHfxFyQ3PsS3g/UgtDdMdRQOqWVGkTp/fc7v9Idu5ZfpcX3V0bi5QgMNqBnBLitkwK7ntByY0
zbYPA2G/u6mLl9VI8g4NWgYHj5mB6v15DI6OP3LUN2cg3XX5IDxEWsv6bpiePuzsP88AL6CWbIrE
5zAGPfFe59UWi0js7z0bm8WxaxuXJHn4eb5dTSfhT+QjqQb8/yKqvuztzL0g44OvWi1hy4Xsww3Z
36Y/DroUjDlNP7kWv5gYQG7A2roW8/tTeg0YrC4124drn6dOwgtjhCBvbTOn9G3iHzzRt/noaVuL
eer+/Sr1oRIq/eWysibYL1/euvvWRPakijdn0Gip/6ksxAmyxk6JQCSkGH3jfwUuXwu7H6QUlTJ5
ZYb1dPxEvIb3PX6rUA7LfRMiu+PzXqWPNuh/mDaM+l97nZ85kVyZJICZM3xNFeVAjgMglz6r+/e0
xXxTqJveDPXbHjW7acg17xuYUeuz0YdTbcueBR5U7+nPbgjFxXIbPU6V0O6Fnqe81zDD/Gt7efsj
ysNkYINdfx18y7OrCvIPMIiMKavAXxdMH/y8M2ulm3/EuZF16bMOsP/xDxYmCs364w4f6qMlsGVY
k3gBIk3nAsjrsU4/kyVFLmQneuyFYNYDe1fDjIc94GWBJjPeBaB+WFDVKRj8i4P2hFvNlKmXgXGQ
tL99flx2xyXrkA/p4M3vjdGhy6r0Sz3n6ljSHBqJuBlKZ3+ttkzZkPKiWlze+/uUixK9luILtO0U
B2eZh/anUcBflngg93bqTBYBSFy5Qj7TQ+hz6RzV3rrypocmLHFnt3tx6TLERzQGk4C5oO93zIqy
BCeYCYN+dBrb0G0lf0B8nT4A5EFO+8o8w8rl/FlhYQgsARnnKTO34sHWflXmeqwIFknlgMimnDz4
tJGCGtMs0g8OVgWTbSRP/jqNeLRFz6K+qRZQ++1IBBRCcUyYBOGcnvtQvwiTrfIJ639bZeXoyPQA
V0HHKjuTPoVxbEINqqDnSymxOE8Mtf8KuV3O6gTrezt4SB6LlBhilbOcpwvmc1qF7O1aC5kCGj/S
VfXb1wttA7wmv19fMDncu7cQAiUu5dtaInJemH6ypf9MwxLgiqcJfo7ebKi5HJyjzEXMseLn/RlY
NhnhReVWZLm967uGQWbtc+tCKlplFY1e3VLojLBZQTFJPlxaJREOyr90HXGrfo9HgavtP1OwIg/t
jk2abjHiYRYvbjS6tt48ockXa6gPDfMzVZbcRroMPJlzdfM/ue6+Z0p9Ejy6kldJ6YSkaI18dGUb
WcLy46E8t/zcm0mpPD4QcnP5hIXeVFeMJ4mk40IYYX5yPPiSLRaW+cMLD3CeZijqccUE0Wm5oyjr
YGiB6TU7B3vmv7P+x1+5FaCNFiWPHD/Z0z84yNm9Nge0YoFlUSOBVWheXdUPvjF/s+YLZMYfT0dX
8jf30DVvh0SlqS41LhhtYyLTP/1XCiUW/S8Oh7p50yneyLU/9uZ++ZksMVTndhmImr0z2XltMFNQ
WHAEmNHm7xaoHiLCa+VUiB60R/Na0G90qhz/xS9SWoYvXJ61TiOzmhZJyZGooWonuMVcXm2flmc3
e/8GRPn8U/NnfdRiUH+MTTgMQpBsSlJJP95x/uK/as0IE1tk/Szs1ztg1RuVGzeAWTpelphQEzyR
t9tsFAMdeb7t2Evv9Mr+ywX14x/7xbJ5ZqDpZMLGF1kxtPHRT7LuY7NVtUoEH9898w0iKhD+Hfts
D+eYqNC9QKAKP9cfhnC5YtyjqgDnR7aGaZTaqyJ9jhbSyUPJYJBCq0b0xZCRzyQ5yZfsvfIu1w5c
oQHwJVAKmbV7xaxoC5uaOeyIfte331l2wGbcJ8zbB8bBAsHzz2fRloS/VpsU13jWYhGQFPC+ocf2
aXhIXDbf93qrPbLBkhncylyY17Zci+UuzOOPSshxZyqeK7VK5eThpsKEjFw351WW3SwMQF5Syizj
1r8LBdAzZbuGgYc3pGp0lYFMcX8BGwwOyXn5SqWvXy8ij7UYzW6cBLF1M8U1tIeKv3pbmoCxbLMb
24QqCuvOyMCb9rGW/fyIcZCOAImvi6T82XiZbGGTmBt3FraWt1ROMJvhvP7hdrWh5fys0UVrO1ZH
cRjeWDpsqZtlBOlVsl/bGO1UjBUHVdYnZt+99209TmnNn/B4gZvVuLYk5F0ibk1xQEqrVkMlzO6B
Y0tU+wEaf6eQmFPbKiOI/eFBOUKsItj5xppU+EK05V/Nw7kyDyl5rcUrACpB20TxBMeGSExrdnUD
uDbCtaBKFAqLvIdTm6x98aw1RTuRhwKkrFFi3qiaL4TXsX5jKEL2NFJ+G9IsoiYQ/AEd1zwUZV9y
31K0WpDkOF+1EUb2z5kzFtcBU0Nc3ZCdN6C6H45nZSBytyx4dylOjdRn08R0PJ1lr0X/ecuHCHtd
AEJBhlpv4++WW0d5y8vRTbN9G4KQy3pAYDR2EfOXn7FdQv1D6xL7hOPpp5fQovOeYQD4trfJ1MMC
BkpvZb5jtFY2lHYd496F+tkjd32uYKgdHyIqVB5u6cp4IRaOZpGfg2xM3cE4Ys9J8ILLDlCfKPVi
Gp4gN87gsiQq/3cm3az0s+as+er+uKJfLQoy8r80DPhERhWU5lhD3MoV3Unws6WZaGIUjTUoVbdP
HCXBArGALS8SuQQPdD4733IazzHVBkblJXVtZeyr8ogoCT1rmEY0wTDb0tztfTNH4VeqaNidCvN8
hnuerSn3KqZYOP+HhqJlrNxNcThk/qMe0B+XnXzfDaHBpK/rdlb70L1Ir3pV/zJrDANbS93lgsrS
3QPLfRsdV8AuR9+rgDcXsl0lbeUg6NeFu9rXoHaYlYub8slSP01RaioG8rojj2Evr8QKH7W6kQn4
UIHg7uHHE58nP+11dFXQbtopOR6kTlNwV7872i75mSXTLROebP5r5nadDSy9YNAUMAdV5d4UNZy0
96RWmq1agNKoFCvbIFhAit/CE1TUb9TooevEN7bRL5Z5Ai4Ll2ABqkAVyrcnIlR5e9QeQHzaLiLn
cKvUBZj9J1BAURxyZs7cMmrOJMxfWjX9MABdjJK1D2ZZMHe+x5tGhsSvMwvIZz0KJm8re4mnPnZN
iaifM7NmZEGMJq5iGuxtpBSLYAUawk1FDIkINezioqD+e2kFKQ2F3JNvp2yeeCl9b1E0G+rgG66W
QxtLoWeq74ZRb7nl2sZpG1etHSg3xeqYenniPxUhb9euSi3HtFgNWlaUEPJHkIt1t1noxTQpio5T
iquGTcsOq2Kcr1fa4Pu7YODM3U2lhw2W5dIbh7Haxsh7qPjYuCP+Du2tJ5/cM/dJDe2/TQPOMWX9
QCencGcZwt7q353sckf340XuijxGMHDgpWfXi6i8H+1e1LUyimufvTOf6bzhvihls6iw70KqJrK3
HBIxNm9dDadcNedVxRHwQgRqgLMjrPaW0clW23j7zCeyeVnSoZkiNlMF4K/AfQ29uImPzwhGdPwj
unFTSYYikuvMymc+CIkKvNw64XDAtnVjR/EisCJEDa2yLfx3szvqoFv1y0+xg+JBg4hhBwnsJy0s
l0cH3W10wdrI9VfamzcCJGH+X8emnUWEJblqUB525duCkVuwSyds5hbIY3zynYk959EYncziaolk
PKgOACo9oLIzZyI9O2YMvz3Yo88wW6Ng+AFqin/W3pChBkCp52NA7M8zlUlw1it8AnptA4XPJoUC
3/HqKyG0GsVZsldgfAsKSeshO403LTVsbu8JD+eaNoRovDAXl9gIBKD9zlpFFEEG+hKpYIVXZ0Ho
FhP8Nl5JBPEjF407TFs7rZPKdW3Yx/S+r0C0gtVt4p722OKa9MX+4jLmVYCxkzwBDp69TbeSpCTT
8SyLBQQP0G0lFg5jJfnlsNgPJ/+Q7vQGhDI+YQ1mE3/7iggHS/IcaxHssctAPnHGrDrjjJXO+6it
IsdO+ZCcH2lJOGPPHRaw4d19vkqxyXx27aRMxyOUdk6DH4HVmH1Vh7H8XI+8rBtr8QbFg50HD5ct
8u76pjvBw9FepPc/8UzrrweMS45O3w/MhSZJCNz4V5AzfgTFUB14q82abYZenVOBAc2DeHUkavFQ
dfhrXwtpH4gKceDvgcILZtrqDKrXYDEeHWFV4mOHu7bCGFyf3EswkfrfCZTs1jd/SIZo3HWHgcjG
EEvGVeLR4oFWvNSEoXOYXls1eRZgXns4QS6EWJ4+RhAzbXs6MNB1aRu6rcO4FQc5iuys4Ol9WBu+
C8za11732LG6a04NkOsxbirdcODR0BLNlL98wayXmdsy/RWbSzyPI+DKIjqWFJZIedU4/QLMpRuy
azVxKpON3K0YdunATANfR9j/eF91QQc6QFPt7QnhvdzMlxtBKRTJNpQbcyqZKhcQPM1vK90Cd5zz
VnG1paC8tSB5cQMAJ8n9ogXuXxhitOI5DcMvOTa71gYOwIvbO8RcaWI/hDhDse86gvV2EL2uTmge
TrGuBfWKFudHt7SaClFzQX0WWrXKsKK8cgruCdQ3RQlzKLs3k/PN4u6D/mFq95AL7580E9HLX0Yh
Yy4LkUuxSJei4bCUEjKBLQaC7FJ6KrWcfPrlRorY1fwOxhU5nEo8Z9IeEIWYdM9YQQjseM0xUUXZ
PWFNxM8AwExNiSVerk4caMWvsVpQRroxYr5dGIgYRbLWecoXtt6ZIufU/8vfrAKte8PTDFitDm7j
Us4Hb1hhE/qQkBfhMLnBgrzIM29LcBhHUb+LmkMVvJx5fahn1w4uUhqV7B9AEJ4gbAuYNo3A7p04
p1Y7JKVTBtetGvMkI7rBJHizZM0aR3GTTKBlLCqYGEQ1gb5VXfw3iUwpVJ7QqQGZ5MH2Wp5gpgIi
kJJuc+zzr+RE3OvjeP9YUtiQtwhw82GxaaRHAJZw+WHNdnKcuJ7hGaAbwZckWYzcGM1i+cHSAtBs
RToEwRPfv4TPdzUojyxNBZVCOc0SOK4cnI3tAERopX/8aZucTkXnCTm6ch5bEmvBZ7GlBJDsD/+t
XSe2jsH2q0ZOynkR30iGmPNe7G/DhJE0D4SzFuc0Ln+5lUYS2Grp+6HdgeaMfe4rFxvXsxL0Okr5
G68bsKe/gxtbsLKjhl+MiEoNLK5c4H9PpaUOPtU/qNkbrOKz6Ey7xbspDkKSkcKRmEGsP4YF55pt
9TeEDNPTtUEQUaCXxQLKjnE7W+Q+IDy74XbsSVjg6QSev7mLkO6JXKjWIW2bwVT7ceaLdFVaCzJR
xHpKl3sA8NXolmRPQpr7YjgnTNYKG67ZsG8ho/GnJPtLxZvN0q/+KRFUNt0M0z+yZ/sYwRUDkB2u
Efdf5SV2jkgQN3Qs3Nk3GN+u/Kh6ucMtUvGVL2/NZCr5M+6NISaBUrr4qYYBgcGUruDG8AiBPGIS
wW9uC8Hxus6zWJvqAQ8yJpLycPsBV9rZ7k8JWDHgvaYAzloJMymKLqqmIGxhoXXxk/H3CVM1clKw
f4zAEmEgrAVA6zgs0dp/A5gO1APMHU+AbuNL0IiAuQvPTQ211H+cwdc/7yiFiOkJqnXHaBw0w+z/
AFQOXn2gX6mzS5DmnZI8bpKcRXKeun1wv8WON26/uwtd4j0i2pw5mBlENm+MvGoPv+aw9rgsObbR
v+d4RQ2yqJaImTpcHZus/d8UVJShBOxNuAR2gdogteMXQ7UtT2MvgsJi46lGeTaw2PtadffABD7s
CujXlnHm6+wGMYZuXMt9aeGpEOAP7iAb+oG/+ZQBDf5rlnMqHa1Mhop9zZ+vkWO2ZOEY712VoxFe
cVRSIDiX7usHF/SX4AvZmmC7P4UDAjsHvOBqhlZAh1OghwSCqFFmhSvxGNkesjMn54hSRNIAZnWi
jxpcg1SFEhDrpXIUoryFk0mVZn7B4beuZgtO2xtQRj1KONwS0qTEnU3e/kHCsbaKvgpQPVB2OJ1G
0itjw3NvHitn8MTAl0Nx/sZBqMkMOVnHjRoD+ijMj7gOXjdOjtrUSh4T32Ge2oO86ZnkXt6J1P5/
XGcxANLoQqapFj9O02no6HhVu2gD5mmaVckOfbfVfZ6ZhULiY+9fK1umGOXRJEFndPu8/mXB2YkT
G64rbcExJMNPzjUPgB4/emHEK4HGVW+2LwuFUAbPK3sFbNnIF+WMI38adiobhvQ1rDu3w4LtECOO
alhtXJle1q5ig7FZL1wHRrJG7EZNtfM/yj+ZlO20/ZeNcDEZzVM0dpanSPaDLzYDQemr/QNtcIvv
DN0+EC18rMAq9fzzREG3IzxL5PH6953b8zGk4hmKY4DfMm+h6M4IO/MkJdSImsz/yiFyyFjjniwW
NBF3k6USahrIO8d8+Kp9alKO5pn+62Qy2+kwZ7WAEpao3zS+CJriScFAd9HJ9slDDeaYcLmNmyx2
BrPV6Qoz1qY1iWTdSKvLigbbsGhmtOhhHw8Q9AuCZiOidsL/vH5dHdm6tTLOZZC1n2MmYfgIfUGr
2kUU7pZ2Dw73C87jmdmBTnN/Ng6UoaK5iFLcuHZzNdbbB6CzvMfGC053mZ4Yf6SQOX1HOnzsyLWc
9tcNK8+dvArfyIR5ANZgKcIVhzXkNc4LjWnNxUUeKmbiH0X2SKE/cEtVsgt7X25dQn4aHrNPzxHQ
6xb0Wpoksf43CEzyCHC1EElcPsgEKL/7jJgiR9TAwcuyCSU9p6aZuz0jCgVxpMUUm2xTiOvxIEoD
FyM5tBGEiWVmOwEFpq9TU4kN8pQ5ZbIzzKVXv0eOZOygx70RD/Prz6ChDdSn/+63sYs4VDnZO0/7
U1fFY1u0Uf16O6qYGuK9kb1Qcw3q0uZnTCqVelPc5l69W4XC+exaSuevZ0EE8upr4j6hbIk1F/je
UWLz7F9W/M1d/4eZQdKxJM8lpUfavhx1z+VD6LXW9NO9TLcL5xrGN5zuFvRunTB+p5ndOOfJ8aUJ
ZMuqgY0BeKQTdYCQ8uLysP5tgqvXi1L+Fso8a/GXSkpKg6Gaij3ZiQ8pbRScQ7Nqe3fTlWPa+o2V
GsTdW6Pz1z0bZJwvCEW68TOkcmM5TX7ETO6pRyWap+v2QuM2PjwkxyB3TbmViq3m4bw0f1UbLAEi
ipxnp4VB2f+gNev35A6yvJaeQWfqS6gJczBHFjEDA+ZabMEzsryjvsE6mgzWZ0eH8qitjrUN5Zhl
WIGuLGuw2I7+blkpUIrF+1jrzT39akkUxespF1WjO5Sf9yNuCpfwHz4keEIo4pJM5sPVXRWHFfkl
xhICtsdG77yfup4fDR4TFVVNz8VKKVt5xYuyi9UWv2J7/TGvQJMFgpTZdz7yA/wX7LCCdXWEaMb2
vBuvvUmNKcH/CJlq/4L6mEfhJfq2OewE/vEb6uIyqVpqvzqT0EWz3o+/6m/3W+6L+hZmpKT3l9Df
sKiebe10FhylijVBQI5iKNZxa3cdNI4qyZZtuEoNCTbQK/JGY7EbVMANtM8RHPK1LNhDDOUGbPh1
MVC6Aegh9y4CLnTqKR6P8KDEClWs4Yre6DiUKcstoe/WhArBOEEVe7s7koLUEc4gBPp+vFMNbE5w
+aVpDILYxQY27DNKNN2q2pqTTutYSrK1TK34gWqU0M6vfQQx4DYC9jbOwA6jtzOcF+j5g3Ynii5p
7oEoJjYLu/98Xj7xXsGVt7PxrWRvoTeRVxIjIQhWUO2SEJNMimvvTDWIFwibNLqETVnreVeaYZTR
BcvKl1Cs2Dvs/S69+QqL2+bRT8IYiY6urzdWcmtUj8mrcRSOFEjvQKIgn/Xi409H/64GM4HrQpkB
SBWQ5aaOu3Dmkkx5jLXvqAaMDYCRKZHuTKdYBH19kKzEQzXpiMkezcjuYoC6Jcak0iODTZTXJGtI
lJNreSZrn+Vwgi8uS709RX+RCjOZ3pAE7RaaR/jwHDvPMiDAHPc2wtAfo5XG7dggNU1zhweMcBrp
zhwY4Bdih1uX3alPPvxuR5XutR7YkyXEdfXmeWATVOqSf0lCfDV7J/rTNFn1pQpOdDC3r+KboDl4
SG6JlepacpNypI9SP/a43kShBxOUrpRgwLsPW+47berwdBk8PJW+HupDxAGWjvSOkYNuw5Maqpvj
vfXXhhPU6my3+thy7EcemhJAQv0j0Hq1aGUqPBpGZ0P3Vhu7rVVs8aMcuzyNikemC6pSlVou0336
BPT2Fyot6qVc2OycxrGHHbOzhsKzGXpLWA0Y6TAZEXB8yuoDt/OteHgoHxrcs6ShICLf/QZ4SmYv
4lr+c09yikL1I962nIOHqH6PSqki4Bo5SYAYfnBuWnx9SUokImd7ZaeEvzb3RjITDDraDvquCq5Z
6o4sI/ByHqXNOnqJBy3Tbvvr/B7gYP2XbJKgDpkUCOYrjc2eHvt39O3Z+1cK3OSCuqYGzwaZItoR
Pr/otwtrq7rYyJt+6tqU/9pND1SWmkSvQY6Xzz3221Qh+hvRFifvmDtGlTaA6jhA4w7fW5nIDelT
JgNdxRCq2iJkXVPKswu+1h4fb9ncxQtM/6l+4N9ZqlAjtE0WlxtT5SjNogoulA1Pm+FsHczL4Ymv
HJbiQRCOLAwsM2sO4u+f5WUJoSycayuepTdOSVBTidd4CDX62O2OvIwLUjr8rXj2ytm0gNbTZnA8
+ZxvLZGfIX1h05YuIlgm/VPb89WnzzOe11gsJMq8dE5CZPuhPRvLda/WUWjOPPu2REsYUG8EGG6i
5QxPl1/HgrSebnbrxiuaXltiwN4Mav0XEOrL603cXqxzHJDpaKVYxjhtFg5XDYe7wopC7Hj6jLqQ
Hdfkfz+JwjMDXqZ/fAfxIKKHu/S8fu5Zi3ExzcWiFFyKswc5vg8MwyG0kVtQQlj7Y/BbL+D6t+IH
i9oNOwyBJxEGKLEKSxmsCUqqmdC3IkVtsqkkGb4Pn52UnKro9l2Yb3Mj6kerPVROilLmmoM34tn9
+Xsr27Q1MU/DcShRRYPO7dKA7D8f5Onc2f2NRnL/8mR2QrB6xSW1JL73E2a1zBKDBlBgoS5f1XN8
l9BV8qcykD6FLrE3lgfzOrWMD7h+CAOU9zu7El7rQTTIMaNlYA81In36U3qWr53imhXIK6EAQ+aE
nMDDv0l502F48fR1Jbwhxi3GEHTLzliWb+MxWWpFvz8E44Tc1xSRSAFyVNfnmGf5DXJE43ttfkas
HsWlzGy16tj8es/xE+2Q/ErZw3MVHi/KC0hIpWrrwvt4ISZXFBkxn/CjjUjzrQR8J0Ci5vVM4IWs
ZOAHGQ6T2jIUFOgQaleNe4DrnWCTDXUJ+CLQnU46+BBeoJhu0l2Y5VBlC+ShRUK+KNTNYUYKEj7V
p74XeFzGXPTqcYGcmJGv8XBL4jVc60W87krTyTVtV4OSE9Pvfjqgk/E+yyEvr+sNGQVcrLHCx4fU
ZbfiF9/wyTq7gLvR0pdbc4FBxFqYmiPiGPkbRWKaZ/R4PZ+SPWKxvq/e36TU8QFBW6LGL9E+5NBZ
W0FKHOFgZ30EKBNURBLKbXyT+NtaeK6y6rqqsyrwHm2h1ZoRA3bRaOBIN63ZjObz6f9a7Sl8a6f9
Y2SHby58wmFNqLhXPvBTHdMVf/S/kiLbpDggF0cCSNaBDfiPHGfhi1O2jF8w8AXEnNSS9ZcsVaNo
rDOZePvuhvUaqeoSSLatjD1Vtq0M5hCLWWwWc/5GuXKi609n8xB/DFkiOvVWciuFwlXMacMAVEZ7
cYSXJw1Et1oIv5KpOTtLHA7PKeTaoiTM8skMpBRAsOZPguPjzIo0YS2sSUtGjvou75gKHLY/iY+g
1R+PugNm4OVb41A+ZqVfrbyGpb9J+/l4VkkDqrDDyVGnPCBOOdg1Aa+bDHkslmx596L5ubFYadW/
PNZGF/0N6RdtUFkwS3TxgNk4tTV1ERisysOsK0KlSlSCvSoe5xx9xCpW6TnQbbF06g5+2dzIVGGU
LGhXR7GxXHOW957RBQwwPsW4OrECz81kO5KtCtC7L8hWmd5anje5N5YnHtqg/9BrmFCflmlPqvrd
0HfaUrRCWg9+pWEJNuzhNeLGvMhzCe2CBTsGJiExqbq3RVi3SXawrMQ4+yaY9B69nZCWAt+dhoow
zGn+ug8rrajWkjBWasXHV4Iz7YDkY6/HzifOB4MZVbGbPxV2DBoFkTHHbJ/o41aXbygc4R3E0LXg
WEmrsiUSAjLd3GB0CzHPp5hJBo/60tlPcM7wP/SW7OG3VkANRpaxP5/LQHPARIQ2bGmNznq93w50
b6ahE7IX6umg2wYqrcGw79LbrlnmwMsKEtqm5hjFwUXQtl+LPY7jImwrwOTGhzthy12sZNKrbuM5
7KpDXKNDirlTjJibxTtmE3aVQZvJ7uS4gYijY2vpSIBq1erRByJPhmn/UcKnClHurlIOnMdza16n
Rz+uZ/BzK+8iphAv0Kpm/7NtOXlM75X+EBOlbC+5G2gMiqRpyOCu+zPwX5TdQFiqYID0Ydndl6Ju
73xj/Jcz5Z0hVTubB0RbOKn+qRFSOzi9MQ3IQmzyB0EKHPOItzXtOuAeAuauP30P1UKU3/kZ6bM6
ZUbE33IS0TNIlH77im5Fe0c/8Z8T0D4kbMXPzLdyBHlPktK+bnU17q0LrEW7ATRBP8S5EuFhXPM5
Nw4cFeuCuYXPavYngnXb1hdhCl5Oxt9LaoQc2S0yVDgjBY5VCKW8eVBGcP1TmQrkF1mkbOBSlHa1
oTVsHj1nzant3oB+OTaoXfjdeDbuzTXS3AblvqDp+ubqHAeDOlwJTCrVQS1jWhSgaBWtVpo1BVyH
ZEO/d+OxYosbbJ1sgxuW3lq1YcLwcca8osYvVeen17ZV2ju5pdASniFtN0sKkTDgN8KTV3lH6hfd
9wU2vEChnxGVOkoJnoI7S1WRcFspcv1d+SKBOtq5cgny0NsFM6KHYnA/IATPfTW47/zoOkBrxWsk
umZjd4sSV6qtPGlklktRyocU5IOKHRaH8bPikRAuu8m8H1uoSimEfVCsoNXYHgtwfP5E2GUG2S9v
hUg3BHic+WIhy/Yyw8ONJO0zK8JjHhojm43IDuOfGoIuCRBKfhVy4qnjKwThP2HnrkevnKjNuGSm
sHJpNmG967I5tFmoxfVsSzTr33NC2nnfs8X2wdcGqGC2gr0q4GRdPHFY43GsDQBcZBKsTiOMbflr
VPItr/EsG7mvMT3n3UmSfIDjj/W4KQ3xZgH1XFs6+G68r3F/2AqYOPbTdn81rPPylD7+OreExBDh
Ks/o0aO3dtLEY2RGYu4ZaQCw1i4JaneWYSF6kdMsmxxqAURf0J1sgozKOapBCjOK5TLISSWD80vW
ctGTed6JIHzjdtnbC6/nXkeCA3hEj4AEmBtMD3CwDemUfcEn6saGBEMlHvOnauiD/tXHi2Rl4DNl
5nMtRpK4UIMRiy8Z9udf/w2N1be5YXrsF1Xk3z5Ur2LQn7Q7p5UZDibs6u/MMg2QXg5Ic4T2NPPc
AUdQ/J9XiRqiN5jWFdBd46a72W+R7kAnOV/HlZAfI89mKNoyG3NX8tkzaMHs7Es7DE/nb8gwN01e
aB8R5DiAI/T+rYdCzSQwyfvM6jyVkC7ZgXYJzFstvZMPpYmQvI8REkVYKnrHBPWn7tCSO2IG4Vi8
EE+Rb9kO2L2SFuQy8qU3zJEMYWB/7t1fJp7CJQndh0Jzr8xFtT2lzvInx30cXf8P22E0V53x+KyH
dVmnebEvjwzeAWheEefWrrxFaqZu7DdKUFjzQWc9OMLjpL36pYI7HRMQrbBJNTBKZVtORm5HQReL
7TksYCPlhFgXYrPdELdPzeKqGeIU1ZZsO7ftAH5mth1a7hyq2zAhgcIZvJmZDf4EmgTVJqilh/jz
LRjIOGh9QD+Hka0Y9Wyv3fcAZ4j+fkpIWjbJQRnZqpA7dROrLzPVmpwws4Jr1JsuHM1eMCVoA+nD
Fmdf/FGTIZLcRlEC8wXBdP6F+9jaxV6i0W7ymTGJ8UJayk/TOjEQLI2JWQ5oyU64syp/BRQ3NJ8E
k3DwGh9zI53xDyIIstM7/zdcQ+Ko867kg3dJ9nmL+snZOWLsFTkq28uIMJpTFsB9zxsp3/KYK3MF
9lHLU6szMMkjEDlRu5HubUXRHLj0VA4jwR+3LC5X2z/7sBIE/hNCyvbizbCp+nFYnI8QqSwEEaTN
T/1eK5uX3FF7X8VlIorfW5OQ4o3Hed7RpR5OyNswePtVNHEqcuhWLg2ryVZ0Nc8Y59bX42WDqL27
g9Df2XcapuhJtEcwpT3kyc+TM8HBlpaIN4mxtkLgKE65ST0hAf/AcaVF2b/5z/LpbtunMzZa4a6T
PRf9IqET374+Uf2D6YvRBmybEUk58Ka1A8A6fWm/153mXr4nIWJvDbJsck2NHd3NH/fbDeYmJiYJ
XpljNZGnpiXY8F+ysM/kUReggq4SxEEbTpVpv1/fYlxP9F4ETU41vEm71X5Lg1sq1fv7n3xE8Zea
D4a9vaMq4sWt/S9u39r0FOxRXMe6nXc/U3BQgKq+3qaCfjhDx0mXfZkBLi5vvRSDodpD+DBA6Xuy
cAStu5Q3aV7C9FJM/yKoppgbLo4/f5ANvwOptnHWjmVzEEC4H193Qi7ecJkJLJshToeBCUyNTWgX
piY8/zobhIUoq/SWp8t4jddRFUIG8dXp5DFWS1fG8RvJSL1wRsuw0yZ07dlyd6oy4yaXIvngtS8a
yDqALuwNuyi5KvZhCEBjFZIVMjpa+ZZpSyMLKOQEYjQt8KkBfYekEHTAqJKBcGpORdzM1WeR7WYR
KN598l6v9BQ29/nr5cdBVgFS7TUX1PBJKYL0K7/CQWMV2CP/vfJv4PBLVl616Op7rb1GiAxZtSGa
Cc0Qw2GMDFGClhrVy7rrritDpI59QJn4BI5W+Lljbl94CeUi3IG0HayMA7wlVciX/igBUswh8mxL
hE1zQQzgvCTHkPEgU9D9PeEnNun/nS2XRVq241pVxl+pAeRHWhDupnfZXiJfYaE1NJOJutTFuxTi
or4S9lyiGoc7K9USCeLPy9Qow3NHbTYk/WQE+soUyV9BMldhk78kpcn65aSIEdw9wQU+C9bEtXEo
8QqSbWbv/9hz/W0x6IrkvRMfQWHL9+uGvGg3Grf6lPGVwyCdlX0Bp7M9XV+Xulcx5ggskubVJxST
JKrKs9NgYuOjh3mz+x397jb0crV64fJ2ggvhIWPp7Xlg+v7kaX6ItpMLOcBXH5V+sqOIb8kQgyR7
SuYePIT6dpBIVyQrkvr5N39eHTzPanbHXO6hMmg+R44SF5FU4Vw5V5s47mKkC3AloL6c/Y+Zvx/P
dUOLDhT+92OxoHhSdITscrgDTCXrbiqEiAh5bGYNkxyTbRfFZyCaMuxGZRekhPpiEzWszUDA+Xop
7XVYEOcw0w9PJSbK/gJOJAYjg7dO/mQpLi5uR8azpvfWZKM35KaDJjo3Ezqubp2P3A5ciOCJUchP
dElbY2gEnWE5U+E8HqENGTzVQ8q4Jk6fByGsE6IIwueSQeqxPAtSzc0FzduWniYwUQNPIUSTft+l
FCe2LuIWmyyzAAJ43OuFmYmteEpoLLJMr/2C2R1DXP8Fi2uO6BER0lfj5vzZlTndU0MtDbNmkdkn
iNGpFLnfx7l8g9ybG7kMK+uwBM94tLLTfQlfzpGSlkJxCNIa6BYynii3Fy9nmiVXTTQAzVi7Gdlt
gUCRccP3tGF5O9Bw5KQN7uBUO7qXhIaxvy2Lf4IkklDIx4K78+q+6uUSElJyAEYovSTpQDEzQOSU
hsN8UHzcJxousou33D3kvgYEOo029vxvhF5ECW+QgOw1CYlDiRf5OnSMfef+eJnZ5O8S6vws0svE
fbH9Sd1d48OceF8I8/d4B3VW5OjNLZlHdnsdv4F8fbAw3SHFEdSC/5nnSK9CQsIq2zw/NChTJv0t
H5lA52ObHqVOZR0UJTugZNmRH1Foosw+ovt86zQiopsfxMl0l0VwLGAHWyrcWwjgIvg6nDjJRYUk
fn9zlEYtcTIn7qpf0jCfCi+YFfR1J0ZG3sSIet2FgKZdohBSrYiMT4BTmqcQ9CpMdu5FbNLbluY1
lZwQDlnmxVbGHSK5mNlGS1X9Jyqcn+iumP5OM6DEp7wqh9PRc5Om2u8pdhXwLtKQBkMGbkGBAK5m
jndfdutVNzqeifjyje/FHrNXn1ae8DTVEOjBcDJlLgD+cqmUPjsuk4uAh7nw2GqQKQ8UwgQUWCfO
YFaRDYzib8905KCAxyDkbVxqTUbnRD+NQacILMy8PNx8mjgiwLru03Fj3B37NZNr6A3wjj131HD0
tqMDk8t2iB82W8OR+lcEDfHekYSWriCT79vrrejmMves8R4/3lbqBH/mLEA3LukoKFFfwB4Htt0O
suOTyciUNxfwuE/Pr8nHiZE5EuOPXJq7OwAk7q/o2tj6JIZGzjRZNgwHDKq8LE0iZwQQlXTp315a
QGQf6Ch0k5Q/OZMZhK0N7yBSbnMUaHsECUnP6FK5DK2ADf4RxQaClLnX1nVNtAat1J+ym+zE+fC9
PYYSyqVuv3bo/+/TkoF100rtht0CEPHn39oH2l1ArtM1CefACIMbgQ63JPYbg1BDsVshINR8JkuG
CTWY8miFp4HczxjTFP5DV6HgfNlWrd8l/PEnJdsBEQHIvclO0ZLt3K66C0iowxvdTbfwoSDgR6E9
RrSjPysyD6RVOQSX/mdPfPbZ1AYMgsVyXkZ2jKCw4UCA4Ie+Si13z2QW9Q44W8f8/3+RcKL+diTz
enm10rRQk/M1Zftgbg6HaAhVAoNvZqR5XCH+f6XOJo7CwVzt+6nbxESpkyHfQkuvkmSfk7gT5Nta
MwizTdiFyb8qMAbV2F2y7oGZE4tapogqw0kHH6ZrSNSbo+C1g4ty8QWXTu9OeZCw9IBl4oopN7Mb
lEm909CPEMkwVHw9pgQxK9VwtgI1vFAXnLmEJsk5OkqY+X9M7bFbvjw6qmppnDwt12U1FfFeVct+
DymPLpgrRI4zYgCDHZgS21+i36Jwo9x6vPhnq5WfBnm8bSAOIoZAS4AJbnKj1A7O0XCDVJjkB3Qa
SrbvnDPRzPD37tUrNt62H9fsrtm1Lku34FZx73KKdx6wa/mnbwxJUkC+HMxYth9ruf+MyH5fQrwq
44nt+JO4x5n+wSu4MI9wRvppR8bt/hrUhxrpSh2gnx6AIM1QtjiEoT2asj6VEhnKF9FCQt2y+yO6
al8d6p734lxoSCekYRkxe6Hy02Uu+4oF+wMaTD2QIl0V/pTH3RmrosT56/N76Velp1kReD+Tg0NC
+T0lhcs77lpvwqHZKE9GkQ9qV/nR3sOiBY9YgYL9gCDdj9V2OcYNCN54/KQlcfkG8X0rlqBp7sw5
EfC2qysbyDgKMK8smI1xG79a00Pm1aNJid8yhrv8PS/3iQs1oOm91sDXayXsMtwCv3xxefcBM9YP
KLCr8hwuFPi8fjFWApIu/ctC1MAQ/Z2zH60SjmSCiExvWhgjPZi10vdFFHjEpA/cDZ25sdSp8rXy
VELHa3tXeMGf90ILg63PoajqehiEHsTqJ0fb8ZTbikIGlxFvOT55stPZs3UNXhCS/S7I+CDjN4LW
0GJCfGyJNUADqHZcJL/rI1mNwX0Sqsmih+GlhRT+4O2nSzts1W8B2X0OT17Xrl0K85NKHR8GrCln
w7om+6oLPtUT/UQsjfwOPQMifthBjakxf7JqPH2UoSbT1w1Ep303mmUT/H82+ulY2by7mjhlXtI5
SDBC3G+uoQ9pzP9nyHERP/rJ+qYzVpNNQayZ9aVOye6g99xWl9K+pDd2uGFR4uOm9+P5B0eb/uxC
E88h+L2A5ezM6WAaPcGk2H2kCUKo51rdss3aCkk1s0RwgE7v7NAnnHLplsyuuxLEO98ZGYnnsljw
G0Ic0qpDZah+J19rWauTlXOUVxUQWoIzFeiEpW0dvpy8NaTts0PllaO4zeu1jA7sH0SY1WI++ud8
a/7h5Tlvmuqyg+88QVgw4YNOZbkPV1BRnLQOlFAZnshSYIZlFZJBGxWJJrJraa6d+imD9hwbPmEF
ERuh1xHa7ZDqEjcAJHgd+20xHamfEaigTQRhIHM2/p+fJrkeumXoQwv/7LVp1jk+qrgWgoeVncno
yBvOfN7BPg5xG7MJO0r51Sj0J6IbqYXOKgPJbDiaBlB4TrVWq8E96mZjHTZadvIUH5rv57zU8Oeh
UF6YfUS1uzKlFlqvycjH6p6liCh9ozuYCqWtPcSm9yxaEg3y8Vc3xKSQVyyglpKmAcNPMcH6TnaQ
Q13uQ+rK0DEtougIScBAFngu9mDAcMCQLLn3Wx03YMl0YflKqNnSKo1RdCP+k1JZp3LUKV4HSgEK
c5na3/FouV41aK+oCJ78i6ycj+EV7i79iJasyEWTYamC51MJ5FtIRYIVXuVaUXNZxT4zWYx4hUEU
C9AFFV4dqRsfOmpOcKF8yrYVGYpF5V3XyN/qhSdzkTF5w0OmCpTL0EH43BF5F3Q0Vvos12lBuuHc
QHIQ7YP0oLFzAbE5YfKDjyJtfb3HtKvQKH2b5crZ4Kny0COasHjlHP5S1JqAOkb3q6o2oaAvfnCa
rwo9sdHTvQhNdcF8xMOWJN7iDDODN8OdwokVHq6Jv+iF9Xrg5J0EfD9vqis4goRkAKoG1t8uIZUZ
PcbNCZttj3VuqMjZ1xUR9sTSLmzWsP20MuNGnkEP6mXnuPEQkMga7vCt3HY1QfMxrWKFvxgGKKzt
2ZILGmug6rof3eNKW4kXWQ9AXz6xpvoJx7jVpiJPs6rtHDE/Ti2ZA/i8m0rK6squDn/mAvbKiqw7
qERKPjc3iaZucteATzVLci3vadfXDdRUA5KlzZQ0pup/K6ljum7PcNmmQMvv7qIMKX+e42k5PaiK
ASeN9ZGJw6vbvkChuVRL4HGQkiQ3hbvFnQ7X0HuZ7DrvfYY9wGHjKzbMD9wTOlJ/HmjLTT4Oj2b/
9uMqjinzIFmZ77q/fBJGrrUyfpD0nRl6RuW8hRjdyhT8JlpMwchk8GuesdK7eLqDLToZnWeC8V/u
nucVUbDyPwOCrqt1tKbB4yiOk+I2ReIE+emZH0j+b4ZtwlabBigxxUHCJ0CcxXf5Beo4sjHA6Xca
nSr8xzP4rZvoJ1clQU9gUGR2a999OkkxjHkxKjSEgrdmoOAIZS7XLHLgxRW4Goqs6njMvGqPpJKB
BDT4Q6Hun/ItjFVfLORXyw9cpGbjfVqPBWMa1CaBlwB4WAcoBqVaGsuAgMzOIAUeMzTKUEkT1MPi
hHInHtbnCFk8FMFlRPwKnBaHAxabSzYqlg2JwyRQWsokCEpd6v+iArTEbcAJX8qBe7PDSyyNf4UQ
RGNPT0DD5Bs2KPAsVdyDkV69z9Hlt5gofpBYw2hUvjSc6jzH3rcK7nz3I1nhmvjt8Bnvb1rRV+R8
CEodlluBomNLQ+FcRBKuhV4RQovMDZ3pUZFnGDIYNEp3kU0vpWH0ZrojzxtQ6BxF+eRPoqX5N5P6
EwWmBuJle2gsD4+d2iNFjACgNO1jgB8hHY8BAL7bDhHhaFHaQS0zRJ/nZc3K1AJs89mfsN6FQX7v
dqCGvdEIe+QaVbcJRPWsoalctRJG0sMPEJG34P98z1AS5HDV4ndQiaXpNTdmeGiYKV95BygOAL/o
YM9ceTBUKGtb+2gYAwRl4Z6RNNU+mdCX5RdB2tQVednqtTBwaBgbhMCanDsQViGphD+wrf5N9208
jZLXvid/JrtvjAc8Y2xgkH66a7d88gVoF34crJIdzt1auGhsz+QzoNILhWXv0NUAKtIlVMxjSqKx
6tl6xkSadIkGG3bqrWYqaVoa45d0zBI5PxNO2tB8dCBYfjDIeuGfQOD0Tq9tC2U8T0uv5kq59BSn
XuFCstZvmvLN7lrhrmqBO9awqArbED4Tw4wmcTigTJ6P+CpgaWhOXwZd1XSEY3+Vkii1sObg4Sf9
JmIeAshCNIZ7MGX7LsD0BWqRPpRuQgNgqLuLeKfSohlgCsb/VqmElmcTKSdAjT/I7jNzGCaa2zys
Yc7hpX3bXZ/8QjkTwJtdATIEWVuknePKv/sWm3VdlGMR1WSjpdKss6X1Dr5dxa4NPxYdUPLve4/t
8tq67EUCR/9KC8W5LQ4hqRaVdNgnRfq6laEBwLm08k0YHRbpLswb2579VIXobriU7CVBm5gqyxpX
n8eP2tCKB/34XpJCzMOgs37qxro5uKVAcL3EMxXSqnVPlIZKttF+ko9gOxP9nGPNWJkHjplsreV+
scp5icXs9OWxEqpejZv0OKtAd56Vlk4yYpDQLeGpLrTvMMRaUNzniatXWrY/ltKw8DnpS+I2sjEy
5lmrhmIenjEQplmYQeCibX+MYTo8r0nGqq8pbkxXSWaiKupjO5AgN7STY54p96WhWPfcIOs/DQ0V
IZOe/AcMYvgSnSZ07OG15qpvyfuaFl3RSPm14K8mIBbPLaWM+dlR/u5Wmn0EBvztnnhX1fI7C8Fp
cHb+hH1WR1CrKVyic5KMUu4bIQkY/0lZqL52viOIIZMDyI8BmXPM/2a/dGSLObPXVaKjK/CtYCOt
WxcQXdVURjsiBmKyLsh56BG5jSjCZUQLAYfixR5+uZrrJjiFwQIZys8AjrEfA2uPJiLBhFslLS2X
gsFJlnq3qh8zT+LXDtc2YYlUphBeooDFmhJqJ1tpZVXzok4+RU2LZNae2eZA4mzly83MRtJLObyU
AjPfRYLngsykGtQpzMxAVE569Iq/pkzoPGMY+1maiLm2fMoSPViZrvSaC68VkBPRsNQEAFx6rOQl
sPUOnILAd6yBrjXFzjQsJSF0pxXc3wM2uFtl5B7LNdpI+besj/1zgFO0zudDrrwGP3j4uY0ikpto
gZ4hCaF7e4HY1nYdSo3ocEfT9GlamWejateGazFolyd/Kd4GoTdBJmsE1hXCeFR72nUFoKoH8QI2
2JtrXgyAvrwBThdwDQNpmOBsgii5XIoxhEdM1lhOmw8L8JgQm0+Er+Gu9S2+obTR0qkdhdILzN++
ThxsMRymqbrLTKOog2HHIAvaxtWPgnHLP+v/K171koqkeWdG9M8NGyOTU5AYJwhadKAcikUDTTfL
XEc/sFAmDbDJAClPHQjcqyxaJY0MUiFQXnYW9Jy1a5id9r5mJRRi3GzWWZyrEaeHEON6Wz28iVBV
Lz+upqb0uvHRsFEfruK+R4DswJ93QOTeFG18Fx8lj8k14ejPWvbgYFckpw67kyBiHcFu74TFaOve
uE5AEBLy5s7WRr7bnNZDZ/i9mGu5Dbvjh+V+K7/TvD2QjpdfuZX47ZucrSZj7dgo67iKnw6E41vW
VnhEX2jeYNskMldCY9jgLSBbmOoStqliROFxG44GIZ2KHMrEdmldLBT5lenxmo53i7xAlyZIrjw5
VfjgcKJzBZSElK4/XBBjboHUasUBWRA0DYTOTnrcq/GiEEWsF5OJnVYmPH+VSszS0h8C2MQrZTNl
ZYUWBVJAnuSAlLHZrNsCINjiAVjwSAQFzLqUkcVEd1mdJBVQP00uRXrM9Uf52hv56g5Zph3ray8q
M5kNyy2Zzpa/YzymK3cihegFGNkVFreKSHM4Q6OBRsWL/Alt2RhZsag+wqHC8ETJeiqNRjAAhtyp
o2QBOHMs+MgX3nr6PEd61GCKxqnWwzAJKYc/hjOslyTlS+i4KnsYz0a2fYJw/T+ezkW/PUtUk7fW
zLOXSIXR+VfbO0bv58Hrd+LteRY3v+wjU+sB9dUp0g9rf7ExNnhdSb5z698uRlQCul2s1gZpex2I
jUhT/JR36MloDopNFRXd8zzTFNvKBuNPm4dTChIL01o4PigRgXwh6qb6CXZYDRIt+WjQUSgm/XZ/
1pzQgLuLgyjTrOqcKdMOvGat8VaPc/Cjf2TSDl/fs7E1dLSZJQ1iso/h+H/MN2J7gZaYCsFdr43j
pX0jrvA3i+dBL4nbWwMBN49DCaIHIu3eEvfsJxtRUpax/diz9J287hw77xAkj3nPnG8NCSG2lWwN
YA2h5MG52DKuXcBoMTC3R4INGSIJz2OYFFTaFp5MXihxwrufNeXO/Bp3eaQ31aP/M4POBcBBBJYx
lqw8zvzwYlJgMTHk1o0LFya5qxMhTPmO48v9oScW2CPJUQEe8hYdWDf2Rnw1Y63/EwafXnYa4y2z
jc+m7bpV/8rTmoc3hmT1An+WMF2dygaPWSlv0E1uCGUHYrgDRigU2FVSo4pwlrTnIZ90GiqqCsWD
Wkyks4FPRyHv+upr4KUJbsl4Fb0MiwPPKQ/tClt4A7Ytqtnn4gh1+ExaGD7X9ZJMhWFI+OmydPp6
tDDQbkSeXnULA3OhmRHTucu0v5SfAhDXqy4QcfHwyFQuSLpk2EWBoK76BuiLP4UYKmKGVv8xFbcz
Cx7QmTKMrS4u//T3bnMB7WNeoX3r50VYawn5nCDGltTW6XqYww91P0td+ZNA0RSeHNRZ/BZ3qRuv
Ee4nnEE9zjKKUKlU4arp9swD5tPrRTmr5tKjYkUeeRct35yWSYDJjdmNkZMizuI4yvyxmgd6Pwni
0Ugk4znyoZrTKxa/e9Vd4T+4s/xYqPAqnMSKqjuErfnc/fB3hOTC2rzHCH4IkYotO41HbpOKmc0E
NO6AR5/qE0KEriYroYaY/xHjmkdvAr7KzPHF2tC8h2pN4KQ1VtqwD417s4EO4MDZz2MXbsR5TSK1
pkQrewtjFOrS4r8VhaIE1SJ1R862+JvUGCMZWHQqZfUu1ZXUJHCnizaqR3iORnk58YWIPTJ9wzsY
QJGDvKUPpsZsKGq6ms7QYzWbjTCH1YnSivU3D9WUbFED+Xl4r3LYHt4aUgolNaTqQenJmv05E6kd
m80DwVzG/ki3q+sWFMhv3n9VH53Sq29jGJ0qcwNQ4uVYryJqZossdUeJSlv3mUjxPDKW1uySDt9b
O2LClFfuiMel75c6podzQTQTGp9cEHnaU+3LoQk/GRMDDufLk+tI9ba8Zg5iLk0yggytGoDLGwo+
6xo1UUCwWovUTbX74OJK/rJVrOxWzTiHY1I+IYWpMkiX5tr2RJZ+XCUKELTE9cayGdLX9W/ecuQ7
Wbbh2qUF54l/d66kCVa9eST8YSLRgXGQgsPpA6mzAtek0BcU1XBWU8T+43mSbZ0oVfLsObwWSc0A
8Z/nbM2wvQ9PuHBFSk1iB3YF3XS4y0i5OhcpC5V5wsYKLIv6ywkWcAA65R5iMaPwUzTjOrwqQmwj
n074V42ndq0EHjRoojpcZw90rjX2jWulu0PR0zNozEw8jbp7FBqBJwYW7xOMdDq/e3+6p6vwbfv/
GZ5ld5KPKVZTM/I08Bqjcy0M0JARtxGy/g7F3pXfx/e2EClbEETuAvKjJs1+iA7QfGsaAQ7Pqf5I
f3uCUDQ3mj+6aoDWPH11Bysr/tO1Tt/jtlUFsUGrhXRre+n/MksW+EAKcKdcW6vbI9hPeCVjwCRr
VFKUWRFGskQ5IQ82NnnXsNFXgXG/Xc7ar+7cPjAqD58/iQtm1YVtuYo6gEfyOM3AZX+jb5KCv/6y
85Pzu195lD4gfnc4KdS6NhseVPju2QJqnToKEevOm3xYkjrSgIHLcV6eeB03YCBR4AVgx/RHWnFR
mAQcTCLBSOJGyKTKzewS2e6aqciIpIp+yXSSZTYGoH2JlRjaTavqMxfQU2uMyTPRyTl/+a1l3rQm
RI4ABj7Q5sN+HmaQZB+H50jPiLvO/ZmYTt/GtkN7aaVZzgF2IvkkBqCN26jK9qLgdQ+VgA1syvDt
7fxePuYVRMEWP89tLip1yLY2X8EvxXf0acaGJ5+i6Ys5X6Gu0S9gDZJzvCLT2uvTiWewxFhlriny
tfyCsNq67wVS56ETS1roladL+WbSM1HfKjKqFKpyJTtp95PNJ63YShDSoJI0oOJ77SeKz8P7erdE
4kVsmc0LHGX+K+06Dmmb/I7EoRsvDqWzGBN9d/tl8cwBMAtWU9GfgR7FvJJdR2mPj8OdfqaTm709
5uYSZts9U+L+71qdlBdrXLugwxb/W0qBoU8oj/CgMPF3u2ors3+tq/f4H6pSuHSxLPD3/eLbhghx
dPuiuN6vT0Q32Dn8y8eN2Lsol7SVtaekCmuTwFFhiCdbKCs5AcviNoAEHEi0Qept10RNzi6oxE5g
gdD6oxavQgWlClBUzA2KzgFykkkazwCpG43P7VSGgi2ldQ6mqqjVT4PYud6GSgr+ShxgUvg9cEG6
AqamXWQt1bNieqdWswkQ8E8UOW988eTYZ08bBLEo0NnhAvAhnKssY2CBAQfsxd3+7bxMXMp53x6J
lhwXqpTZ4AjWm3y0tP0C4rFQUUchxJ/Vd3lWylvqg3EtCa6BQstJQp7yPUAS3KaAH9YMKqcHg7sJ
UF5ZSS78cu4ZHFgQR4NRj0+3Jt9fgI7yhXy97Y1aBHAcFdhwzoI+mIlo5Oui/lJhwkFDiXv1zxsh
qfPvXJ8rMmC6hDLk/b34xEE7Bpnrt1OjKj2WZEfUVWaFNwMV9fPXZRU54ugfHocf/mhpqAQXGSXU
4byg0xw9i8Xus0RRcCeuBfF9unXmE7nspSjfbbq6VcFXXR6ZaNKgxTQEYwVXq5qWpXpCwM6+m0qT
oN/58MByrz/lIyAbwVMYOEO3Uc1ki5DDLKgxwNAEEyxdYCfUr1fHHtPeD4Xpug3xWUBTyHZaMAjp
WN26ND3hYelt8c9YoP8aWLuJZPF3rQL5D9szJrN67RIPt1f8sdqRn5vA28TcKDDEYgv7EzHaaGeM
YN5LcRT+eoDFXaLjl4LDgBS0SUhlh4ZQaqsEI695AWRMXMwJSu4+lvFqRHfia4m6G+BUT/bhUfx7
yxed7/01PcbWDJOo3oDbqAPMf+/Ki/4/EO7SdjVSlgYky4os63sN+jdoyq3txXSy9qbqyuT0gGQx
NjdF3tS/8zcxFZWZtqsT0i0KguCWH/5jKzZ71XNsydjgEIN5gBnBANB5unS6kFdL6L8aK6CABtxp
0qdCfpvM3LX/3UFd1WuyhWrMSXLPBf5iXXhJ95TEjhmfSWF7IGyNPGoGBYNSncDsAbjtsknzpP8l
KBL/8Lr7w2JJB8H+XMqzoSSZWLOfAUPesHcB8Lyjlyae5IindzNpiKp9gkA06VGH121WHRQYWY4e
mJE1FMW+q70jl/AxZsKFiFHH5r5Nm0WpajJonf6/xJ57pZGESCuubGTuJUJOkVNljkQob7YLAkWI
+N6r3QnAynXLDrlL0hGlR6QrGyZkws+f6YWWLY8N3lODVC2uwvU/MzdLzTrpd9cZLeyjEcTuDboK
Igj9gyGfPoaJUcXM/F0rAeB0S9pPeAlumnbBx/hKv7w0/qNX0uXFMW81Pa7PT+nxouZHmyjE7zyM
lJjQAJ8R3Pz6yUDt6ne0l74emFenYptnvYLcblUNfeaWnd+uU5zVIj87/RsHrot/kcsPO3KoRxmI
Jil5gAwRS+ozuwcg92dMu+gkM+O2IQ/yjSRlK2ZV/XiMEnV5Tg5MGeTToZs+7okjXlz0vTf+WEy6
18RqgiA7RXjcAaIMNaMVSCFN+06A8sIRh09T7dddCwU6L8E1CygBEzvOY+z3hzdeuw+MDShUymi7
XTg4i0Rt8uk3J5Cy8O1FO6CY48tg5D/sVmMQTq5iZIPmfnEETPbXMfOjbln5uX5Wldcv5h22vvud
RI6DfuFlguLIv0fc3NGc0PBh+MHi7fnYbaPzKEO7NGd+LSULpF7wjdERznk5GzPoMDfCQZTG7Sh6
6xM5ycSBn63r2EHTqO3zzziq+f+4SlaFgi9+oKasMNpo5vIfPocGuE8RBYkK4nuSjKUlmxxgUoO0
jHOTBBvpfnssDLJIgEbbniuC1+v0g/OOIzkw0CyypF7+E/EjK2MW4G1HPgqhK+ekl/jgnGXNjoTj
NvZVuz0mZmbGcYkhE4sMjNGzNTdUaE0Ff+Qf6XQfRBoAkTE3g7Y7ZYd28TGDeoUcKK1UcFa+E4U/
1iO0GK7IWMxRisiWabQXqtbjkZVp5qRPwM4621Fcq9M8ebL+qSRExDAzGA83gw6qUYtOizfMWJm4
VQUR5+ruR/f5zM2WagQbXv8PCR8wl2MsU05Tk4LyUe+QrSVzXgs/s2pBgmus4uijo+qsy75Wwf2J
K3xwWeziwYyG93Kh/yGLkHhBhIdSZtxH9L5Jef1j6FFJd20FD+2rmK6kWIqAQijqN46nLgDUtzpW
u+xmbM4/ZCfSTcJhZV35Y6qquSU55JuJTbOffcGz9MP2tjGNVYVbZG4OzHfFPJPKN9kn6pqQXmzH
EyFNTfcoh5bCK+rdbFirl1MGpWemPkS39eursTOHHndjYHuZAIQaF7ist1BYqH4VFDCECOvvD0kf
+Ps4RAbML3Ggiw+VrAD+Bie1tnsJyT9rryhqtvef/aDU0oabxbM+5s3iOeqf2DsOoZ58x7emcunw
qcRKse6G2fCpr6nKv+LQ1mjOhRNFxmMmuVqmnlWtXjmOAD1YOEsznn4GQsrV9IRYt6tfDGlPy1pO
Bqq+l9PK4kAsOZuR6EHsSOCGJOuF9QkXEO4fDcd4s2l+CDCbCZ2KJr0Y1F4SM4bXrJQJ/dVkU6iL
2ObtfOGEtKOm3ibwSuU+nNkcRVlFl5V/5XwTojW+rgSfz5l+S5+ra+HAfk9A6kC3U77uep2Z5+LG
lHoByO/KqWHJmCHMf9HacnylM36c23ptzPiNyrRzTBO4coY1qcelKhbfXKAQJjo8NTwCUPPeBeHX
RoVbc91aaIQsMGAdCO8tXqCZFGANoIQoPRdhuauVZh2uZJstZWBWZoq3QlSgNO83B10TMTi7x+Rt
IR943/C0tBO1WvXDu2NMgUuRup+i4qIWTPOCbC3vcO74N8Ni5NBdGN8513tMiI2mhcjqIWsjDut1
ivvA95dd4bkqqhbTFw+Cc/HI3ZQMRm0jwn/noZuoRL4U1FoiWySagFr81JAtF/c8VcJpKiGVGZU/
aZF0n9/s4NcHNFvfpodH5citgdLrVDIJIoP3NYJHHxMDwUavMepK593H048daMkImkzqlDzVy5Cx
TwVDWxhSJj3IFD5riwqC42r/K4ukLKJcVgpAPRaGBDIv+5+1yMqVODYgcsgmZeYZY/Lr6K+/M+Kk
v1PFrLXVSIc4r5AQvcfrXdXK02eF/tdS/l4kOX12B69UzTsKKW6zD7K5ydPQAEvPngCtOBJeHy9T
EHAgU6O2lAJfAhZCBh9yhAN+KynS4ijjksB7kVDJunJ9SHTLa2GOnGyn5zJd7aYEnQ6TUPB+wWEA
4gsvcciNG6wKEuxr6JL7/APQ+zY8t2etedZkK5MQhd6Ui1k/yjGP+wkabuPbUOJ0+rqaOY6UYxcu
Gzn9SdwrcqI6rXraz+13XIzlqpIBX4cU8wdv2z4/qIq93xheIze2VaN+1ZHF5uPsy25MmRvXxO+X
ReuBagvGYX08ZQ9NDXqJk6FTjxu5MlBiPf85zC6eLgzmmpSYqYJZ/qERqzH0vwo6VumcD3qvkzTk
S33vE+jqEAa5oJZOJvmwlsQv6Kt5j2Yfx0nWlXRCaDoVK/yodJbwmta6bv9TcXYZobadAvWcPdMZ
COhqFtXF0gqpmYfLwNt6WYXAiBlrdaRIf9PWSzRRVbtsPP4PC3XuTUMTkZv0Qd7+JyGW6DO1J/gE
0sd4jY0Qw2rtUPYMC0r4va7/L6/WCr886Jz+LBkxYTb6ZN6EIxAHVR9RDqF5JeRH23dNIDhQ04ij
+mDdqgPQMOHMrCgv902BH9QusQcxGqIElUrwLBmeieFZaaZYIOqs3uaiVv+N3H2tZHi/TJFDnaw7
qAVAm10G5K3z5ejfBjB9VWaN/fn6MO6n6jGuD6DNQPgSxpN2YeFlTKLe3vTOo1aS3em8rW1caHXd
ypzgO0eP17WBt4SxNPh2dAh1Xm5+8JsaZZY1fJ5wR28jyu5oqipIeJqOHX2NJzLVepZWlwOSM5WQ
AaX7od+9iqtqpNb8sQl8MdODS9Hx/JVjMATWB3w6alRVyyT7hxqtJhpHMb9HMIsbo1UaM3h/0hRx
jA1Q1Xk9ilfeb861mA8TBetqTF7L7UbayAKDwZqKmFI37kmO5fOvw47yXLMjqGrzjmUPfQHSX/qb
E1QtGiaTlHgNL9lT1V5kekPWNYPMdgb+P3vzKBhvP1A+d2W3Aarzk0r8Btf5mYbP8qCzBGzNC/fZ
H1V06Fd4lt29x/n76WIVP6XjyhO7WqaT5Iq8CFSLH4REL3k2Ep3Qft+OBfOdGN2Dv3VpRNg5Pwey
mvqeUNuZz7Dn8bqDsip+gnjbC18DUK6xe2aZTs/r1cAGeGX3nZzWolXlxIISmCvrmlXzQuYsfzVZ
Jwll8249V1PDKwzuR8/5s0k0rKWdDpycObtcOeIzjCjAe2tciseeSzDolnQIwBO4MxG55K/QApl9
Xe5JJtUoU1Xui347HaZyn1wnkCKtdZgun1eWeMzm1hiKYTwHpQ2jRVxE5Cgz9opSXbnDiZxjOzfS
gPVwmtTna+XBZ3BT+rXSg7/IaRZY/BFUIIA5wQ7v63FHUpUsKrtWSwVty1668UNMduba5QqWwVwA
8t9iYuJHgq7eEvqCQKxJGz5DWeePKuzxYFMxgpAWlZOrUeB4ou8LC5Xen9v52AXQf996cX6vaVnI
lbm4S6Uo3g8PXNxcoGYhl89ulob/pBPmMsbcZZBmkDi6HfCdJmFgduHoULC2dSfopTrCk3QPjx5o
l2atpbsicMQXcZUMJBr+veozY01aJTy6lEw4t0FGxKXpkDo2GG7qNuUsdyLmSRVQ57x01A/2ijfe
b+iLKPgGIIpsMmV8vTDXw2gZGRvNBMogITug96rieGRz9wiEorQaDOdIRLXVoGKPdbKOdu73V6Bn
8HLNJRL52vt7tXkdyxDpuCMkTyQvvxLiV7+BBA2/L8kYet1ypemtQ4YkthNrAf17sRB1TqKGyv7K
hwuxawD88D8VANmRr9dAGOHN3eyeZ/cmwsKmjmVOQLtpqJwxF1BWYsmR8jnp20CkEOHmHbUsWfL/
ZVzbP+V2FUaWScF01veL67k9vqgtgb24Y27CSdAFHBu2wBteeQBob9+JvoLUZa1L/4WkDnOTctfN
f43CYUGBOuqGDKskULgBJScF7eoQ/vC0SIb5IsnfzA/9LJbXv2InwlkRrfi66TL1Mh4GICnQuJbc
5cp/xH7EuvpW+seDt1klMEDX9BkZBqllSsDc2P0kLE1OqPtsPoJeDvHLDnKrVlAUXWi0MDCJ8khJ
qGMlMMmyzShx4zLEoXN1BEn3poMazfi1UwOyJNxuJETiIGi1v0dhLOktj5KrfswbHOAnczQWXHiJ
6IY5kw4EpvfnQ/+HlIs1KMW5AQoK9JKkvHHaKOmZ9HN15O5cIB1knMEMNaBAPh3qVH9Asv2IQgQj
Ynv34+cxjoC7fpyxES5Ax7JyAEWUG/J2XyQmSJ9YtXpMivFFAmxwG9NBoYr0B7ve/f4QEWNs5DZ+
6voh+vk560uql+cLZ+EQSAW31usquSB80ci+z1YmCIp3Xejt/xWXVKab0+NL8JHruYjAgwsT6Kyw
0Okg4pEuuS4uVi7jqpvyIuLlImAakOARrqpiAbjXiOkZ+UkzR3hw4U2pzXuum2PpkReNWzeAzXte
W87YNq2yz1wzT1HKeKRIaK5RO9zdn8zuPV/KT0ltifdhEblrdy0OzOLyfxBEJRuk8BQNv9P9eatK
lT7TOSovQZkHMndUneS1GX7c/sEUA7vGHq23t/7GJIqgIA84ILVcfxEUXMYfpWS8hN00I3yVnZEj
Xr39V4VEsOGSInZ87LfOhnTz8JDsTPx8eXT1V4yruWmpHYCutF1WDd0YHvp/n2iGPu6GDTzc95jM
ETvXrqR/lSnVk0CjTt/vQ+H2cCdjFtxZdQJWvrY/aB6aqd2rGNZyVLZmb2/Hv9TfSqn6rSg1T/EP
MFcJAV8snFR04c24mOVzG/TebKjBVzmBwLK2eaehuk67OIKB2l+CnKMqIL6FscJjg5VUDmVGvEgk
waz39F7stjgs0biPY3SIfVPlxtGFOvtOZZAr1kmjHyv4I7pbF5ZC5JQtCl4RBZaNrwUcXzfcBDQ0
cB2iypCv+HS8jvb0CQoAba5kM1ZXKtQsA+Fpp2yIVmHulx7UDDwNmqd/XeMaG/QCgfjb62Fx+wsl
wZHgEMdUVft7ykx5RZp18sItapyCjpygYQCTeXP78y4BMC3isQPK2Y+bcj9kKyE6PvfNInVJuwx3
mpjbleyH4eGGE76JlbaHbFKkO262T5T/6LuO87N31gNbX2HC9wqES9FWVkvAMgXFVPYZN6bCSKMo
LueHDqRm2q0MGmZQEeI6+K0XCxUy5wcV83foB3Su1ELh17kmD/V8JibaqClv0ENcE9QqY3iKv0ob
GDFjdaTpackqtVuYNsgjjZdxKd7jT1V3KFWS8kCEa5q//yX/WctazDfSWRzi3GTSrguSVwcXKRw8
MdpZCh1aeLQEI8lE8LKmMUwyxyypKDyIQOlz2W1e387w10PlFYynUC1u9TZXBHBZGJYe4nEZCxo0
uF2c7y/f2+9wNS/GCAizabDuTzb5TR6XnL72EAPvzz1KyRWrwnBkvVFkz4NDYsmi571+cWZ3no8m
3uoOWByOVWUYVYXmSXeW2Dq0p5irzJME6j6BVk/HrKPgWS/oIaEZHJh8QlYsmNyEjnmw3Fvgce/a
rnBoqt9QxQqgQ1vV7u7rEBLSxn9hUHnpaI7ZDMRk6AY4dAToSACrwQfzLAd6opnvqJYkKNPlClFi
rsADTjBs/FQiTW9Mjbfdd81w+lCR+a7H4L/eoSnal3a55vX5zHO0L2Ifzb4G51XSFfE6jynYzjlj
ocH3UXJ/PGKAgSIN85196FAsZM9kAktwm9qJ3NVr3d5SGtfq0FRO/hO/LXuxQUajXl8Ww6sH7uPf
UY8qshfcDxuaJti4HtRjs65+elfP2mZRQe5lvFKk07yX/QkWdMTLcvMn1bc/mVM6nSDv530GTIBI
NNor0v1NBOJKLztyESGmZEAC8sMxhGfY19GA+DGgoXdhWF2Ts2klcC3D+bCtu11G5/XDcU0RX1t6
lMepM2b14+q2SUpm5O60yFH4LYd8Ch9El0qCfLIoAykleBa6en4OtVuDqnRAPdgxWK/YC15KlKAU
3zxi0xvIwrSL7YUY1bURSwV08yaMA+9jSTUIMFjbLK90AoJm7J6UqJj+YGf5vLnl+bPqnyrk9dhJ
DCbf97jMYgEcpnl6E5sTmcRTGv5kEgP/xvpGNDePq4TxVZaxBbv036lh6uRaSNvzlaUXH9yHx28L
/ddKYSVVOd8Iw6WshGz6AHmHMcJtjN/hZ+EYlpP20oWCN0KBOGPjLiasAQzuPWrxX+UWx+9skiBN
KAjMZR8hJy2W90Ny32ZBUj340fzQnuI3Zj1o1WBKlBmycWKfb7lCqAWmbcSVoaBSpzK+8wvQWLHO
fcUiuzbsPLW+L9AYh02TSyT8w/jyB61580rxov6X7/yrThlgbh258fwInb6DXeBeejp3TM3abx6o
ndH3mIInrDBZ/Tl6BECld2H3maoScum7sGpuzHxgj9dyC3H+bLHCy+xU+F+d9GoeZTxNplIKVYLu
j7FCfK9PSuTFYdyh4T5X2SuqhYlSBxsubzJgcDrDW7kXBVYwe8knaTEnfPLZXGCC9DtuRGVH16DQ
8WJfg6lAGC+sZCIMfHf6xsjKIxlwo1VGrcrtS6vtDRaiTLIpLrjFMMp2G8lXeNXwxRlKJNOkf1pY
bKkzlSANF8zFh34uN4mq2gQ5XW44Pc9Rg98m1DU+wP+xM7Jc0EeS0S2p+8s27qKut/AcjTgVpYOZ
RUb9YTjfCG1rZviJgT3d12Dw4I08tJqBP9fzxgTZJbtArELQcBMZL/Fxk+/rooxFJUaGb0yp+Jv+
SvAF2YhSMVA6r+JprP9y1iy58u558PVd9EbrAbKe7XxQNTdpf+UPzRYWjDmoQwUcozwajXCugXtg
ERDFvl9Y02vH6RguvXnWcvMyVSQ7c6QjdymTt77mNZLT8VUPNqCcLdP8ykmySG3iyd7LAa5ObzeE
MFpqq4/aul9ES808K+uyiqFuLfdU+XYxWtpy68296oJcaDaTcWZfXtn0zAB2/9XCi0yRQyznTzZu
XLyjqXXVZE5v60KNDAj/MyeFy2VBxNE8OA+bjHSfMB03jHM50oYuZ0sTxoVSJR8a2tW4WQwMSi68
hB4oWD17+tCtQPTTXJvuQjQkY6nlfrXVVkt61BEZ0Ntds1s6rykmQBir0KM1Uq78D0gQcdeKHVWc
1CkYOFDXwJ0G3sfajn1hyhz+09+RV1xfwvgppMAc1f8R0CeKf8YWRGJJ4/s2PqkSoV6P9wvyVjS2
Wj+dE1cOPSI/V1UWkdWMRka09XnfZf8gb5Im1ltCMMkno3lo2X78yi4LNgqzFRpxqJ5dyX8Pz0BZ
xuaVW8Y8dRipj8ukgp5dkRydhDEYjFo3pGnz2eM+kJGTMWK1brO3weTiZOTtOMEpz/nvOEx8A1ML
aEJx9rTj1Rs7O6dxoHFp9Uucs5Rg2kd3f1cejiZWUpHstcFeuHt6ZblVH8JVvmQN4gpYPkn7G6I1
QTxCEdpcx+uQvn9jpJmu+MjlmKAJp0fn8/eJEraMZ3fzQis+Wg8+tSpRwJh24rpsT5oXgFOjvA/S
d/91fBWuf2fab3c/oKF6ls6r8EvAYV2tQnL1rJh8bf/A1SqI5QJf1m9+qnO5jBbCUdTw7KRNl9YU
Dc/P/d0w7v/8Sw/ilX7BEGEWZ44/2r9KViraaPTJRDy8yvADU/C/wgfk0sPpplcaokN1eK1l+/Ek
E5mZDJb12bfprIYlCqm+O06gIiJ2uirF20CxLo2xwPF3CKAWUS0LA4G/V5atRrX9Y07g+ZX9rlkJ
NiLrULWslxWQdr91xGFQZJ05bVtZSGaBLIJDdqnrTJ/71mJ+4yt4P/Gmz5cSgoEX/yxY3oc8ZyVZ
iiJpKqojtrMVIVFGX1XXg0qunNB9voQrZvgOhv9ZkLtuhkm/LZma7cGpaRHfYECcBpwa1TvpGDsf
OQt5/3ArMoaFmkItg3e+rwdoZu4YxL1ughEvEwNB4W65EQf7wuqD0YQuCK1gOLs0+9o5BR+SrhkB
Hw148TVNIlU38owujLBh9N/Nz7BmgPZxZjdnhaXC0cOHBTLOPNNUdXm8vbamerK7q0ULPcDJKN3h
iSEjpEUviKB5I3xSPFGgbMapAT7CYgE0THqZULu6m5WESqtOhZTb+a8GDSJO8dmihJA6I2KYIap/
hXLfRlbyAb8C5mEas8/0AF25A6iNZpCPJat4xRJ+a/gowbWGPo//7slBe8xAby3O0a8l8FOCYc6w
BsBnWZQoP+k+cu7wqyd0mF8PdEUYwmebfPHZoX6FqeM75G6yrvF4+LpWxI1b7+KnmQJuhl3x/vY+
2cQ04tXqhRZ6hjjctn57XiezHu1iOTuHh2g5ohkGanyEYSNC4Z63h8I0fz1RGK16JAlbqjcdyxAR
G57DOL+3KWXZPQ/pFDzaDR6ep8BaadOu7HNHO3gHIPoXrm7dJEKkMLM7N6YFVQBvdDbzOGM6Z4L+
4TyCPhqFvTF7ne+wDInTSvCrZNuItH5NqApzUZ6g75acsl2u12ewvGhE8DW5mTBFDe4KYXtdW2cK
reyprO20pKV8V4flT56J3TjvWmadfjPCfpY/EVS1tzf7fHiGBTUkD5kCPFGj6Qqp8LFnnTRugUSg
g/TdJMzsadds2ZBOFnyCb/umBEMf3KQ2tN/uZzPvXYtxYCgvniag/PsMMVYBwPvi069CXSoECBaK
9xBqBU0zcMlWxj96fZzOMnDb3nW+P3LBq9MJDgc4uiCLcvw39KfoSiKdMAgdBcyyZteBGl/Ik6lu
CQfrsM734ele2wYnScnKB8DDZa+xc3L0RaKeKM7WxikkgmLVSpB9cJVas4cKeRReqoOdlQK1SGqQ
8w3FadGHxZ4ow+kOPnZlEImuvcyCvBeZ0Vj0szKSoNUuBiH6HnENi0OiWtdFS/BmXF4Hb0rLRFbe
Lm2fjTUhWXOHUHB0Z0eH9bZ2EMDehKT3aEaoka/nZMTDSKF64uOj5oUgD+hxViaq4a5amJF8wLTo
VJ1evYLGznqzup/r28OT99HrMcDfgDV2DnQZ4Vio62FKnEXmhIILWIS0Y2GLyMfDqo7YKj56ZHwm
3SLt8sQz4dNLHLSwKOV3tbE6NwZxLv7cRm3pQsGhufLoOAsDv0ZWr3bvfSsgHN38tM9CITnIZWG2
/U0RrOKE0ecTCc7L54wr3FXr+LHVFrp3F5t0GqJAAjJ/IwSKiGNUPySOl1fUtdYDoRJWqwZpDDnN
FnDsRVKk0/M4gVAZDxnhOBcOerTC21ephn0e2TVTtVIIhfiKoWvCuFcppwti8ATq8xHCFoO57PuD
m/Sye4SaPzi0oPqJXgrHyaKDnssQkWfsilmtEW36lghPwVhTXJzsMMzpk+CB2hiS+QZEa6OWTYx0
IfSZZ/Kg2z2WkMp6QKYCVB+SpFJZz5iHE8RrNnc+b6WAJVi+HR+GuFFQYZRt8kWEWXeLkFQijsMf
RZGZufuqPNDf7Dnn1EM6Oa02MYr2cyezTs5sdtHkAjlw5DPijdMLTmuFNUrhyObgmHVd/QHW06KD
0qcwigF9vollV8okx4q6b5OWNgaJb+PM1Tm/UdoAOs1PsOFLLr1x/OfGRUIdy5eeLLC+DeTS2z2k
x97PySQZFRX79Sn8ssHCJlaAAyHULACWYw+E8x3wWK59UhELM6d0JzAkx2/JIo6iuxgvXTVn/0wy
ob+jkdU/NTUzBbqicyF8rT1losNOS9g+VnOyMAUqGZyFZzxI+mpCFXqe+WkdCf96smVgtsT+9LGk
JuVVXO9mKRVyuqzTLcEapsBgKntD5ugEk3g+CAotP27/2ay0DEuXF9zPRH/cABOxP/rO/3+FO/Mu
9b47tMkDC/0URqkPSWEqaqO+0KbBnvXgxjJDf20NFLUVSJCSBTWRayym+NU4qkHyKK0Vywphzm5M
wpzQPvVJz3S1VBe7Zumdfy4iNql59dkFj/aLxtrPudDQ7Fc4uWK12+EOmoXxzEK177tbmZCASatg
WM02zg8Nhfa/BNcihtvAFdu6IO191Trzmf7x3Lij83eZw2WQmJMkrL/RczI3hd6dO2SbLI5JnrdV
MICuysEUTop+lrgbrGQWBg34byazgj4+aQBuOMWJH60XAwfFM+IRQwp28YwmrlKc5bj/QZCvDNKt
QrnD4mNymMYjmHneCKdFwcCihavqurEk11weu9Fv0iVkndqXzSZkxbjTQRW3iu2ooQYMUuDexXRf
P1Ws0nHaqWcU3Ub2e8RaHThBZg2hgOt2XBkS7JAkKVp46TpvyY0IWlW/l+as5fOf32SGvgdNLd24
8VZqkOztfQBpSJfbzNnkUSBMHGMqHJQIWZJjde/0XNR9OztU9VsAJUUg2/9NbuRGLtKl4jgmh2dH
NwX5UyzUamtIYPtu/PrH3/2DQM2tY4V4jIX3Ux6Ctq4apxt617vGeE2yG1ZAsAf+thHX6UfC6RfI
nsHTQtF29lrQGEAxZr7CA9KaFzuKCvJ1hNIKxh3QfFGV3LxpCb8kKj9kZ30W3zY51acaj5lpV6Nm
6IrzWMjwTK4FI6d8Wu20wZsXllFzUDa1NfiXlrumdcsVjVl1R2UFby14gJCdC4iYbQdQN43F7eo5
q1sQYhTknWxHi5bytixiRNyEv03OuJGNGXP47dPDUrs+xmJ85+hDjYcCbKmnEjnDyHdE7tP/JTLL
kM1Gla0POVtKP6UNbTVKRrn5IWYVR5csO1jkHGr50Av2/IVVIQ0k/UDu6f+1cUgVmxtO/pjR3lzw
afdER0BR8HnOUwzKF59v1WeLPMR7nJo5HxEVaeprOOzd7VhVWeHROlOZXNP1YR3pq/ZqlKwUgqTi
RCfEbxw34HhD6Av8hbaFYPABV04tD7dVyCdSOnI+AE2azmCHHH6tn0KBG9PTNKx4EQ1mZe2n6w34
00qU40zxYiwEsMmSsfdp+RwCqL3dyW51Jdcpf3pVswnoiNRsSB1QtVclCcXDzNSP7MhvTLg+SW7s
VgwuwkGBhKI8OEL/4F2S7cT5Gs8AN33izMsNm7bezdDDrqWCi6cXEsqFJXa3OhdgKqCzkS3lmdiE
xLnW1yoMfBb+KOEsfEzXZZoHOV+KkQuWm7jEtIPHeBYMYMh+OJhOrElSpUTzBgkhdR+AupGLaNkj
Yvf1ww8JrKOXhjedOePEbnRQ5ISkNzBzZTdXHSIAUJ2cxsxVSGZxagurwCM+v1AZoqV0mruVbkzQ
gMQod52QEHOflvwzmCjTvQydwrWaEHd5ehaekOXEV/wkeA80BTqzoeH74Q7VvNLi+OZ6Udoog9gj
h/ZyrcGEhVRFIKvjBnbCUSNwgb8TqwhUq2tA/2214zfocobaieldIPX2dPzEYGxjy9edYzgu3iA3
iuhFqSuyLtmmno2QJzXXliEWZKSzyGvaAzomlPi1HzZfxlPZruNiL+ksUmm9ncUszTMFlNybi6D4
D1iiNL+JUfQlpxRQvgQACYMClr8ae+kcq7kB5vMcIF9ORionkuoQVTOwgc+xhbmCOOMcuOowBybZ
TRqKL9LtlUP6iL3NA+fZ2vvig/+GLdZ5NWgcV3MsYgUokp0OCXXWY7EPLqagoPVVvZjjq5U22gz1
UKTiBI+iL+V8hr85hI3BdByMBOp8LvaqtRxgJN038fs/WPhZgMd7/6v22SE1JoxKYD42MGVWFMic
haHKDDXd2zOYs+gsmKqDqfmRD2tA0Ps2RwnD/7wYHKCbmLk2ejOQNw4cONJsbI8b026iQil8DPmu
sxFF9XUhCSODQ6dgGC6lZApyyd5Fm9KgJngxHw5jz7FFwgno3XFKT2pCryA7TYqY2FNbv2/GgSUK
jO1caV+RWn/7hSFrriWPqGyitRH9hwlMu06UHebGeiDy/7b7LkhieFtmM5WeMq/g8sOChnphe2NZ
Dwh9+klpqBfF4BkuYmmhU2swOQOWqruS0LyZGdIOu/o+Jam/L4HQuR1wZl3XjOYY/orrrGvsuWzu
Z9FSZjIFwXr9tX9e6SyEMYTDx1IYzq9dcayQJvg3uPEsy5lotq35a4JVU5sGnaG3WzNhWVzo1yg7
x7ltXASHFNPFM1Cge+l90LPjHGBehnmup864KK222VLhdxKneQk2cNDqrYHKpPtDXOg9lVedd8ov
mj3kk+pSIttKetLY8iMtjjeBj/jfl1JNY1zOQ3axregn8yj2c9PDUIuMjO0GegKwUzNUo07tJW29
D+yjUQ08SnuZJcrZlf6g+xb+w4VffHWhcP2x63AqqU8hed2HenAd5ctw2Jdd5UM2KsLBiPfOzbYG
BRJ5C8ZU441OueC3f00m9ComIKbvdxYqp7wQWk7VaMN7KppPbNEeyA0L75PVPKW1MTzow0O96VCp
0yDm4lye1zR1GzW6w+LwkkZubNVTNjp1fSurLQ8isoiqyXU0MH8YpMgr7Pw2oe/yxDqG7JFr+B8F
9DfjfVIKMxtXsFSvZtD0epLRdtBFfVjTZFZtaxN2WMDVHWFXxMJy6kdAbv+yXNpakRbPFGaj2QRa
/3Wc7J2EkLUn1LxrB89zyYngg2KpRp8n7cgGySvmxLKMAHfPmMGE7eym+eZuYyqG3sk+jOee7gCq
ZDtu5tIFLC5W55neOZz6pkE1VzI9ltSon5qwT/PkyVQno0Uh/mcaPqRvDjtCZ2O25dc1U+LzB66z
VDa+CTBDT85Zb82fa+pawvFlye6GVpf1VYHPPI/AX5BsgWkhVsuDYBoUqcY/ZgaYArIiJL3OtnE0
E0I6nn/ALV0+SWKqcAuOWEvEiEU8IEA5v6oYUYwdcA7CrnNBu1IUBhOKZhFFTHi2lG1OJz3bqGJj
TQH6hM6X83S4TgTs/ziFnCpp3t6De5oFTy9b6nDFaToLivZS7RLOw84U9vSeyjH/utsoNPUpQ8+I
Jl/azETGXeNYzS+EUU1kydtqA27t567O7C7cU8zxJGd9XVc5lXqushkzALgQyorGHtIzmujf4D2s
ezqY7kQii1VpJdpDIea9TKFZ1bCkFJFvdkhB60RPOi6kpjSq0XItjSU5Vshl9IedVVEododWIKK0
xyL9Y05YThf1ZGVsHeJkRKg00Kbu1OyxRMQPboP7s3x6VbcVE9FuoqxmvnlEMxvKpYn2LYWJT6AO
fW1TfyUL6x93cXslzQWe9AW6TZm0yyGHCsp6hWDABJXtdMUwGfx723p38jpJnNN4+n0OPy5ER1H7
RKQBMmNCCUW/QQ7JIzlUFe56OEbmgA5UXEYNlMd/N3nFcVRgizOb04xo8Wb/UmDgmZtxPjlaM4ni
yuVJGfS5QTUdZgmgU687bMzKUp1wQgWg8hOc+PN6dIj1TMbdS+mf84W+b8ZxWUGlA2bsi9aDOH3s
aby7WBgFeTl/DELn+vj+RUt4AjPfn+hROjJejPs7oyo5ABa3oZcCufajFnpgCd7pCnK/0mbZ+i+1
LKIiTPOGHuSE/oRdSHNhbJXAOpmjL10/VJ9mozKMH6sx+akHB9kvj7oa5WJ4vJR9lUGifNaArenh
4R6U9PErT0KeCfL+DLgrnv4+Q1rdpCLz0h11LLH4tLFJ6uM3UMF93QutVRTQriuEzS4zI4YGtBKg
4Di0rQfSmj0+FXngWI6sGFQPZePt9i4pLQHrDJz3j+tLxPd9rPVB4GiGvGV4FB2NTr3XfmRJsr0A
4jLnbsFU2CRJUgHDFSFsa1LDbYEpCtxJqSN5bTiJTX/n7rRg8il5LL7YUlOh37GEpSK4w8z44bTB
2GnwaajiXSyB/1TM6aRdy0q1UQeVkEShc4nIwEuwQJa0OyJDZ7ZM4Z6ApzpSB/HFwamlslIXS0d6
cc01dLyWma9l0sS/xZKfoP8j+zW/p5XgUC3JYNkAzS75hchGL4bPDCgbngfpQrGRozZZX3vPeQaN
IgFLWKpkUCuvYPsQYcuESgbQ7mLmU9j34Vt36S34fKEe2BkEKl2uusvW/fpti+ogEezUoOmAdr1N
M5YeqFN+Z9FjNZ9GxfYBzW8+l++xIA5VUixKsHmd1kA2dexMdaDVvtA6WajB5seONQbYmGIODkMO
ltCFAH9JcVkb5UlxxRTz/5nzWYHKtIbpXFRnhHzud9MDHXe1wS4KHC2KgO8eLDZJwSeBXWAGPWck
PhV9YIyTNOzXfw5cS1yTiRG6uOlNdZDWDkqlus4VWqcLv/GCdEkchflx7/x2pBYYXgAAG03WUCOu
xCetiy0QQFpzX92PFRWkk4ywXWbYvoqDkR5cfKwy2Y05SJtbRqNowVnpWC0kAnJg/2ImSwrCsrU0
pWoDXen55Wj3I3a1PFuRlW4/lSugtAwjFBUD26eEbKmbzAKsD+0z5ETjuuMYaQpdiSVOMijmTLsC
6Pxf58FN2+iZ3Lsa6s242fPaIjnDs1KNU+yxejFRufiQmus2OLieN2BptOfxedBnUeUmRk8sT7op
PEGwpTfnv2EKV5xdwVc06hUNJ7WykYDmiW9vpCoM/47OJ53wE288tITLLtMsm3JimYctZVhQn6G7
+8YBcNo/oHb47d78Vw5Rtxhp+9nREDu4gOhvwpVGDY5AF1XqtsVdlH5q6kdmrvXUqyXI2fJ3QvnY
XCInujS83mTzvBDxb1Az5aPlfK8TAftlbwvnsY81g6gf5yxmt5R1Kpv02/eDENYClSlNiIpPoEMy
c5vdP+tgN8UUdzqcuFvhiwhl2MDyPdeAeJXZDAACyzT9hkH8wHq2ElpA+OWBOS+boGx4ZKI0UX6s
gL3S3zhAV+J9nFpvUMrUyEY9FlzQxCofCAjdsGXrlzXaWFyz6Jz4gRsm1t8RQUxOYMZaBJAjoL9A
aKD6ZBH73G/D2lgP2QeIkA3M7DXQXZYT/uqNTJR8XyOrcau8uhac1LX/eNgBnPIiOiZEsHzkC+7F
KDdWU9zZQX5tkm05R9Nn/c1NGwTDKSwDfn/M9p5awwSJw4HzQz6kwPwNxEwzMuCx5pXtMV3CfyHm
o9gKaweBSRRUGfQQ+Zl8QvQDEDSrLbIp4dw5zSEwOcf8IrVM1dPuSgD1i3rzS14p1mA5hW2g+74W
LO6nsUsU/LisY4ZJFgU7EeaAseAzIf55aQe6Yo1ar/YbmY4o2rpohd933ly6/pVIC09EiB7aGt6R
/aBaMduFJPxCwDw/4PoZdubwgsfNBBMFVS034lTKlhjLVbIEIqk57C3eOMpfdsO5AiivfdBGdQLL
6ZfQHIvZcvGTDR+0cbXt1Igd08HvTh9nYDRNROZyBOSOoWZzPVLExMfApjQCrvOXn73YodKHPQjj
TotR037Z3OupVnv6xs/q0NTMXkfR6YP7aK8g+Y+v3WYgIs9BZZkEBVSigxni+TR1esFPuUpW090k
tCDs4xrlhb31iksgmAj6BfzGZbcH8iLSzTgckrJ6NuySyHqpbQmsQ9SDLD61lKAY+hiVFSH+zjPp
WGoV9hMS6x4SQSkhJ21t0M0sMaBLhv+9potS3X2GzP7Y+nKmjPbnytYdC+25ZayGpT0TFsXvOINl
5ZDrsglKb1FUX+4OifieWgTSSb7PZFin3j31Sh5N3YlWuu+fQd4vjDMyj5z8TWmDiLcpgpLImwOK
YDbeKTmIlhNWoGJFENGaT6jPE1H7hjsMWY8YyC4gRh0ytGmxlLKGE0WM9kZhka5kDBJTVjWaN+9D
gJN2gXh0qDwVHzk8nXmes9H5oJdR71Gou5yNQCncAh8/vgAyZCWYzWpBRC+JkTLFD96e5yt19Zkf
EwMyShbcb9Qk85zMcTrFbzK4PFSOgccnGpoKyAEx5MJVbbUekE2erUsFjq+2Zj3BhfSb/v3Mf740
zOqS42hQGCbp6Kur8J6f/pisYAicTNjP50CCar+u1OqmQ8SPZSOLE9bgj/zRwovLsRx+a52HOj9r
38thwwT+wOWsF3M1Ab7tfckx5CQR2pkLU7VTmsto/J3qiQ/cfsrKV9rjZ2P2CfeD7rM6CDTAmKqr
VBkFGsri9qjIpQ6Dj+hB//78UJnhe6WcSCO+bnKy7h8lOZuFHHqPRDhF/tECilaf83zT6+ky23C6
qCVFIWdq+7cpe8IJBq5Npn/0nmp7xwBCX1spIfs5xWz0vUHAcyxBrxkl1RSGjtNWWGDzyd/dKCxj
IFgfftHYAFochqEGbOveFnpe8UgeLl7fmFuoyE/y3U7PDq2NwNVQlpAVbyoIRLMMXD1DAAEkBo/3
Yzt0lQk4o8q1QsWlttQPSy1mrrZ9ecg5lA6A8xvlveqkDJIOgkKIWL24QTGQCnRKGURnKZwSMwSf
Xuw/cbN7eMrorU6bOv5TTGWQjAbzalnC1wXXOVlFuYvdgYPPXXM1tPaHLMwAHqnZwPyJ8SD5mj2Z
am5PDHcrDwMnpNkPUx7+FZEouoCAtJOsuJwSZuNJ3p1NrCvwRQ4UN3xOcyCzwcE9g9xx5HmKAKYQ
0bJEUrmqnZxQQj5OW9Yymp2sAgNl9b517CotUoYe7ljj1FhAjxLjSLKghyYx+0iWlBtLcT9kU3QQ
LeNf9ruweAZ9qJXw9gAEOXy0hR7BjedtJKNs//XQXs48I9LUb8S9RHqgtMQHfnJZGW8HF5PkLgQG
xldzVLYLB4/3wHdCbZ/KPX0vh8wsE68sb0N+qZDOSV4YiOTrXbJj8PhwsZt0JP7Wtw5kZF4QtbFf
iFU4ig23d0ruS/bwamMfpeNjsp/mQHZR1otGe7D6+igae/mQZEQESkFLfehqMA3MdO5NmIpDFdiJ
L2Rqwd8/Aj+NHA5i1Bn3ihJ7rfN6OjYL30xos5hWOHUbFRNkNGxZXL1+88o+08QOcWYSgfyUqQyF
2eZOugYDMB7xzaHbMy5jdlK0dP8EneRe6O9dk3x6Ch7wZzjYvLwKj6YLK8ubodjRCaAwfKB40HWo
7P7kl964knfU5sJGQmCPPusCbz4sx9IrlKaerH2pYUWmZrDtHNkAOxna4gRCCsQcpuwyqRYzpZlB
/G4spEXFWtTaj/BSz3ULEko5rwwi/NDafuOY6pA9CUAWPeRTjyj/I/bH3GNU0Hc0fG8m0mkhdZva
tsHbQjpZWUrcPvFlnW7Y91ZD8DWaawkSwMxcbbo5Lt9qdxIvfCWxWyi3P/EkW3zMdaqZ6caXJ2Jm
McuzUW41lE5Hm5g6i6bFSnx3bQ9aPVizBvCS4ju0RuJp38Z8VFwPcpiAUqq9aRD6F/GpZSfdpUDx
y2YyK7+8rNkUJF6Cl6yLMpMGDd6idw56A44OPwzbijQm/XyFOivvScfd9j4Il4UQ5mutynz0ye9l
jCXSyDWgFnH35I5dQtmK9/kw+zaQOV9Mr/oTwHl67+RjrsEH3E6aOsniH44TEPECehnLcot1OpbB
wiE+PZm5i5CgPSC6sQQFbrEqZ2AVcFveW7Doh+vz1E+4p+rjV0m+3nC2JQ7NpbT05ZqW+8dMZ0L8
DzHIYWjUyfGuoEGbmhotMigLrhusod7JVb6EQHZtyKaQi8hlKDozePqTz4WT0wk1iQrQgcJWH9Q6
+DkIXnyKzdaxkfV5ywnShs/yIWbTwpytWlVVNJa2XhUV7DWtTEOcIn/70YRoXvHbMT+2x7fWMxDJ
EJ1YLUQPqwa0Xx90cINDoTw1bSCxOnR+/FkngIBrNlSfZqNRVSb2kTKSWwyzlGiTFAWGKpfUw2Yu
ID0UzZyoQuctiRe59yWZg0raej8rTUEY9Atc+YNdMYPTRqWrS9xubBsLrdgviOtv0IEKVrTe2HM4
wipastzGC+xsoFLzoJpM3baYSfsaX8QJXdwu21IqRAOp4y2bFv9af1doU0MEiUoyWaI9/CRMk7py
r8M3yQYr1L2nFZ7zLZGuahCwAXeJWlA+WCz7S3qemXvUDSQ8/M6dRFqVVwxLbqfPS86rVzIKsRQT
tlNDkeeEIIU67bIQSwryVSkOC72EZTxHG+3vpZP54XjWXMDIK8wpxIGnR2d3AOL7wvrSvR8RFfFw
p4nhmpWeSJhCCymy9DSk8yJBL5+zQVeI6FoWtFM2xWc40bc50fsGi1opViIhBJrx2FMLPOkd5g2g
cJyNcYugNW9zBpLvW76AbUNAV8I6IVV9WZIDESBfuCP7hZYZO8TdCQyUnwf4DQ2btqOimrc1udDu
EWI7QrimNqPoA0T3B02S0kV6vzOZju/7cBY6BOOrcBB0LG4o5Z0CLrrDBD6W+HIkOJ+8KrHRZQc/
Gdhk4Cp5m7UoXJTZ0Q/0B6lTXbbJAm5sFAD1k4LY0YcB/VSOBWyJg3JppnL2kBZg1SZT8WnTQq9J
T2nK5J2wn/ZbUzTwy49axKnFVpd5qNR8ilpCOzp2rgiw+On9PSDGPI1sCY7XC6qek6SNicRFobuW
211v9b6y8beGDQ3LRKgXnBExC3pNRZyZh1VOeyt7bww7qDyNQgzLlf01WdqJwNHxJPbOn3rGVLHF
8QSszvSH/CMjmI3mIb+lG5PTnMK/otxaMtzgTMJeW/YHv9tWh9NUREEwpt6PKi3WW0Y+ne4JbKH/
2Tsb8Mqnugi5QXiJmFXYYq4yNw7jSAqSRboMermvTqtPILICslwo8GXc5rm3DfJDoSUEsALEIOEP
yZQK3yKdhw5Pg8x3pAShmj/avsIopEnzRlidvc83BsZoYBlv8hPhDKFHpvqmVrsTfbpcU2DgneRU
KP6TJVkZG5GatzCI8IF1JCkmoIB+uitdwM4jhpY6h6ktjB5dQy4jH68FVlCQ584vCj+jXj6HVk0W
GsK+diy8Lkv54xYf3HNxuHv/EFziWhlkdyQEVbfHT4DgpIqR9zxugzszQCs/8Clm5KzSP5SiHWUJ
tCwoNyy37uuOyXGfcIJTY6/ehEPv+FTMC6ZR7A3a2WQ7lS/FTaELNvDFFMuwmP1lwqo9Tvsxekrj
72tdG1SUS1SCwGdvL2kmchzhexotqTEh4a7WOcE3n42dYh8txN3HDL8qknp7g/3E/nxMItV2Q19O
cRC2dcNaCVzh2euhtuvr42AneFgSNS8xMXC3StwS7J6E0HVlY4SPtDI9l2mBK/2n4o4HchZf4ev9
mC80hSSDvwFaBfYFDGVI+TogTlx1aMpOsiAUTgFmmIhf1aCNJfwUDpKDDlm0dfiijvi8TlImT+sO
xRKGLA9EjlW3HXGVZJ1b+dyLq++mHPdUIjyYvquaKHNRplGrI1h6Zz3VTUiQXVMAHbPzBP757Apw
uWZnWAyJryYfwJ+KvEf+N6B2IlH38pX0KIYtWt2xAgLoE2KVF3e8alz/S/JElMHrpVMhBIBHpWjC
HCmmI1b1QSD2V3FqxDE8k/yHKWmze0lQ43YSQOj3lpXxhqVSkftIIZpOyoYG8d+Y3oKNDJYxEfEk
rzS0TcYgnyZAzgB+L4BgGqcvhxvHLjUVsp1skDqQiv1cZ6AKJc2W1uQXZgIyGsmR3bQMhlOYM8OT
kdwDFA0qR8pX8VDXP4wbBwI68DRRDBCiWCMU8TBWV42vg+E50FoFOAoOX+o/uEWY+Bno22QKAYg2
jcoAMH9tk7qNex0+XZzGFJxF0yzTLSK/dVcP04Za4cinq/oNA/uboGMrKA/kO53afI4kCCgoAw/V
SYyleBEBmMqmF69hizMun228rSh4JmQXEYNVHaeU4wMjRzaymqFpOwnVOTZHxWmkyIhcIL5qnI4H
iONGBOITiVwdxp1CU2x+Zv3oZVrRZmzM3s0LQnJZv6ScilcGY9XLQb7YUesh9oR1tMmMIsNCVDkQ
/doCTdWDbO3z7+VslRTG0U6wew0oRl1JW9ttF6iS/jWZkCSlMtZOeJTAePstRm/M+vvASjl8jaYE
Hvr5//Lh4u/bjKx84De7YtBaua3XFgUMLDPuDTYaSsRkltX0d4RB2sczLRjlDaJ93G0R00dkLb8+
Z8CEQw+a6Yj7xFEtF3/CRKN+z1ue3tuXhU3MfIikCUjqSi9tuBihjvbGIjLlvP6i2VRgFKm31qp3
klt8ikmg/DyMlSkbK+LKZXVLInskqvQouXIMKdkkt87aO7keQMP9gvN5Jrc9+IUq1YHkyp38PxVP
sU533BKZ700Ix1SK/DnK6oZkkgqJF5BhT9Q7qp4OzhWg95vSM5hD9x8UvvqV3sf3UzcyYl+pkUwp
1V4LVdKMKn9zicaCw3cc0bRRVnPPzf1+M7IztDe/YlCeEI3GUQ/RHgm9nUktbkEGVPabeXGqDrqN
g42fyQn+6klbDHbj0meuhBSuA+u8BWAOAYyQRj6cdGyMs5D86wYMcPhT+WIno/Cnc2zh7zG7ZgDg
pxNkP4UuXvhayWJsDV53Leunocrqwlg57opcfwzpSbj7p3cxDXV3JY9UPD/Gk5YPkqpoMrL/GdjF
q0aaQRlSrLcOzcj9Q6pkQQd1KRLDCRumsDzpb/3AW0nIlpME94zrnbwOAHxXT1krtqK3tfDgwU0X
Ua9k5LGhyB3YBoJ+1XmGvmi6pwDAKYNoiheGP6+iSefuPJq0xt2B6ZJ61v7Hp/NsSIdf3EOOZBOe
2hU+7LZy/ERgnSKbJaMDPqX63w5wiIqkXGFlIbrr+N7wYG2SSqPFPmGcMzpmMWgFNlAirA+gAh3g
58qaupUAYHrr9prrPAyP+Fb9V2+5EyXgYMqOjNxirnMcfLjje7O9chZVUF1TXDONpGwjZ7tW193D
n1Xgo39/iZDSxH96Ec6DO+cgyH64U+jU2yn3UDhNlbNRrCySIK1xrJrIw1PKmFDnoT/r5Cpjb8Pr
TfZDm9I0YZmu/FYpm2Q34Ruk/2qqYcBsAwvICZkqmV5zySQGq2QQjsO1tdI8w5FE1Ofg6w4OOUlC
8NKYbt05srOBnwADgNkQ4VUbWFxca2XfC5CHk9Wu/pty2wHQXOUliUpSnKavVH6oqOfFJ6H3Y649
fBsLAf8rqR/kkHEYV222Rg/4shdW7ZmWM+jwWEJnbNu5Wet9ZgzBG4G2QZzEettVwK8KPdwE5ytg
FqXcbZz5skGRaQlyhV23D9/umo/LOHgtzfdfyz3WwGo0XXuTGgYDPk1a9y6yk2g1ZlwajsoQO0l3
cc0S66/KHbVoaDVQ3G39zZptJEOSwk/mcdOj1zALhNxVpaY2uNNP7HtfG+Rn9QWimeeCpTE1UCuW
9jEPX6rYwEbWlN2AMP4e5cup37yViA6UWMh9efjs9rc26Nh0UXQSAM7P07W9xZliJUYswa1jNiXv
P5esEHFkIjC4ihWd5LMEh/WUIMYMCYiyg0gpw3tQzzXWMzmx27F3YMr4ezQ30BoTiHOS1u8/e2Yk
aAjPZyFxGL6Mk9dJSXPqkF3+W6joTZa3Z+lkZWqfo2pd9nj+eNb1xDG7DfXJakWjHcPl7ycJyJaG
qIEs+f+Pp0F4YmhjOEEndwB391ZwVqudbMeOiki/jUryGmsN5cBxUqhQCw45TyvE9w/o3Oy2Mkfl
B2ib+TEJEr6VlYqWjzG8pQ3dHxncHJw85mkioOH3JpafU+z7PzNcx7fZgodnaj6isBJ1TjU6aRlv
vQ6eZCywzh9I25PCW26es71Y/0h2S4nMBi/6B0uPy4pnJf8b+4q6FxSsA8iDtvEh2tcvoYBT6OE8
bfFtCuu3g9FLcxutXea0iCIaYUxNUoH2D5LgNjOYg48SwhUAnSm5UQE3OQ6M/rRs5ZLEqpbUiHK2
uz7qm/QCGPbZ7eYa5R6cdpd76mRaFRZ1/pC8N4MyXJe4rGb0TsI+kUkT9l9p097cymT2iFYvpzUt
3MmFtDksK7kuM3FHOx6LbHOrI3Y4aOX9RiQofoTxaIYzfC0NHYH2IVZKXYKVd+Q5zU0tC78167+F
x2QvzPNUMFJXqBgjCS5XRvE6RxS/kvbI5wILLk8tLVLAD2BwrTFKjHADFCoIZVWINYtTTY+Wj0M+
+CC4DUOMz37cOfleEDbi69vqGTAQgXw2ThPigl4NMiIjrg3iMwwLEdjTrFqVkXkEp5qHhCh++lT1
owpw4YKQ48pV1hz6LxwHPElpM7g/TpRhcpivnkPKuYDNNt3LSt5+SaNqAHkaDBNtjWNlO/Urxx92
+CpyXNihNlgI2Sd4I2ngJJzShhmtj3/ZibN9PPpjByjVHZWTtrWOXzX3aLVgUUR8gXYh0IV1heHo
3YEQAfLkMUltntQMLaSti5uoF6GHUxklIkfbOoX1tbMgMcU4JxqSA0emGS6Z+bVjn31vs38Sd7pL
avTfnSpd1qagiQnd6isbW44RLUmFeYdzFQfdSsXL6xqR+G66owZ2DD8dHCmyigKcHouLSe6N9jDw
9uXEsNOh9CLXSCVN9kHzvC+S0XzSjZS7SU9SBKH/Kqn05eOozcaDMbCyNLCea0IbWjdXWKhhiArk
7E8qMfDM9CauAiC1q+Sr/ftSnE83kxjY9sPgpj5KkcAMu+yLh1GMt9gxd2K1ztPzA2jKERGDsbUg
RONU5+fl00xkUYiMVG8g6jkxa4oktmjso676//I07xOZPC1fLr3RGfRchyse8zgksraBiryYMNWe
Rw8RmvrKIw0qhtPAKCSiwY+goyYQKHG2lkcbrq5elrCWDYTXx0o0iOv5Ao5aubap4Rjr9xRJiFe2
v62UiMXINk2h1VUjuG/ncGtYkEnFZ/Xnbbb83VX8TvAzQgK0utIeDbUme9gAlvAXmMwnSZv8uxeT
SX1yNpccRhB4gbu+1PJv/UcnEZRrdERJzvU4d/htmEq+/lF6f2ynm9RPr4VCMETlvzDf0Wuvvu1M
xPplo2WGFSgg6d+to5S+KmD/Dn8X5nO4IWCEDDfab8LCC1qEAr7ZyB13j1rl4FmbEjPVbbCl9ID0
FconM9olMY+iQcCVDIEP7LxCGOAiXmJaKk7x6kfkV0QBf16ncxg6vDOy/e24Gb272AJMrGpjdX1T
ULU6tyEp8Gi/Uu96szVMEh+g7Vf7ejGj7NbTyn3Ino931gOCOTCCDafGblqxMP0+cV3HXA0NkAZg
+Iw3s2lnl58Cb8vtWcVxjM1GkrQ2+6gyqNzUYbr7D1qeDMEGhbiAbH6ismGFOl7AJHgEv8EYW/4e
18O8ygLBkNVZdwoXP0TmG/+YvkoVtQ/s86a5/jxgHBqZToJqUC7L9bN5Nc3I00bHSuHCc0WH1NMd
oPXcaHzXSIJ3hGDio/o7DPUyCWkkGFTNwQO8zGApPpLgEOhEqDZYtnhrIgRJFdFW8AynEGr/bRXv
pspx3H29Dy1qWQILvmXO3J9AnoML64DVCjl750kNIgoILDdzDEUEFQQdG9DQduNOvL7I63t9RTvy
8p/v43RGz2m5pEdOOHco3FX0eTxkx28eifzUlvWLmyQm9LAc4JgoGGvfp8zNSEDN6BJk/JqIQpFK
/OGsWEy1xPknfRTizcEEeblVyQ4a2+Byd8zFed4gc/PMc7nViYD+WDGOJ8LAD6S2QuFbQERHMsTh
ETyrt5nkc63/Uhs9SLTLaAvhCUn+CQZn+Qf56m9tyC0cZRUMsDunUkV2UDRI8szga4sKu3/ubsMN
q3/HlUsIqKwRSANFO2UOfazv0amYfwRcNP/FWvkOxWPtc8b1HI+QUtUwDX1khB34/AzrSAIKU0yJ
HWMRQNHP8pfptcIFZNg2yaDPZdwhKOyaW+s0FivPaGtn0B4iONebA9oMPk9HpQQM2HmySERY6k98
NsEvyYuchzQvYDUHplgTg6tP5JpNpNXPCMAOvYqlLqXatonBfurXfJl+K7eo1hcOoFq9M1EtTO40
7jxzCBhJ0o6w58h+0d3ZamWKuDaU29Kopg/BqMjfVagFNCVicU5hb7YsU3EjIEx+te3K7Gi4O1PZ
MMyFHTqTnX86VfBtBO8eVJEfOuTZmS9vx1XJEe3dkzZQxAQgLUL0y571msflxWDSbmYLoezEoN1d
fl/vAfRlvAC35isG0oMPPYfGy999PTxvDEv6XYV82Czi/Dytz+2dQvLaAQSvCm7n/lFi9DXygOos
86qQOiJYr15Rdw/cxBmRyKd1PLun76EN+z5t7J55aYEsFrMfMX5OFI3rCGMK2JtZUhKyf4nQqHtB
wBfShSU8K4mbUIHwmTduTTNsETwgupL9BC+GZ+1gRtyvI/Idyv83iQrXNBpUIe6dlmgYPcJ+Zxvh
RCxDs9FSaw9VjXjqpaDbpzu7McFwPsI80p+u2886b2sdHawL6NX2/7s1xuGx1BGfkJIj5pHHPYrv
lusFb1C3RyUsOJu/tG8kq7gvYmCCjcWlJF52/giV19Z17+kERj4ct6vbtsA5emFlipewjdYqdLN/
YxxhMrlekBAMVBY1+6ZeVmA1BXQXoxmAoHOTAZpTqO/3Lr1OFV7ab1ciJLSfx0cRXi7oqGrnOqSa
VPAvcga5Cpn+Iyn1P1DUtEXyN2I4ICvLXPEQTtlVExUI74PakXNTN++AAwyhCCzqKgXd08MF0qWV
g24IZoWjdLvoorCJ7lYH8ZaHG8lORRrsjEg+c1ftEdsd7bYxTpGG2ooHR9UFNwXxfO9LT0iWUJ7T
TeBIGuiLM13HQFPCgXT8uFizooLAvFbPSJmENGo8z8Tes/67LcJLzM36GT8JVZ13ABohxN7F1pmL
vX9ir9fb5ygKlFZIrEZkTjjA2meje+2JXMRj1FxruF9w9IIH7HKSNEdCiCT86KSKsvhIVstbv9lV
45v8IkbqqodDbgfFH3rcHRtWoHRl49VA8Q7jV6ldq1TBUDLPienKlIN5+RQbVCBfiMqPe9OO1W4R
mcCTkQJ2t+0R2VN+qO5vkYelEpYLwkxo460+nrCflrZjpi4ydjTFhf+PnAQFtvFvr6i0tYxf1Ejv
YzVX+zGGTur41btd2PaG6PdP4Yo6mmxzEdJ+yzjk1doQQlcq3pEiRoAutnvGYHkIhOn/nk8Lgl9L
lf+scHxcbwK/rrrgpn0MQ+LrKDQ7omZRqE8l9NlsSP4POMTOVGSjSgKo9i9+z9JMlS7Z/NpmGlNP
xmN/ESe0wcnFPyjsBFwxA0AWc+8AU9a0mhZl5ZUKojcTRmfhZiznPrZwVKFUNuK1aiOAZtt83R8c
Rhk6otiuPRY+PLdeFwZRIt8nPmuv2PnsTTp2gOx/pJPNgy1Cp/++WCs3WItKqXIDcVy2Qk9T/T37
E7tK96HiL32e8r7Yhf6Kkvkq4oAedNWtnhqM9lDY6Eono/qVq+ky4usSTWS376tbW+0N6j6cGXYu
o4g3dvO3gR1MDNpmyd6S/hOOYG78crRfkk0zQtoWkVYbLfPchoT9BvKYxB5fFK4T9U22c+JK6IJA
bZTUq34F4BM9FK6sMIz3zjJFZmD1/aH2syfkbCjSvpDVWsKKAh9/pou85HftkavJlA6fqeE5Hbha
nit2z5U1AOjCNJCWwrsf/5UyqGl2IcyP9JUEQaZIAzELaxw6qBwhrx/wwFEUhN6ql+kFNUoJT7XL
JXwvZTs0oAB1a4EbQ0WrCXfRKyQn4nlIyxnypmtXoEDHZhcovLU7mklHZIALgX4G5qnnYCEpv2uP
E/5pm0vCRw6ms6ZM9aQqBj9J0XMVq7OrBb2RtY0LxHKWjRt/zRPfDhWyoaTOY/s8NrNJdGxxeJB8
3IrHFi9WQrNqb08Bdx32I0ZhL3gCAJq123eukpxfijgZdxNQgwpNoWqPDL82pDiYF55JYhpG6Ks/
yIHYO+aHwUeXrZ4Rltd9DTg5bN00ybP2ndcxzfRnQjicSDkwyK4rclm6fMUMbkYEwBbJmNliFY3n
al0QtGnxKr6ojaS9SI0m/BTaVwn9CbjEoyzFtR/IcpH3nORRfs+K/tIWQ2WIMf3frObh7Kgcock9
o8zr4DycVTp49Sbci1bV1c8Z+aZuv6Uz7lHqC2JaEAIaaoCITAh4DB6k4Je0l+JG7oQp4pvTQUYk
NQYxQcX7dcZoQay/2Lo3qLSmQNbnJ8i7lHtlaZy5Yn+gS0Q5BiV7Mn/60UXLV+KxrQmIzCTK1dpc
zFlF22xLSYHUGvXrOdrAZ1Taz4tLnk0Ku7smk3w+3A2AB/++gd9Db4aXvN4LiUM7KPdpx2qsxTXD
+9v70iQIlUKeyZ3YHhoARp2TdBhk5bGSVJczSOBqv4+mpzUsWZx+OaPKRiRpObw9lrRcot/vdCPD
C0m850NgBmRHYG/ck6x5f/tod33IZMgHCK+9Wwjv1Bm64SVWLTmI2l4MFxV0Llg3UFGkFVVOpO5M
sySt9LM44lSxD2/2dqCVklw4VW1ofmi/muMn1G1KrHblDAD7AXDwvsOYxe0oKoUu0Ri/j61f6Mov
qKbNGO5tSiwjxAUNjynPDT1/2co/g7nOzREbcmYeBMXv/HCfTHK7jAPOLEcHZfA/m4XytLauprHq
OZYUTYddEMVMLJVUiMG8b0x64Ak0aY7e975s60MjQW16vqi3pbJgUM89tt1eWUcVvURA5PHd8flL
TaLe1pyh+x6lvLcmGwggXCm2K+e4aT3Xzw8Q0sASzXlRWpoOR/mByUJIVNaAdYwzfCcjW3cWyUHK
sRY++TYVVOY5if/E4oVRxhMicupeL1ts80RDD4gXe+uxPSIOpGSiPvInB1SvzXpgio7DBZ/6+5/2
Qt0x1r/hl1nLqZisAYIDEaJMYdeEyTfcKA2SUnUUNz4ueL44ZbBdjrXbmhK27JR+WHaoptWAGoPv
b14Lw5fmm0W+gsBx7TI30S/fnuS3t25KurdMnetRjiabVdyyxRuhSANZUemdAwHIbrZqB8lPLfSb
XqpoStk4AFx7huOelz4Sq1eRkQghpqzsTtT1d95GjHtfox6CW0TYStjzQV7RjXuMNLrdV3GnhldM
drnTKrd3UCWNhanJJ65S3/lW8BJ+WoI7CbAKPy37aNWCeyqIHEA3CB86mWMSBjVON7kGotpmSkQ1
5zwhNSPGIr4sx5RfmXk0oEIUUbiQ5kPYet5LANhEekaaBr6dp7AxcjqhLD0JELBzaWVmmxpbR8RJ
3OA5kctxSnVmOjU9zegKXLHzvAE1JWIOagwTj5JAXY+vQfi5rwukjETRcajFFhSrp8TUpMcABxt7
ErDJwKXSP9M0aqzGx/aeQ3T8Flfe/eC096pBChUgTu+GdogbOk545QyUVqYZMUJM4QBv29TMW/yB
JfnLaXubADfREyt2xuELedaDrlYpArbCYw3obwbJt03Y+dttN40uFX9beiEfCUvIh1F4Dz3N2fY1
OmzF/bL9Kta+aKpxdA6mbFUOZRJBDYEzPvX2Up4TaaM7xArCvt7dos5WCSv6Hmr5SPMi6YGEkoqv
NhyfhOLHPukc/Bcb3Pzw5xEKDNXAPxLsyWTl7Ls2hwUqfu38rMlKBTwlrDYdRRlpEYhfwnQ1DYXY
EMDF4A/A220OHBrEdGlyV/e9IZfizcnpeVNp9iaGttFf0xNtHfuPixUowSplDtCjPFxdXhfwY7ih
0WCm/wSZ4YPpTcpREwRwU0AdiBSEXdbBY3aGyISt7MPRzMECjETsYB6nEYfyUmHhN0tNuHs7yiVf
pCzqbc5u1OD4j+8=
`protect end_protected
