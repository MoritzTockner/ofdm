-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
DL24FPfwn8STNjjrlbAHP8k3SS7VeWAtSw2thNEbvvpbL83f5C8mnJlFec2Y9U66swADotnCKga5
tydZdq7VepZZNy314eVm5wXRZSaRB4pp6b+k59RM+cI1F9lM4m8rAfgij6RSvt9JI/biUjJX17wU
2dzrnTixQ2cLT+8iTGBZmixgQ6sumJ/toUgGGa+feXg25q2Jy8+YrJg6jbKdD6HOopE7vEI4g7IH
h+ofeI5gz1EXTkOSk5r859/hQ5udJSmQ5kwqJ01nk9VO8i0ppcQ4pzwVcfU/opvMd/SI09Lwe2vE
IDLcvuBdcWUux8rfwRuvl/CgLw6NZqep44h1Lg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
dHXLDsmeoVoLmYa0//QMb5PLmOoX3SkaeRfpXzGrMQCmIwhBecv1vyxnVSaNEu6I0N2Bvb/WVMRq
SjdcOFSsZ9guwjv2NYfA8rNkP/lpEvi/Kwz0YSd0BFLE3Ho7ZdOGy4DuUmcuHxIaSjFUFWPCZiHH
rTV/O/AKCyU+rPom1xgBAgIY1NPUcNvP1szALVWuSbvEplLmGZSkclza92OZ1UMPoP1LBd9Mpq6g
VWvBs75c710b0lUz6mZuNIRTIekwI6MXxvXz4dhXCP/dqQ6nrI3QQiORYkhcPMQf8FN+OkG3L9FR
I25XCsrgbvR7ZFvzB6uTPtDKbW9O9Av+nsNAiMKIAw3ZLRufzmeLORVRnwMeR/YJC9VydOvvLovC
nNprn2mZiKScIa9lgdKoUwBR80ugA1sWh1lznCay5TodAkRwNcc9BW11r7MsKDpHBe5S2VaDqA+a
AbQNSKJq1bHbUW1wB+reI+TQmcOI3SoQzZAWsHREPTvPIcWMFxd6PcdXMvvalYkQiUz1hwhi+FQC
iKHHyZeoFR5ivDakbJ5KP20+KNd9kf3QLALyGT6QrNih3P7PFDQ7ZuEY87iFK4B3HVHAR8mUdWDV
FL153CaJ0JMX+dgwS4raT9zMj/VtG7ogik70DK5c7bQ/GsbFg9B9KnFHXWCa38PTekM95XgQeRkC
x7PkF7os3im5qOgkyV4HHiH+vFWOlJDJ49v3slow9h2kMqw+h27TYWlHBLQ+QzGLsNtSY575g4Fa
zLCksJrE7uU2uDW8hGZ5n+d5iUMcK3ThlUbJLQUzuIc/UzUMs0ej9TE4n2Mbpjjx+xx2ZmhomCzy
remKx0fL+GJVSrYo9s4rAlULNFJUZCACPEOkreNvZdJjU1UVlu+6YpEMSC8bNKTsd11a62x0rmlf
t7xUR6fYVv8N4ujo7d49Q387ZL8vbnJQhgl5wZlqLv+S0j41AFoevgvtCyWPx+p+JmMsJm7Lzg05
wKT9DB0NWde+wXT58TFCTVDJe/dP75S3IcsqrLZ3UnaEi/75Msee0AR/jQorHMZZumZxD1FW4a7W
7Kw8FcUJECS3CSjloTgj6Q8tZnUUJiFRjIJRUtvsWfg4x9xlHI+BZyhL/c5mvBR3tP++l0El1I+4
Eo/3s3q+9RrzGeGVR3lNfC8QgQCV1vpnFJBbxspCIYppqIb/sivwLs7NRG0SasNWp/8gZM/FBukj
u9JfPWiP+1II1/Km/cA+eQeswZiBZu6nC9Q3g/tPVK6olvFAHvtZKDH6eA0zmQYb6u1lGtkKYmlN
i9jpv6rdl+VwHabLHjzMpahdMsQ2NZjBMthnXmLiyn1keZERy+nMfVBl1yJBxN9ObM6oI1F95uMO
gwmurr4QG0EksPiz8KlQgZ+uY+mbl3VUMYDH+/9P3KoiFGgYqD/Kue3AdOdqHflp1U5gwroYknYp
BjwFjcrlP110cOMapOHsRFkwCzs1wpHqTBM1EgZOep8NwSA5Od1RjY2IMOyYr5MjhQnNnwXRnZPY
4DTDrY+080iQQuBEKGuCGR8xoMAHEsi2ETcl2bgqW8XWCpqWqwxOcGX2tyRs33Phs7XoAFSc7phO
DasyWEVmZ9vdNwclomF/yzmaqun9tig2qViuIt396eL+OTE9FP4PoGLOb4eMDXn65hmBjz8Wlen+
8fbGrjsrBCkfgUkASG6MGm7grJUYswqcTzblzdNn5ACzdrV7CxX/3uFrGPB10+kQdumvRusYiOcD
fs5soPD184CtJ8/yZo93mubaRicRwwLVcfNGK98N9JP75a5ePyZ2ofBTyzCD0hwFT05OlAMN5OcO
zSm5dmBdJq4siPlQCbyTWs2ZcYuCTkonsxThNpPbALfh7Orlb4CfPM4ozAZEnxkk0DjFw3/BaZmN
C4gVgDxRhTrcU+VVadWa53ILbrqRZEYzvKULkU9pOQ6xHXE/1f2oMbl6NGcR1N2dHjekGyIgxy7V
UhpemXiupVSmMVOPgUbjYNGpG3Wq1Z1h3+XeDM8QovmlhNuBT4gXcVZFup091YIRosbxCFqBV4Hf
4Gm+OkRU+O8IKHPCyC2ImN5so9jPtwilAHuyacto2oAcSINueOQ8DSujZdCblEo0w6NWJjxx21ph
kere0OOsAay0sygQz5INvYnPFoDsBcdeXdaeyfp4vtcUf0F+qJAcxTHxkKzqEuqKpmCBgGo4fz0z
2r9LRSRnfq080UKhM9ZYJdVlYZaSat7pFF6huerQAOtt6NztKkdR2BkIZwGpgIAkzQmWTXemJTGK
cacrxQ4meEtGDsWhTK+JRM/uqNPm9UGkOaZcnSmWoUkX+3+G9wNZ0DgYR/8lh2WnQI4rpZRMBvH2
ObRME25xK/7ZBiPcg2hE3V5amHp8utog+xpRUudU0x4s4OD6nWDxa/tQTxxhiz2DYzO5ljscW1/e
pkPZgHbc70Cr2hcBBj15cOnuqSdRZeKtDoDCCaHO2JkPwYrPbdGQBQgyshOLUwI9UverlBPu9aPA
BbIan8JXDBcWC4U2ijJ2iJ0pOWGiJgRfnPUQdZ5Yg8mbk+8R5tihfUyfFrh2iv30wF+XR2elYt6i
Tmm1OeqGw49E8YBfwZs36m+vsQWk7rL0GoB3UpqSKEy/dvcfqOyxao9klu4DHdh1DEHxIabrzBWi
LJ2g5KdjSIIag6z3tq2O8uvjaIg3Fffl0T7hgJ6RAmN4CheayDxXTSHdyu47yW4fs2+PZHwCIwP2
CZWhiM4MkQlpAgDusWQYafOIbIYy9gmH4C04JxdJVbFOV0rcxv0lFjhv2sd2E7it/ZdHjCjz0Zj1
QskznU6EnI+sc/bBmLiyh1EOWfd0r+rQ+otptapUjdhDfBE0ZPa9XlzpWsnNWC5A/ipyzOzQkPhZ
rfUNIluSfc9ZtXVeMEYA8EEFCyOgSVI+6JF+CWKhpCusW8odbwe22EDByxXen/SmKR0AJ95UDGGy
Bs10WDAhIEaL7+llqrlOAKk6Gjx5Eo9ZLYo5T+loOIw9OpN0ytCxtuQ9oNX0h4RzMIx7p7QB3jX4
iZ9C/hIvxe+xcjQBkalnlYq6f/SsrreKwXBfA+lwcrm1Bfq4hUwSDxJvnSCeqC9nFyDEo0zISMKX
Is7cpjuBVZ5uJqez9hPTpX6t+rNHLNW7mK8+fqIbhhTxuOGOWnlNnFA12LSkalZ+p00X45OAA1Zm
chWjhOUs9KQqlxV5t/3RmVLHLMH3xVlVTm1gLBHaqKVhWVmmfEznRkoK/dGy66p8/0RvQQzEZtjj
trBaivdsY94bj0+icYV8oqQ4Dgg1Owby3iVbTqRJGMVYvr3C8OqFBVa8ZlyijeGTk1tKVwpHCyPe
72QGv2MVXwq2twP73colKQfI8hxw7zdWWBLybMQXHyb5L1rD6dpkIafFPUxP3pNMFb1X/w05LccM
VhfYle73XJQkN1LxhO6mOeiMSuz+BOiHq0JbIZATFRFt6YZwxaX2Vf0843bPp95K8yTg8g1PLvUg
57g9o+/pql/QeaK3kqfSjbHmH3z4uWPKuRJ00hlGvCrUvNspn7zkEqdXZX2gFm0ch+HrFlOYw23k
avCjeQcUKBM+I5XtjrbgBFIXLkoj4WXql89YbiR4kDEMCZirtEy74dErgGu6i9vcIp5DvTwvV4bq
uH5VCAd26rRXOLmD9WbOZuea/BEiu8c7IbjA5TI2AcXmaHERgUdA5vnsYIkenRDrowPpyHMIej3r
RB54sW/ii+DvVS74ymMRrFrRPg06mMG7NFABwme9ZKq8rqduADrrhhEBRMcoTcrg60sWYBH/mSl0
+0/B+Zb1NGX5rQbBz5T6uCvTCtWagldRa0GRTRXK6sNpe4im3ZKKbhqpo2lMtZ/T24VMVvE9kQ6Y
FoWXb1rOYT+oXydvt7O7mOJVu3qirkk22LMpqYaFsc8+CUIZcSiIiaVHIa64Ogqnds49wzp8L8cg
SUokYClLeCpTU3sxB9qW7DQGwdZ5Uu9PVEDMmPitcOfFTVB0b7wFFc/nQvHum0hSZTUN3sTkkLF9
vfX4Q+H29n3nyHd3+2LJvPKDqiNYIGq/IZ6eERD7DAqPwVKeiMSYt3FFvYDLX9mdohJW7LKg+EYn
t+e/enEVx/sf4CcI45v26CXm8z21foUrYcgdfK9AQ87LF5cRjf9HGLUyQZ1LfJdF/6dc9Hk7M3Tw
acrZdwkR/c36oYvdki38ibErskmTNW7uTeK7Ze9MHQWnCB71xL5aGN6fjEXVH2XxfcXUAY9OXWhH
z6bNnrsTVKfRdXvlvvDrYs1ZdEzF3Z6mhWNBhuZBXPWWzyYA/D9AvTml+3F1u4q7KVgC/aHhmTv/
IPYqXwJw06HWKoxzn42GijkJYT19p3jYNbAzsZuNPP644pdB+7VUYW3dVXSwLoCVbk9KlMFf1enl
r6Bv9p1stir0PEo/rOPmZfF+phx1HWWTlrhlgEf2McAp+iR9b+pnjuuwOPQPKEhsJyLbaa9csq+L
++fyF1QzWxmu9BY1IiQwEPJ4y8avPRj0RSc67UQyNrYSMhybdUcrtVo2gHicWQBNuVrsABP1MO99
37v9e3U6HBOaTXgvhJf0SreU4BOAgHfQoV7fCpOv4MOShRJ/prdVy3s1v96S1p66YIQdn/HKalEA
ax8ZXGwWXXfVq/3HcHpyaaVierL4Hoyy+ZyB5ITDhw7Yt5NbIzIf9VGLY/gwDxM+OZeXGGEUJiCI
UTComYmkFMlFXnFx2AOjE97FEo/m0GSkcK7JxLQllOzoTiulRiwwnYlTP2dNh+Cv1zbjkIsCTB7D
WJN4h2FLgWftRX8GjCU7dPv8hVltS9rkIsF+k4diJmysYYpV+TMXBRVB7p8rgM+7pDS1Zo9/F9bc
J3096HyPzwMBsR9HulbyBz1EmO2YRxdTf0IrYFcUlGEI1XaOY6hVXN2e9o7ENPQzSyChq4Gsa/17
kQEpE/4mt05nixZG2qHkTQcHaX0OoFViydtwCn55GVMSTu8LWBGjEE+ZuwAWbleIqPkIvEWgW9uf
i5ZRjJhc9AsFQmCkVlkFc8YjOZJYh774TLsLoj1ViYnL5E3awALvzq1ihR8CdCKXEb0slft3pgxA
jn4Z6FNDTVujoAahIqBrDenPzPa2cdmica2jATgM25+zMDy4z6mu0FtnnGbDbBBhp2t5QQN0cMW0
jQgjDP6CD3xWyYcRrAQLuFJJS3fw0anzEXCaKzLS10RLw+BEKgtMLj79I7+nExOZnKYn08AUlWy7
EzTFabE43zk/OE0dcsY5NSLau5UyRkfGhRiTszBrxdytFb4nOfP7Q6hULBYo5cg7VpiyHm14awZv
2zk9SIJxVxOKO1c3laoOaZHqDfYcNjFmlYKgXGQT2M8npoFOazjzOHLgGYbQjU27VTvpHi6BcfMC
V+8Up0npQLO/DFD/CPmaf4TsfmyStuHCh5zYg40ugVEKJY/ujzOPEJ/+PD8tYtJrn40dg8pvEe7E
jBufcDYX//SZdMQDqj/BiOJtVmUdJWp5LzTYvdvpYhPz1hAcH51bAygsZJWvHbiaqvHPM/bSxlwc
26QFGLAjZi+rvMoQgPSeowiLDKiEmEP08vxHsq/6tHA6fczABImjv9dtOqo6xqhwcWiHE2ZsclGz
O45eltiPoDcmGwtv67usIyob2DtVfi4YsFCDFgzQThWKK4AuBWsAfuuR3A91ly7aOuoY9y+0R6fi
VBcr8gU3QmJbebMRp3wG8iMWQQVaEhCYNXdqW1Y1+cNlP4CTymnYVlCiEq66FPl+Y2oeHEI5kMb1
NwG2pN7ywOzVAFP7cp6mgfgm45gVTOSi1RAVBqIXcrXzlGmO6tmNx2F7eX/hO9mj5nGcE7gYqIGz
se4MfBRXcI1IMrKcZmd3IBo+2y7B3p58syYmCCORVCZ4dojEy895sdNfNhikhmt/6t5pcZ9OCA4M
SUsOs7bLNkijuwjmQs9Cq1MDvqenqVjhkxUZ1PdNZOFwZFKXDMaPKCragQIWLZjbp0KE86reJlKA
6TitZGTBMoa2GcnCbr/5KRFY8k+SdFP7knqVqXqkwub+y2QknA31fR7sq62LjC5WDKIhyg9DgVOP
hRDdijbNdBvisevzqlYT6i6U2Pdbj6ff+L9mXuPfF8lQWjH14SBXUKK3+GXOFCg/q/c8XGKslrZb
XgEa91w4a4NGkX81VvJU0itfSscM+4m5CBIm4ga3Mk/P51USbVCGacPBvVMPi0xb8CboKd1pEuAE
wUtloLQJfeTq+sQyvmBavJ7LrqpHKYfBvZPMEkh36py2Qp9F2OGQEMQmgEWTkUr31fmnYH2QRxX5
8w4pdkPwDwPBxq9+wV58+I2tVLc+QpLBF7tddmr+0Nxhg78uIk6TU3fCMEQ5gZuPG4f1wti2bxQj
KWGH6shtwlxb91fvoNEDCIH+eHBpYD+H3MDxNLMtPjoStoMq5tmHSDqQ42OnGhLnoo+MC2QIhh+m
U9YkIvdQvSV6b9cGwm1DTKP2dcn0VzYTYulLqTXwtbkItuQzeNk7vtiOw+0SZeIxK4VSHvrty209
8gZ7fiMaoCj2msR/SUAf1jxueVjI87PgfmPVKJ4noNtI4aVqnDx2PsFBMt9JJrIE9GZ3jukTtS9v
O86vMQpofi5vKsCzO9ULYfkm8PCMZVPG3suZYGyGTbjYJg6+EKg5jyzzlxTh9ipdqUsuK/nFlv8E
S8z6xIdmS8rn5VtnmYUlSfbZjFgxO6Q8DvPUWQiIBLqsWAgn+PaUAjMoCeKefokGWl0MXdKKJEHH
/qU3O0p0aokMp2aaRweRq9eUEu9dplL+U+L8SCSiK/EeAfznpAmdXZOKCcM94tYUYg/VqhDAKp1K
ml4NB709R3JBJneLaTI2zuD3VXX9ptZGz9FD8+FaHrAmvzdxNn5hVXtXJp0i3xwOWrxPIq610vjT
R/mOU4+aCCx6G6Jrsj1NfQlPuAwHumHpWzmbfP+IE7vlbXPs2l+6N63CmUS45kpOcommPXo+EY6/
T+H9rZ5btvmDmdReT3njp7qDOZ4TUI32TJ2YgYWIq1whEPKiHYYuNpgvfELP9gesQwyaSbSGljC3
Jo58ZzVFki0Vwvhr/u1aVuMahMWSs0NKMKK/qqRF2NkVWmqFLhUgUb6PiCLpgsA0nDs9xGbd2OV/
AaJMZCJ/HQ0LE4/WCUCQDeaNiVkVVo2miThIe1TnESjBMvGXdCMZ2GZYHJDWWwM0POaUhQ+PX3WU
lIT257cfkILvhUWns8SXIwqaTrNY0YVDohsjOOEz382y0qzudQgYH9TKGNfSQe4Pmt7JvSTFTvbw
7kySfeMRA3FaWC4E2ImEMMdUtivlVAK5ZL5X0UIfosd12iRprky9fpn9J8pXShMWqxfdPmjQMbID
cwpjVWszZLqeevcdFPkXk0vAgf/v5+EGgEf+sRGQ2Hcz3x2TSIea1BRBc0Y6jr2lrpQhx3EgUpmY
NUwk/GxqUkRWwOWOmj928+sAGWnV4XLXtvYskz9OD4jJuRyhKg7i7eZgU/q0TV//i6NVds0VICTa
UrO/NSie2sdzibUUXRojwi4gaiHLMeHxY0vQaAWUDpR8L8dKIwInxa4iE89dZcv/aKfXi6y4A0PN
z9WtKHoQZZD6JAYWvK0aAJXx2/FL5wY0Nllef8azitesB9fHaN4AYuVqAz+VS95Sox+8QcI6iNKL
cW3pSiaKkLf6oEj1dWi+DdRZvz5pbZCcIe2Z3qX12YQnG/3EvwHZL96DgdT+G14MyDkbvo/rkNuz
ruk/Iypw5wJ2VnhBNfBJQv5OlE3uo2wNBh0r3A3a/1MprJ57RP7otyqEdyeRhtDuAcrUGWIWHU+3
QjdafU8qlKboy0vLtGzbeWmId13fMkAwXOS/AAseWbUZbVh9kpDk1aRPDN0cCEoZfw9F6M/3UeT3
EFsi4bBxKNkF+XKVx3UFhES7+B3cutOrMYr/YEBab+PXL4VcVy+R0zAk2bf70IYigi0kc1S3AYNt
d10Ou/Kkrh+Ct+S/rj/1oH4k3bBWwYEPZLQBlJ43xJkBp7nvDIXJJDjBp0XI8keDmdQWwKyrNnWf
2Jwz5QfrGHlKBUc/KRFO6+oz2yVEt+c7r7yNmO87CEt/Jbg84OhZ9f81ZjzItfq40uN9pNxdthGX
8N1ESxZ6OJ4uHUpnN4n/Bg9VtwU1gIZbtz0LVlUIbmlOAgUH6he2UcwGALtQOBqMjnnlilUKbWPr
t+MBXdMkkMq2IAMm4zIRQzeRKMYogcfdx1ad0nqGOT0tJNGVgVNJtOLJxLMyjuJn3Kr/j6VnzrDA
YDUDRS1tuM1qjkszqFFkyRJzcldwXiFa1kNzSHmq97cZXg3d/KECiV1OZljOzvzZt0OtSbgea5UB
+8fMrIe6dRIIcBG08qR3LSEG+Bc3a03mcrys/vwWuuqTpMGKq/4uaFZsi4siFqIdkcGTxUQyBzMn
c+7L1ziYzzyk+6iDz3UN/XIqLHf5X/5bksh91dEtg/zS9TwMhh8DieNVJ9TUTYD5/rjsngmzmO1r
f1yW2BevUocigikZeobwCkpIoKafNXkD5UyzyLnXAvO8uvOtrmKrwiytOqkBiE9qTQ0p2+jjujTu
GcVuQ+ZEJqesS3mZ4KiU7r0DclkNvXXPz4r4c7lmqoxyR7b5nggCaGEVQilD+TpGu6FNK0aquIH3
pgWwuKS0BA0bXyLMcoE8kDb08CXvgr+8CW6h2Kv/DBMiHjgOYg+OIAOCN0gbdMcYvKWBRO+xtYCY
jI6EmvgzFDp5tQZy28zuBcTyReprgyc/1+UBTF/xPUZODahXquGGSjiyHB1iFgGbapcwGdHkOGn/
z3wOw7I+CF5eQyTfvk5/QiLziw93CEC2OgXWeMl+And/vwVOdFUwJGXRxijV+FGdnlOTX1UJAVBY
MZmdqhmYuIOA0BCyiwbfZ93N8JvDbCCDcbNY7u4hlJA4UTt53hLRLKdE/YVKG4BY/PveYPPeJA1z
TwbcKk2TslB+lBaKjG3QrGEPFL/kaAPitWeljV9oAqkeqCneefftA+eugPEGwQ/zC1yyKld8y+Yu
lSsQMPk7KrUs9AbufLw2c9W+I2Rz5iNPd0vnPqBRElGWuEF/rp9/rVmygPPxxQzqVwVtlWIJWiDg
5QpDn9YYTRYtMpAdIaGpOpjxf8vWLtmkcL05ULg1O5+7OHOsqsDl55yVbJe0NvwBYRiQW9fazS+8
Fy3sR/xUL2HLvoMCPmBIjX8y+Id6KRNbBI/nIYmrqtiqpEFrpss3w0VjZUmC+nL+7Xd50joA3TbQ
6dXzLj0tpwpnUg0QhHIgYK9cpbpZg+VKypv7UAca5Md5Kyu1djWk2kTcgeDX4Sp0NAELOfCeRTxA
BNvU+UMHiEd2pdXv5F0dQw8+kt+B7V35HyV2XnJgP3NGW9ACoj7qZMA98xABMKJ55wODRrLzazJA
zVBTBJpzpPEASwrBxMQ8H3NTBTVIQas+KHz6eYW95p/y+X6SR9Gj3R1ktZY2Fd1ZrQG3jkBgKOHk
Q5x2SX6GONAQhzvubf5Qoj8/QIfH+60S/X9CH6lJV3m7TXNEU02SekfcyQGM6HWmeK/10FX6c4GG
DxEg2EcS9qq9VFyWxO/J052MBwVuY9Jv2LzKIikr69zJWGNL9A+G6xfvL0qsSIJz0lX/6UtuhZEN
RGKBp2JE2/3PVwMB7M6oWyndUpy15kMGIz8IfzURCcs/MvQUZUf5RNfi22vQTNqKXWxgTnghD38f
GNzceeFeVhT03zXPTjO9HxqDjEj0saZs5db/qFEq+mutghIEsQuxGNWkFQlg32SmFNy1nGNPAeMl
KMr1qtUy9xYkQdG6FOb/beGZGMel0sroOKAU0NBe2Air+H3vmCGfPOXlBT5SBPeVGPmOII7cMgNR
KUccSdlPmX7W/dJ+rqQY7Ze44y5wUQwsu+y9p7p1Y29As2D/eCLxbc/BrWbnYVs2AtvSp08YrBYX
G7i+5gAhINErIb0nwrbVyeqsBcQVca19xGQqZrKkzstbwQCCkyeQY4Omrsx52QIWwdq137cteKyU
rBsHKtcUyLLIK0EUgCMc8TcCUzmI+v2KdICGzQI5blDSSLR8oznFNImI/TX2d/PqccJqwuXYdFF5
5BOeQi+zj8YIidXQJGA3ahLO4+N2UzXYSVmLnQg9OCGMwHAng1Zjv0ZIJXgLNBbv2bPHTKRSjWBs
oDhUdACPs9VLiQg6v2CXmDCmpAjJuL7zE72P1qZWFIWVAN2kzHpWyVfqamjiBPRyBapi7W1IFkvD
I0Hcwrx/EK6p7v2+enpR0VzezR3AfyMgXA9vF5dPTNlNSGrlUpR/V05BvjPiMeNh25z2ZCEMvW2b
Sjit66n5fcCtbmqWB2Nkkl+PVTyH0oDRL15PixSCRjF7B/z3uUAxRvVDQQuMQ8XMie450et447qp
KKV/MenWlt24WEXg7YIjB9qI2t7z5xNanbg8rp/cJ3C0ZdJ7jDqCO+wBuIG3x9ohC8iBEvwd2ozD
QvY7KZxPNDC1PhcocPevCiOVc0m9Vq5oXcr/A+PK0kmosNZ+nNQRSCSeUvVD34ManpCKk7CQMqki
k2OKFhTcoOeK/YQao5swlyWiq6ZTyplSgSkGfUxesHefWCDjQeFSWZCL7s4SwvblG4AHRBzXLRKN
gBo4vh2MdiT6JTkADnCLSjT7Rtgk1nhOm+3O4FsRWqjAMj7xFyu3qhqGqAl1RAMwaJfKgsrl+GTO
+cnPYnxcU+XDTW1IfdHH9JbNRlQAz/DyUx4nEP7r1NDNVSonvOX2q8UcH6Ux69bf++jvflZjg8u4
8HqHK3wVSZtjoQ8PK6JoLMIgCZ7E+mUlW/QRZgvK7ypNMOgbNg/YaU11BGzfkZrsEtFDNkVnWfct
WMgLqdIMfcOIkBhWlIBzrxeysM+QZY6gshvUFIjWqzBwZquyBRN5N56gshKt4NFvaAbzJNf2QuuW
sfLLXHSqihJ7FwO0Bk7jZVYLG5bvg6PfDYWrPyY55h4LHHQdYpkb6zDJafny/SMsYF19SJOInGKH
MZLiGL+PpMeg1+OTc5s+dnVI7i4p2SdPReW5ik0PcE/aWvBKyaZB356AMkrAu6tJK8XnQKCAcVIN
b4zq6ItzO4rQdtewqn1JkVhqknEhk5yZdWmwSkoE0jOQh/k+oCeBxjTJqFnxTFizrf3kBZTsH5hc
vflpEGCbS8bNYHvS5qF972GhC9Hgt+38CBSrGH9weXK3YlVaYA7ZGPXy9/lNIxK16AAl7H2NA2aV
qSY3dve8P87hKQR0xzm9rtx7kr6+VRaqzn4gecpkBgcSN/4QGY2tFn0AZJBA9loZQ6ys3k8C5F05
TxWnH9FE1DOxzVjJnHuxLTWSdB8IeXB6pZDULYFTV16Mnb0x0XHhKWmg01N7i126Z8869+ox6I+j
MCiPqQkLF0TkeebiQYG0wLZ2ZACgAblLjTCdJyh8HC0HLkK5Q9RwX1olGs9SHwTl6iru4Qjv1QZc
QYnFYxJQunW4P/bgFLAjHUbFN231G8Fi4L2ekumXpl4oLYC4PE8naYp40QoGWq0MLYFY+EGGJbKg
FEELWG0zQ/3gL/TLLsv55TJALsaV4GmPd+/QIlKjXfDQkukRyD1Dl+XbxAEXlR39TwEqZkLTQCEu
niEkw15z5GNoXwcCQMie0iRVxladmGm/exhv2kCNYrwBa8F+9HWCZlM2cRV7y7RqXNv6rRAAm90b
EN1gqMsvFJ4bKVVaP4CFGBjG8akYC3b0YcEW2VPjI55Tfc8KdUPMlc7JOz9cCze3MC4n69kl16jt
FSV8oWPVcS7HOEDOBvpyV7E+Qht4W4YLbD350I5NwcU9rsq7Ke/hbGs9sKX5o2m5hcrmW8wOvMtl
LlHnEGzsZaZHcLenBZoxsXsAQp3eFYbImheXWX1DpzpeZ+gyHsGWhb/gSgMHy8UeQScMz3FLtzaT
hzp1VCh6PD9B655VBxNJ9EbiYn53HwO6id6f+ynQvKk94n4nE7oanOs4nEu0GIsVnY32BwCNLF1+
Dtc6nvapHqTnxWJYc40/P9KSleZKO7IRxsBZSXSU7HcKYFfslNfPvvuSO2gpGYN1IIOfJQ3lLn6x
McfiKYM4AFcVo1eHI7axaTtsffWt3Fjlrn8KjdX0vAayJitSUhpJqvw3+QE244ssmiXmc/vVYaro
qktWn/umU1A9XyDvN7OV0bWoIz/vWcbKQjb/GbmLf2KZgmvjE566dPKyVhSwraUMJcYeln6/0r2l
anunyAN/cG9+Q4rQRzenOH883XCUfvQ1z+rPLbSsHa5ldSFmq0e4WgX0FBAkHMYxSHCqzRWgvDMN
GRHOZsNhNZuQOwG1K9qNradZR67AsLVuhTM+o5T+yVs326OtXC6OyGn6zk85MGimP+TqLDOwcYXE
XFVHWp1fpNu0eWKK1bnT0g3tstan6igpZhvgVwn9DDzvCQfiEtC3apGvur+KTpLDlEfoJWspnjmE
VG+6oVT52b7RD3f+vykT0xxW45mSi3TufJ8QKH7fZeNJzpUGE6KAcqIR1WRQFu84xLrO2PYreD5C
yfp+0HbSfxXSCgGHDUy45fw+Juwja8ig9IUiMth0gLyOWZAExb2DvcPFd8smku0WVbahj6GLJVUg
WZ2ks2djiN6tVWJxD5RCHRRNGFf7O7IG4ujjo6qx0gD/QgRSyXUqSL1n/7NFfwNk4T/evPkHNJb2
UM2ftBu9wHvUsZ8FbMRb0gXhV9aFZAHVkZTt/bge3Gxj8S0Ozl2JbxDo5K4YSok1vlk5+2mgYoqu
LLg/o1Yn1Y975CQk22v20W+F70nnr7C6HpeTxOnYlSGNdFlRjWQbJXOMOwwnG9Jq0usmzqvGrv8I
Pq8xGZVBJzAPPTFvaBlV1gbdBKDNrqVUzbJLpqlVgq2VUNi/ssZ0UivTn7NRfN+WlDG+w4OFBWNV
IGp3A9I0xVvS4s0df9R30OJrHceurEefGhxLRru5+pL1aQes7GckrpSccHMm847ZfisY56WbB2//
LhVt5uZ1sz1F/291ARlsX9CGAliJBRnOTeWozTZe2o9iZoIxAEeJcRQOxn2qEZ7q+F3XieD0RlAr
P21hCyce+HOMJSGsizJ3MwhTqqtEsyGH+rYTY5Cfx/M0HMvPqhPG0feSKswmfoSgBs957Y6Oj9f/
MdrhQ6uSbn88A4rv1ad9tMOVp2A10MBmP/RsduPX0Ib3q6pVVxlcoPKNglnfM8R1UXSZZrvel/SO
9ylqAC3sUswTSCfoURSZzd9NDJ37HFndG7LQMjffuCL9KdbD0Fc3cCoVMw5fuNsev5ioI/jM0R10
aHyPKpriLbcvh0gHp2ATWkGY96kepVKGofC6Q624MybiqIJuDdOHEpNDko5GhbPw825HnXS0hWLx
7Q8iVlIXiCeMaKSmoZg00Mmrepx3lM8ApA5vSjuH3my+t8eZzmcuXqx5IdxAbQOeCo4KQn6lLCjc
KKEuyrZSESl7bklGRmVvv0Vc8B3T8J04QgohFgFRwdNnsCF2MNSf3Pn87zANYVExxmZMiEoIM2J3
55P3PLdbuX002BwXlX2XpU2dddcdY8AxBZm89OagXF9phYX6p4gQpX/d6y3q6euZ/zo3c0Ibuqay
kRG0KZetYPnzJIL0q1p0bn00N/SMkJgCoIMOzN/2ghZkEPqGZmeJ4/6C+IDeOS7HcoZgLx8V5beU
wY7iEhXTzoEWaIK4/8b+gllpnsO2cj9GAvgWijvZa2Tj4jcd4qspCX1+PmJqFdqwLn6CvSDBCR/S
mD3/WGGdXfqFAdo4Nhy+WgqMz4OcKsb9+zSI7dVgfb3OTKPQltY38p3GJscVdSQvODLcx966DCmv
zQe7aHqWkgT+F/9xaDc97ofz0HNz3Ujzu98zkZtPrdtW5YHoQW7Z2bZGv1GRcem3I0fsg2hf/Ysn
+kFyXrsWQ/Gcky2cLp5ojEidG9L26sSiwZRYx4eXiOl03N3bREodZxhhjp2LCyuv9lUoTqz8UZ8v
ep81hNXEYWD61s9i68d9wAXBAM6pEwtaETbKH63KbtLyO7Gp0N6VHOUchCmIC9x0EVeh93ERam6z
+U5kR/lrlagCP9xsSXI30a1zXTOX7cMEYn9HO8v6Ct9/AmKO6870mavWVUbALMWxlZsC9939gqIk
ynEn4GH3wBSkp/1i7gNl9ZYHBEC9dhH//VXXUehSm0ym8PIDfc3IbjEu/vTiOlFYhcx5J8dgLkle
jxZQ1442+0v7TaZ7/uzx7fQZowpTP/u6ZIAD8m77nIA6ozqIX3ZAPRVCPU5e6bykiDOOV1RagahJ
B90LB44T98ncmOBz9XXo1rVSfjH0FgV5FTWtXxlKlMuxtzH113LagN7eS/K3E/Pdp9YrwgIZ5NN5
g148Ss/lEstcF0CnP1X7kIU9dT1jVvPfXaFVy+xW1NcE0nUy8+eUBkAdXCn5jj73xU0duZa0LV0a
rzhYOgQP5sdpMkoTUsl+dukZG9d4xF5Asn4D5hdMstLnnWbnulG2ufqkO+6gK/0iJ1mmUFBXhBT/
UBDfpncVWiISN5JFLveT3R6raTL7t0yHG+roAjZ56mZS9U3NNg9QRAltOFPVzfH449uM46etoIxm
ZB2p6aNO+r5G4ON227k4HDILryK1NRBdmaC6hQs1r6zS1MebJbOtKDvE4MB94X1oYGQDkOm8q9t+
dbDmLLpwa4jwTkdPw0ig9+BgMBmNMrzbj1mfIAXzHTvcPvj43t10kFTGDn9sVB0v79ErWreUKjTD
84N03mXO6ea+6dDZAu9Gds0xqj+Xpw/PaEk7IdbGOe5L1qX+iB1ibXT7nrpXWv2mmvxLUStNse89
GQg53PFNFNCR+NUnhRHyKpLQfr/7ZtmW6cDVvBOxS8cRmroChFiuehvMzVWwYGXgfe1+HrgPPD3l
D+c5ZNnWrlGZSAVy4O6bX4Cw69QIFmwFbXFX02SflMFgwLYalyg7KAL+nHwe4MegMof+0FtZsXO5
p1izCYamxDwMwYTjmah7aiiYRhLL4DivEsEmBsiFvR2RerTmGC1jK+BpQtWBTluXvYJMHklX3R0k
XO1Kmg2rzfB2dQIwss/+gORTjq3N690wq/DCrb2LnJhNtqjH2wAE4yC+4XvSmALYFq7MNfbA4aqv
feNoZ7ffbZv+0hCzPxnl+yMdr9yHdP+y9EM46UM62QAwIYMD6k+YjEnUscWcbUs6qNE9Yw5gxOcS
scuuNIevVPeVr/JvvKWe4pKLgd7yA8yfI+x93Bbsx/bx3KnbTMsESQNFgknMqhgKvui7uTzvylJl
rD75RORV/sh/dG2KK4renIl+q/ootLSwisqejLA1h4CRCututq9LwX9TUKAtqYFEW6Pn8t8/fJHZ
1KcBq1ZjC9jgF9KTUDPIEllHW9FJUT59ax+gXKwW6sceB1Mwzu9mQY9GNH96peI7sixJHpvvLO/q
KgYR/CmwFwrF4ZsK+e2q/m6R8mJ17TOHEkj9lrJieCulhfwGxIiJECVW5hr0+3s186BgGQf7Xmij
3DYv6HAu1FcQiQN03psBiZ3CEoswC4F4STk3BL5Aume9DSttckSyZCNgdNQFYWPhVqyptVGUA5v1
AoFUSMmZHNKT1R/OpCAlqGtXUvOrzaAJzJyO65DjyVQSTfbNzGt42rqxT8CUC+d10MtW36vUsD0c
SKbtU5sCkkyPitYo9ba3Q3zAg/a39LgpB81WRWjM4cLS5dw47Q3dWS2Yio4TruUtmouB5DoHU23Z
ABpQlWLO6eiIbMu7ibgAtb8QmUYfSKx3113NLvBsIx3xYRzyqGwIry2uw1NWm1bgoiIfCHFmy4hA
IIPqxO2ruod7JH7nbbSMMQ8DYUsORq4MuaZRvt6uH10Wq9sSzd/Gsu19SfDDOBExL/OlCGJ1bP8T
rRYb+6qkHvj3xjoG6hoF/OpAe1/dvD8LwPGPDaTDOGbBp7oVtqC7AWhD28H1L46sILvIH8qx5lPB
BNDNez/sseDHZ8XVvobLfHshpS78431bNVV21c53ULS6I541OR3d5VKbVvmXVUb0pz1tlX7DpdAc
KPHt4f5ZgDlJLtkF3pYhVkbL8UMQ14iaBbaVRpUby7wH06WAms91jhNN8+Ek/RL7Srz5nl7rafb7
T9SmnWNUf6SPTKqFIHvNkEbrfaiWkxTzj4IxImGwNz/aJsVgDbvVrjMYR5azgX6BHLe+pYQag1t7
l20k0WZAKAJnhs0RlKu+sIr2B/vjW8Ihpj+4xCpQQpwj8Cy29CtEoNoF+39P/7MmWOVbVd8PJoog
RmizpVJjGEtj0RC9mHp7zjDGzv5KlKGFdnEtS6MjZUgT1GlyTClrZHVRz+lWG+TMiQakEgcv9/Nh
8YoGgKiKreHM20Yw2jyNAj1StpBb58mlg15mwKrtS7AIhBA0xcn/uh783NpMcO/9QZ64tXUvXa8Z
MmDr3A93DrbEuyodYGX0s58twap6+w/B1apeLfcZ6M7r2y8EarQK7JDdq9ekYYxJjSioL6FIak0s
EB62W20mzxNg/eCRmCsuOjejS2zmw0OQ1R/Uvp9NRx5TucBBMcGZq+tTs88IX4Kcd9A9NNIER5sJ
5qpElS5Oq8/igr1va4N4y2QAVngjuTCH/qaA/AxfI+dNSp7IsGgsWr5WE7U6eAA2nwLufTYFBbZ4
ZnoM3hctweUuow3nB+QUWofgksXDr7avRhmI15Wk3bUwnLdDFTKNIbZhVyz6THWVIFW5hsEV49D3
LHGVRofg45LZZc2Bb2Mtphh516zsVYgJsS7jhaWAse5Pvz86JQbryNXERiTRT/eHmrd8SKOb2wYJ
kFn5I68pvfLePBrlMNmkU0Njwyp+JKbJVNifh9KitzpBdosgp36eRCsSGxBMCZzKjVAxMAdbACc9
n8ntS9OFOB6i2TxBcMaERW8q+nLcDcWwORh2WuRf/26pFtRlN8wof4Aph6bHGLm5BOKatK/j3f2G
eP0yrGTMgGvVZeV1B7fqIFiGAqrLcyxmSJXB8FpPSiHbshta8KHqnovrpYumIi3zSvV3sOPp1TFW
h2IVNodb5DhG7YqcCAiOBOC2Y4E4mN/5h3r65I/umN3/e3OmXHvO6v/DDngE6yKLqbpfeSniK2TB
f1rf1bCvjMNbQPhJCVEud5ToChBk9m1N83MOFyhL7EeBKXTIwTsMUyAeKfMOEQUWlrbgq7KzusX7
8fC4/kVhGZORUIuiC8vnmwRytqvGGI9/rNRVZsg+OJFQ/9Pfisb4zvRHE6RmbNUiPVZMc9RUGxdX
RHk3CxOagJp0llXzc33mmIvSTTAouJokNh9Tf8JpPhutU0yTxTmLwGhejVVM+ur2fJx8VSzv5oqT
zbdTlJIksbFGxQTSK8mfNEdCPKiWmiAYtNfZjQggQTkoUoH9rPEiiqW+bDCBxeX1qfxrSPl7TfO3
8Lv1VeDOxd4dVgp6Of4NVdJjs6SHkIx+FSSRaV8LiToeDM5ehbVBhyv4qRaoDiJXab1YpXC9j2pZ
Wv9EwE6Q78WAc8AyogNgbU9q0qWWFGH17SFCfajvre2Q6KLqmZMAuWmFg8Fv/kaBeadG8ZeMJcsq
y5aLoIEKLH2iePhWU9CJzDCT97Vp5hslKtxXL0E4tG70qCRztOtnDxXfCUDb1Tr8t93s77Xj4hd3
6byHKqoo8cJDlcIeFvtIueHwGdGp/SuXYCrVEgyjDcAbBgYYsNqhjAZrQgxa1uXRkGrWI1hjI7D0
CqU1VNl9GT3rC+yuo1HEfPu6r+b6p05tT4/p5Uadp5VAhHKqa7h0rKGVVpzbBxXyl5EkqIYz4PRL
hJt7+8nanxOs2vgJgf6nZ/EP6dTNwMaIFKIfk3Cz5Up5MudfpL5gFzt8MTwAZMt7ep2kE1lhQkrl
oPTripkvoQcrtskSKcmPinP6ywXhHVFOLtnkey+juxRXcjpLXq0d01HSLoA5pFHzv76LrRVBks25
lW0xcr066CZ+NQKEzj94Y6+b0GUh02QuQOAebjIGc80QvIZkWmfLIluMvQ8ak0Y/h5jQnRBpybmW
ZxDfKor3016VoFD1eukMx3+biRM+rA6erFErLdNdKMbqwSGtFL3MSA20Pl3i8LBIvr5v+dIPhhkL
vu46lbn+Wi48oSxRKFvDByVkXZ9VzL6/MILgIuMRtPm9iPq/Bxd5fi+w8g3PmX8ol4F2aGOdJjHV
ShvgD+ExXrawEtz388Hg0RIVHS8WFKljSeqydG/pcaCr9UQtNFe4PpBPCVf49YootxAvmPBAHWHQ
MNf/HJ1QLYcvYVuow5M/TQU32KhJL5XhsLwYvLGjchRbR3zjxZXldhI08rVut9Da7QOOZAysamEP
Sv9+b0Zxs8jrbKHGQuaDeiByjTGgowlPUVKCMhCzldGugbtnE0G7+ofkc9g1YJenyqZlmOiohP8D
GHXmBdhlLT81iFHQel7oS72mUZIh8jD/ld90NkJWYYHLnx4ILc7ux4wSUXhRWJh4pSUSD/xxu1Hl
heFjDDct9z3pST7+Ln2IvULjs4dcTAdEcwAF7z12pli9jlckUSBGhwNEedjq2kkR+8iNQsL5kDir
GG42tUdLvWR1EWqBNww4X3ifRX4uLNuQkP+/g1pWRH9MJG7skww4bQFq5FYhzFwqkgmHSxkQKqPY
0jKLNkB+4BV0vN1sbYQdeV95rDunlVpfAyzQolFDnlqQUrNHWyMEk1UpG4sQIgjrX3GMum8m3UVl
KXgEwBtv1I/4h4i/uD/CKfxlbTUidMfLPYD/gbEDweEvwaTJZ8CNvNrLvyGTwIyn8q1sSFYnep91
FFrsb0FZLiz5mygKr/+SZP2QJWN4fhJS9VvMTI6R9zVzpKG7qg0GpSf1FbPsr0KR4HIVZMCTXqUu
3wO2yatiyhW0a7g1bOcGyQ28k1oO8M+1upbViyxmYV7nCf2RAaPUEXcPUWMt7VIQhztKzA9/VYOR
YKZKyZTMb/W5ZWv9dZUzfhLOfM2Ihheg47Tjk1ufFIiP1iMmranT/CxXqLIpCZ2jAxoSdR+a89pM
Z0EXVVTb8dUyN1jnwe1XAiCpCTFO+KC+SAFqE/smtgSqouN7OHw+GrYRdzeOgRD7Oh8LLo6boJJq
KLoAIU3Eu0aAFBCqCC8+HCQQDd5GLhGNKYxKAiF11M7tICPpmhR4w0LN/RjWGrx+oqjXNyOqdZoC
ObBgz4Q7Pz51aWAPsRUtIb1Q1l0TtzQrFBEyFK1RJpIMz45Vlj4uFe3EAGo5ZDoaeTzD3KvSAs6a
u7epz+v8Q/U/PbudZ5+3k/iG7KG4mLMMzBWAAnLdx7ZC93m2t0w4nYa3d8NLQCB8kxz2GOZp/iRq
VKwLRsjh9j4ceNr0SY1j+GNES/FLAB+HIaCtiJACDminGKp05iobGhZkNNR3V8u4i1AYh+8zGlQ+
WMNNwYseS13zYBd5O/DkwmSOcQHwDZNrhnuusFPrPizVtjqHNXRbgAQEj5mP8l4y2pHoVYx+NfOW
KC1K6SmgtSMi8yRbm3I9TdnW9waluYcYcFB5iQg7aDqpYvudHaWlw7kzmfiAInm30Mrr6X84eN2p
7CRXAu5/lpQSOgGtW6Ww7/3xNaJjz5vGM0e9UcSag1ynpRV+hmRGWWAU1EsHrvb0tbaJhn8Kjq4g
u6TmMfnB5/qqpOpp2asv6NBC9cOJ6bJM/ZnYGc1Me4QgboPtpcl6a8MMbo1Sj3Fo2uxIjNXWj6bD
R9y2+61XTNxRrmtfFxp4RetDUAyzmCRLM+2aDfMlnbD0+YwV1ys+lb1tbIXMrD5BajOsqeZ96gtA
jujtl9v+XF7j5ou8UxCbNPDRIKp15Oi8b4+Pw3E0xe810zwinqhYJwI2KnAWkhvB47Q75S5ZND0v
L5WYuO2VUTZ2081VH2zHI+oM/rOHU9/jNJPFYYIAivYNhoPV02JnDj56tYhA0UMvUvzuuaW7v7DJ
BqnIsCc+JUsMN7zAM8QZsJ3C97rG/rdAkOTt3CT+uYU0Edkyh7FpIOVHxOV+zfEToyp/bixRbeu/
BlILusAgU4xMuFlfxmH06M0RwteV9h2sY0gejiEAKxPuwS+IQhKwHyGCN17x1UVp5upI0fCus+ge
wilDjehI3AE30yBK/GJwBuVnq2NBzoYik10HMV4XwkSsToqJlTt5AaXgDt0MH2Fn1pug2TTyNqxB
EE29zD1+rLvMtOr7Pm515am+fSg85dYqN9/ud1A4S/sbofpTyZS1trJWBZWJFfTUwhULE1BTKCfl
uv7jTr08Fub6aotKb4ixgMdEoQ5w49502nXa/YPntivuWJASut5/2tVBh0GM9ssDDGS+U5jGeLM6
mjqcPKP3ZSCuXuSXD4ALcTjOAB04ZS8H9IOq8uxRVNbhGFie285P3Cs7WTYR763U5p6Vk6uFbm4C
YbvZS7gazYu65ylsakB/tEZg/Bb12qaYSnIOh8dPyVLjBxfZEfMM7rNP/MgJNHqoQ+5wcwtpSM4j
BOaqeiTA86u+FLOeFJK692VS8+pLH489CNIBRiEQ6Px94I7Vjr2oPRv09nVXETulLqERVgf1dUEm
AvhUusU2BkE3tflcTPsCH2ZYlKR2fUSwlCxUIkNiTT0s0Ux1QfRb77mlRT8n3Wu3knBwM59mpTRy
mW4s6HnXgMi79hsFJIEBQ8ICXMDVKFmzQ4vRCcAjG63k6cIBt95Cga3++WNba67ZH6iXDu++PVJP
XaAAt5vCKSMaNwmvqQ6sihdc+91E80CW5C+3Wwj26yV7aADIiY8ILBYYhtJRus/UVlSVo+NH27ZB
VgrqufxOaimLe+jxRJ5R1ApLJksW0DqOz2/HJUE6A6//xau5NEgKMPR56GwnNkrN4x3RcXpBZJ+H
Qimeu3qNpg8vFNKL5vR3dFXIMFvyF0KhBdcqSvbuUIJJqCbJcYG+KbqTCKLjclyKcVxjppv3g1gd
gM7ug5KhvJVsgD368DfBmo0emPQ9EsqAEp0X0euEfORzzRNlRY0tzuiqbg0WteZX26NHnmVqYxI7
aWlKWdZLrHtfLslWxbVAwae/t5K32BMjKx5mEp8QlYLIUTGOuv/GItL94uqeshIjJYJE5CjvDIWa
XgrsvB1H0RpimxHy3/RSMVZ2js9hUa9/ri5XAEG8+yjEOpd7LE5RF2B181HSWsBqcAmsUo+QDBp+
xq9EB0rIhBVhWWYd+HtPLx6kMEnoWR0kMdGCYZq+PVbdoj0OTckN5YhnjUfbKFDfhtUy43yiBH+/
LWTwNpWU0qvQGma/wwJRGaEOGfbWMmKRuVfMdYbLL8qcilH4BUML0XV3Z+dnhX2OkLYJau9qFOw9
3ubbnWmlhCyM31jOxugyd1qr7QgEQqiniRyhQzK+bg/M8sD7Yly5lcOYtRPFA5Butfi5kz1DAp/y
ct+bcuv5Txqi4CKhoN8cjQAXlPNWp1alvvpaUNIm0KjUiFcdvpjfqGgUrUm4bgsfsWtc9iCcy8i4
jFLHNN5zeufo2H7/TIQj6a36RGd4/1t5vC2HfD+dSERcFxbVVmBJ6c+JDd8bYJrG4cdNp8SoyLls
gPQWPVrP7oKOk/CsgkZhbZsAH83egp6kEmrtCDjRa26xzcMBN6ofzO9jtiPuO2BEpeTYjyNwTmcv
yUcZ5ihSrXR6gOWROooTIj1SsQajZiyt16LaYdgRvjkZWX1rGJYcolb2Fv/jTAYJbIWnkAcT1Mq0
lzIQIdxGmnXH6jEdhQ3leelrAdk7YAkphDBHulD043BIq1hVf9RXrcaSIzLoJbwfjM2WLDOZkS4p
6ZLudTiuyRP2sczdfDGsyWJeCBqZoowG1gUYvMAkCrJp8uaRhG+4dmQL5OmrCHrWmpIeY3ndXBcD
yFC5JY88+Wkp1VWRCncn7cEtXcxE7jz/oAUCL/scfD9N/WdTciN5yc8McG2IygzcClvye8FRe74o
QXpZfuXtEa60EflJo7wNoj+6LPO3dHO2ougwrFR9v6sPRVNRQSSnryn/5pK1b09YNRLjZKPGNRYU
gVl2gXv1dyP4DlolVAbuVW/vNCPWQXF5Zxo36q/yEIW+BWn8SfD7N56yYkOxJDOVSIhjUpa4Shsh
jtSol2c/fUO+Eroi4VglinPppOX6X100XTDnbqQlyUpSZeSAh7Pk3CzpsraX3fJPhXLLPj6UFbgu
9r7YlepeHKYU/z9eNtqaGjQMOkmyQhLxhqzkIGTDRHyAGhgFWFt3acxXYh1a+TRUPpnY/VGDBSA7
gQ9EZs/Ls+EFeVIIFuilXaoHVA/Yzzp3bei98pGBHWJi4VV54Vx3ZErQ3TOgMuEHhnjggGFtKyCr
LXzrwCtQlgFPly3eBIlpVEPaE2U6go1YHTjp11zCeJVhp34DaRsdDB0CytGMZ3pXU82V8eiAzbnh
pBLpswNDnIrhnSqj3fHAR59+uYQ7lE59DtqElZH15LkKBr8LqzW6ucg0N95QJRKQRJ54Ni4BdsQa
vr8yxsfMcyE7ajKgupcF71yop4e9v//RT++oPTS0p0Fkk+6rbaQwyhRN0zkOtyJ+5OgdT4NHLX2X
llb+d8f0o5HIn8wgZehq6KEaJF7ZhiqA3oPdhoHE4OFyuSTAD+kyKbGRghnPNIW0pYEpNUlmR8NW
nRV2TRTLL/yzWGZAPqLm+wWzyzCvN0EdsjGBiyaT2HNAYl+0VyW+AeOcU5H0kHoy7jvh/mMRfRLR
qWvoOf2GHjHnwLEhZsOZuT8IYks55e+74MMur5VvuaYapwHzMagOIDzEgdr7+NVBbHkA6YnAuHRg
0m4nNZni0l+RK8Nz1dE/PcfNTFNXJHPaN7F3/lP4Wt1cM3tSHQbfyxjJgFmI1LNQo4Zkjep1ol6a
FpulaF5NiQIcx4NOxrDbbg19+4h+xB49ddRRDCRF0dBzq2UFp3Wyz0+9TKTsd5cxwiF6RZNGGAG8
XPCLGv4a3uHc77fX4PUodOfGGLcBjLHQITJiyWKHZ+ztjyZc9D/COuV+iizzHgIwBn7iCjcsKbBu
G+V4AOuaxWtvgW10XhQpJEFaQTsF0nZqBstPfYJOSW595mXVaexywTqw/xNbTryJ/9WE/I9uKq1U
mDaNNS0pTla3/cP1Itp7ACgS+MiiAnFiNstyN9NoqR37LZXBz2aSNuvQeW8u4C4JTDvHb3ZPQAO5
gQJ8y9D+1huHr2GmMVf0Ttk+leXfWWWAave3NGHF8yLXsfpAoPnp7SUpxwtDcnBdYnZF1z6ATer+
FJ4dL7tp5wansMF7sqgu0ey91CH8AR38LqpzzqFvamSRg7zZ/v4Yhu3v2cjh5TJCm3b0+00kRH+d
ZFRAgln2zUUZ/Qrj7uA9V3Rfes7bNJJla9SSegCaVLWLyPtNL52eCWa0nGEaU344FRZBQ2LWYfc8
TLtYcSv3bxs+QS+dp/xelHZjuPnZFcgeFRzqJrM1pyEvauZYSwDrDLT4Ks8+n9AxwU0Jk+plVZF2
w1/ilpAmc+k2nbgbLOwcQxo2ZfXTU8f3f6t0reILMMN1hw3RSYFJYdCqGV/4gDJofvEURzPWEbvE
L9lArkG7/16K+LtAVlTq2dE3Wr0m0fgcw0Rkmaw9hYky7tPVrFs5SzoUW7yH5obTu3c2VRxVgelG
6fhD8SybIPyzbjh6QRDpf88EcSuQ/Gi6UrF0yeG6scMuVAWdTVbX4cNn3qbsAwaj+V0hN1Og9FVD
6BlzcgqFs2LNVXvIoViSqwodQU6u5lY97ASAocwrnsoGu02kZ/EvIRTYNdLHu/j65bKH4vtW86BF
4uDSREs3/DvXB9NczuygupQ+PJNdhZeIyW+v0HLvjF9nx4YKCQXxFDBtf5vgw5ku3bsUPdLvM9qD
yGdrV9kbvfLpz/7fDBkllMbM9jReFjKNpsRdKh5NJJA3MBqy+koOtfJRmCkVxe3RES/i7+g3c2Cu
y1p7Ch9oVnb66Vv/Ny64OTosFss9qdAqhEXTseie00ZHBrnC6ClKJ3m5rn0sMpt4Jt2P6WLMHMY6
aDqWciNHGXcpYTdXJCzeSoyYkCXOd/UBpnxBtKX2L05Fqn2SlKhHaxK5C/9foGBsi7LLXvStTEV5
2Tx9quT82a3oH4SmWyt8HCMJgeQ7gY6d1cD/8oxhgxnF30QYErG85hWCEub53tcuhMm7K9uScYNC
NEAA0RfN83Y76uP781CriFga48gV9vDJKiWkyDIqu1zoBzdFkmADRGvqElNXmjYA5SjULSh26HC+
FUsQz4fvE07E5iCtM34TNH1Zb7QCJsEgy0Zmo0tReB3x5HGEGKl0p8614ga6hWJeV1rj5HD23XL/
SlYFu2VzqkK0zBJfO2dWaQm2ZpNJXadPxmXzXRktCtrMtiFp2No4gJfWXQCLgO8CkCmp6hF/eQfw
4jy44Au/dbG09qAekB2aImNwGd4JdgT3OLt/t357GPkXgdsB2Y5eDNsEC3Htfz/l71dykyVfXTx2
tUHrjFNLZgT7kqOrSw/TBTXfvg7gZHuaDLk6P3Py0WmiE8DKKH2srhWbSMivHBqg1k1z9QYeYnQc
ETNaHS2dOTD3t5l1yDTXh1CqrPDkSeQTfv7d1b3r4r4GhmCgouSf35CbJa4+tpLMO/ujuirrAJZt
KX10sT2t7aN8jtj/1AdaGPed9KqvA3JKJvLt7JP6QvT3k8/IwLdRTY2mNsn0ldaMJDwGCYYWqSXK
gXmmIUjKIo44fNizvgPmpUyVIgwAbWzvAUWeCaEdkf8rkuIq74sz8ASAGdmwwIVLditkVKb/IP97
roQXQmdZ6uGwsaTCNHMdaIoCW/PEzHTfi9sOawPNniqW4M6JwaEH65H26HWyl3exQnZc1dl5N458
Ua4oD325+sWWcgzAJ3OjP3Q6xExnpeQ0ea90l8epo4O20SjJcw1QTz51M1MbWvcCkHTk6M+NmIJT
7GAEjlH5d0GB6i+5owlnpZFRJtF+6bw89Cp+lwMDNpnnw9hijsJtaxr3gxbvIuUOc2FdtVhILkjI
eLwvEoximxj6phndKDzpbiadKLj+3qVTlgWfqNCM+2ED/S91vsHs+4StF97WHQ8Le23MLmG3tqjP
IMQv+Gmr0/nU8omnZ6JPTBbdvRJ1tgFA/1lNi4959lqUtpEn9xTNXuh96SFJqfGELHTzo+W3AaWm
J6RTUCZvGttH7Ib001sHwwyJnleqJKbNV97DvgI7orQSbbYb27SeSFRRY0uCRcKl4dhFaVAcj4hE
NfSf5LuXm6Yxx075ABo5O++G+UbOOkquq+RDYpSXYLZeajQkL6EWLd+khx/DbA2vKJpuhckOidi0
e7KeIiR/VnNhf4LhePzCDX8V3wMSXiMVquYTJb34XSKA+278lr6vD5WPW5hLdKLMHufbSNuVqvVS
qiDyRE7FHqZfyVx545bvPGGek+2+lb/Yq5Tij20AQinIzt/mCKEXkb9yWHTAhX+qE9mxgPtBOF0n
Y1yvB2UfaNNFZwvXNZNpKvoUt79rzxGu7rZI+75JUUVvV7Or/E/vlxt804ipdQLWl62+qymM8+IE
1YGDx7DB3eQqixF++WjutR29Hvzfj4Nej5o45Ztv3IHk4qv55TU1vyAvU7d42BI2kP9UIEhp7hvk
qg3W1TWfLtf0tiuJrvooZHD6lrfgpuzCJmiMQHRu8GSm1PTiZDFWaEu5zvHwh9CBvceZ8vXmYj72
PjYD8KZyes+fvVstFJgFfYpMdBoiK6jV2GzCjtSl0tt2D/PLZ3U1SgHVJgJYtGZImMfCwQ8TKNNr
rYUvK/qQSKrzQo5m+0/Uu5VLi/yFMnvZ+WapxE/0I3NNR6XcHi1XFQSUacBY1fq9wuQdBJAQHuZF
vSI4pwVwpSMrCXov05eh6fRQ5S2Lsdc/Qka7WFcJyMVRr3JHeCoJ/iJ9mBTjrQZKjpLuvy/xz2HM
6mO1fyvfuhco2u/CzRf4jOofCSK1eE0MWcD1A1hvZPngj638Ziec3VJLLDgBXtL35OnOpmh7FsVx
twk99z6XfOwtBc7ddh9uTt8a3ogkQ/24OMUoMyzOu0eV/lgaPO3MwL5bbYCVbpl1U4VXCIvf/0JQ
C/v3trlO+hJzKfG1mUiNKhaoVR8GtcqDo947WNtY64090IHevjjCpvg37YumN1BFOHhlUE3Z8eYe
wOk5AEO9b76rnUj+5G/mQhahR6IzuGL4FCvXLKkFNA10TcRUsFsZg7RceDDw7FehbvFf0f/U0tZc
oLLuTZdLYzJakPUCMEFgE44OI4Qj7pEzc5dqSm21O4XRG9l8OWD0vTjWwljA3NifT9fBS8WFHl10
2uMwEOxwCLwJ5CQxnBKPDCBp43d0elFEqXUPxf1yjGZzNkhLrTqqattGFsRCNkK0sYpaDEu6nXRW
kjXbnI5kBqQQpiwvQy1x+YXAAYvAb0MoZzbW3i4WFNF/6fAfbPxGTP7DDhsPlCOoY8U5U164BMKC
OyWsqJfwtP0li4y9m3QjiFnQAQPesZKL1VKyjuCTgq8qP9rVUonIjaCYe/4nQ9abLl7Rh7pBF2Kt
pqHIhKQKoJS/aO3405LvVzrY/9QFeva0LNf9XMvOMzYZNNmB0mXMnjCN609o9Qqfuz1vLuD6YMwr
oa8PPeSphlu8Ng4nmy/JXsT4SVq9v1cmz4hmCh024s5SUkX4+JEdgVqVlfoeA7wXICMPAGY33H8q
aytDfJCe28v5+gEuNfdBorKZvSESZN2Bm0SB8zy8WDxs90FV3Ljh9QTeMC4OiIwAvEyuHjUl2i1V
99eRwbhOjku2gBMEFrd5jVTkIeZTfNcgVNSYdQKlRhV/qVGDRxBVDJzxOCZmUByEt+Qmhm2AylW5
RvJ2OwhxHYAbI+VISARiD/xKhTcNH8kReRuU/hEqZfkilk5VWcf1UZSrrzRc0+BD1nux4kzNxV8X
soridwtT0ZQcNZVri8fF+qJDlxd9fyfDyvD6pQ9xIGs/V3Y3iuHEC66aZG0m9XrGNdDkpV5VGsQU
8+D7yufYk1QIPUqAOwN3pand9chXbqAIoZlJ0rECOPDsrXwzeUrtpEvQSxYQw3oVdatCwxuB4iVt
/yn2s5lnzkBUe/pJ4LV1U4wqXDYfQxH4a/AnmiETmL/EZqRPcyC5iRrgMf52QVW5rrMDp3Aki1Mn
5TFoOVoL1b3By76rPiDcDhXPS2mzy31e346g3KypMDxur/MMqzqj0CrGPNnKZI+p8YW89HT/5r1Z
M6zvXodJeikcFBjt3mogxCaIStZHNNFNsns4P6J/6bJQKetxkQvOfi6CnHrKOVKkZH+imAE7ptEt
1TYaqXD8FkjrdaDYke9Kas70zpW1EchNC+GKi9luNBC/cDjq/gmfYm2LXRPo/EZCxO2BerrR7s1Y
rTZNSrq4XIkVI+7Ox0i5YYPHHYdrgL65ydo7IQwCGsPiyTRisjnFfSF2/JubqpYVA+4KwhXP2HpK
CtPLEizMhaL0Qt5rQveLQpfDwNc8oy3eVqpHAG6gbDc51vpk6z5QAzA9mNaxRF+p12B7ppOFvTFD
EJ/PGL0x0MAUvyuFb23r/Mok50QNWggEAkzqZlLlwKUvS5df9NQrrW1N2Q536ETyrZM9egMxM455
M4ixtIp0NgZKwS+5uaq9HNqJpepIXvXsHyHrqaBKvxrqsIbToqQCU69tZxVs6T1jNWaaXNZ0zrUS
vskyDKkVj8RFyT2mvtX3Whlw8fZ85RGDXETB8ZQoIjpk1ff5GBG3bWZVGwYsOJvLj4qrr0dK5/+n
+NQuoOJh33C8xPceKLbhnGf6VJgBBdLJ0RTwhBrrhxTFH3g4GOgwbmrCIqN90t8/rTes5OSqzIjJ
TzAB8habJVfc/mV8MvJh1uj8d57VbCwztDIHA0+MvNHjhsuXpauScI2X0Bk3zP/MbLjZ94G8MUTU
6tH3D0Pb48g/dv1TnAnRFHFLlMjGTz5q2bbORZCPI/18Z9ZQHvJGUxIx8tLezSpfWmwnps1D7LWo
4pmLP9Y0q9T6A450bSnfIsylNObTm9PvSs9BSqFqMNEbmcZ12AAV07XldcANpqfeQHr8hFHH3Y+z
fT71JVnCVNlR5rBpOg9r1bW8V0ft0PBEmFPN6cXMXAKQBOcGallMMcTdt0MtddmvjjlWUV6RCFl/
t3Ss8SrAiAZtfHJWZPogGCyn3vYaPVMl7XWQUQwuxhHsRmxBr13WqOgDQcrtrs9e3NlfWdiTFpXL
nebrUbB5s3Uki4y04mVtHXxu4KJYLPtImUpABZlUiB2a68hqEYo4Uj7mtMwGg6+ojcfdq4EGls6f
6Ym2yZdedhEb+dSfVTg6qpOemk18Qixxn3p4MW8QTEvFgbVgkTYkXJRjIQGscwcDQQylnalUZwzt
Ixx/Gww69MWlQwEyX4m76R3BndWimYlPYFByQTXhg1XMxP9e060scvNgmSiUHJGgfwbwtKfZGNMx
COe+Vl267cvlmHm0+Fu+tWk7p+GpWcKGHLDbFCw/D5JtIDP7EwVI7ci/rDBfC+yA9xncAWaf8kSy
9REFT9CPFm4wi+FTyPKR9perEPH7covSowbtEYShiS+v3exgQeQ5SmY8pFCMEwR71nb5wzDzLqtO
rYweDjE7Buc5onPVVGQilKnFnBPUcZDvHNzxGBSK8NkzDw5GEBlkpH5DhcOJM2k+Z4zYWCqQlDgj
PHFS/KT/PRqY9qJ3bbsG+TOWzlMxCDfV1FsGkQN5hyPeHJcfvP0cIUfU/QopgvMDK/rZYDy7OpNV
kyTUo/0xsEJIDsD1m3YxGMydjAYzQ602uOFGClDL+e/vQAEXY/txyzazp0MSQzjjcJ//NX6TTrxx
KU7aqI83okBxdBNapmND/yfO7D1umlawHduH0zoLjSOnxKlF6TFqwjirn2vjNTMvZggJgxndHFUM
tHmqQv6EwnC4pINg4FVCPAOhijcMy/kR3qxR4sfaOl0SiGE4skAdurz8yOnflwbi0q5tWYW9GDO7
69O6DgFM07Y1IJJ+HexGKTeaGqSR6UNi8G4r4nNcSgcT+QkmRLXLrCN1eos23HP+unqU5TW4g7FG
e4m5wfaR5Nir050ZxMaY4aJJ9nVuku/Xjo4ViweIxHYDw8lAu3StLROVaThcCxWyIssrX6iQdAQ/
fUKxctCU1PCaDKTLjlBV4VMGylxGwN2aqsLehahoAK7zjAsU6OBrQItNL1FQZFg74xNKz8mkGZ2H
kIEqKkmk6FTCzm7JQMERcu3C5JonIpBFp+NCWswKN68Y0zsn/JzcTwrRmLf0jKdmZVg0R0wGP5oa
o5a36pfONP6wzez/jT+dQvg5dfs0y72EVPblyeuj+WWJqmof/TcDdys8bYs3KRVimugIJeGAUhQW
fJb7LacyIf/fd+aU2XeJo6sFzT8Qt4kEOcwHyh0j70Lq6LcJIX6CYTWeYppOFv0f+RCawOiBd+tF
RhJbnlmnQ0bwQPePCF+HzQOPsReB4yEaHMh+7uJ6Mbt20UCXJdUz7GZn0hiE4PP4iUv4VSooKgm/
VOUTCs8VRt0FK+BWxiIKmfvnxOCCGbmCnxAdKVd7h7S583MWQ6NEZZzcweBwPKwm7nRfV1jB4QR9
3HVqN+gPLqEieHPO6IFpk+gVEiZZheTpahEba+76aaPSeH5+14noyUlcEIoqlzyLWlkOr+phGBP3
incR9qKrpMHNN2MqZZrHC6wRRA2jUSrACAYJmS+MQb4BBWAoABpwCqdRAAIKjrxgYB1INyUBi9dG
aO5R6sqmUaOpOnta8drnsaIt6cy5qDKRTmHA2EiBgCRj/k8cRksZuJD9kTTThUDe6inH0qNIbnyD
lBIr2MjqB1t7c1sJwDg8OSKOsO911cKsRgw91boiPIpRASTewvGwXaJLy466zGp0Ys63TE8QRZFL
La9Zuaz3/GWoMYYnV8s3tttJP1HsoPZLJ1N6EytHqI/1/gW6w+diNwO6fpQ15aA+MZGAT/IoCHKG
UNYG/qhgCHRnfMwUer/SBJVD4BcDFdEo2IZxagqzk/l7JwyN20a4NhBcdP2oEkRNv+/bsmYHtzc1
Pa2q2LYsJDQMq2EgUPIRIFpfAufhdXfD6P6aiU1Gi0ATNnFhIX4Rz0TLTb/HZg1p1vmFG3pKqXoK
SCOe4fDi7FQkZ51qzBSP0Z68I+1kd56oIqdVHztvbI1WX29o+ab9/XNH+68ri2Y+9hekJz4xovgd
hk+HYp9ypvvTE6i8U+DhGWRm+sty5a6UXIymkirZxBqHdWqhiydJPPUvBfpi38a3TWRnn1CkbwA/
6xTQMlYbIXFODSQtx6i/d6+CjLtfJ5fFnwGs/wC9YJ+xt6/It9I8cKdAsG9Wvi1GOsnem10JUoJI
LZbBJ1lrHEe/vPqMRR3/n46+xau534zyIzU7yI+pAR2cHU7sqsVCyPmGSiFxZsqofzcznow8eiA/
VEDnouISGZ5TIupp07CsI5q13q0klVQhnwx6xWY/CfR3Fc4+6/a7c1U0bON5yuajWYCgVK6OiOFi
lHNBZc3ZzfXWXHwg/yW7wEFhOS47ttVh3JsL4V1x26fQaMe7A56fW5AyZeJFGJfQ3+N+sh/h0nkj
0hEO2dwPTjvTR2PZLhcxp0YvrmIlgn3rh6lZkM1AKXmGzQboo2GLM4PvpoEFFJnz7c5h+e6Wb+LV
DaA5Wo+0VQlwPO1a34RF0cjQrazP4T7312pL33wLB6vcTILEtR9GuXsanoP+IunOf68xhEsHOTjL
Ar7uqHJc/mNAK3XaVtkvtYlx5vbECjNdP5+8hauLRy/VX7CVx2MABje2wsw5egdYNi2oDR5Q3D9/
U9K1e9fY5mmYX/Dge9sI5r2XQetU//fqWRTuGLBOWKMAYiejrcy6YLoEuH8XZiE7uGWdQfxmPZCr
fRwN27KQgSGSzCh1EtHTV4m8szjDgxlrf+lkAOvCjMMRHmZ2+eJ99j+O+xYTHJSR54ctwP7Es0Yi
6tQUPGrXhg5FF2kErFi0XwtT+1gI2L1SgbUZxidHPClKBuv5xLcZVK1P0Bia8yTtI8WCyCNckwbU
/eEdjJk8NTPBYGzZTE5ysXbvWYlRM2G+5G/DbBzTtaIaN+MXwoQ596IvUKiucCeMSONw10OmxWBN
0xvP4C5dZ2wq0H4mxM+s+5YWY/v0tAJ4r3TB7eiq6OkGlbVNDoM8/BKJUOFDcezvVDh7chI2V579
Cxkc8ZyotBqRSatnfbggceuAW1/p03CaIoFBSfTrEHOiWq+5sb3raZPIFqDDOtuGOahRBAHRmuHc
ysgrv/256uzLsDl6DdpHS6D3o0JFR5b62hmEvgb9VPJBzz3QWB268cXcaEcusUofxiQDrOpJNtFt
hWuC9sWEJiuIrFjByKpzzTxr7Nf9ndFSveqnsn0LajSQakqSLcwrC5P5VbrROvRSyy9rYMULBoto
pssqz2JBZl7xqSJTfv4Gu6BT/nDaMORE3i7swkml7l+3qIWlI2SMyIXq2fgwXSY/lJDU20iLL556
Ssr5zAUwCnrGpXyahUaraUcmxum6MGDOwaGxhMLdoG9iwbOlXDY6wKtNUwsRldt9Nl2f+YLpOUea
t8f1sExvGLjFj7PMae0syuXWRlZs7MR6BwkPtB7Tp8mKSYgxtWcwtUcJ/gpNJBk8AljoIDrGqNjP
75whPhMTHIh/23VJ680XhPLPiodqjI10DtAIOpbn1JP04uwa/eV0A4wQ+Bo9sRXXPRZstQl4WaRo
v19tlHsaneR5z35pnWhlMjM37GoRCSHmvThMn8YpRZWRuuTNeCE+FBKc4AN0mjHXmNj6x+JSo/od
VtgTzmqK4NsCxAPt9hpvWwdgy48eaWrAs3+KyZWGBX82VqHddglPgKEsck41PrEFRNF/kOxY96hB
KcxutGOl2/ixbTxiPq8KcgTZmzUHUfjiH9sxak6mcFmqMb2ku3RXy7R/RLt+gvHEsxmdZBzpCR4l
vHBI+0maHJGBzavJtF/c5KxrlHHr2YZQys3jNspGyN7MASjOaE1Zx8ub8Nw226iU/AxU/DM2BI+N
/MmC2LU04NbtK+eV7vzkG8OsYyylSx3/BdrjcTQvFwqpK+g7LsFfMBUQrK55YOTbq8wfcaAWZ4ZX
kMmxVJCvM14CmdS5SJSPV0edi9GFPbcnyGFCrWSU1apD+r+SrDnlJFpFjSFsmQD5ZKVmBGKOnBDq
aftnDrENH6LzPx4Tmv37AmuaMOGYLS7ymPa+96cQRC2DDVz71UawQr/U5TAOePG0oon1WwVz+42J
D3RLA6F4qFhfDhPvUnNp/SRqP4czPpDFc0siSjGsMadz3DFOcjDXtsNFkjSDVh1CXPwCmZd9V90H
6UGtSKolLdY4hHZWuWJRjrtXmrEbwMHD3vnq7Bz0aohETVMbkNeaBna/k+wtAfI/vhDRO9s2Eo4Q
wKWLYlHeM/EKIq9njqD0kZsKFfSZiSN6gZYQrNEXx8uOwE+56fxjGuaucPicwvRCTFdhxRqKnMoq
sD3eeJbteyOm7Iu8GbXO3H8mOwQQ/glOqTJBZv2GFQ25HkUehzz3Oznj85QM1k69nbNnJ5sAm1jH
sjGdlkLm7i9Q+g6i0FEqriU8YjopCiWXgGYlv7AlO51vfc9OIzXbpf9ipxs4kQBYlDrpYVs8gZtT
Ok2dkxy9QkWJcWON7g8t+BMLChtvsEalTlctNLcL0lFDFmTPtaM2DsMBIFEoEm5+dQaAa5g/o+EC
uf38tLqWawhVYg2nrOsJ+kJexSOuCkSuThv4UxFfvtL1H1i1F1urt8AlfeHob5R99X+YPbvftT8u
r6wk0c8qN1X6RTefjTMQMS60QSxOE5aNMRS0D25dIubpFIZ+/SBaYLAnvySAQv1zH1Admj6WIazg
T1gwvdzSyM8Aw5ba5u9WTehl3ZawmljgqfifbM3aGSdfI7MRUEkjmw3eljSHWPpLga9CpV30uh1l
G2ghUlkYoAHBaSbnR6eMJlmIwXQEUdmrnpBiSIDjkTn0YuSRbDnLTh00P5Vw1P4UcawxEJEd7Yet
jIluIFXQPGKE2N2jSU4JEbC/sk1DW/Df46Xg8bFdiKmtSqs1QmSeQulg5TAaNkH69OJaNB5zNd7X
hPRrwvv7SyLrNKshvcpJj4Ik6V0SXFe2xhlTj1TrR0puUPFIF2OLRad68ve0afO/v/i/dRkeAopw
1y8xVKDRyWIAuTKlm9YocMPvOioWSEUGfhN5dlisDzjIptT19avKo/ma5n66+/bFTZJC3t7XHjBF
sU8V4wLG9NBI0/Bn38EW/IHjCNr2adMFH7GydC4Y8MWdYSLqDL2nnn9TA+TC+HKtSV+IU3wzfs63
0UzAywXp0RcDu29BY93K8j652k2eJR997sZhEB/bKhWfgtPNHmfheABrAL79ASs8pOtF5nukozxX
kAdVWBUBboKSMGjpnqKpoZXSD+/SNfOQdOPgWjnGTUEgd/w3LjsYyUQC7GYVXRMLGzLZTkLH7WHa
T0w9UFhUuJwJEfU595K1Id/RzG8G3jf1uxosEXfa8/RK3dW1Ejz/dY0VWxrCxY6L64jlF3vQU5QM
w0WvsPt+BUFsiwELN+QWWKbHqKodgpVQMeYGwkp7xZ4E6dimI/0gJugAY6wCAyROM+9+jofnZ07W
ClWkMJ1hX8A6iyAfVLVmMXRLves1iX+B1vQzUb164I/Ow9VcWorTSregiHyS/GjHVgyUr8Qob9a/
TLNGx0NLC9lDPR+0l21tTb21axBuq5YbEtHronRu2GsNcUPAOypt69AyhwHMODrOeAZ/Jea5YCeI
3PL4fpY/b+yZ8s1C+6LNdEQheX7La6KId+IFBbOOjkzn8QUeDrvdVQIZz2jJ+R4AdX45B1Q9iQUN
tw268qVE7YoVCznDo9ZDuhB+iGtiCOlgGqKK0P+H7cWiVQwenuaIdlVjGGodAeozW9wk7exg+4rL
tTgs2t07n/ZPR4lY3KrnGpzkD2qGBxkJ/XfJ+7TjLPLOPRY8pzAxWZGMo/D/AtuQVe0izotjWXxU
Gd5XEAdzes302ViU/Qvr/vXJE6n0rbqpWRx/KnSs+W8kMoYHUcYJ/8AMIoHLDj3D6dycN7Lh6a6m
8OJmrDELGKYO1oVLdk1O61Pg2j7p/JXW+SYFLcOy0Pzr0h12+7lpIPkn2HZUWeyA8EsokWUn8eLY
MDiG3Ij7tkzDa3Kn2lysL8xieNU5KLAaegQzFqGDRdqIV04Re3Y4FTskVD8SFdJwcwIlu8ySgXUL
bJdLimmhE4qnG10NYm6mynEqYD/fCgHXm5KGccBkjYha9b8adx3Oaakse6/4AuPVjp/ylbZrdySY
pHneKy+NJ/XEUQglIUzIJlG49l+xlrqYa4u+oh62CJlgx43lOxKI2a7vzJwarr8BAAGAbKOfMpED
52gz8mK/wrG/1CICAmS3Lr/m915mJDd2sdFlupybwxy1D7ppYbj7K10PyCiX3TzcIUU17Xbhf08V
wrwZqCrP3QqsWqSSml/cmGYXWRYF165N0inlawUzpCGu0T+99KNVBj+Frm0nuqy+fbhiOriJn/vz
fW6zkqinB+kdt5Bj/IJQJbPYzcGLN0+DGagtGOfXKfpRRAE4Lt9Y9DKnzmT9cF1no973TQFzgdUK
ZTv4EUdsyMhIEn+6hNmr8bmVM0ir+w8kppnlHi6uspIdeLKQfQXJJ1GKcLVZ0jpe1uQqEbXLUASy
aXIszlKbFIx9baepU1p1q+OGnmzIHcVDmhCr2/jy+b9LCg/9qWuDr9DwQBd/tMx3HQNi5cSyEvBk
zs8kUpleWogY3mCK7F7fuGKxGbrsw4nSpDgzZO9SIOxnbyXv+GlJqV/yL1be/SsQ15wQWECHCV2O
bT8Z8GyJl/Az+UaC38gCklBgz0UYXaNNJmD/CpF8b3lypmS/PztnwduHp6Y28oLb4ULOPWxrkwYv
I3hhG9zDD/erc4gD1vVkABtsmY41gmApUhnnC82Z0uenkX+UTdqN7h87Ke0fNcKh0FYguRQQ46fO
6gone/c6MaUszvktmqYCl9x4FEEitbdJTs/n3cnOFly1oHiBZfd7Kr85yYKiruQ2QKCQyQrQvLu4
B5QFpzHqoIJTZHqcjecX3DUNyc+idk4TE5EfNO4bVcyAQ1HtUkOWE+irqvv2uBn/VUKhAUyv+ld7
GsieLXH0gJVIfPAFrppExPu1LYa5tAj4NpA40476dpHxJ12WpgWPrkr9MQkeSRrQ8jBLnBUGvqD5
rGfVZMeUYmyzlZ5se1m+85JgcYYxHS0YQJpJacE17a+CL4MK65uhAaxkxdeAJfdx4S45IPjG8soC
nTBnyY3cyrxaK6ersgpNpIDW8NGcp5Yb1PWe+U4f0VPJOFlwJl3e+gqELD0al/2lCQManF2Ygd1i
tMgt2Wyxxko05yTd2NfBYdZiyDvioXWekS9Mw3j1HLdAxE4+W8O4L6zzt4leJV41m1FN+BdXt0/b
HdctX5cwGDm/b1wfKd2ILakm6jGuw58vIzts3XH/j1EH9JmQkv5Dztq7EXEY6IaYHcWbLob8BfG9
yXILnkL23mdwhJMYx3qD4+DdzEuvTJbtRQQh+NoSdFr2xz8L7300TuWxlPXUu2urxvnVHJWClDlV
MDZxpP7X2e7SYWCh+ma98p88g771MOgWJiLMHupwVhsRlC+lhW9uC+UcLi+53gx7h02zXg/l2YMg
Ck7fwQ6c7aPDL8c3UZnxDtF6QcHI0q42kRm8u2ixnfiADEjTUjCBnz4EuGjBwtCRPZvm12qYzv88
N1sAXAyBQFQLAw2cBFq0Dq6cscnnuP9ciFdhJONvtH3ZnvHuH6X2NlZRUKSW+Q3FSlgA4Bj76LiQ
hp+Z/7TD0ZsqJWBW4siIUo2yp1AkgaDECn4qB/n6tay60xeL5GqrDIMmwMRt9l9QssFXTMeN/iru
MGbbm7GF7wKf7BbB2EjnFvhAFPAkFEJtpZRoSfU4ex9ptG9vx2oiSwN1kAIoQS1s+Q8KObR9fzoY
LRnEFyKGHL4zlpmk+cCfZOk2Pz6rp//fgTyflp4eF8674wuep1kACnO+GGc7qfpXEUCG1nUyYlAM
+IVIM9hhsImLlGwlz9gSXrRR6vtJdgOh2r00K7gDoe1keYAyOUBXyM2SPD1R/4iixXQrQ5duijv9
nGvkjLidSTKMRSuIL6UioMZeUVNVfqkNCC4yvClpdui90PVnvZ4VEXVNlb4kZHzQR58NDx9K8lkt
fl6ck7GV+NMesz+d6mu3pj9uExo/RnbQkoZjGGoQGelTHUsZpxKE+SPI6Cj1QdBrsUjbYHZr2v8y
7ZoyIsrhOGCtRHTk32uCZOin8ztyw+Q+A1QdxiOtnH1gMtTtr23lLgtc+e+qmcuPW1Y5/tpF+USQ
EclCH0ULYmcnMsnUt83b41RMdANrYFrOl/1yDTn9lzcLCl/M2A7Ary8qnEeWXeVV4KIkXpDjXQvn
nDTPZLjHxcNm91nJDrmCpNfBgVsENK1OUBpOrw/q6dYaV0kSvAGReINs/8ZGMcM50enjdvo5bdbP
w5w2BwBCi12q0uEu7XJ5vQJ/DbDGAGHoqpOH/W2nCrf2WEw6CloqP4KDnv71F8pDwANOfSwlkqVc
2oGgaZhl7weNuVIIgDwIUVYJY9h/TlSsf3FJ8fUmp2l2wg8X50gQAEqJ1bnKHZP/v7Q4IQCjFCDz
VM8Ic1BmBoegbhWvTwlk4aUSi/dACTYoW9D9ObHjjv0UIWZhY947tW+xE2FlyuEPh8OYm2RVICsH
5U+PLsoKEchx23KiSp1wimPex8pM3BchjDHUQvseFTSV6Z6PvxoiLfMQCwifSL1+hDZTER0Du1TO
T48rLG3NCtvukPK377ry5fRpyWuvdQTRauCjHEyEjav6ECeWHHtOHVwpz3Qsd2ug65/OS/gLgG2j
v3nUIpDXVoiai637B2LMWH3xisURUk5XZtdtCekdD5nIetCPFHF+bUTLX2Bb7etmY1yZKJ2igFdh
E+2MARtxAP4CvHnznsLMQhs1Zy4NrtmHlNJQBjLAgmfQYjOqDSyv6nsFyQxloRzYOqIiOQp7hWpo
2kOZlUMOHvobUsQTuLubaJ14uvwmUUafWAG7Hfm6qVLZ2aWFiVkGNfZiosSvpHjz3Y0xdTtnZ/rI
pjSli+UHo7RjeBIqxVuBWXGKcWv0bEzSLdmHi9i46OTZgM8U8Dx69dShRli1BsZV7xwYqD+OaNcI
LFsTsxId950UFm3l4XFz4Z2sYtD6JHen0FkH2zE7rzhrdMtnCcsqePCpHDr4cxJ8qOGERANxUcYZ
r8DHEEvdBX27xmvbxgZlle1TRUMyTS8C0idZmlJmY2Jx4Qj7YYp0j1PIjGyCZZvPOg28dd+lUhJY
kplU/H6QxGmSxEOSOoGXWwK7Rh6D3x1ZrXtmI+lfINR7dF/9UU9Tl2+gtD+q3aEzjGaG38LY7wHH
PIb0X7FrfqB+dp2LWFXJVhBZ8E712K7M9ztynplRMV6YAJraCSja0gb8Y35QGOv6AlVyNDoM4UBr
Eg1w8sjulBMk+hY+9va21GMc4XBXKQMqyV4eyT9QJVTnsXYSQODi/0Cu/4c88zLMHfcn/r1nj4YL
9cM6HXOPedA9TGR2Wt9ROduFQHpio1vTnJo4vyuVt4jehAdP9HAMjtU01jY7uIRmCyxaKED8/6dV
wdE05CK0At4tgyPfKzlLUloyj5zS6DCbpH6ASGKeXIjmnH5rcPxsDGOFCg5LB0GBqP4p13sxaT6K
fdU9sOM/CfAwf6yW5wN/gD1qO7dEDDEwNlsqviiDuuOWqaGYLxIZBs4ilA2XQqL6tymmTJo5Q7QS
iomV4z7bOfQ9I9U+PaXKY21id4jlU9FLlcNvPIw7iU3bp8dkDb7saKn+LzqcR2WrXAoGHkIRjSII
2clmZzltJkSP8GSmCFkRWl3xVC0ro+9Oz+k3ReMc4QPrzGCM9bA4CysOXu7xqp7Cc3caqeSpFBev
HGhSQBrGw5q4jKF5lxgGe8oRQMscDJ6QdKyCYKuorJtWOCQu/H++Dpti+L5Y7Y4Z+1yDaz9HZkkY
UEm0uLfbCS/8A0HlljQvKjuBu8+mVrns3R+OI+aDA31AZLdCBvotJiaSqIB1TI0lyqfts9JETLBz
mq4gzoZS2+AndK8m8s66E7CxKnBSF0E3hiQqPs3GhwgskY6EL/fFya8kdTnOhUxtlWZMyuXo3Jmy
zWO/liPxQQODgW4VWAiShf4ZReS5UuMUep3R4Iu1vLsT9EqvpNaszzUKTVxlOb7CNgbzSBipUwBG
JqwgCXtZunSXVLDTGduSe9Vbal4wkmRvq2LP8VtI/zyDOTtPXe5ymvzT8T682+WiX/N6BjCtz46n
/ivXu9Y6SpS/yym4vX5L+F1NS6yhAw/Geyv9cTXmpLunFvIhuaxoe1kNCQbQCfejN0UAqTzqy+tO
aFzotoJeitfpRYPAYd2VpHQasQuzA7DJUQtw/S6bu1To0mswCQzkmmlpc2aXQfsUpmB5VxPBweF1
08vdgH22+4vUmiUmlUpKLhiz4E62MywE4//igg44LZec8qtUPMuHMRuKS5PxhfLVoOYu9l5ZVjsM
Z8b5iazk39Wj+6VS9WJ1WWNWqHXtadBdiBYwDRO0Q92YoSqTQsn9VH3y3QRTNrLLWr6WxljZQZzC
Ntih6+fSksgYTpTtUhTkOVbifHP2CGKqVkwehc2qDWNMTYJfE0Dv0xc2S3Bevl0epaPJTvbxxF0z
zbl5fnhkoFWtHAoOdUmweLoBNZ0587J4CEATYqPiBLTmsfc0ihlzxhZBIdKh4T1r8cjybgXUfWN2
9vZgnggqByF88iSxA4GTjCdbX9UqnM9WhF+m7b8KbwnYQYMooHDu7FLZB0zw5JfyPGY8Wqcg1bKx
s03H+Mm3j8fKkYFI9i4rIBwPumRZDU938YkkE8tC6xBntgt4GZ5KcRCymXnPxtv5JFr2cJRfBZ/6
C3FJFSJ7xgcO9SrqFx/FdsXnKBVgM3XQ0Yvn8BFk11rrZNFmRR/b9eqIvW05utFMJW0HlekOuKwb
EdqNT3EcyxRSCAFWE1wxoH55HeZLHDzJ5ZP6oElVAer8WGSsVPX3OiEVv5JiqRV8NOUOLaEAw88U
m5RNx1AKLY117c2n9vpfT/JlDSdDP3s1g+CRfjn1CgvZ81afIDnF2fQoBlwp3XLM4RAdy04mW54g
eIPmCut19zVFzYX5egIoiyyW3YCHIUXsQtzZ7y/b5uuPzpRtEELqW3KoG3uKH0XzZdwKO/5UkFPY
wXxkdCZIHWcufrYsUNjimYq9JDok/UzRX+mcpLd7ZBUvYEf0XPExSvk5E5CufmvpLGFw9xeYyXwo
4KxpBnGrOiqE1o4rBJzuAz3xfFckz6yr6kMzWeUrGVjaNLxy4wRXtTcb5TgXW/62LoysYWqulMqc
sVrirBmoQOYRcCZbSOTQtANaTRbWLnbRnLXAW9XroA6ZW7dkaD66yKomgkRNrEz4loWkdvLyFhq4
Fali1Gj/J2957mOG5bZyf13Ta32UCg1UwD4ILt8yTFvZrczW8GOvLgmL6dLkH0eNcfpJ/1YWLuTj
aOYiARRJYfhC4fCwOv7np2YiJKSuggZJqDXGmzlfVY8prmMIRTS5zctTUDoeLFYCj4IA+YwBNvar
3IuwKYlqOeCIEs3sHuZHiSSunIS8qbaVFboXvPF30Z4RcbMyWbRwoAO3h1Q1RcCKfLfgRC/Z+zyD
zP4j1tHHbvdjnnGlGIgAnDBvVrJMocWAnLYWSMl5bTdMJucyA837n/zIbo7qR5fCNXR8/GNKvLdD
8Ym7MJ950kPL6gq4SQwmGcm/dYTOGGK+ONOybcU3J1MrvM2m9W0aC/K1IjYry8XgZM1DJ4jlTo/z
VFjXNJs42eXsBbfG7FEEoWvNnzbhwf5VorQdQSiuzZqzM//ZxZ1Aa5TShzNKVBsgCNP/6sjb00XT
5Wt50tN9kLMd9T1nf7RSZRe4hjqv9gOcVfxc3iVlgWNsSoTrGlq4yk7Axuc/ppd2wZbGGMutuQzM
1ra/cvwbcldPSds/ucQOJ7PMtDhodhaoFO+henUJKCYRmWk00WrHwIPRrWAPc+U8V54sV1R90mhu
cWXX+AHE5Xx5h9c3GoeqA2MBj19P8AeZynsmhdpTM5nxt+oJRXI941lqat6wU4yNvtlGTFKbm5uP
ii4izacQch3F51YtReFvYFgaxyXUeaI1gCQ/ealR+8NUaizgl/GdqpCKtHFMAAEKtkF4ou9y9er6
Dz4FMJW6CceZqGWZBqfDP2UNud+rNoW4Q/uEUi3ceiHyr9KFbNJkgEI/RI2556PUg1DNOVstt9ex
PG1b58+LqzoZCywN/F3ELbGqj7r781BElove7wQQTOzDfbTOhApDxzXKRpw3UpAgX2lkhJktO9yR
Rm7viPQ+V0LZ+bqHFpZ5YoN7l4SPcuBNfDZx3AWaG+neI7f3MqZwmSnIP9zW1vT1GY2bFwwauDq1
yAb1GiDe54RngYUgBSzYwsZp+5GchA9l1oULBIKVw+eEsSHJVymfCVY6tctHJN/BQ357TU56DZps
0sRynNELyZcM/uyUo3Sxf69iAZ/+lyiSP3EOVE9kgiomRpGMkPxOGEOCZztjbUMrkqC4QfjcLWb9
1Kgp88pEuUieDveOSmLssNxmJFPJyWBoTP06Ia9FZ3EGs8RbXaxXbxj16kVh2mHaysqYzPK3rrNl
a+xved84i4uolgPPQPADAudELlbWEXVQHZlQGufVN1XVBwPDOPHCBmjNSpnpjJGO1fL77bv+CD21
kLl1DI3xM8UI/urcg2Leo1d54kZR0I9TvD9mRqqTfxan5g2p3gnwkdYwxedpHDc16aAXx21+eZS1
2czgrlZY+ImB2Tp/E1ngh4qZX6B2UNaAuAKzDJxyRp6Lsb9EVXBoFBZahISTXF7CJsPpWibu2sQa
HEcO1t2Fg1p7icYJEeOFBDu2Cw6Cl/gsTFHmtcUf0BwCcJ50EaBgfttasz2/3VjxK9R0asJ4xcnq
LttwyG1VtU5nopNV8ABM905u5/iPxnSQIujwjpQjNcduHLy8MVi9q1z9LhSPeDLKxYo41Yu3FGJ8
2rcdkbihIaEdEppnsYes4xLt4ML+zzl4HHxB1DB+ZrlnZ1ZNhcJhVDHZVBFOvqx0whxko82zAfp0
HGsWuwBjT3wEFDdPCphCnMPVNt51KFq2sB0+fw980eP4yE6C34MIirjo+2uVj2NHjgGdFMXlQpLv
k+CraWXnUoeQYZ66nR5RN3jHiQ7iuEFRw3BjU3YD0MEeghOaGa0P6PX3yAm7p9uD1IUmODkFBXFL
1bX+AcfQDtuYngvyBVGE4kF/e0+4hj79p89S8acATMg2EOY4cH1jsroadZZfpRzYZv9/UrocVj8+
QRpg6ITKjbjkmD+erB/fKPlG8HaGYdf4tVsLC3ufSasLhX5nEWHNI9ZxSTtLBW46vGQLaDkAMIDY
d/VSYpYfPu60OCh4z/v42D/DP3kON3DDME12DVweGRK7L2sfc2dAohGpTUs72AzyqiKjssmzgQlb
BXHBA46kudpkd61WJudj4mvwNkTJiDOrRYZI9lh6YITcb+y7OsXbxZL44pdGE6Dc0PnvCTmZyCoH
mezittXNBxF/NzKLegqL93C6aDKyxCtMB2h7+MgjduaJfXkmgZrRkDZDnwfT6K7QhcEv3leWw6Vf
TEghXHxV5NI2KHKDgpmereYUf3YEIJ5I3iJ/lKdCPsD64v4H/VUVe1PKgBe0T7uELObfPlt6CT1R
F7ptStPalk72QuTcdrhSBeU9SWSdhpGWEO1XmkXwnwsJhDEFb7YO1fbanEIm58MfM7PAGivPkvzB
JSpBB98pqVjdEHVC48qDmSVPrdrnHPepM16dm9Ed+Md0sJbdi3CUhSp0/i1yjrerX4vmOublShd7
HbN2RX99HKCrfODtX4QPIDPhHrWB1cKsOwB49vRimSMewwKME0y4x72Yabqv78iqNb/mRoSCIALN
BDKTBzDr4SS2OFwGIAGXoDyFhyYsuHVJHRuwLSOBp/ax61+HWlLQV1luooSAaNabe7EdrnpErAit
z5U1sbjyBWx9iZcYhYHkrmPdXDiuHCsST+FnjT2g24ipkMHE5xZL/so1BXigE0DrXeXejoCmo7Wi
wUcCm5Dyzgq6UP52vNTxn8oLBhRxUzd4TzLI8EV/yGgXOUQ+zhqpGSFDxxBjFR0Z/z1fbelxsYyo
Dk+v+kwuIWJr+boCU8h1Ze+EcobDJQByRSmCNGMRZ5SFMbuOGhLDszY6fxMr+YBOmPQolSuiPKfN
whav0YuC+cFUUBb3Y2B6omdpd1VteEIcsbxWFxz6GW9J9CZWOVvz9wVHQvJg1ToCYRp8RBqpBqF9
pvKpJNDco2zdaAjkcYnx4whRoeZzRt4VS1Rlp1sSNdctOVzXm9Ufkat3o3dlKCtZfZYxe2ge0x1x
QRbsAcj8oUuYmeQdcCHwWtMI8oualrvPA1LcAK+E8DXzG4IcoheqQpTTODPFLmNqKSRqnFlrwsIx
h1RFYiwvaKi2Ce+H9pXUs1e1l8rR8t9sGHcRw/E2T07cD51CR2tG6vktnX1dqZxySTJW30akVJRP
FLAAMMfldf+qN+OMv9NDu3qSGgj0NNW47EwQtg8b2b/gteu2Y3CwHJ6PKA4QaWbcjIjlKBQoQTQ7
3lmIBClHG56fRNkBueBVVjX254XVTf5kqnp6UxC66DjAohXZGTD2kg91qUdJcrXK8h1avj3nJCJd
cvua/x3ioNNm4CYQMBznqAQjWIuDCvQznPLMmE0T1fEJTeBdiXSZxgfAtGlyQiLzdz2D2RkMs4ul
QT3qpjrwHgUsk2KjZfoRnXdvpeFSMnlB2DNsGeR7clN34Uazyhb++gIEpy4Mh2oqQ8LCfS5+SPb4
a+cplZKpPKvC8JMF5kf+ena2OYH3VWiO8Ppnk9wuTPUcFzWcdUsMJoLtXifv9VTlTQCCfGZRTRTy
+YThZmiELR0Z4w+HRdzlwjoXhTeoIab43cfTDt/ydOgU1wyCq6z37y19gBNUSWEpRWqZjk0eBbLo
GUz4pJUyCN1ainYoxSUONGze2x5aOv0Q2evhBXaw4rIZjzq4bu3CxfQYnRrcgY9TFaQGW5aBN2IY
9PpZGR6Gubxs/1V2qwOA605hLGu8ONiYdRMu3GXq3q2LdroM/u3hQ14tkT6oOoP6DE6vvz2xSJoT
vjKS9A1FQyzJUYk66Fc4NFv3SEi8clk02UpG8DAym7pX2vPbHG/baHsunKus8pSX6HzvfHfIvw38
lefjf0j9hRLxXJKcuZfoePvue9bBwPlw/ifA5sNMtXnxbpaySPIXgzzrZDECEtf50JDdKGoZfyqr
PGsLGpf1gU4Wb4h9CCHpj/C9rSsXZPNYTtUtrz/ssned21j2P+bh9hJXXHBSLuTjfQ0ePQMD+9qT
Jqa9vL/UlRZc77RNedXzlwrx670h7UlHw9+4WIzZ5T1vmz8uiYV6oODY0nrnx/Gb4KQNWWLQn4U/
MKs5yOGi1t4Umcr8f6uZqT/34poloIZJx7WWncVZwZtMTDMdX72kBmtLpG7eY6W+bxuk2NM8aRGO
vHqhATJQQ1hAP1Ykx+i3Le1mw5HsZswR13T+sxPmrGi9YsHVnHaBu9/ssD6ZJdQiSITLT4ISwl6i
GGTJszmv+X0Kx4KS5rcA1wse6NhS/fnKEuFEUu0gS5/AxFAbovTYL9PEC4QJ4NAyh5+4h59PJy5h
Ssxexqf98VL/FJGZ/z+Ue8EQW2Ljrrkk3NnKQyAYaUXXIMwp754fkE2etyKhozC4iXi5XE77+uDN
lvoRMqkXXPQF3hBeaMkeN+W5oS2tyKQUS/up6wQYUY1ug1/+HlaKjl0uPh5+7SYzAU+eN1g1KXJo
N0DQWhitszo+AkKGaKUeRiWY+JLX27iQynuqNG54GP+39BsVNRwBwPFQ/2IYKoUluWuamFLlNeeY
emW2bn9THX1ckbUedRaMQw1GPFcOWbST6KyhZQufvNJXwriASBzunt+p0dGiZn5qQ2zmSRqgPN6Y
A1UwAcGz7Adq06mkmfGSH5/dAiQcXxI+J/CK4243POqVEmjTlQlRSGHTK8CEFCwOGbetuAmX0RzK
ZveHLds7EFjQmVQUsK6pujg260q2NmW8EKEfNhas3jKtjN+8sXlUD4kx3bX/PV+BRYGLgBHvJmrF
vjqu2l3Fp3fAxPhculcuKi82/ZYiaxrx3/wD1j6Sp1wdSNgZV8sfoYUeZbH4ng+RxDNw6niwWPwZ
A1TtSaxxLc+rQsEOLj4OdKtsLFlF9ove5v+SDFptPMLCUUKbZySnt2yHECvxEAcfAUOGVrCeCFXv
a9ZPSx/ntDAhNxAXgrqehwueRiLK2x1GaqFr86ciFMyJE18laGFJmSkSppgQUxObutt7aeZYXRro
dudkkgi8WBWgKB/0kHhrJF+8tnlbIGDq3qZimbdpe25OClpijrsAH7wRE+byFlrpnv3Jj4EKrBqm
/+l6sriFa+RZGw+Gl7AlakgqoqW+c0b1zXz0Tvwx0y4oKUzqzeviRJ/58sI6K9iJBoDeVE/5VPFs
9Yq4sKEYuB1szzSZrA5iLAvdUlsjclHNqdhg6Tvul+5cWwSpOFndQPBCFKGMg9jMwjfAh8ESAPFR
EK/GMBSq82JWA6Ik7fQYdemeZAgUbOsACrieSXwzRPv1OrxZGuu7OF3TSUXcDLK7/p3eVEGyr0oG
GxTzo8Ouw+asOmptWDGy1NiZFVXCzA6G55MY4VjsCagoH7E+pCpSKNCOQfA79NAMzCidJR4uQZ/m
+6ctWEUJ9xi1mwpolx2E3cYqGxsHfNUD9BUMOrWcNc3iMZl7/+Bfq3iYLEYBjZT07/6FI5EoNPsf
yO7ffBIbYx8+28xf4ZxvBpB8JV3lO6mri7QueAstGdX2oi6HuraFP8KOx9FNHhh7Wqcn86PeNAop
UbjS5KltCMA+rZYxeBEjByOLLrrGwb0GYwP3Qb12fiscR1X1Y0kpXiNq0/CtrDcmAEIjEvzXxYAi
Ome37SiB1zC4k+kiNxy5R5h1KY5+rKc1clHyD9W+/ySKhvUnid3RrGxk/YArgx+ST0yvSJPOi4Ec
dQI+dCn4JHM+xJTH6TjfY9/rIS0dBjdWuJw2zOchhOK/F6dVgepCMWSqfVji+PvjgxX7ATSZzA90
4AQBXuh6W1v4d7dNCKXHqjWhOpSY+wR6tis96kMlUVEt+KOdbXVSH73DM3v+3H7n6yrAyjNk2xhe
LNFFI1RTEAm11AZFaj4wggJFE+TiB9ZS2jmFXSq3/pLdaDYZjDohc83MRkzS3myx2zd8DAoSCV1x
xGlTRQaeMsXNWtWYBGpYMsoH5t+szpYEnfFI6MrANSC1bIVddzr+zdGoa/dGxDEnn1kgQxSE5DZg
+3VzrF48Lcr0RTsWFIHKiB9FI6wPcPVNb4czgCZ4FhH5/+YTVLnQ4Osp4Hrw/mjyIGJjJxCmajz0
dn6znqkKscKiEQgdlS0NJ1D8By2hVQ93IWA7xUdHepQoV5XTa5KfJc/QP7M9ojubdcfAleeDvPyx
89hOFulu+0RmQGldNJB1a2U9wFevkC5EqLfpXTZv16mKputppTNim/SzzPv0WshXUrTvwNICd8js
JP5bfjVFP0tJPgf/y2J1KNFJ12VOeCihwBP2vkgfBOoRh4pLOm5wNadTDX8Be0lFoC3lZbkVfTDf
1WnAOKCpKxsgjH3pEm/ekZpVa18zmcIuDDDofU6PAFS0vqqhLDDv9CTsfFJp1WqHH8KEsljv3+EZ
QZvz1vlAG0NerrD6Cle4CjetwLPURGOHpVlvhKqYe6OPDo80irhIUEmpMlh1YMz/mdeIZJrJ+uKD
mcqfERwvK2oFcYT663ursgL0zUfsHg1jK+JtTxS0gU3ythjruhFadoHW6eAubzgqPQKI+KEK6oT6
5HtytYM58KGaf6kWg6u8zhWGddj8hXHRyJ+MCIQ94DbyOx9nApLwCmdMZ8lKA3ZAEcIzUw4heDGl
7xIe2oO6bWv3q2b6XihedicSsAbuKFGeTqiQMBUuzRm4BOpyECOMnAmuvHGZG/10gt9mx/DFkTF9
1hGQgUKwzgsJwIk2lTZdjG6HSFSAMY8rBG0Uty+8f1OZbzGRrDP52iaNrLpyVl3LmhyaFYQhzx+8
18BHybEkjhzt6jrzLaYvX8gKZuDd9VyXtXzllaBClTd8WPSPcd3j2IswvQzxdSuSBnOmRDMhmLI1
EiLWEYUmhnTQijHyH2U08evFeZ1YG8Iy2uNFC9IUjpIyQKifmkQPE85B6ryzcxy7Da08M/VjAsH0
yfJLSHoZxsX7griCFFTy66GcOZJzVyguOHN5F/bXmsub2Sz19vC6O0rHEBYGTiBepd7YjCZxUXHu
esDUtHPwLLz1d1uG5Rgmym2JJCDfM0gwcnWeGsp2N+PHknvRft6Y1YTOwHLRWSOL383eskaJmN3T
rrA1ZAWJtsi98/9PzoatsHKo6HNp7xHcnEqbPKl0niIfQwQam9BtU6NxCS+6Q6HL6RBxDIpYiKAt
jQv3VGiU+nrhZY0i+LlCa5GNZRo6JQtILMxmXm7tcJUXAZl8TUL+t8vyciQNLVoc/ecy8ehg2zsl
Bd0q+keyTGo67e5GVHVWeD/Gs0TU3SU26A/vKEE45VVmEkpeMSl8bWTlkegba5MCpt2nGXQdg0EH
wv0H+XRvPLewtFrK7N39brewkYWadfufI7+BWfJlgUp99RXDfWk0QXxM5lvmxSo6AScxCu4MTaNl
8jELKysAC9BClezK/Rw7b6FdqGrmtJ9eemNF8i2dFj2wiGCMVvhqrXptUGJ5xRCDR9vi3a46A970
fyIuhL8w1aAvJHTic7CBNKQSgeeEHr/1oHMy+0g7X84JhdS6nugr0XJ8yXN5zwRLSyakF2NGKULL
VTBB4Fh30aIA0XlQobZBUAsa1pqYviX2DNyLUq5XBhbc1dqH51f+ElMOjwkU94MvXMt31byJDizr
Q1B2b/4n0i7wpQ2ml9/h
`protect end_protected
