-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e7aFd/CRbsj4igh2lwNfnSXnHph6nYbuFPbyU31CGHIdvHAjQSvZ7yabNNNnVc1+CIQFd2P36cZK
msZAmf6PStcJe7BIa5YBwvDJIK27wosJPRnuzwiITuBXp6mMcTTTY883d7UoAxksNYJA99d6vkRS
2PoehjD/Us4u1qbQBXSYGxAnxGefSo3Xb/59vQj3kGeaJHXjOt3m0WtGXhsNo2udB8ZMD0xw9xLW
RL/uHrKXUJfsEr+QmfPUkSLOfOX9cgHEkOLX54nULxU8zP4WLCHlObvjeBaY9B7gbtUGybXJfauG
kn7wPkkPKG/u0KTy4SddL0xtsYWb7/LVlW9Cog==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25264)
`protect data_block
CSYFxkGhusXSrqaLbcn0ybrMQfwECmGNvH762Q8VcAuIBNrm9sSEYC4+CsB4x8J29ok5ymW7FnJX
2Uo87Ud73Em086qnRr8t0CSPnsi39/sMEJ92t6Tjj0LH0XjZLBY0T3+g/VvnnY67x9SKgxPnqoOC
e4rLtvF337k0gFvjMreF2LI6vitl2nlRiwM01xPQJsXSA8dQECdgZidMqRlh+ubaTAWYw/HEYvTn
KjKb2Zwd1NZ+/XZlofYgOQwT+VKGVmbzMOEtlpddZgsPojZrmNCzbLuJu17OXh8bd0keoVq/bhBr
1xzmSVSCEAEiyfcC2T3sEuLLeM/pLsnienzyuWJl3zUZpTLYESkPhzdHSdLjRLpBGbxQrgVgilAV
zk8dN9UlAf+r5z1JTbcyyvxbqCAnDW9ZNSBoHmM9kfbzC4YxXIfPr2SfHBTQSEmflkh7fY18j+Mg
v8KEoZ5+kOpmFI37A4lXm5DrLcA3N/Qkck6TsK/GfH1xCIsUuYUcn3FD6jvQpOXctUGU04gsjjUh
SjFoJ7ErmRgTZ9hG2jXY/7xdIZ9Q2cN/AI8oFDRi2lZiDJdfkNvX0/L+Uh98sqpertJ/f2ZSZjuo
qxn7Lwf6pGA3QkLLot8pQdGqq0IoVuS/fD5cgT+FMmmKtdKpH4GYfu0camRH5eARo+XXrvqH/iq/
hlTpm0jxTUvXhf4PWKFSkdc9f6DLbAzPFc/U4mHscWrqoOxcl/shr3oFLUOEPjjFQB6MiY/0uFpm
7lCVZ3oT2UHca/rJHrthNCGywJP76T5pSWvCeHGPMdHlHQoZ9gLGUHBc01oBa+7z4SUSyunenlnO
B+otY024Ti2i0I+KiwAB7uxd5IljdeWb8mzuP5Qyf7H505nS0epMXzcHmp2kTiH1Su/C5rJ3ps4e
RapJ5Y6eVSXgVvsLeJesSDuaWDva89i/DOSoJpu8YWu1uSa1uBLfwHA1TiS1rLNgnG/E8MO14UEc
Hb29jDdRt4bu5pS1Ku2kRUky8CEoTsaqqQr9evBmHf2F6RkrDGR4e+sbCDljGZ48h1aIi2pw8y2L
qNBeW3bIDZAnrgsof10dXhWVLAuSgV13dFdBlMDcZ14njq5pD+xTxV2ezuh9XdubcydkFg01QRPT
mdL8TuZMmCxIZ6M2uKzbQs6AoCCj7I591GBP7oUB16oL/sBY+j2UR6mp4QzgLtHv00NoNdqrz12n
S/Fwi7rW0LU3ZJ00cXCqH+mCdkuZNWvERMa2ZtwLOD3FNpIdeI93J0UOj+5S9daWpK8QXY0dAhkT
IQtaKB+l/HF6jyV9lZdszvhP2p8Y658ZrQ5R3qD9EQ7+P+y69TgqHWDE3vBqHF9PWS4aiqJEbdzB
FB/qDwCEVYI5LogfigoF/NrbN50RX2Tqm7sCtM6+m2RB1cu77neT3bzRUKnedXrleYCdi6fyczQl
yWm/89byMCcZYw1jKGo4X63Cpq/+AL9L0CZVdO/3LXqpZYrTMEQbHVR8e4bWQI+eYboWEx4RuD24
LazMxh2Kj9Lhj4u9juigPKO7ia85Yo+wi9XVAocU0YbM7uNIBXVwD0xyZYHbAgoBhep0ErGAU5nP
xCGsSUke8A1YEed5RntPGSXfY9RIpxmAmViLDAKL6rAdd5HvhROnAftARxH0wHObOcKJvxhbi2Ey
c3mEkgNlDZZvttyIAPUfGQcHvAzlnwl6Ysw7dQmr741duch9bGdeNtn61SBEsTBwz6mNomNO2UQl
KFxgeGN/l817A810CAQpXsqE27CqwPy9vbUVyE5o0Dp9uxDTOMAYhGhfFuRuFYTiNVTgaNLLHWyN
Od/Jshc6jIogSeNl4f14ZAd/wlSj1SIMWIxPXlofrVEQANwqtgEOprc1FWrrCHL7OWES4DotRvlI
QNKcRc2mvG3hRVhjaYP9vOk5pob3hjEozL45IerblVPAcUJeDzEW+r0k1lu+3JWe0YTCuaM/J/71
ZDmBpioURDKcRVS+oWMEJSv1kPCLj88pwxE3YJLx+7pgEJFAxGiO+tz22dCxwP9fNwRj8GOeAPq+
RYHbA+356PenvCwDhBRx2+oH7wVHcVcpPJN8WnYlwEiG69dsfzL5vZZzM5Nb5yk5Lte6up8EaxBS
VCJGOfdJg9YhK4gRcshfiNx3EQ4LEaRLRkDjGHvwC2Gl91qsxstJTU21vK6CoYSASxJlzyYrFjmK
DG6R8XMMv7l3xxE+m5uF8Nx8OdUeF2eyJBHV2C5bSupjhHplII4bzC6PK7ElJKsSCBxd8ZgvzbL9
t0QcDd1F1w9NWAWqWKzeqF4nZQlL6VptHlKvlKoLrnGm8J9yKdieYDsV5JUdEILUVb/PBQVLFhaH
EZBnDA05uoQUUsxSqNQ63KTLMrWuExBbPyCTtMPCTB7JresCliH3uR5EJPLU5fw2BtS0ECH69x2b
suIbF2Gj8KxGzDdgKCbbFFxhf8P+FNp8PbOSdKmPDRg0zWDqI4IhEQJOCMuyudBedFmO/QfdHNsm
zVJqUe9UFHsI4kOer6pXj041QuSL0njr7elcF+ii3L9nPaxig+dgEtc/PPYXGD7IhMk8jo0d5Fie
6PA/99uw7vj2gP4WCPuC9GFWWZKc5SlYbf0OwzP7tpx/Gtd2XcHaaY7OxOAF5fHI71dP8+ikBV+E
/nCv1nJgz71wtpDKU3llcFIxj3s/ltCD+bSDYrQyEs018piC4qaKdRbBtefZqRyFnb8KVhPQY3dr
ajnOwBmoqygTgnw5CGry+NBRMZOiDRZM/ts4XLmvXyITpwGVyDKM7UHaqyjeCTwfChZqzYHTWEI/
/AefQ3l6hlzPskkn5YnUj/wejSIu/ypDiRFBYCCNc3hV1r8UNN5dNT80Azj/rsgoyEfbPhzM6b6t
KaFftmdfuBShwl43ZhB1kUovcgAKiMAK1adRRAanAnvIvet4q4194Px+AzF2z3XNoJWwfYg+Gphe
Xvf3cq9CwF/ghPK91jW97IfjFO/pV5CVv6uJlJCkE73P4hYgysBfEho+1hCERGgnT26oIUxwt7Tm
UhlCwZfs3y1xbD8Znx8uYk1olFPDEkyFmsK5uV2B6C9f2Kfn6C6fIWy7gkDYvdWk0aV2KPUbFZKS
QcCQ3rNHo4ndW66UoJZ7lojYdni8YhctoWyGciJl08TrPseyMAN6w40qZHLBYADq5q+d19BWLWsS
83oKB44VZHJA3C8sqYAjTwAqL9n1CuPX3+Jt+ToIWKymbiSkNwlk3Qlst7G6/78GHYH/K29Nzc6a
GoHzTNgSom0VIEQ85AbkxLArEEIHEnwS2DGy2e3/0R3XInyXXu9tui4hmFrbNzVlzfxHmAE5YtN7
irxc1RYGbebGo3Bg4M6JcPjgucuBkxwgTB+YwQKHQUXb0fVg+qzbWaMUpEhvgnkWftGOdNxl7EQH
xU46UCtQ4Nj250aEhuqqNShY6Rcu6PFTPiI4nqBLOr5NlA7tJZHfJin+oHHOSBarWMXn2phw3qVT
axefSrSQ28ncCXmM4Z+RxI0aqn6c5UMU9jgQcqYWkJ92TyEh1XyUZWw2/Ax85j7xp75vZItG5Y0H
yIUsNtp+ZeWC6oGqEfCSVIb/i67dB4rY60dI9J2M2ddB43tfN1WhOAwGla0hv3EwFji0fK3ccNx2
EIU/TbGgZCKPRyJmEuO9D4CHG0ey2hBMwJUg5NnEYZyQzg0u+JdfoVgPc/aCSrJ2q7zIYo7oZVxJ
T8XM4DdmVIbCO24mbUM9Ovulijgl6Q+Hw3TyKqSEAVgDZEjieRG5ia9QPfed7/sQrSoCgQW2rJhr
jrT2QLfVqx+PQAgFJySngTQ7dhurNtCYRhDPrmvpwr60TpXanPUxfOPBFxlDwcFHyocwnU5xsh7H
IQgFrTM54Bg7EsFiWQoLakAGR32ElsPmYuTiHmjrF78L+YN25fxhgahYYYU7CPrgR3wVBQKR8E6y
jwZ/vKSgS6yv3mnu6rc3c59N7+iHoPuWc5LFptb7bPDa0fgn1hwkbc7t+Au/z2buZKLrpMxTqQwo
PBPteMDyj9vDicD7O+sb5kWeVZHD8OpdOy00OwU1y5/RPJ33+om/2Usz52tGJLOwjged0ZhA2oCJ
8hglpTkZhmxwe2uXETxn1BH4j8aWGw/QSleq/uDQTrXCPO2tmkWjgSDTZriJbZ0O71Klskqfflyn
pMmTODAa2cRHMB3SByl8Al7ypEQc3j7wdWQlftVB6a7ilkIaV2qZm/s9vzXWNzMS5IHaMgpqUue3
ug0xXIjDSA/Vcs6lKf/kfAtc8duJVULnXRn+4lkDsmb3L1q63Lur+D5nSLLo1hYmk/KZQgvu02LY
M5OOHnEMlaTxLVzs0nQUx387X5g5sR8EO1j2eA/jt0v4a5TNwBVQYMRWwzFyUmhhOZrTXzLPyfrb
0xLYedUIrRMqCpP8FBeTNSNc/m3EvU7mDWJR2GNmr1KKuQlIr8MvsCN49r3roL2X8WL0NCvdEQIl
MfP0h2pRgwlGd5KpdiPtDaFNMHpwf0dpcqiAIU8hMfdq1QJKWDYFNeqN5YuFD6E1d5jr0a+zf2rC
zmn93jkj8+wkjk5uGZUqkOYu7dzU1MqaLQuJwC4bzUbkCov2KdfXK/+Y0Bz7ARbgJB8dWILOyex4
tFbga2Hn/0FIaLaQqzH4j+JIEjIQgvDP+OcKufR+pLJNbZz5m5qCjMZGoX17vqp1qeeRPaQVi3PI
2ECsf1979m81ECIrAfZCZ7F3WltYNG2N06a2pOON61u3R9JxPU0+tvU3ezuPInn6H0eq+DiCO8uR
2QA3cHPtk4B0g0xpS3wRH7abOXcD7IE6SBf6CJ6BUnRRRGvG9lTgcbyZ/iorz2yDiTECjVbDmyqf
aUiUO//XscfsvltRrDOyHtpSheCX3ExeZFqnJwAV8ANf3E7aQmaRSpG5EM+Ew9ssWW5+I9mIryiW
mJE3uLt5vjYJsur7hnu9RX9E7wUnGIFi88XxdDjDITvKNHgZCKRxyVD/HqpHbSDgPI1pgmhY4k3S
h2e90zrDBvduN48tA6whK5yIxG9fR7gl9LxB/iPaeYxDpnl6ajbkRQA70/JbNVlHh9oZlywR71jS
YoVi8Czlrjrw387QqxZH1p6SuY1m6XSwQkDMWZ5tkGI5Bfnqx2HPV2/0GKaoK61r7MiMz1rk2YSJ
Wr51PE/5paw8VdrOfY8mfE77sfc7TImWiKGGwcQ8o4j9eJVEIex3S5Ct0eB6PAzL0ywnhZiJSKu9
b+GWavnXz2f5T3tMN9vp8uQ16GFdYLZ/dH0/WQM4f2kg9SGPzZdbacIlIyjkNIn0FjU3degv1f1R
k3JoENdIxh2uPmYwHu3ukyEac3La2PvMNE+t7mnksSK4b8+lPKTfYcxydDeB9E5hbTqTBm8ws44J
IpgU1VAh4agFE791MvfWIOELruHd2hjiAFC0IK9EGhJg3ML12c0q53DlO3OT8YAHNF9uSkzj4apH
afohrkPyt9GCTy6UsLAQ2K6JVAOVfaULqzr7/qySlAWW3Wh+Xup8x1YmtHSSOlYHjGivElcTikSa
CW1xNHW0nCsFQsBAJ7y1SUj6CFZVQZ6jv4ANFGJf0Bb5Eh2h054WJZV6AcihWp8S2qv34UHHnN3m
+JwSD++x40MkHyyTjKWDA/cLrRrLBn+CJnyNRtL3UGVj1RybWJ/oAjGCNQhAHLZ3WATqQogVbMHQ
6s+MDPwrMQ0yC6ssnNl/YYFH1x6iC4yQZe1O0iC4RyIwkUKRzAtFwCPAQT0T3lQmYVDo8Aj3G0TX
5b3yMd7r3Wh/3teOxKox6XF8Rj5J0+680+YCVk9SagUqOkf60A0ilyI/SyC7ROGCN1XcVf4hwBEH
F4fa0RQi//AvrTXK4KnFnVIFLqCx0K6Gz8JyOHdyY4hCYMO7v9bhO0fVGpM3ty/A8lE1WOI6G5tt
u9VpZMnkTyclEbV8/nAIQsnTjW1HVuQHP8kK+XNUoyrSipEvQWg3kuoKQhoqKn60tVzO/ZwYCqpD
ym9e2yA031PnVCgJhe8rJoYJfa22hA5NPsgiks0yOPi0UlnwlANb1S4rgxa+GXBRdl9YDVoG7uzA
0vdwSiCMwokcqxsvPoa/fxF717jMA7I3pNYeoXkktIsfibUL9G6I1L8uyIrZDerUZRubG37cnf8l
u6tjAWhuTUh3T/OazeLQGdPoZfts1K3HWO+lA9nB1dXFp6QoY+aqIGvo2v66PHGsc5kol5xEeTdz
FyVLqXt1GRNzjOVc5oWkKu9kUhp7wYXRnVrl7f4xg5ZPXtGo0HHlFQClVd94T8IakobABgzjHWta
IeT/WYZE5pi+tOgj9zWyesobLVfDMA+DAXpd7v3yTdi5iTIyQftGTUu5PCNf6Ao1trnjSajU27LR
QFYf4IwwS79KBNSp4Jml9RPEelZv3kqhfbAeMc8ars+C8ioL2Te6bPLvEFzWTrntiJ7/xSklW8aV
iyE5CEPOx/9wYklMugfGictYfqY4zsaIYY/df0uesrS0jsnGRyYxzxpAGjlfX9AWo8rnFPoxBtKc
zGG06Ar0BgGOBREWLHzow5LKYnnG2BGXG10R+vhj39OJ4LCt0+yF9A978IX6Ko8fAqW28YHLCNe/
Gj8WnaylaVCyPCmarV1CPEH7jh1zE7pPjM/G4dOokmiBJ9t99sXH7OUmMrh8uIehvkI1K8gUEs7D
Kn/FxYh+yqGqiQ2XkSbmI+FUKwjPBpUlT+8wXsgAWOQYDWt1fVgt6oNnfH2NN+EI66m3oecd+Z3b
4aquHPNmMpnjKCaBbwCWE88RPMdq3lS6I45idJo5Z/yp0epv2qm2rb9U0vfje/3PxFP7ISXhQ7O2
w2aBG5rin9Elk6RMrKbvbuVGic1QhPSeiUQno6Wl802OpKN1UZsl8Y40gCyCEKnXSQj5GcPxRKoE
IqzaP3mnUUik7U0vsowWwtUhWGg94SNZ7HehGzWuc8nE05UM6LrUeUA8Xo1P4TmslGuuFw9GoA1L
WwXxXw2zAEfDzoCuKDWjI4LNVaSZtMi3suzJOLfpC0v2OvGZQsv4A7V6FQtsrinzgSoHa9QfIGyK
lyL0JucKd+VTWvlZTRRAVevkGThWqOURizp08+BFojLcBj2ZN9hUrOitU5yYFlnITM6yuODmy8mT
CIkLDBqlmh+hDOTcDsXnfMNGtHkQmEh54wP0Mbx0oUqGSp/yy5w3VlP0A3f4E2MKaMsQQvBbQAh3
oPfJc6oOk9HdfZjljOMvmSH1t9rAjAW67LZoNLYaz70rWkEgmPOymw34H33llNuH2dAE0s44je26
d3liSTfN9XYy3JfWG91ZOUkgJf0EZfopP5IWENdCeqzBIUBbHRRt3yaKcqq/IalWc9RRiNY2/G7n
p1jApEA2EjRnpZ59q1p598rN7nxof7mYVDY/+4t3XFF9Lzh+k/DpCC4VKOX3fUsA2cy+wRgDcZpo
wQF/2SJXtst1/fdpn6sNjXcDEdG7scijtuWac5Aj+7tKs/8gBnOwnQOVPGMrUONgrJVjWSsrOLKy
qT3A8qZDJ9QIQ/VNjxxQSRC111Dy9tlPKpmfnUaZun4/Q6AGW7+FrCAAO8aFifnP4O5gt8SGxd6+
2wE88usdVuSfjVQczzWYdsaUzg8/DUdPw6lyzgJOx6yH/BRN8RY1mU1qLEU7VO7AeMc8iSmJmI8P
cEk2Z6KFATXwsVWxGd2otpPCjvoSwCH5QMkRG1zNRusNqdibYO9LtLgEQK838oBx6+A+zzJdjQAK
bK0pJqoJTPSsB6mlLlyrK9vJWdUjto+i3Yj5yDg/Y/L7494sOD9AGPubUxGqTDBoYkQoOMcnr4in
INLe9s08kEOG+7OFD8ydal6hldo5t3RujYIMs/J1AERTBzXAz4yS8cNDl408xwY4nKMhegUjRrlk
+dFsBJvkB8fR0eLTp2yb7jOLNeMUl5aeF7EnHSiMIMq0zAho1lAivt1telq4LxNpSuymFADMabee
UhE4a27oAf0zHzsawp998ZYyko+AOjbyvgbxLd7XhRaFxj3tkEn+Q66gTtzM5TzRzC4yr4/qHAKr
CRrFppYU/4o72Wo/Hvyd+kmpi0y4OaMyoEXxjWtbm1wjbfbUTOkaZnf/5+Y343ExPG/UDJVDRKPh
AVUFiE0uv+CS+V54Og9xLdIZqqxeVeK/j+qDJ2Ohbs7spFgEO6DADD4Z4ZkHsB16ccYZSeojEfrl
qm8YgU+cqhFhNRW39VUzLIYv42F1NTyGrhSSTtz+rx/aEpJ927K0aemYdvfCBHHsPh71konVh9xQ
gbRFrhzemJbNjk5WW7BUg6wOgChPfMd4ptiSPFFrNoJOum/jVkX64CUGZmRj53EBAJiIEqZTaB08
o7oNFREa2whS2y5xCsxw68bnm4qUhxvZigFJ5XVUR/N4LkozDzRH8/IIyeaTJAwEz8BE/PWbWyLy
9ElShDkuiA1US366QViaY2pxJ28GeRkte94eCjC/2KpeyzHDrvtCedj9PToAMG1HCiFWMHV7OCh0
xo2TqXEeVcrDCRbyx0k7BCsz42lrux5+rhxLpTCjPg8oIbjNgXt2nR2QE6yuS5h7d64ds+KkuQl5
BEHLxD+nZmMUFgUrOYiCxkBH9lDtJTWYwo6GxcesrP4e5nE1AabuvUUJDpMPMof31hdVZioDSVN8
uwnghWzuVAephvS4Jnr2/cPzda3cYVwWaYIvFma6IZgJs2ox8Z+iRtVfpTh25OUNBY+W8FO4c2Do
Uae4jiiHo0Mg0dskmiXEtPXrTlDcpfLbP205LF7o7Nd7m1Xb0muNPkg5VoR3GgPB/APgx54k1qwJ
iY7bEww+DBrGiiwNF1WfnSZVVI267lhnnDqS4+lGseo6eS4QxnNo0oDeANLfUt2PoupjtR0KGpD0
TzTDab+aMHWNJ0wm4V7SmHeABIoFNPzyiTt4UFdWWa/SErmN0Lu/e1E/9hV3DHJZ6z6yslzowXtZ
so6Z6SWJRhFs4Y/JwTbf5gQuxqWmAqRIREbbOCR3Au1Ls+pwr7j0uAz7lcUAzbamMoZaoU3CzMZ+
HRpPkswx/KLI/3ILiacFr8KBY2Amt5o4rF45s2nGUdlR+ADuiULody1DZfFKsaTK21lKRUCw9se+
ykxseDboGgR7rdgK1xm7XOIP7spNVopFp9jJWtOh4ddENJp4zBijNCWXqClEOL2yf7lesxXMmPoE
4h9J9sfvbOoU6fBSfQI8Zj4MA4nMvr7RGAap7rkKCDlwIkbM9SkqtHiOSoZi4aBZYtbkdXRd+EeU
yYyZTwAdCCntLQAtXWey/hN4PCbfAustT+rExfX091+vdIOoeED0xBflSx5UMP+zOjoc9rlgZDMS
B5vOgaNl6nGNdCBqLJJx1IkTJgzPRwxibr6GiRNG7rPIaP/lr7BIwQt6vLWrcfDrDPAuy4R9a9Di
OvXx6De65e6QYYZnmiHH2lJm4sUuwUipGMZT41eQ/ciF7gLFCH2upA1MqxOWSFQyE2cv9pR4URMY
koTCSfGMhdMze+Wa8qSbzP7EXp988hmPQXgTKUhdQ7DD8CY4hx6psSoWWtyvKAzbV1/sV4IxxA2H
fSlWMNCb9I9dX1LvLoMmvaJ5guZ8yaBv1IftlR4Ngdt8JUlLLpWAusF2DSC9xGYj5zP5OCErS0li
xyBH8sLAZc0UNXG3auwnzpUeeMdiZSMELJLMt2O/29ZAmAhm6GA+V7m0TYajUGo2afzzTExQPFYc
KTZEh5ja7f1g1vv5awFuq2P62VEu+zWvc6povlEWJefghm6vqpOJzzdNFSMPbyBGeNXUeD1MUfT/
MU6mB9UpSfCEzAU8jpBGIz+EYgIL1IKlHNiCuMKeK1vuOWPIgzZuvTt5ptgy4g0DHigBZnCE9Jmq
ZxVRJvjpoTVyao3Lp4aqOBLLWsrB2JEyKohei7uHxj7GnyjbWuyvESK972M7ippYbBaeVqpMjTj9
ZOk3EuTNnnjmk52eRC1rC5pGHlp4njXfLVdKt9WO8LlKf5n344S7DLn/GGCj3CYRi0oCXYqzp9tE
pkS2Z44Ly3XwnQejq/CapuyFupIrI/GNi6piATZN3DanYb3RXb+UPrn8yEjTAYXbrOLcyeDr28LF
ASLfQvy1U2b5MqWjZ533SzQYy3a5B2o/J5ecaWsfERHnClPXI1LtXznI7o7gjB7CQI4L3+KHmVzz
YohW2jSN51qvL1lgFY5n38pYKcwwKaTmyEZx4+DNxN33S635NBTDSCKJ7soTrUGWj3m2BqzZtUBO
CZJRsI7H+QT2+pSzNtXhiDgNGtWn0iTuzv7Oozsj6MQlQu+habLNwQ7otrY/hdYSFTkUIS23DUFy
Op9C63fimcKH0GhEid8/KkzhmlBHc2+opzvUiAwbtJbjVau6w6OGHkEFubt51KZqnsXjU+ufLSSm
dd5dBqFwHQSBc0ntLNjdlgA9fKw3PPEU13+T8I20s2jNOmhuzjSoxFALjTRgUMuFEmvvkKsDQ/A1
b7Bl/WgbjINTfhjihi4Urp14qa1xh/Bif3faHUI5KlCRIHq4oVmVoZExl2mCBah47B2dieajVOoy
PsuoYX9NaEwFrKMrBlIGpQOhRpz1a6Ia92WdTr+izIu5gvpsL+ZQjb9lYzg8ZCBjZpg/X4o6g7n4
2+s3xkBvBqoYBHDrCoO/uDWjIGwZRBZvQ/8htq05mKi9DCLXCMkxB4ZjNhbKtEteuTsj9cMSQDnv
8psqheuXxOr3bXnJaMXU+GVT2KuwpWy28H9/9bjCoZa+nf3JPaQtghaJZRYomvKaAmj+Y+/KG+c8
47m2N83JCg6jKAW9IPF1sVOSR7w0q0Wc0jq73icFxhlENYQpt6iRu77FXfCoNTh6VNTeEqBzxF/o
Wv3TyjCM1hdTy2LTF+jRB2rXYVIQtl3IIxlNO0X8tWhd9DawYAroMrClyGdYJG40A1vtAtUIMqIX
Pm13bLvlQLgWl/GwV6/XEQCwzTNsNfjB0KpS4Vw5PbKa7lvVXEOSqFgDL8H4Rs0AIZoKx3P73fDb
Cepg95XqCTRc1sSQGSSlWKamxa2RrENIuBjfq8jMsjYJYWrUtdNwn421X/ZdzjPpcvlfZNSuU6hR
aSUC8hnETIDYpvrorloth3kER7tovO9iV3m9E2/B3daPjZEQpLwJXxeYYrjW1zT+09YQatf3M8kt
w2m/IKNRVQ9G/S3bo3NA9cZVoBxRNZ6uMvW0eymCxo05IQbGXyXf7gdh+OdNFrNNUGo9TZzIhlEh
r4i5KSNfjLjpO1wDhQccuBIRTz53lv+8RfHJA6MQkR0XbRrDHwe2zJqQaM+R/cMk2BttEVwVAUBD
H2i6L3AhAOeYK0EHHI0GXDad1DZ17mc00AOCIlMenBMBu1oxiFl8UNUP5Pu3c8T14keSbBOY4FWF
R0Zb8nqpaq0xDQNqiz9P0/aMcyOe9XCbG9wDnI8Mc5z4pN0W4aTlCv4MXJmt8XNI4MXXjw1BCpba
e4Onhw4CsA1ifwQk/gZYtvDlZ21CphyYCD6zi67MzDMg7qIkKfUY/4wq6q6YVtYyxT4EoTEPsFR1
OxmElTdnqBUCZX7KtS7eFn/6TH22Slk9sZYSMn4KFw4U0UxSWlMywQQDiitVtEaww0Be07qeVCzD
0VgBnABqbxMjuPnWdwJ6CkH7Rn09QEppnwyOMZjq9llA8r+qqsqinfLcpNcSOuu7ZxrczjhmULjA
JqlnnUX/egh1yoRfGiuafiCvKIocjW8nAMqAbYMnW6dsuHCv2GqOVHX8rpW8DeW+UOE1stFyvKZ4
mMAmIkwHElQFT2qtRnbksI9CW00iKh2Sii0EMX2NcH6TAC38li32wHeseJLb9wRxZdjuBjDySTqy
JV2pkorOdSKj2hTFqLjK0Q/AZQbugQ+D53HQLNEoTXX2JsLM4XUph4bqJvDZpfziolghOAWDVJyN
DfzqYrbyxdvlC2M2h3SQCHL57BKCEYn9wd/9VaWVNCfHoDnev6kl/EGuoVa5Lvd4gsFcfiyToH1S
ZSozzqEJUiTg8CxbY7qfG9KlbNjMJ33OPZYKTzwv9y0Lpkbp1lNdkvdWgIS8BFXFE++JsE4QEd3v
kDkTyKVyVs5qt9vP819tl08J4SY2GzO7+Enlo2hxSFAcPm3GX0mzynUDOWOoBhuQyvNaRvif6oZK
lsVG52R1xykHjGxXxTzfB6L05Tfw67BzCbZo84EZpZRVg0C9DkIVMA3xPJQmI46Y+blfoAW57lGa
YYrQNwL3ot+oAwSxITaUSs0Og4OIr2N4itEDDQqfVU2ozlEy/rNOjmfAD1SVXV704f7qRzLsA3kW
fG9JqNaXOwbNc/SZWVXefXhX6sNlmOzNBAcgnaWryxaU/Ym4654JXGPIrgP3epmUyFj1hldCJL1E
tHKqpL3XVr8oI0E4c0+26baxHdJa96Har0Me0pvgKQE/6/k94z9rT9d3Qwy+qmnVn503sj1H6wL/
IrTL2KNBQPXO/KTryLwluPIy9SzT/Dz+FVVQQPjfGG33KOkooMlvjtHawVZSo24rE4nlK2wC3IhF
fSAaqEWbGtImvF/IxO8dzS6DZFFqPPGpKfUQWRa3LvqAUHEVSr2vdAA9OH97J6ZcpW9QioFB5tLx
LYqM0XcAYkUIqZeAL2Ybtz3kanSqDu/8UHpiM1IViAk52LblDVvyKLgP1pPo5nW0JWa1TaHWTta/
Ki0996xJghV531xe7z1L63GgveH4X6OkeKIXqkwj/X1/vSU5rrPXGBJT1/zCF9SmlfkM8gacEtHM
sDazUiDcUZfBMWwFC1w2qciHmx9mzx0N9lMKpEG+qmSkwLLQjSBLqzrNuyOB/XV0nJ3mnN5Hna/V
KVo3YKaE2ycsWGbBQ9wyo/cvg+iJBwSxGououXVJKFct71iBTOp1h1F6JpRPuGaqtMlB91AX3Kuh
mGU2ULl6ysrE3A+DFUEgOmt8Nk0sm3B/ZDcZ5uyEIob6X8PVvRtbxpJ0G2nAxUHZqiXJUzNlJKnw
TWY5d19thqOuSkxKLU8TCqYnuFu5B+PEiAqKjymim4wtBX88CuLB/1ZEbn8nG5ELvNufzac9YtMj
jYm3jPtjiMvvmJb/bAR+G6YBYluUriFbUL+dRNPrtiPonW9Uoco0m2M23qK0yVsKExkbTWX933mc
12YnqPDtsAMvFqlEcZgwU3icr33Or8TCbo9jiAm75xzvL/MNPApZlpZj76ndnGJzH1Z3Ym/QzFJz
D/O+eiMNKCxU0PwMfnVOHl12HhBYBuFSAGuI0Hu6fkk5bJmNnVdTNL581YUntWOnclDpGjeIhOOU
WsUz8wHguXAO5ZZEYggeSAjXITGHfkjo5FqbrH2YCC4TLP5+X7CTuqTsns7JtmsHY3+olyQaRyT8
Byo8Ml//OZgGbSutPeuqZwd7lRX23SNYoZqrZHZCLIvBHvMTQk2a3Rnta0x2evz/HQLLf1PTtxzv
ttXgE2gv2hueE3TVJatuBz/PtJZZtllEuhXH/sEveYeSC2OIi5KKHjjEZaG8L7ehhAP4fVYAqE1/
A9KCCCyEMbtpwOXZgPa3jzADT2eh40p2jK+2fC+VtcJ4AMivliVgrXmara35UuB5/WlEjG92IxiW
87b9slleYyKqDSejNYpRnn+HYzSaWNa/LibvTAbHws5RM1wzqUI1WNy7O3h6670Un2OZ65704Yj7
Dbz+l1EJWyQfK7b5CvmPf+DapG1CUmqqi7jR84aDhAxMTuBwXX7DyzFndJnsekloC43LJrWlRDz/
zyPc/DzU3YoPpSekB26C3r68bZ7WN3tulrRBDL9Qky/g28/mM1UoJMl1xh9Om3HUN1VdAOjfEoca
jWqA00g3l0NRYpj4F4NkWuD12cW/BoykCVAiJrXqvvJpqIawpgmCM0hycuw8y1RiZb/OcUv2SWGo
RllaZLFvTH5oF9cJ8n5tPgv6OZEQiRFCFim7rlDTCiASMj8RYbV6lYfJRNCCXt2aWlHj27Ib/L6F
ELvOeaa/JJzgfNdO6RD9rUaYf0ZmkFJyhD0aONA8Cu8gA44b4XrBZWrW23A7i1Y7yXD72HlnxBQU
faJC8vEwCp2Pj3RuLSuOWB9Odu8j0+ufnLPLA6Ie58t5FXjd3baZlp6aUUZ0VxTzC9jz5VlgG1z0
gC5METCr3awx5mY0Ork7IvXAve4eXvDRdxazYt0s5p8bYX+H4ZUuzBHRhCuNVNe+kcCrYBbhmZx2
13uz3JB1xfbHUcOeeIZlclU/5LiwrlqLVcy2hiA+2wsyXek/sk4PwApEuH9u4tcm+kk+j06PETOu
R2Ar10uElI1Zx7c6EL3PsCIth+d9IsYI6DdJCFxP8M+dshUxc3oONbvBNw/D5q6X9gipau3zbEHm
rYGZWzOlG7rH4Hi5lpWMYE9DatZJHd3sT9CxjJeLZ02ckP7K/KXjdeZIT5PfavCr42goxOReuDiV
M2p/Yer9ri+gO/vUToXKqRvdDg6vbWdqNOTGcpkwIwraaKGrCVBsAeVFVqJzw02BHaDpL9ia5C3A
7Z0ZXY55xnQiKWKhf7fM3dk3f9HKKA3e2DPf0X5pZ5VnwI8Pnidv0RcpxA+xLSY2Ro+v4QZTQVTO
pgyLnUf7Bc//p8T/Ezx5K3VZ5oPr1Rzw4ISKUSKVl0D8pKrYKqU9cPUeTtBIfjHxjb8yXIVnoJMF
w6Mf8ohnLeUT6q5t/IDqbKBoVab0QeSzSVoLZVPVZcNApoBUNwYeEcYpnrnGgQXUvwlpVVXV2LeM
5Gkr9tgm1BDoKGs/wn/WJTRm/tR58uxfcgxkT/WKM6PfQNkWfEaFMselYrwfiAShlFQI+Yf/PdkK
1x2N3u+ckGhMTeI8m2qrSzcMtkS54s8BTMpE8HQM/FhMEtD24/XAqiBvhM3BxQUARaJxx2McwJgC
aEjSjc3PWOjTiybP8JFr7yTyiYs4RCAMjWAXTzmkDdJDhUtnknzERzGMR7ZMAgilQl61KAO5romW
VOu7K6dBZcii+5KBDWQY6oxXj0eCN6+JG3eEjHxtBMwN+6+o2L4ZHhIf6d7A/TIB++vGP7dHlMOV
mT5lydp5cgkNzM8HJZNJ1ah+evmamIHxVehlQemFF8kYv8DPnVg8kU8vdFisLE4BGIsMfpt7W9tJ
3UaVsPySJCKnsRJz2F8Xr7GcrmOAEtWp35Xs0AfjKdpH57yFTo3OpC9iAsiXNJ6rWcM4ij8/SSmb
4aGtblIj/iiyXitcQXRNQFtpi5p3U2s6bF0hZCQasPz+4zmEedIvvAHuvn77d6rQX58Ax7I5fVGv
DEjfYoq8HsM6n0GpW8hGzPN6gvRikqgJ+a4wBh5/5jsVuro/gJ3ApDCtVr4/xDVWjiew89qj3vyV
8RojayZU5Z9NOcuE3ugW0JggXPn1MGKTD4zS534SLnwDE4ewgSlmBzspxySR9ZOBXUTwtPoRG31k
clTNPkU5XdvGnMU8V2KGqAQp1F6pkaO9kC6tG3BLkSnXN6cJcmpdAlt+EpsqpXV74bhEr6d5a3iR
p1YEXRTBIpsCWgUufz/dD/U9FJDa2nNCBVePUEDe5TusJQkzSJWir5WtgnR6+QNeiUNjU1olX9fa
yA1pXxTztDwgYgx4zfJAbi781CG51jQZXFPh6wPi7j322kmfbvhWxqEXU4+eif25wRhPPmuonbKo
vNGAt5Q9AzDgMWVhHCjjC3SkVPMoQ0bn2DLBG1VOBO5peLuPfzDYc8+cuJcOuZrryov3I+IuGmoh
9znyubSolbHwT0yA7QEZPiFtI6S7iRe6ygsoBs41qM6PhmOS6uVte7SCU9uSKehY7V6yF2EkgoqO
LB+cWvyl6sfaiAMcEpyzEvvSdz2dfC0BMz0MXTQHAmbcKRVW7hBM42NM7D98hb+QEkFuAo0oW3p2
2Qq8f75VcLRtsjIruJcZXNyl/W26Bux/HUDbJaQrYMX34P/4oNdlRteUdL0FmTqtgCWiAEdZRomg
TYT2QMqB0vgohtbneLrlthdSnG0PnZwB3WblOUIxJDGdgdn2uVSZAWiMTtb1kYIe/Y+gaAOOfMKr
fatmHWPyVk9yjybCUG444EzJqN7mILhBfJ+gBy25oyChHqpA3L6z+t27J/Ob+bkOrQGs+r71SOlA
efiKfKi7mOGSTUd3pP3BrKkutdrvKIKxhNjDPyld1OGDP+ms3spvzNJT2S4spAU9YaOl91Hlaphr
gX2KayuoOLHqusdS15OGmTyriFyC98nCJ3Y0eH70iV3sENrYCKNDPaWtUErwiOFyEBf/AsVOmJgQ
3SxZd+g1NP1ayAktr8J36NBVBbEqS5ZbdqAEHV+jGJoGnSSYXv73ifi7Xvqz3Vb6+bB43oYPmnxJ
XqdS4u+9M5C2MCU9ihmwwfsR5JvkoA/Sl4W9947mLXbl7kdiseS9bTYCXlHLmkTRCC61NWC9hyeR
tF6MEIepfjDWE/tYPN95DN6gFJlK0+RPMv/QypIOnnX4wJzFI53iHGuCXV5X8CJmBLVS1V+2JyiJ
Yx+2vYAxzAO2J6X0rCL5SdOJ/dLXs8wWsmcpqBwPLiza34JCxyIabWHjwyYH6k+yY5rjoAxKBweU
Kv3TjZpxwe4aVrcCcEq1w4OZvlGP1wY37Wjbex/+VBonwuftXiKrWJTzkUs1ygUmCwDMM+/kuD3h
0RKtaYfHVOh2B3QqkDNoqCexu4VI5YeAbWYbfdbto5FK/0ZZy7RikkV5pIrJyFGf6eS8FNqe8Q1M
BG+0GDzJ5ntQsK/tb1W65Ajjo5ibso5azMVceSFBCf3jjqSJ/S4ce6ZTdpGkTnXWMANOt1kzhShm
hCB2ZahZP0WTw2UQHB7nGeRnY/KCQjBKFs0BRqzc0dg2donlGnwoSyXRhB//AYuefNGx7XuYIJ2h
f78KPmpt3EFtI9KeMvhUB2KpwjhHMNsy6S5KVUVixVNn2ZV5HNFgwPr8YlOguatThzz66G9fvXBb
PUt/6f+YMkNd3i7ZP6vHyRqDVTG2xB9C6bCF51ZcDeycqJAfaFtK+JcYtK5bO76OMbGz88rcRuJX
MOgF7xxfjmH2N6Mq4/1JWBF5Dwzu5mZuUz3weW30VYRF0byXW8FSqEBO5LAvU+206u+CkzMeUVXP
Nv0GH2IumxCQLpJJrvKgncs6JS0VN968CuffT+azjyDs3DBFIv+oE3mAo/51oEVEjKkhoK9GHuMg
lKNQ5igMcyNm3+vefwbcxybiiBNE7CgL+XuEp0tBsebu3RGRM/54WVmWJBJOybwNcuGrruCA67Rt
Yg96BWbqC6QShKLM6dgQDUK8KTm7zR7x+CGT8QGZYMXfrA5stQ7FS92MmDF4j/x7hG6epKNZeAjS
WlXoi8a6adoEzL5gXjBfieF8G9Q0Qp/ikVmKyTcorng9imgqhINI9Ujn2/wr1ozShWTvdcco3EHN
VpAZN9h4S0DcYwcOrfHHunx0daQzSInM1nxYynjurMjBAj5dnc0pfL+qyRwFG+ED9pw+Y1/jZhMb
1O4nq2dofcOBC3bxDOKR4FTxhgQPrON1bp+2cA9n/7OoUYqubHwq26TpRYadhr4wrRFITsYInnHC
w106LxrV1/SdJYnjmvCI2ktFPEmlgjRYGmH+zy/QvXjCaeT72EX2lkupqsKv+0FYpBBJMsWkJ6ay
Xp9DHVjjsYYki6AJAXKqUVO4Et5pEfpHZsa826bNTNGnVgsphRd1uGXo8b6K+V5vGVTsOkvzL+xe
6ssNugucB6rDBc0l29C7zkN+ppRQn4g3kynGzux6EGjXivonksMFwaxQXeJd3wmD7k8S7N3Afa6S
VnDotWHhR+bfXi7Ihndo27D52e4M39kyW4lWBeZ0sYZhnIRDDzkVYkEo9Ev/THR0E8S71VqfASxi
dMNvaoNgH06okxEw6M/aiA2f8WkpGLQYgaf2UGmKiL+EiPSkPrngKB+p1A1qJ+ERsGNiIqevhtvD
ce0LtH+9s8tUKvkH+C0j0r7WQtOpQD5TmHf151CE70+j/D9l6FNaugU6xTGUEIeAvjwUybPfuu4B
LAHJoEhk/P8jaV9XctA6UioVTac7HtbkM7BlNDMlIc84uX1LEkvNSoOk6ZPCsLCrX2pcKsBYX9l8
8+0YQAzVZccF/TZMFQwipUjDtIIKhu4m3bmeifjApsYzo/ZohHz1/jFSq8Pg03SV7ZTvP/LaNRkn
YqUPZTmwxegxs5ywbaQNfRGX/YUoJMYg8wvjKBLBIJy2Wh7VWv9v2iRDeexKS+D03iXMBCvy7pBL
/GlgT2/dSzpiNtPF4a9IByw6V3E7yWYCxWPwS5tqUAL3FwqfTzU9fb1gWqB4fVfAMzOKVdNcb8sp
82Qo1H1V3vozeurNLu/kpXbRHZ8XFEYuUpqPZTb0F+CTouWkyo5VSjBLl24+aWNhZf5K0/K4ut2G
gx/x4KQNETXl5/9OqALA6gPUIsR7namm4N1YmjTsRub8OOCm/Gua1/M4y+wBGg6pn06rqiPfLy59
wHuBi5fOHrWN1Ck+Nmjw3FcuBH3nh0FZujW9uTWYtxzzvYCuER6/owxFlQJq8Qjz5Gt2qvm/R4Lx
RUN5KdVjX51xml1LqW71kzL/I3C0BB6GZlunn+Fwlc1v9Rz6j0WxPsW9gO0nMzMZyJHBRKH22azv
lJTXqYz+DIBv1WAvJtF60TXiezhtdem3XmisCht613qNixjXn8XP0BPzC5brHlQOoM0N0F8/IAKK
xlXGBx05eRpQJBQfdpYK5KTrLyBIUNcnVMRFdGsRgDYEVgUfe0XQuw43HQ6XbO6L2c+5lmztQP2s
lZeGPn9fGJlDq7cvt89U+CCwHMS7KniBwOKlkOxwHNwwSivxN7dzSgceea1qaAy8bcRTxK+4koOA
CZVGhbaA/8d/z27g8gyKpsegUKpoC19xpmhU8QZt/zML3tMYqIzV/oMm0Briop7Kd8jenDmBs4J+
KJb7/pFxOaxyOxt1CF5Ed+uhE/Az7xc5rIcO2MvTVGv/Uz/yCmFoHyC+W6BjG9Ifk4bTpKk94bUt
0uyZhIwVvuCKO5CHKl4eBU9u8FAr3GAG2IwQ5yaLixCbP0c/GZrDk9F8aboFFuD/CaTRuYjlgVsz
K2iJsOd86nCJvsMCxz3n0w/ma3ELjokMh224XKrjVqdUD/QfMP4brL9SwMZ1ymZAjaVUAWCFC7vs
S4luMumGVPWH8XYT3pRmnFfqm+owJ9olsZ3SR5z7iK2wauK1wClmlUSJgirj8ebT131kqHyep0iU
Bn0SCuEWJUWHROBrylFWzY1+I6BcdYMcbkg8biv2e3ubSEte3EGHBejR7Zd/Ox0igm5usAZQp8bs
8yBQ0wxqr9U1m3+7xTnfdNNHwW1g8I6w/Y8bhK8PkAzm9MSzmupqVZL5n7Q5OPNilH3/fprzI7vG
KSGRhz6erHzrHVNa6wWgxrkWKa1rTZX+/rCOGbS5eOzYTGA021BDRq2c2VyhnghOC5HwY35XplPQ
V/s7+ZEt38T1mzSBjfZx7/joo7LfSYQF/guf3uX1cWX7I6K7d0pPGEPUI+iJoK/gYbRg8xm8IL8u
SWo32lWYwb+/AIyL8qH2GQ9XTJa0LLnM/HfWBhCtG5GuaBTP4x7gc7T6cT5BO/tvp3UtzQV8wJKj
OV/RNgJL7t1BqVzTSbo2FdLKIBp6VeBwVgERQwdRnGpVHHqL6eOl3+g9qQtXLgpcNZMOZlajSyPR
dEhzKsq+lb5FI19liQrOJRwRA5i5EqhByuzfELXvUHi05arlS12wdC46a6uuj9agvC1TOXeU0TNb
fsBhKPrjOIw13AdgSL24QK1scc9ncAutbxstuEISYpos7ploxLmIxQ9BFuq9SjwAumdolnIMWEU6
zFsqFvv2+wGdJlpANP3MVlGjtW2hIt4E8Sti9idYjGHeNKNg4Z6sji6zN+38l1nTtNNys4KXqGzf
mLuo0tiuN/guifW9r8KkzXsd5O5td9MXOjSQhaB/XRA7yYqBpc+aW1PIeyKtUarH3RMQP9SQWGsT
HYJO+bsJT1ryXMejnZOwqqDmEwqTj/Z5mJTmuAvaI9yUlENq76nSwMfmGsigZII1GEvcRQ7xEFg1
SY5RMivYNaNbiU0JOwUL3tdVTmpnKDN1tGs0vBVVQe+KohweUWpOsDwJB4icbPL+lhvJYU6Quowf
B/EqzTroIAQN4oW+EAjTv6cRLEa80ZLLJb/wIUt8Lf8sF7LW4hEOmFQXzcK25Ft1sJXhedZIIcoD
g4ivN4YlJNdqUlWHLG+7DZfINGG8CzdeA8gEZveJp5wL7WzPjbVwnFIpELbL5H00ZYy8tcHzTjXG
aZnrqD4N5wcccaxRHTgdLUyokcDqSJY+AWq0N8Yq0yIA2+EUUirjEY62QQmOND4X0Anbsj95pSZz
c+aT+OJ9NfhF6SW9o9+8d02vO1UDBbZ6lcNXwC4avJJlRPj8LlQdhaGh7et+ekWTJuy6RKec2NdR
JcRKyhEsi+b7xJvvgPfunltCmaUatcfvVANkWhLwl5qSSWaOZ9aMD07rWUyViZJdCb1rmjO3mTOW
02dtkV7BMuZtNPUf21gboDfoWiHzwO4tnIO8pihlK+1PUTpg7IsmGPLCkeqNR9qWkT5pQCZbmtto
hensdZ2MOGoivE14FAiDK/6UFni8iAB6Ks5oES0jKsVEnaALuQfFLapJfBmFEtuPyHcxYCpo67ja
NTb7eyx91jUBXnOHqCdT+wSbZAXdSlTRzTYp7tsF5Qb0pOvZ8JJTC5DEaQ4FpF8vFMWihqeDnZC6
RakvAeESwix17yEGE1UlTZZ1Vwbon4lIAu6S4K00+1ISEMJO78GSCZyuFzt8+WcY4ZKYAji/X+At
AxBShUQhZNmZ8k2ItQMFjizi2500nODiaDI6GteNgSwoFq+jGMObIuZNVBB0V6DawX6N8QEoOb3Y
+PZmLaMnsU+OOaTx7fu6/eDFU+cqqCBxRI5xUxzgbQjnQyEO33ZFff8Msnbpo8XC9Bv7DtHXXZbH
Hv7TohfloNRzJ8YzXzUvW33tBSGD+SG/XytDp3DnaJyLlGyoQCmiwd2WGVOupDmeqwek0Zs6YT4X
jr2hENIotoymQ6ruJQHERLkZ2viXb3808keNpOfkH8cZ+y/bMOsIEjvgLdwi9Mo+XcY8O2g+PnaJ
nkey5JZGajcboO1OOrkk8G7lRx1vJEUii08reoLxamcSy8588/1CgR13VPTXmW3/Q6mKiYnut7yO
HM3bb1MIqwMwgFVVL6wtlcXbEWtg/PF7vXXA5uihYw20MOde5+liAsZvxB6/tWQT0WODScA3+TM+
tfXTY6hkmdbrB8QlhFy29FPmRO/kcAZhIkwHUtcfzAkqGUXer0+HOdYrhud+sD/wrRV46i0KCgND
wyeoSMko1sUzU6o7aEiLTyaKRi1FF8rx7/iMOJniyX1yPKQS6UbBJoT4/jP5A1QvXhSAerZAj2ti
1GwUt4dymnMYCBo6KCBnWnTMbD7Rriw4ftdGsnAyewIfBPmUGIW/YYplFSgO/6nt8NBI6/czj43A
vqarVX6PpLE1SkJDoMAZ/JZplRhx6kdR9VXMzRznm3iKtYhjbg4egs0yva27YKKerhH/0HwWo9dT
/KG+Ka4QGZKkpDQsoQlC2yONyg08iibKcYOvbROiD6MNnOgBC0nmACJpimaTne0pfvvnVEbGlx+2
HxfUxEC6+oaO+F+fUcw9xNOfu0Qn/wyuoYaWn/euuAC39rokSqxgSnPRHk9zcAxioORE9nmyt3Bq
hssbDbQIvZ/1e5lMwCraKL05dNNlv11iL9vVhafVUXTGyBdZ0zXUzq4YkaSkRramD4l3xIc10cxh
F+2y0O7I6ZOVYvFKb/L23e72H9o9bWZE+2MjfHJBm8dZVJJqx4A294bKW40q1UBkLz3ZgzkBswwX
E+GJM8l91DaulPnXWrIi8wlCZcWAeHX6qpZAAzr38BVouUelKAGW3pE0Y86TIWUnYSN8/EReeiss
qAQ7dlbn40Z+esiFFsDi2mngLnfO7YeSZmfjX22IGO5B2g6uusBSdpK0clx3AOlmPbRutV6GrnSY
PRClSEY/B+5Bgc83cAwJENhnH8q59V9RM8tjhWrlw2MY0mtuEflbt3qGFI94+F29Ptac659MMNQA
fSryPheqhKXPJkF217viuGSqiksO6/4LeLhIjnztsVeN5p56LsZGPvk0dGEUrFlFxfg2VdOYfIDf
75W8nyNSArxLFRJfLI3d+KInm7XOFqjWhUkkpOcJqEJgwGYaet4TCmBZnpx7fh++p0S47Yr/gEju
uyWLtEmlscumVmYZJM5m38/NfDOu6k+XuR9UZW9DKYQ/eHsxjCwU3kjpLQMbQTDzyjdLUTMhgf9Q
8fHNTxOunNRxxGkwum+jv94IQ5QlmErkn2TodnmzxQAW/3NjLx9RZcnvH7T/IFsBBfEewduXrNLS
p6j6xJG57EUY2pGAQkOZXnbZz+hr3yhtFHFSwkfA68V4OyT5pcx/Lh7m5k7GP+Ug+EObonM1d6D/
IMBQA/8bCy5QZYMmr+YDYS2ThAjjr4pKgNY6IVvZKLUdhy0Jcj6OVNKTzFfd0uYC/JhJ7mFvfP2+
J1anh2vD3+9th8aB8Ag3vRgaCdVtkbJdxDnXOsUwpFo+pyH75rphnQrVQriiiR9Cz3UN7YtcuwFi
pfvxXsYiWIXsbLocECzbdA0GzQxxMFVthTA/M6Rv95G+Wyb8YKHtAIMepV31dRuRyhrDp+BCBU7x
yR1RfbpifwYCKZB1Dl2xYxf+F/9dJTsl0baldZuMYgMS+h9uqwaLxkrlC1b/VERT7qNx3MhIexrx
Cx+5iRpX9hE2grmK5/nJ+RfY94W1hHCdyUzApAoeVRe72oxXpYwfsL3URvst+CkcQFnRGIfujyzP
Y19RKlCkckfWSF/FfeAVQmzx/Fa9wO4Y7Jdl29+wktxQwIFOuECtNcT4ArE4qeF1AD/pvBkR4Ogy
Dm4f5IyWRPfEPBDHpYXRbioUwzOoeVOxZoYq7tuGc5SsgCTPaSQzjNn4x6NreOB+9qNzrhOwygH7
bMysLwmrNzbwDvkfXLnedXb2yqkwnags2AFAa+ADDamkAlvfAeGHNKetoP749OjeHRY6dnZaVas4
ZVhXjJKfjnw28ZqwoOBMjfrN0X82BkxlQj6hFeq3RZOUj9bJrf/aWn4fmuGiIRi4OZr63tvW4Ayo
oCVBpNUFwDsc0QE7asdO5ORB23g5aIDe4ER/HRLFpdH0tfYgHaYi+ceeoKvQjzr0cmr+y3+Tk7c2
TDCQpJ6bJxbbnLwS0uiKs4cNeXhIS+J5rIA+CkqC3YZdIDRxvwULRtVWcnnk2J1XmqgGXnW4QoSS
fVVgA4QPI+RiGZRGCx84vXonh9Lx+0qL4k0Adv88Eij8l3vYiUpLFdQdSM3w2aCE3cBQ3T0TAN61
7IC3NOCuR2elAAGzBIwX7p49x68iqYr2jHpzBV5H1ovDOZbymStM0OXBFWzc6xNSAnt6h8dPWsvs
rMw25QHSCQyQCT6Gi+0vGKFoLVk64gJ06QdXemepVsdAjUcQWnOUT9dZ5cZexvOh4IGC1Y3Z5JkU
ErsTpwLoPOm+Hk0OAGYjri8wC6cPhJ9kqwM8sCKPqlWtwr96IReEEM+zOr/HhNiQy+/zNXlicu1c
zhCcpEcq+bmIrSo+k/F8FnblTHQz7AnaNbbexkzis9uqZFi52c96FfKUF0xiGo7sp3cSlwoPuiHM
tnejpgQis0mcZKSTvZP3mqSXwhJ8rjOcejkd6kLLCN73JKar5MeCFOV3v3vGxfPRcc529VbeypW1
Eq8snL2501WxeXbsaJJqW5Zv2ZAEQdaqAekNkvuzJNdTylX9BORXu/xXkow4buzIzKhNhMxokfFq
Q5QvlAF8B1CD16cDLtL7Kna4xQzTLvv3va2uyZs899QDfJGMFQ8LRrBkk/MIWgE2RQ3938iYmZL5
mFWVn7hvWxIzuYS1z/S9CrdQCmy20R+xjripCn75T2S2UioACfTTvabUStOSxw+Rd9yRA49o20ns
K6FYpHskGJZ0cBY0DV3ixdU/VQ8CoK51xd+BlxOO7kYMHcDNhypLbNAk7koprofoEsYtbKbPaYUB
ZUNVeOiuw1M0aq7hBKlQzZYjRpa5vZTHDDZKrvwnurP24wBMg3e/BFN4k9UoezKa3QMQb3DWl67P
VfSiwiw0nkB0gdev//5k+ne9fQRvS/1tjXe8Q69XtyHk9kRwosyPDFPHu+IYGISukKN3dvco6Omy
PbMoMuXXtYNRoBFCv1lt4sMglkhWt+4XPYKGfvpZH7ZGSF4HAmskB+ZW9SAXrNKWCHQbi+RUPYZp
819UgbUpZsxA9fYAfUg4oI6vt3FRgRvfFJAdeklN7ajLrFeXPA7dqTKA2qDk8L0M9cxIfFYaL7Jb
Wi2ojbNwTTyHnesKbOZnVyE0oLLn0e21Gvo7I/98gMOvDS25C0vNHxJZTc3eyPJrQkR0tlH5o5Cl
FVZvzbEn1qo7nHql7HTsZnUG+njWdgH1uAzm92/FWJXYDkN0fAiKuEZb6+aHKP3RbZp/npHNQ7Zd
kWNh2MS8iZ6DJy/7M9nwRXRMmgFipvr6E9ywkMNm3jhkk1U6o2aFK/yZ/lMs0L8psABc5xj0Lpx+
vJ00VWSg+Y2rHxaDUs0OEDR0L4Ivp8xDEhMGCywz4FhV9+JbIenF76li03Ea45uHvuANYzmp39MT
IOoQJ9Pgtk44MeOVJBUxkPebArvSjYSPpTvXOzqm5qou3FCCMJE3u+RknzJoEHi9dCmhcz91NUEQ
qBuAL37cfoJ1mKQcU4oWfhAHgM96B4ivo0LU0eN577srG05OVN4BZyG9I7oDqoM2gJRbJWZXyjjA
2fRcacnERYjwbYUrwS9E15JAa+DCI54A6lNa7Tetl7VFQb04DIuGT4KwKtMTj805MzgSxQMaSVON
mhYLiNvIZGTdAJ8b5vVNbzI52x9PxUMVxyiIH06AwVEPOCMmARsguE1p/tzxViCnMqB9trMAo47Z
KgdIwQhEOnm7Ty1S4q8xfDcwbF50nhyO7RbA2QvBLNllC8N0I9iDmH2zEr4w0gxcYeI1t9E7GJ6m
g4vY1GpsS0vMQgPxJQ4pljLqpv215m0hhZHE9wGvZuDcMIMAf8TQq0WcG04BRP9mgx7q9agQtYg+
NdP9LbEhrWJtDNm7S7SFp/QKfkb1Hz0Kg8SKMtI++mmGORCnZcOGMQx8kBYWrqH5S7svsdthhuZH
AXCmio+5QYadE3mP+LfOTyfSlYrdWpocAIT06vNQiW/qhU2jOWJer/Kc+ovFvC9P8dtvDW81T3DL
UuvSAJpH6PEHKpfAGiLgxw7p5mQTtYsnPUvy6B61jLSLZt+n13ZJ6zNSAR9yvkppNatwQiNSFi+G
S+JDdQqvp8UVkHFb7i2RnTRNv8HQpVPlAneOADrgTUJEVFBmlyxoSmNN7YWJsNb9lQ0M//hyOBJV
LXuVuqwB9rlnqWhEdmVQyQsEPgfkxuUWgAD58rrsiGgpDZ+GiXHJQyxSc19BzjexaW0sQqUZbWWi
kFSK+RNdBAQzVCaf+eDKWnfkWGT5EvW5pJNzf+AgZaMWQlQPI/LMXEnZ5jw3bxNJ5eJcSvZHAx7S
EvEf1FuQmfeSODjfhwCfR/HKEjsSgGXaDXlDXHsuMWsiGrxtVRxoaIiwDsYUbTiJNRL/r/QF1BMW
QU605P2p9KoNsJa1C5ZXKm0+JqLujcPNyUSpYrFxYSESdoJa71zKyVx9tarFu2+1aqgy95sJLaa0
Qater3KjdDfh9kmAawlPE7ZkmHKRvkMSidYbTlgOtjz6cGhh8YzabR/7lqndsr7ZlRA+HOXR67iP
p8y4ndcyVEznUIqtZnL6crwCAu8pz60Ow6SJWjULkdTNPPOngJdsp/NlFrdBKxQFuqUwK2WnqkN5
M3HQ1cH0pNMxYTuJSeHVpzQt1nv4H0NMr5K5vVShR2Dyd7wOLo8KDvszsh52oOSGlSsCTyrWuQsk
4iC21y/deJydJERUN9uxcE2/am0Z5/dlwCnzcfmIRJOjrgt1a1yUo1jNc2f9Rx47tC5skxS9f7Qa
wcEte3Wyh4/rAx8CCT49KjRHoJ2tP3AD6Tl0Zjzy6EmU4SqLnqGAZMQqScDJboyY3FMqo7mHB8SS
aTYLjTpo7NRvfNlyOrFY+02MQ1cOqZGUnh3KhoI3kfIDYBNpKSeJ9Uf2d+mZPQjTPjO/PNJccVoa
FJRTVJD42nU2+Kf1QFxgPTAqfp43Md3gxe1E9hlYZbyiJrWkN585/bUiDCeibaMqwvXL/87rbnBg
mT4uhmtQ2CETVUeXA965ZodCH4EeM8kINXqdMHeJtOOwFeiHrKMEqGGX1z1sn5XEsNG7iQxgnlqb
QDBTM/s85DvATW3ziWWRCH1wqpVqGRSNKBjAwQmy7sInidQOeUf8YT/TKnnEAA5W+wjm5eJF/nBK
EtykDiLy3PbBbRxUuasXyw9dS4Nl/tF8FS6afUDZZhX+8txn41d+4t5AYmHPtjioDNO6a7UzQe3E
uYXL06GQNSIsAU8vKzCiERXSMnKqjBSXFdlOhHPBYllspsN7YhneB8T41NWE/PtT1I3lEcI4wnrk
90sYDBcHfgM+rS5D5Z9PVEm+St0hOSACclfHOxvp5F8HZnIPuDcuZX0njtcL6iCA9lVfql1ox3Ep
nMRUlJsAEUDu2kLYUHth9x7qgNIduavH8202pcvmu+ORIrPIg7SK70f3qqxeIIampMf+ythSHBBt
To2jV4VeOZhqqRqmG/JXSs1bBlhVx/J65aS9kHHB68GaNGzhrAnHmi9W+k7bcqGgDYd4fzJHDQaV
vZXLvXH8OcLMRp0Nk15gV0C6fQ6u/ZZQ8OGCdz8+aTqfs8s8SN+ni7ZeWLrfUFisI35gfV1I6LvE
tDinukvRBIvtN022He3fZEg/rqCC76LWNLH6eI8nBnUbb8Lvgv0oCZJuHttEOe7zTSijt3tGPtqt
sOXdVHQDS6YZbooJD81KH82yzuRfRBHF4xK2aMW9RtBJyyWlve4GAaH5ytevNWT2I79FNSToGuMc
z+2sCc9hi5Z1jGAGa9lDszxLeTRVGel/Zhj23XNGds9X3ey3P8Pg0aySqo/nNf6NOasM+4QIdzJn
JRFFZ6iypx13qIAlIE+Dld0AJ1SqVZH2KSfVw1B0xh97Ra3Z8t+4cvYclzsT+QEy6CCPk63M5hNp
N/kKm3kxGZSlMvjcekJG4CyH2DjVxEiBLfQlGeBgx6FmpqgAbbkB0d+fBv8OQSz/sKoRqToTSdf5
HKZaxLy/GiQgW2RB/JZ3ZOBYRtoBCTNapWb8Occf2uaemlwxaWeVMbCrHegQpMLdowdpvfTI068m
JVGdDNEn9guarYJZUdwWgE26uO/C+9iqQtVPQRrqZ4zdwOIXEQ7s03ZBwTdo5Z0+dYRUA4oNWlF9
wTTHlIoTsDAhZQ919QHdCIeE2r/nImKLROXTV6wnKQvUAc2OZ7yNY6sxRcTgJifZx9I8RVJ8Ad43
V9Pd0DGir4oUyPtZRR3hZm+b985qXfNwkd4lkJH8NCHDTTDfJ3BZnoVj4mFn/KxSxmwdpDDOgIYK
na33Lfb36iNZp97lhwTWH+f9RFsjxsIQb5UOLxdugP6TY/MZeWRqhGlHmZpWDXzeFXDE5phwMWAW
4HZzHE9HUECekxb+X3NpdbNfaJ6W2hw+6pIRPeRweeeDaacgejTh8sYpFTmvIsNjI0OKb+CZVF/J
gzd+I4KuYjzKuhLdPeQ44GPjDK0Ggpz8sgoK3RayQftYGEOEfapecs+GkAQl+X+4yUrQhgFRAJSi
DXmR771NoNfFYEU0IAs8Rmpe1BV+x4mvRs9RkWwDeac0Iwlw9xj62jZIJFIMm7psh/fq/faAJzcZ
d/10Dd2KnzQFJByao7FgB2yO5Ox2feR8DcHLcEyywZVwIueTEpMiGWDGptLSOmvgD+V5iAvOYuES
wTuFLthjY9eVYPI+0tagVqik339zVLqj67hE8vpWI6N/9b/VH9FIxFNkDryUdnWPXPDp9wuGbe4C
9+9Oxq4ggLAKOgmFqlA0MJqSjkedtU4XGdEg68bk+34jXSpbyiU0MCpPF6evOoYOMBCPMBzLEbCC
MhwvtZANlDYeim7Loe077uRX/orPHcNPspKcWdVVJNUr/5WWRnaJ0m2JDjtHqYPNESmH/z+PnHXK
ysyP+fQ4aIciUNOWTYz4tx7p+lei6QNKRkhi8sXPN04eHYdLMMZwV7Yb2ifpMSaiY2iOLOm1cb3b
UEQxxCpjt+rY43mnbcETM+rPXuIrjZSPScwWnEgEFHzTkfm7EQbTcfLI36njrIGBSFxuLMgLoVXi
p3jQi+ceL2hL64z2N+CA0JCmWmThJ7jXnYJQas9z0doylZnshCu0XggONgpr0bGUBeFvmT1MqTVl
UhDxoLh4oyErW40kWzLXzc4Q9vk2UPMEflhGrrIhqoUSw+rp9+cFnAbZF1WwVXFhm+Ro7xKY4utb
uvv7gYYPCk+N+GJChBiTOvZSB75v07ElnrE9op/8m2Fx8OeeVQZ+8jDvlvBNf5yMwvCun8a6Foyn
RppP6WZfeVNAiiPRHQCyH0EJ1zoxk4Tw9cMPWM5neAA1/R6OSd/qTO4jytjdAwBrB+992ylP0PLn
blVa8LdKJJPAvUgNIwy0946GjU2wZ25exijvN+lffxCTfQBRuO0Wg0JIxP3I1FoEIdn1lQeKzBoB
PG1Ikvv8BXfA1DCr0yG2duuO7P5xSHCnnwB6zshOirqRf9Tyj4NmQbNAhEdhw7vcG8h+PDr0S6vQ
UQrbtX2dHEvAjLPc5zcmi8MdKq6tvbURZQOmKR8ByegPBTCwxgy0IVRT6S+pqDggg88HdPb9rq3K
bGZZk3x0pA0qqoir/SF4YU1npp5mx7rOkC/wREqY9ys6SPtWHLUuXokKadgt1MhGsHPS+tCTqhnx
TS+8aJ75rgVa01B7YGJbmI/osuypWrLKijf+cRGROOxEInp3HFrEj/9pNcjIb+/xLO9HQdK/UQgk
LW42a3ldrliFUnIDCaFDeTiyooygefi976oHICN2m6T8rNwZ7umyCY67D2T0QfOP35xExjHxisPd
/f/0SctPg6BMIvd87eWYaLnjiC4PgBGCOFEd4TompaRX4zDgWryQiTvJFE2LeSbdbfjXFLZDWTmt
AaBJYxpECwZdi4b6wGqs16OTRvvwq/naOet6xWbjbdxZBoWN0sU/ij+Mcd1J95ZroUif7Pya7mFf
hyY8Z4OvA6uVk7d//fu68tsE9Y3KX0NjKyl0UEWd2bu6YZdi7GfRqUzWUV98hncFKzHzVxWU2MM+
2wepAEkDrzMInNzSkkDBD5J1PrQhElXP+DuVVjwOuVZwX+WnA8hZKu8IX3RdbCuP6dFDle8fr+Lr
IuQlgEeYOzWXd9jhrzl1VVcd3WTmrFEa/iiJ/QUUSvmCTOQNj8Y8WtFWReXBdWyKe21RZmwPKG4O
jAKSpY02hEw/eFRYn3AtGhHyKe9mgFvrDQ+EVrpYjOLgwDW4GgOY4GhZF435wysXEK2tNN1P6LI/
36ybzgUVWuuaBt1J8hgnpS3JCvsTrQiOD6gI1tRacMr8ZcJnT6G13VsNWGFIjMft9GDcO/yZ5YCO
G4iqY95OylvK78bL1FZJteyNgJwbDWiV/tEKqDOz3FLbfS2/6ZX7ZSz1UoZ9Q4lOuurY7PzhUPCT
1gzmuL0OfzwJ2b0gXyTSkR/E5zZ8kWjz65umTiNS0UtX/mpSvBMKCuHLS/sdfd4KtDRNrcXyZnnH
ZCHbAUam5Lf+JHSOpc8jjd8i7tEaoHXRiklL0l0bYm/ZMSyrjxC8R5GiBfyxpnbRJ/QFccERH/Un
jbMbzuE1zprsspewhkGCyApIl19dggJt1ws8BodJqSA9hcf5LNi/uGH5Bz4K0jREcd8p+jcm+30u
VQjyzxnChu/W4/n2vltWGsYiUsTCTvcr5g+2RSi0kSau3feLc881hhRhvhvrnfTj0Q7G5dNQnt3B
qxt4YtjfEH1pbHG7Zz9jo3Iiv9vPrmdITrUVIPvcahDBtg/OvCTUcG3cj9dEq8j1QkDnDGhAPI9w
lWLlBqMNZ6Jablzu6wY80aM6F64OynPoGjiRrbTdVK2j6XE3VsZQUQri/jjMfmy0OODFr1KuEuej
h+cfe5TAUwFWRHfAlrRuOaQ6he7genpLLkaTLwaRseyeowMFoXDwczjGVjttkiISWt44YDlzaPx8
uv1C5GpLtbMTmwVrUqBuEubjToZHPGR3i69AR8wzgRh824x2dpOMjjFZ31CpxpZRDyCOHXQXD/jE
KDA2/Q/yNt3vKxwuYcjejNXeDZaFQTUjKuCHvBM/W1s6xj0GS2FgE0TfUvzLr7EXeAeSgd4tceXY
WI2Og2aheNcYK/UNsrKC2SDErII5u0yUaBBPOaVMSLagHAdquBInbGoS9flrP3U1PcSliyE4n4qx
gievsieV7y7cw53FHGkD8H8zqO2A1Nux4ec4CiyFXl1dX7bCkDVJjCCmAvkK0GYqZVECt/PnMOZ0
PifQkj87sYqII02xZ9Y5aQxqZvRyibBgBh3JRbm3/bUGjcVLoKGdo9izLmiqQ6BEdk2h2bpPfIp2
z7FQy+iNRZ0/6RQVzMXkwjzYmOEInF381rIXWTBGnF5QBtA8bENdpVk6FILPAn/O7D2O1OOyLNKo
7Z3FYDWW7dEeHR4Tbs46xOz0/8tkBUB7OEqhXdD/RT4AbvGkbWjShjz5ncKWQoUjaOGnYYY/H/pi
Q/vzCOI3y/4UXKIna//BJ4uJdjCjrqrZRO0oRil6ZsqUOz15pqABQNGKbl/xCBpMJcKSv7dQJeta
WFQficqNSEwiFN7GcfFfW1gFoGIxb/3Bluz1oZh5tqQ3xsX1SGg5fIHG6BRrsJuIkWXkd5h5Wqug
/NLV9uqPhCB6aD3mL2mEy8TSVBr+TMT14yIZZC35wfiS3H3ICey4AWdpWmjQhb7YxO36lEes1bXt
ayY6GiXa2WE/nYbM8jO9B+GC00hRS07/8zrz6QyYN5y51tMgK2Svn55LrS2E2Qlu4xXh5544CMnL
LzIfy2ILtza/atZa8JNIGaqbg6rqNbkfWziw0M9J4/NEAwNHpLiU8pu2rOLOBIISNeq0/DM1kOex
IfDlOKa9qB6fqdXojS1npXCOrMj0BFLtk2XaPv+3FevxvvR+2bhe4h/vxxwKWOXOoCNhLho1XOwM
0vwXOxy3R8Yw0J85UMC67OLnt4nftE6zlTfBC0HbMNmqw0Ebbl/opJYqj2fus+Ww8zpfK78TVQiw
6NDDUTbKFalbghPJlY6WrYlMR58M2dqXhkhql4+ME5+AcPPJ+ZqzWpRiIeEEBSVL+QIvCnU2fwTm
z5sd5BUv8csx27jU3zzqWAP7p1dDk5tNvbGF5OnLIDrK5iCJeHRX+V1ciB+xx/zytmXUy3NCVq78
LjVcfrOfZ7lp5r4+qLQGqHALJn9R7Y93QeQjffygOgaduEPGUqc+rDxHcCNQaEUEnG6iPivx04N7
6hLz0H6DVUXR1UWJl92Q0GxMlWu+aRbWmVEPMymrcAMaQowstAwW+tolaNOIdvt+M+/vzssU7ElK
wMqF4Z2DEKIbTMIroprAeQqFWt+REX5VggcAeIIUWtEOTUqg8ILJFw+kAjjHkDFCx7+YKc5CIABY
TcqvQfIvH+Q03YCFI6I2qF3P8kJWhVzGI+Nnh2nSdBf0eAGmrWGE+8ZbpgUIb3TA0ZrhHZIyXj8r
ks38nklo7eDk0VdQNRLJgfpJOh0PmqlEM1I7CLtNm5Hhy8NfcnNL65g5Wle6ROfWBFbIdtShbpVf
yE3fzhT4pD5iEcMsIdS32Qw9z2Sm40PK3uJJEuMihMONu+r7FAinBcvOSDNKyXjHufPlUmVOt0CQ
sEeEZjzRWmiZbqAgvsxf0ktz0XLW9/RLAe+nZQFWnhcF0751T5M8JZl8C43E6yZgPYP7OO44afc2
ZBAA7rSLM6XMPIcNhI4h7JCfLtvCybSItV8MmJhMTw/iJ+hpYiJsbxxfWZCUGPIJrpqD6nXKFhzx
tniWtfkh8iGF4nWDjoNdCXGh53Y1crkQr/cqd7Yk98+pB0FKOKL0Z5zA3hN2vgD25NwFklkfMNBO
bd5wKE3Fv267hD5I2NX0eAElUmJsLNsJBlhJ57E95irvb+Eee1vGXPz/Uep/NQsPSh2mMAxXg7V5
JMMvitEF/OTR1s3hjEFJoiI46CmwYEDii19t7Wwib4ewBoFi1cGCVbS09jrISzgmF0XfowxxkYH5
Y+ctVBuB675Terq9BgWqL1lD6l4B1U+CkEyS2txW0UGWCquFJ1cjwUdcjYpeikkip7lwyroDKSG4
X1kjYSpMZQdltiS2l9KP50n3SD6GxH7AtlFwEjEfnEr7VOm3dU7UdWWjsn3qS8zXLy2xEw4PhpIk
nJk+vFZyU74SfjYxjFlUd6aEnry6bPQIaRLGWN313wxTQuJ/JnCFNP47GFzcVktqTZtFTVaKZ13n
3j8YrwbM7K5VFXzkmxYxMfVH4v0l3gfS+H+J1x0qzuBft0D68W5GPNC6p8vRBlBsf0jBRsr/LBs1
g+O2Z1DAYTWIFEv+jcqMDdASsEUIfBW9ZLnxQW9Oqeu5ZrLxVw/B/Bf0br1klfoho4oPcWZZezyw
lSCZ1jF0nqXwJGz1SOxrNMpZh3bS8xNYDPFopIIyar2PO/stmRvjseunFOk5sH3oq4yyB38h4Z04
m9wT+BvCXmzN85IKP/Z9brf62aWTAMek4vnBOMXqumX2Y6xWJH06uHfH8PukW+YB48RlZfO27q6K
Xi8itfsS81tSV9KZM/6Z1cztNOTsynRRaFVHfksVKIkHbS9PCBxc1J0mr+mdHTk6eyLwhzuz2UP8
QV5JBBpNSEaXS489ViYHHYpBIg9ulHL4Qlf4DDP0b+g1rqoyZznlR7hjpxiKYeEFPRo75/xa6tjV
42kMnHb++tMiigbrIRudpyiHNd5uRJJIjh2norNSsY6k0gVoOFH5SckvHs9iqiwCaP4SrtGur4Qh
wBdmSZPbY0Tjm0SPRVUIeqTeaqHu/EFA49zMzUv5ogpAmI8JGfDiFx2UuRNO5ryb5rn1OTmteVzc
WgLvlqwtHyLyPT8D7bShJ3vLEaOoRu6PBQmBQn+IaPAVHRAVfToCbRdp2fZW3XvkCnRq2/0BcDfp
oPS3ddbJvVSYXkJZWy8LLixQ5q7vWuCR7iDNnV3NAqNA/pIfIOlv7np9cjJE7q77s1CBc6lOL7tN
4bz8Pld8UpBc4pOaf5uqS1ZpbdudZiQfaWHH8q7NB8pR662sB+h5Cl4fa3BeMw4vDAoOD/J4rfWa
8QYRfWtupLuSV0d/MMBVltpW+ndo5Zdmon0EU76bjilYHRI4qdR+24Zm7/9ZPQ9cxOodeBCGA9JX
2VowKRtv1R6IWGNcEIZKPtRCnIbCfwbcRDzp0zydXpIQfPVaecM8jGT+TKhUVOUd9hFinCHlosY5
hviNsQExDixa+TI+hDsSs4fOmWZwiXmtvSHS6ZTMzNKAycXle1YZNJUcjbt6IN8BI3DMTB1gfpZS
e7E/7yYQkZtVBvTrUg8ahdza59wWcSQpUr90p9ycIZrTQY9GN21J2Jky42XcEpX9ROWBTuaT8XKc
439Kzjt006QZZibfQQ==
`protect end_protected
