-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xR37czgYlY6lFnMmA3E3r9N//6KnuvVm+brBCQWxm8JsdrlkSa7hMhaShM3NoUsVzn54qhbvkBgd
yDW0nYQ7sgDya/NPv6sInf23bA76XLnSwuh6uVMHfFtuzJD5ip34IFCqXTHR8CrF7zmvzbPNGGWS
ZYxJ5jPabWKepcmPog+d/nJ0gP5dQnsAjUusH88iMEnljJQm7rQMqSMMTBzw8uGeDf4iEt7/JqCo
QKZP5+CVnaG9kXfnUx0hvOYQGO6oxupUs1qnVUifwjAne61Puc4qLMPiEedYJapCwrZSuwd0n5yC
SSRBRD37kI8sYWVBBVgky1i++KORxtst5QN8Ag==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
0njqtb5gsmWIFgbwLG3CiYySFNh3i6DqlDc3hsUzb2GszBS7FokPwP0x3vfjJ7KOjtujgyNtgw1K
WwW4Za6elg/kMBpFBaCsDIq9CPmnUaCiX3NHuBUvopW06aBOLp27C7epFyttmxhr1mSVD82iWBjy
1pL1XjvFNYUoxWD1x7dXesCcu++fyH8Zek9ItSe/jrOfCiG07FQzGDC8qQX10xtCI0Ztb7QoUjC5
ogjqTfLzkus9iV6pTc3a5JGETFXxp3APOxy7kz7Iyo79Zr4kQjPZ82pvgOSG++qSjrx45LHIG2lF
A7DMjsLEaEmiUBvLidugrRyUZR0RP9ftlt6i6ict9NW+QB4zhjPxhe719fcZVqvGEMGllTyLKFYO
ISCQmBygj7vhdoOsfMVB1R3O0O2CSDRqaO9W6b1siLNUnk7YAQsXO13mf/YHoG8gom/lVgBrI4il
D2KIAEaAGjiohXi33CbWC+8NywGn4WtIcwHaaYTHto4lAbxkQsPjWOJfeaNqqigyONUepkdDNEnU
P7NSzlpYznuif/YMtGRVVwNY+DvjWjhESnqrVKi4DPeAGFZu1y+pzGNWALrrD3+/QQIZiimUBM6I
65b44oGmfK1l7Db3qKOvfE9drLedTLSWIyNRYyAtO4t6IDL4bhqp0dFsWwqiKQtRCjX5li5V5in0
Oa8Mk3Yo8gaCa5RMYg6tPQfQKoDDdDxd/+tNe+JQGCCXJKtTTynOH8WZ3K4f3JGLPIhMJhPCi7EL
2U+4VBoM+f74lmTHLVHx1o5MFkciUCt7rwpvluGrz5ChUaoweDGRrv+fRBklpFBGWKjrG8/6MRz6
0u3ZU/f/EiABvUMAo5ynhcfw5N9MOpX3zJOIJ1tS9E+n17m++hjM0OElbK0b4xwtSuHVgef33Mjo
DoDnCww6aQOhcnjWqdtS9jX7GMBoqzNKo7aQy2JHTiorkDZunZpxGuWrXyl3C9Scxq1qUm74GJnE
McS5h1foOupHdnD8nYSxZwAw2BIoQKhRHHF8Uqt+iSXElpTiXUo9GgTcLHJNqn+WAJhutXGlqwyB
4XIA4eGVmeLQkFPwQ7rtt1iITKLGD2/S1aUQxIdUkX2DdlISP6IYa3woocN2RKVvKnFrH++oLmTC
BJ9khPRJQrSQqlFIBggCwRFje5qH5+bmDc2OhZKpjWqBX2CCnFLxD2KBLsNfLqIkzGprpVvYsVGS
RuN1ml6WuyB8jGaIItsR4OOZXLalWjmBv2WFWqLHtSueoxklLE6Q2HOcBwVYEgiK2ubHMb1cj5dw
GNOPdt089e4O3wLyCHVUNpeJPNE1E605j3QMHi+OaQPMUbfA/mJa2ME5Mnuu/4/LTg+blJM20L8P
IcipXCPYWkzplLT2utNGItWKLIVJ0OufYVuIsNfNSei3h7/tNJwg3EimosvK23lQsktIsjhyE/O9
8PrUA0J0mE2an7ph/xyq6cgjyMKlrsigJGJrZVnpjXEBxOlGgY7Sg42Qo7PPZppo1Atki5ZYPMAI
Z2KyGbZwnmrbetH8teOG06UlLZFYhVamIkfsE2Ntv4BLBGDvkGV0oOctQe3QTKOA/w5aCPjXNR9a
Piv3LtzRXsUSlqVPhxH8iMVNFP1By1m136qAUcZrdddPxgRyZ1XgpdXD/URZW5lj8M5IAQFcOq/M
qFCrw88uler4DpT/rdAoRqQ8AFhD7BxFssOiv0jbTLwPrD6NYcVkmEtSwdQAauuCLAbq2wD4wkMr
dmlCbTZKFoKP4c34rTOPbG4FjlFP9A8sMUyN1CxBQgq0S3hfbpzrA2rDZiHPlr0fhNsIq8qh14JR
XE0GgEbBYLW9V1xOiLNXBrUYF1lnri+jxvsOo/OgbrPY1PhCRz1T1VW3PW/4eQbHmv3GeOfJ6mYd
ShtNTKWnpDvpzoDsRKvYkjBCTXJX7JSG+wo+9gCOdQbu2cyuIBw+PAn1rpX5bRB3q4EiTT+iqsap
l4Uc89V/Nf1uWJHC/KKnUeV8WNhdAO+GVHl1bg0FGNhaj9kZ46ubWQ1ElJOyLlFTG6Fhv3sOb+eg
y3EI01HOIM8ShM0SjKXRWelivKj1yW+Zt8exnVM3yzcapwu9x1zYemgEW9DgocBpBsFX8Qbh6x0J
oWiooEk9/hVYJGlUli/P2diYcAVbiVfIQbqRRjSEL7XqOPui4foNmTvGNHOzw0K0beCfdfOEBszL
oOia/kajJQvKUpUDMvV693oWtk58y8VFpJHZ6sqJbD4M73+ax/Krsx+6o6tDBwJ4P3CactF9M1St
L7R3/eHrGVwxwgRSJQ6rgM3tVVO+IavZzDBw0XeJ1RCZOVpcX4hA9IChru+t2lnIRDXPiTqFLQFx
YeVBR6vcfvTwBfs1aUgfue5Fcl3VXmksuxMryYSSDQjFIZjTpOcOk4J+Xvu6em7mXLsuA46N3Hic
/1WzFYFQa9CNQK42puL8B+hHMfP0QbmAiDePDtNfnIyU/TDKbsfM3/lTE9nwCbCw5u8wR5SjPFZq
4JVZehX9QY+jV0hd+E0JPl3g6cQ4WzP7Pzgv34IkNT10+wxlipbm1DzpFzuXkmaP4T1eUXKambNC
HtAzJvIHszmflIKPdoAU6OGvVevz+UQwhr+lyjWixLR0eNMHLXOa5uo8R3J86vQTH4Faany+kByl
4RKXw/yKs2TTqtbYpZw+XI5WtIMNVsaveGPOnFkEhf10hHg5ZOIvHIlfIRJ8/yLvNPnhZ7OcOEl/
XK9Zp35DIKmjaF5yZaaUkSq4IA492OVjmhicA4QBeIfhKFtkty3p/oXqAeK4+XpPHVlyHnl8gx2h
bAeIJgm+pIwtMiun87abRK/kjMaP8pnkgsiDK0ktwGm+NN1wYSMzt6hLEOtb4l3eogUkx6FNFstZ
0DAGgLTuX1YaPyAsH0saPw/L3F2SDWREvhgXSe6P1VS9Lq0Z4Bv9TitV1ml89YSCxQAUSXJ5LT3c
lbYwlLuESbY1EsjA9JJ3O+yh6c1P7qF0hA6dfhc6dNDpTmMc0gsnN6IK8hTqkUZU8+rgtz9r86R7
PPSl0OUuBEUTNDWNGn+txrULu84R2PRt1rOeCorn27ciG3AAaC8GDucxkbf1iKZM9Zvhf27VkZQA
9XFdsh9lu8d9ti0uupI5Ipgv1JxhPNC/dam5gj7YK5mcA+LcyUATUZhGgUD/hJ0knnsLkTenR95W
2XnTjttWF6xP8NGU5aDh6MionaRfTfuKZLYKbEkTWzv9pM4QpkCM10bscArPR6bSE+WO1D5R2E5Z
JYJYfElGkZmFbNl2I9SS/HqxUNfdm0flISKFwvlq5JOUkRSMW3D/NHGnsUqsAqY3zoRtPxgJT7y3
ubPNYEqNlt5XwsvfdA+U7n30utAvCZoF4uWlOJVjC0nxmKjOuEeUN+FIzLAvQOXlkzij83Z2Ja0Z
E5qtis8mCLGFAK32eXZWygS97QAm7CZWLTK+kFYa/dQr6T9zq4PNYXU1rJNxXpn7zhjSr8xNNAKv
ff4dvi165Cf/+92DTdpqgR3am/C+5gCM6n/hdJ7/yp8gKtTZpniyLZvByHEoO1eK3J6zeuCwMWvr
+69Mj6f+oX2P0fWa0/im33g3Ei/Avfhbf277MH8RNWIdotr+433c/AiXSmfiPlMAoF4qJea2ynEf
FLy4HDgDuxucF/dfnZ9aMMe2oR88Zc7q9SuSoAhkX/0bbfeZXOP7eXw9dD4UEdDTAnk0DXXhVHEB
iUlXyfa9rHkSajGzi3fuX15QfHEs69rJqHRncwbZ1k3qCagLGUEn+GbudoHlKCQ86VJIO+k0QtKy
DUb9i4p5ofcS1wFosz6WU30Ld6lxu2lf0lw0ztX2Cjm85WK4x3yzdKbDaQnj6qEiCQnYoRZ+46Ao
SfqZ44Cecs9jzMm0dVqkhlR3PSDhodW6D4/2aKBZaeYuD5K2BuY3mNZ5q48XXpTlZ/dmNwqLXg1T
X8Alzt4tjj3njvumBh31VvObb8APp7KShK+hdmGAIz+Sc4sDKIHajQ4C8nnOgrgZ1RSimg5dQhAE
eODccJjD0aP0upDAKO/wG7LQalcunTvO3oe6kj/QA6r6WJQgOia5TKBQYvAtJcfnVkkKApBcno+H
MiNi8VInVzNlH6cVUU3ouoehfNKFVG1wC7ZI0hc3j+Y88I0puy5R82Nlhh+7Gf6lS44/III5Psz3
wGSAZk3/EFDDBniXeE6casOQoTC2T0pBdZ55yP4mUA9J5Dr6LVdTBokqZjmLcxVL7Gh8DUzKICYa
vATaEqQRjcPlKUiLjxCTf5y5a80vzJoBbBkMd8J1iy8ePfHVY0vzAYB/oJJk6tkHKa7hKcpOfVA5
kJ4+JuoyZZEnMieNk5JLe4Qi6wP+oj1ZBUaD3H4bjD+wosiNr3kapzLDw1k0uTu4bAX+61Ex9FJW
UmUoV1wgS3l/y6K/Kjh5teg27D6I1HqJtz8vhYczCcG/y4bB2lDWzGBv0NpOlkrxc/S/tDTxojHI
8og1Njdm2YNw5G8Al2p18xc022Z7KULbc4ljcJmHC1zCqlsCp/VsHTYo6uUajxnxmIFmHWzvLXVG
PQ+KwHvjF9wxBID8tHNo2PaHDQNVEQWlDMc9cSMcgSBPs9L5qaCfA4t36I0DK9CBUv0P6e1m23aS
/WsR4vehfx4UTsLp58kRLWADpcNgON103rmRC/B5dJtAQRRW3dwwUIO/KMIRW349fece3k3wRwi2
LXexbK93dgXkU5WIiA7vGtrCpvRjGCC4np8/2v1l5mRpNwB0HB/T55cyhTVI1xvqvGAGthgHjt0a
gm5aFkN9U+JtSZWb3Y8yPeZ2SrdeorX8bpCzuip2VPLWo3yZ5RTNrsrSUy+oRFTskxYwqtoZO3YG
75JTalyn4qOX+21cQlHLfiFT5Lg9/XrbOI2nkvfuxtePbbRxb5UjXCSPyNobLuexbrNvJ2ISSj37
FNXcfHsHLTYnsl/aNvt/6P9uWD4wkLKlorgA+gXPzerem/skjXum/zf3RTc/b9TupMWB2oDyViVv
T51C+t8uX2gE7y0mmwAL5oGvrGrHHK5jOMXgYK2+GO01ukVti5bnr86orRjFIBXztqJBSxPhgls5
P+vul0uUn6ccBUc8dwqw+Yi7WHjsHy1X4MmuxiFvGCFwhDw29lxs59mNkaSVt/AZZjhRO5hXOKHt
B4OkleqZeZpoSZcnTTJo+9AMSQHp1Gwe2r0KACLnuMQTy6xcFbBpn0NVPP1RgnzmilY0aJ0CUFZx
XFuH+izNQiwUXn1y1+i16P6l/dWOlshgbMaigJja+hnEPAnjrGJgqABwTBN+ZD8qMC7qv107V90D
p/ooTHrE5ulX4dlyXcACX67bzsT10+v1zyKkwneqLDilJndeDCT5/0JusfIEC9LU3bfUduoeOi+u
pJ+3Qr+8AQZZm2Ryy64/Z+w0MRM4Kv156X41fj/jef5ssRJ7r+okpMdx9p+uddxIXuS2J3JWLYPg
/ziNyQivQ1bSGu5Hw0PpjvJqVtwI4bB4qIGkOP7IDW8HUJneL1UpqZVsehJ3uihnHc8crMNUDEcF
wZXWDPkY1J91cUCIR1GBuW0THBTPEzDHejPfd04lLsk6fRw1NvtIN8RQNv6m/3XGfUM646kajuPR
fxsM69Q5OlK+xpQiACTkd/tNXiKdmPuL9TiBpy/0lnaWMCcjQ9vlAN7s7UcACQ5zaABWNk3vxau9
Is0bOnnqZKJ6WpIOvr5lQJ1pM7w3Dicw7tVa1pusz3g73dIREFlOlZyk2Z1bE7G2f2Kpm+9GJ8bt
APixitUNQRpQc/p9Ke1XkmPZdU3Gtjz9VhVoTiFWrkWDvsYHT/43BfeS26v1TsTd5Ihv9omnqAc9
Dm3RzUHUPyP1S0XdpMAbvj1vOWeTphzDosrgxd6GcsrE/pEE0H9kGaRwdr95ULocX/9g+J9ozF/p
CIYdyVHEpLj1OPIVTupMWhVuEJuDRa8eruFjVmZDJePpCC7uPTq4ndr8EdF2M70/P3Wsv4/bQGrn
Fy4AZILyVArHxiDyQ7SAwUC4IzloUScygx/2eIh7XDgHH1mZj1wIrgF8olf3jzKFJw5yH2fx24Pm
QcGF1Pw+d1IGzUhLYFKEDNS8F7NAoWaLqyDfCBV1fFbKyWiOMrrwjH/sxV2rYixdoawSgffdCvbp
hzoydqFiQCGZP0qLWDj2BrrAJHxE6zKzKVUpisPIOvRKeZqA4hnVlSeGpzf/n3hjtrJP9g4wBLfo
jxSl3PWKphcJVj7pFMQukjkjMuwg61yNZBv8VbxiKKdu2W38bG2KNnzGqEZ1t+zRIVgm96W00luJ
bzJP9h4zLKCuKBEF6dAdyMqD2oQfqRYVN4Jt+8yI6T8pesln58i2KVl/8xqsSCFhEwJxDWqHoqR7
ZzEWTjxZ65/vbtKEtME4EH2n7Bw0wLEVUjRNMpHpvpMha6eQTM7tkFLulmqE6lGhM81SexMl7K2U
gHPKTxqVRuYLzcyk/EwzCR8CdJbAiU/k6/UsjxWQd2gFC75wbymMi0B3snxg68Yhl91WkQuFgSqm
UTC9yky56wXUFTHeOZ2uiI41lSYYAfOFMWg1WgHzf9qTeMJ7xp+ytCtvVfd4HPnPNl4mTO2bMsWu
SpMVBrUDstZa7cdb/PZgKgFCz5uX87DGoqSW/ZO1tBNiXwSwY83Vo6tNjVFqFt3CdZdbqkZImiSa
HX5creMTLnyxdEOQ/j8PDwpquUkbOkmeeLRFJyu/X8PsMsGuUGB4hN5qOEcPj8hKNkfZHwyRDUfB
nBWlVaP8hJOBN6pS67I9GfOpQ3+/Xq5vZEzlv/VuEYNOlXdMI9xubFbUv/hf0Th/k/WwbpmVsKYu
tJG0hyQrz658XcGoz3mvT/tY+n78dyzG7kyoeNmGsu6yCTOJrlWcF1Pjgmd4njwV+1poYJfxObX/
DWeapr5YunMA699KwA4Qvf+baeM4hpRcUzZ+fKn/LU24Vlj+Su/K2teXCdU1U7geGmF0EghhWoTn
4dDpW7zGsMUcAVmxK672vlGWY/GdEtxfDCWoAIVoS0v9leFjupM3fngBhsDpKeibXt5ouOnV0Zpc
azy74wNGECKtNPDZ8GKP8DXRFKyp66P8BZLzIneoajJDHSG6XWFIAnenetHhHMgAEtW9kCuqXTgO
M/Uh7i060oeISvcwLswbGtrvsBOV0Eh7vQHArYK+HZ3LP786pHPbnXHotpmRmQhybRoe5zTeC9Pn
LYvdiCF2gcY4UDE1hd6DOXg/HmxsrTnGYRzA9CU8l9M/2htiHq3tjmoPa3pWNBY7k4hH8/vrOdNy
wIt2W8bHAYwfEYOM4qgSxk3aNuzVHB9+Jd/TedSvEfw1r3xpREWnxc0CuTuf2JpunnPQvqNwRXax
WWih4vWkuRd6cbW+t3QvuVGpBj0fmGIPINN5oCMI0JW4LTzwASkt+Nl4EXQefDCsUr2CjoF1U7SD
rr/RnCgmw8JYeTo45yoX3ktQJ/ZaLid4YUaFGAwY0nKm1SEH9Lz0j8Q28ZnvQaMW7HJBcxkGiTHc
rIHrXhGb2V3XVf4tGuFwIf4UJsIvKcYAIXMH4y7rNfpy/aby3XD01+4mOODevIG+K9kfrVK04KeH
m9JlaClirCcHoQGdMt3ScARNaGR/dN2wlD/zqyhypX2Ci0yv414p6PWaEqTziQdhYEGG2Hdpq0T3
ImxEkpi0TLUWYmVNFtG3CLju7JmLGui+UtyosUW1hzduSwz7m5gh3rIuRRY8F91uSzg7/rEM/ptf
LniEWJri9BXV1dPw8xuhcAG9+ec6aOkJk23mRpF7jzXME2T0g60nrRd7r8HCJDhnFnRdDD7BJn3k
4wg8h62URhvVQFbsL2qglcOx3hM0ACQo72NEk2BRkf2KR0etapwdkv1Rt5gKJSz5fzL/9R+A+S1l
f2eNIOWTThkr4E63amH8deNa0LlyoeRl86/4RSNTbNR5t6ggZh7PJqB5e+mX2iMg50PCLxQBAD14
B8xVt4Su265Y+0uZtuet7XsZN6RjNcWyhDURkKa0/bJYgHd48dvl0LXuwctwexLi/0aA8ZeegMG4
UwQ1lKaeAO6kFdGElLm1F92pMhSo77MTnIZWnOvXXi5K4gwVLgj/e1RYkAT1rJIEVc80xLjgTfyb
3aPwW6umqbvEG2vdu9T5yHjNxNpBXppBTWYvu8Mu5LkSSiw6LVwRStn0Yt9VMLA7lJgBiOXnrfZL
IsT/RJ87o2JV66gLWv7JH78PCKKKPp8E9tVItQzyePZ3jQ1OVxMxpBG8VXND/0j2vBNTDSH6c2/4
YqWr940eOj6Tqilgz+AQ/Z0+o6L+l7d3YQlMnRC68iv2hZ515hLboMNdQaWvK4Ay9K9rdzLrVns7
T9nbas33Aqz7NLTg1sdKf9oqmO/u/SJOGTn1JEGd7uWtKoRGIuRCfGmXXUHb/FqT80TwGP4e3ce8
fkgzEKaQqITTv8EzL2TuTDfiUmrXDgXUcaju3VW9g3Xp61W1UpfCDsFoYlKRYB/XyHHTlswhJLzN
5q8wuFTvmospLJQTZejbtIjIKfzRSgL+1T6QjjceufgHT869al7CG+0ToylbQZn1VVww3gR/nTw/
qBBddWbmnKsAyU/gvrSfOQur461kauMIolT0B8TGBwSWcCCTJFQ2rV7HW02T/2ZwaCdksQJL+IvA
tyBvYMLD4QFbESUg54a2nKsfZ0WyCEmj/5sRJZIyxykwyycHIq5tEIWVbF/5K+POvam3N9zCGi8Z
aGESqyg+aI6+oRBGfhFgHv8q5YDwHf2UbmC9G+7FyvMcQeD5sZnX0OPu9SkoUrHrmV5FPox/Y2md
x8VCkmwyVf11rN+1/wCe4dctjqzzTfYiPFPq0QQA6RyIZ5+ivBPk3t0G4IrQgrbv6GCRsdMi+F14
PfvmoRKBhk+g7jbJVTR07x7zI6ZIMV75b96yMpRYZ6F+AXM/Pgs6TEO0aXu08rx1AmsLwo0dSUzw
b2qXOjxEGbPlAvVTQ5vN/r3dnpsBFN9H2Hp40YLZmiNKHCDczgkA0yMmpCHXGRk/4ULuSRZPHbMp
PkwREquZLDj4Vyu4i2TRFkVUl9UOACG6F+P8mSEB550EJ5pj0LHtKJPOp6Q/aBBRRyCgJmq6eENo
NSwuZZRCPoAXxxNrhVTbuidxWb22f30KtCecn5jPgJiq7KhRyuwOpjyH5K7EXaaCg7kLsrQJNzff
KTBKXZAMcEQh038I+x0AfZTsYleOD+fdx1Q2kZjqObbBMDWuWIYM5M6uCVnHQBsl8QEuofEG2SaJ
GNWN8wEDgfSBaxkC7TioSskbvBYQ2Fe7sRgynd+h1SVcitw325vNiCTYtB3siSVoaNNmSAKv7dqC
HO6VSXhev5ag4KS9p2tTwkPCjxzquc5APqmkY5VD6F80KKYAor+HNeEj5pqD/vKaX6mv241D+Cq9
bJnacLNCr23O3/dNamvzPVpkhITOrEkfGv5vyXNITlCmV63TUchp3zNo8nem2k28H0v0oZ9OT2zW
2cKrazApBwDkXnSBoMAhQ/dmYilM3VoS7wAegW/jxBKE9OancOcVWgpRpcxFEUjS/fn1b/4vCka4
rCl6V2JEwnLufavnOxvNsfPHaJ14ankCdtqhWnJJtLwxtk59YsRiLCHS3WGybIEFVQP8dDXBoGjn
d+F9tDJCGz/7u5Vpe48leirxRYRH3IV/0xi+/tcuzQBYzpaAdrjHD/hCSr/DO+BM7xy3fbWu66se
/E8/3FYiOS6DNFVTf+/GHcsiBK/xu1w5ApEFyjLARnpzXghqxYJ2Ue6/zzq/N/Vzj1koa4FUKqCo
CG8SxK2PLKUtj9id8277FrSwrs1qQLaB+3vim0NPWjiz5f3h70O/fJGZXta3M2YWtK0h3PfsM7Nx
GM1MQybj5u1ty65DkoJLTho/pZnTV/ccVby+h+UNQH3mnV2gEASpTvqlPVNTvgDv2JKNCbsKoWOm
p+rkce0nBTAlyZnsu1m1RSXYaNA3RWqX5iRGBAQedu09B1xrtOoiEKUtTrkguGdSg2QQKyNWkcJq
4MD9mdrV8QK8ThFUl5IIehczFDVGmuHpMYhp2TnO8calxbFTB19tbFBIFoWJtg50dzpuRgKYUB+K
JHwFTuOixFFaoOendXdwZAUwDZIQvo3e/2EHJmmWONYry46n4tEvO02zE1CRIa/vHOh8OFZQGNVF
NdMWc700xBzcsUvSDaFYdCemFYIGFeSVlIunpjr0szd69SPCiJWE4w5e6QwYRRuoeMJf86yxCl40
orXn6emYNUQ5BxoTpNQ1ZVdBBpJRnloDWBrIzAfBMqXS8mflEjxeBFANmUbIl8fr4vcKYagtUH4Z
bjItRfxoNGMU8vCZD7LriyGpABFY+TeebfcsL+aJSF3gt6UIqAaw/Pjqr7kQIi9mesXg2dX2bnsP
F2zu5vSt3bkA+1tY3XfXQ+nan8LknipuHMcb4nDqIslpHBjSuEGu0wUlx91JS+OnqdqbZYAKywas
HEum/S+DzZUd7b6sU2rL7UbNVUhqAIYnCVhgVCzOugi/MN6WeBOZwUzHX3xgbi/ZXvpHzRXqUzUV
aXX1OOVhygngyEBYDeynfE/NuqKXjbirY5qr/mKrEgqT+y8HlZlYPbL2k0Oxs/XpgZoAfsNmAWhD
8wRa2i5XCDj1dRBysYxUsuV1c1uCdhKwJ2L28NS8IPyw9hcTflmT7UFoFyX+lGa1yZ44uu+8/zP9
a8OgzIbvPvjMKocaXt09jwrNkawqoPl+H9RsPtY9/d9AI9IRkdxGepVeLyLhA7PqvVsdytszgsd5
oc/eBv6LPOZMLXSjTCRvDyzBjX+m8frw8yFBjw5VuDc10y1IDz7wAWakSuMlNa2jYlIvJsDJXYlt
vtXLINCYe8lp+5nPSgUh5Xpmc1/quiBMdJvvsfSy+mNqD95hdbvPvm6KdWZ14JB0+XgaZr5ENPBZ
Ppq8P7ZyMEm91VnzEDPXnGDwg242l+8gq0+mVaAI/p/y5u3WddHE//dwihFIsCVuWXNFQdFXirte
mIKJaZBHapckvDWEoa9nf3HPMhmiO8LtWyrDwMSlzWCw1xP2KwjeQXqM9GbB4Qp1JPuk8QmvB6nO
riGhjWx7dcPSYfCI7/q2L+qx+4BgR4fZPwmZ0yIYWFc9S8OSiUvqW2HroteqMXO2bnuYPrZYTRro
MShgIYZPVpCfskaM9BAEjOPU5idU0r/ne1EBP2LYsnmReGN3hm6nkfOcsW0Ny3gXKQTQN9LO2/N1
w4kniTZNks0jLWzcxhawU0vsONg8Q03Rmn5G9oO2JDJDl1ejtjsIIE++obKiTLZfopH4ZJUpn8c3
bbLNH66CdgU9mkQrUCYNXISBVfbEYmupcwkOcQrYIv9q9gIP9DJFdac9ARfNV+t/K22w6Jdl/6aL
ar/wKKgG8bNgs/rwXiEL5vttxuPwVawXnryQVS5aoNmvROUxJK9VeFJpxi+ZbsKMtOwisaI25Xgh
BolNbNDHRj0FRs1t47rKhGOzeocVWmacYC/1XpDuNBA/KLGltFDzInKWMVS/UXRjLXzXrzWJ4tNB
0O7uJAobwRuVIS2r83/ZaiWmudzmlWZQdFIxmYb1xJkNLdyrrzQaF743RTmLaYtjq6r5wBjoKGUH
BUr8MSzzNjNcFIVL6O+p/VPfUsJ5ea+6ESABlz52i/fVaX+MB+/ruumvkSt3SN+8ktFBtKf62AY7
5pmB1Om+pmQeEFPEo+tPJe5vu3IM3sI+zpCsZc+12egUAjVa3bFr4MAH/l7BRltziUJOfab13Jx0
llawWoL8LYINsI4GZx+vRdVZsxk5FoIT/OIv5yLQUJgPJ3oEYNF7P0IZelzK7KBo27Zli9xzq2au
Behz6XFRdkqkCl5VeCIVg24rJbyeIRorM4c9FAUhQHQCaj/wCAU4xUeqqDt9AlT5Eaa7dnDP5kNT
7oNyi1WJt9R1TWcYOhD/M6FwIxvcKXfrnXLkF7pHtPlpuTLJEqAGrufa1yB8pLYB14eBMAq2n67H
N9PiV6d99wPNFdVF/HgxzmAcPBORfBWZpoDr3DtsEYblzPghM+krRaKz4fPnQObmmTXPK+EkfhtH
Glp6hTX/uIEdZVwLSFZuHJsjvu1KvsEKiYyOICVHt6aMAYnyBYrn+lNTtI+G1VgbruIreqWedUAH
sf4u4xtHyIYx9cw+JOHFcuuegzLjF3H/st41DnDkYc4hI/64N+UrJG36F1EYE56xE5RIFboNRyBK
daFAllSlKOD5BoXeonhQ1CsZ9YYK1t3RbTzrOcPTfPsPBGh/bfa8aRXp70A2u9MK3ueVLp0L1q7D
Am1dCiZ+9z4me8yl98UdEM/0JMQMquIc7lotmDAxSj0KPDXcpKMXbpMK0UNjGLYKoJV6TTZvjeNr
M8HXYEPql3L3IGXe3wgzOBWewf3pV8iSd89p2F7/UM3CSwu9vojh6OyEvS9iTsTPGSkB4AI/H9yS
r1ALC551nz0t0sb7y+f/NJ7hU8SZsOpAoRMvMIJ8oEA3b2CnbItBsM0fcGWj8bpELIxs7yPvaodj
M4AoWit88foFjNt2AbpgWMG+uQcYKPq/1bJG63z04X7SJptlQ199AmyrI9c8t4DRGSqcqIzEqHsM
OLo5eWDB+q6PfAeuFvoEsi7hJlKizfrlI0x39p/dQT2CJxn0mzIW20skKVV2n28bCMl6cGfi61Eo
Z1JefRmaJxD44idb2XcCGzNInUKb2WzEJZ1q1mFQFHGW+rZghakg0q+syq/2+VJzMhIxAhzxRY2b
ES1VUVlzntQCXarsyUhh5gRusGXuzws8hfmDkNTr3k/wG82zpKgkfxkABuVHQmKdyq328khE1Edz
JUNsiVVJ3s7hZXSgGSdrpI374iNMCmnrzcy32vAZiPsjovpPn9Az7OP9Wo4PTEJPRoyGAhFj0FWq
1aU8Cenh5Ocl9+HvUFNgrlj4JZmyqgYfnrIVfpDdkh/M2BPrd7x4bZDDd5Dnzau3ne1grIMKisVb
+IsNbwO9K/nRy2ri3PL+dqjNqOpMr/rYmAx+ZEhSWONyn76rQNst7XvV7hPERDz777FPVIFU/wdP
2yl/xetZ7nVWIH+t69Yjh+BJvnYXO8XEZTjX87uH1VMnDS/5Gtrm/hbjmH3wmTc313iQsoKGwqbC
9bDmUfwknU9kdWpvS7Ku7sCCqou8lXX5ljWF3GB1mJUUMBjPXmLHZO7EeZ3kCf6YK5COuz3EmFWI
ykL/ROcaH0K6ZxJyTusAsgNGYCKwsSdddNyapLnm36bLtvyvsMVq0hGHPGhApBKMFuzNLuhcIqEb
GNCtYQN396Df0msJtfoPobLUHfFxSeercjS6Uwba5JggZ/8DPPGfhrLTwoRzbeBtqlHchwIKJoCI
o9fswqAGlViSnj84TLhaFFMUpHyuZR7eq2816vC4UTxe8lmTGICqomWM6Ejkv/q8sLkytrroa8H1
OHfFw6w6LZSs0HqJ9g0adZLARmZnCnHgwd/96P6MYp5alplhZzdpBoF9W5c2bduZjxHoSRaI2Z2d
ODkxUqrSUBzyNn6yQJ8Y1YY/dGHDkrAPwdD0Gg9lg1zvX0/GWFXLykRVmQ6VmNrT4UP8VBEiIZgQ
HrCUVbk1362kGMPvq8otkTOZpbZAuZluxCGsS3JwqVZ1ZQv3Xc+6ze/0Ex7WiPx9JSBaRaR9DIDV
/etkJ8KBDl8VXVqbJhk1lmxc+7g4l70msTGlYv0tSxyANgL7yQHbHo1rm0XYqD4H/xlKUR3C+jbE
4Hr8avWi1gosOaoWrd6HmfufGdcMZbFjvvz+OPbjCBgiXwlqTf4dj62zvJre6OyUzXe2UDhDFd+O
CsL0LbdgKHUZg+rjgNvCJnzuKSUYVyLxjhcCmRHsSRc3ZWMUPgZm2lPMFbJRTEbMyeipr0FdFJVp
Doe5D4ge3of4h3XuS1bOY0VsCeb2YmayaiZrCzPRuWVQQ/HCxPpX45fPwbj2j70l8CKDdOYPiSDL
nMtf7t8mGPpXAs8584GrAg9JHP1o+gFf9GsZSOSA7FIVkDRd/Kw/pRuFIMX5F9wu2sn8MGUVYuM6
VaxILasM1nFMonzvzAwWkSy7TaLfFKS0x0kccd1jDDefHQpQkI0vbFnxhtdLv2QvpmzEGeDS0Use
p3Gh5wR5rOonHhgU22qNhJBZonHQbVFeV4gQtWiu4ZLh30JQb20eLLWulRw4QmBK80LvadylPU2y
2fuCiyR+cDouETOxq2d/0/AyRsZV1nW9RH9+Ooa2F5Nypju29dwmMCxfuZX+oao7+J/+51X5rXgj
WJRE/we19Wd+IONBp2boD3TmELypuwCO4uYiY79dah7IVJMKWwdJElDpf/CsZwrQpcEL0tsKP6S0
Zg1DBBPqsZbgb67vI/2gI74ubyL3mf1/5X5+yA1l+9XyYpW78qL3NbZ/mFlX4e/f1vCEPa8Nlukl
IMA2wnBxzVahoQ0yNP9ROeY831Vbc/twtFzSL0pxVvZzUatKt/ga1g+1BR8/+/bVW3sryre5GVAF
VX0PIO9q8mxi5ZH2/KdieBNnLYO47EkUe0alAy8aDrW68mPQnp/XgXZnBp0f459cu+OCqp4tf3bb
iMYIqYdOp9toujlxiwDBsAWol531nH+r7DSfo5ykzcr83J8J3CBoFf7750/wuz6VkzmYV+ppoEas
qOAy1gnApxUALBvboJw7BgrpKR59gr6joQgEjk32VOg6uPqpzaxV1nkdUGigRzFVNaN9zVIaGU+V
VtYcD9nlHdnE3ywUFQhtRZO8ge2cxrvB0v4zsAkDiOM239Lxv0N6EDY93zCYUtQW/Zm2+xpjtX3i
e2gkIZAjCaBBnfEFKBj34K75i5/aDSnC91P/+dinUf1Hdy2FnCgNfd42Pis7oFLXagnkXdMTAbKA
QoynDnqv/gm62ozfDtYeOS7VYX+7Jg9NMxX4LP5K/TPgwN/abhMi1wV7rxfeOHqLbgYJg2R22DsA
kFzpSZR5/1T8HABc9qDIhFvMRdBzSab+qqji/vk2310HXIYblCitNn1Crjp9AZPkAdT+0u3Ee1RF
0y+N/Eb1iS4zYiB7b/94+xOUj6uQPjVQgSG6guAoJMqwtIpLZkvislHWjaEr+EK45bXvIPPr/y3c
xFUw4koP8aZaAsLQNnU1smWmR57Z8s2Ri7kh7CQp9fVJMSp3Y1/Z1K16fe5/WlDoJkulKXxOVOAz
ubdKvA+4VRTadE0qxScxlHHyLgZU1qxjKYxS8FX7zTU5Nv6oDN+ltDFfvJPAgM8BYZyi/52BiOY8
krdawo6fkVTwl+7YgRaIzorKpUXLvmmkso94GWG0RElRhR2vMrXo7sKjidYKE07rReTrT3AzrGfV
5GoVThcsuIwNSPrRiMrT3QWFc23EvJJ3xmoRFQsDx2bb8j6gK7hYf5l5FgZMgmImiQyNxB71Oy74
ZkTgnsOsL9KR4sNQZtIu5BgyVkkEQgvMYn9zjVLFblM6wGA+Pt+yxbTj0ROQ8u2NG91oozI/Aa9v
LfqxPJpkCmYxKai4vjMzFIaU7RlSn0Z4GlGSzWEoMsOS/qjtq2Hvt2C5Rslf7P1cBVCLSUt/owZF
kWQ2CmXdrpmDefRvrHerWYtEGyidFkyAZ2GYO/ZQ8frJSsLRWpnJBrm0O9U2oN3vZWTVUrC5LE18
lTR3KXDYUVJWlNGgvjcQm/o+V487S/Bd1PnBEBme61B2VYIIqo2bKmQ4naN6S67inWP9e+h5ZTio
uFKyUeXcLwMwy7ePTk3zN10EZXK8PrqWIWHCLHvvArmsKF6LTVjLh7NLgfF4T1uHeR8i+dkzqHgR
q9+sw6amSrtlKYLS7qTGNTtZ1ay7/Pmbu35dleyAAdLBhZBraw4dkRxfLP1McR8MDj/URrDSetlb
7MhsjKxG81Zzg6mfXvjK2IE+hqlhOdGU8unh0MMAHwS9MNSFFMxfJeJohXcV4ozNbfbhIDVYf+sF
9ImO5BNZ7uj1l3PtQR204MubKHEhv29SRhJPSWYNbxEbxYiEPOr50gsp4jY9aCcddbOF8q/rCR7G
Gt4ec3jasrVFckJVA/sak8iCUmkeko0++WBKe+9GOb4jBBeLCf5GsCtsNOz+E1dVP3i0i6RSl4LY
7REHTRBiA12xuyz4AflVOIhPskt5+eFVutYHN1LtgNvmaa8Ngf31GS7T3pHROJvXY2lhmlu6gcwT
12+Q64gLxdBldvDKuhmUUT+Bb/9IVd74BP8Aq49mPFNUFLJq/esjnHk11GdUYgpY1e/hcsnrQOW1
9dRWVkJPahfOSA6KHrS3FS79E4kQxWFNYRu0iTxhjalQwedg3v8UrBByhIpuFudEjwO3O0weFHRP
HsRSnnWSjJOHBS9ynCja9uPZeXFi5iw3aVrZYH6OzgepWqqgzAYR8BYNNlCohii9kt+7uypfIlFn
9GDPOJuiifBMJm7z8rlWHNyP+q+HKXfyjC2Y+fZKgxLBdfXCXn+to8FmGZTXVwZU2gqSmf8e0xnd
DOvrzNskFMI46Iv2vi1HYPzVTdVuWX9N7L7RxciDUMBarZOKY6QbHr8bHujDNdpb5Fv9hc0kzajg
VqZ/VCvOuitRI5vaPzgMLEAv/mvTA/30uWk7s9hirNcjQCD5UVEGC5rqsfLciQZJyS0H3uFz+YPN
ScqXpB82pKscFtZew+OW0tOSQ7WaDaN6DCClFXe+y+hnDr1xkC4U5n58W+KHa/EHchb87iROZ8aZ
rl5Ad7MMr0d3mKC2jH7GI5b51yhZ0d70p3thXV6AOecT0NTQ5ebro753hnWqFcOyo45IeAZmZtfG
idesqgi3VUIBRU/BBn2Vmv+AFy9xFphryWugoRZDCnh/Emgj2R1CfQOaudAzoZ1FxuOH+1Ih6toI
c+QwFsNDFBUchnbBJPf+qBA+Qu8GlGsZeY6/uPrkaKd17vh8GZdMR4No32vf0g7Ly1DEW5icnInm
98dRyuX+SvcQfVhPXW68xONuDvUeoHjoDinY7ru5w800cbg6/yYeiWVN8sATnPLj7aMNGMjLcQkF
c3uNlDwkRp66HLyUdrP7+21jWuKnuW2NyMSPlIgHo24Kw76eyfv/HmTzrGxlBeKcF7ZgYAXFQ2tV
T8mhCBnVeCFUBbuS4whBF7aF3/axfl4iBAn+Ox6VcPDB4jBwfo3otRvE8s7z3QDnWjiSLfKzOpxy
NJG6Smt3d0OGLo69qCdOHEH0fttRvUnlW8uqqqm9IZNwZSLH5tjiIwQDudmJ9ibCf9w1tHw+aKPb
nkxG3LPEtqhhjrxySGEKy7kr6/chuHj1aqiNpVjhQ/p5bdCGfOmcxxATEFO2x21TrXJm/vGzPCvM
k5favX9RDUDQTHMyu9wYA575jqXRykY8sT7KAl3gMSu4DwA/F1S4hg4YjWqS6kW6qbbZQyE+jQOT
xPVe2g58WTT2IiMyX8divQJdW4me6iSt1NnOdb+bggj1HMqgwARcw10GzepZHPUdtG3jy0IOuxWZ
g8VVcXuKqTPS145tYzcv6Jo2ISt7kLd8MVRkxEZVTld5FZ5BJhyXtO1wiRG5dAZ7QcXR9s2Zk6Sp
RStrHG+W5/h1s7kAbsaYrde3oBUV/nQScd3hlgieX4LgvUMedF9BDupmebCqrwvpihrdSijraxUL
Ch4Rr8V/2mmZ9zmHGbtG9tMm93+q46CiaiB6GerXIhxMblPrgP0ETmWEfA+FxeqVPfIfBFzWpneA
XJre+4uiZse4WrXPbjtbKgFe7wlaJKkfFqaz89zl3nS2XMfdCsUu+yS3Px64QmSsKSXRVmso6oSh
wbGv6hUc0xPhRSliNvEJ4hn24dw2RKklTv0yfbrw488OdmKJbl1BTzqMHjhZkebeNcNdrial2PeY
Y41HrZU1X+upgVWvmmJOLUb4/ua52Zy+JMRMVUjNnoqrDGv8xBkYXQpU0AQRx2HfKguHgW03gEZh
OORnjCEucdZOtasxUULspaRAgi3QB6VfzPiSLYMvs0nuMc+yx5fkHsdyFyKAOL1sbjPp0XRK51sr
V1egm77pSLVbW4Gy/8OePHOOJLKvp8Q7UUQBfVZK2dgnpI7uggDgq7zFpvZDt4Nmao/AIPCuD4mx
HsiScZE8MtNjems854l5acue1G3M7aGGLkjA30qCSvFcx4Kc3OXHvdM87tlbDDqpGEQuKeZS04+u
cDwYoj0F1nvmI4g9rPbRTvk2L+ZpPm7xNizMEL+j1zvzezOkBVAnnqh5uK/SqFzLY5cR0B7qd90W
P0e5uLFNUjiV9YN3j+3ZKTwMk4fbgU46WQMjkIyof0MthK+309ph7xMTPT3UlAVZbsTu+gH768d6
XP1x+P3dGzzrt/CXr2uxU1WQbV/Vogf8QFHPhZOSmujQX8x0gbbpmw/M52e/AoSQMuHCpc/oijbW
I2B+mIGfmudssUdiUlwMAaOpvucxIA7WIhjLtVw/r2lsP+akn2DpPfs9YTUvG2xS3EGWcrHvDb6x
bGo7QgH3aM6m8YHKtWiwct6i3VGeGEMDMA9SvDWNLyZ1wS7qGTXnG0uI9eU5qQ7zQgRhihlco7kw
TbjhP3sWmR3P61u+ZamJrUaVNAqOCBJI1KtEF/IEsZEzPKcKkpvbqVH9s7gcWR5YcpSplxQgRSpB
c6rB7LaUGeSotT5gf2ee+jY/9xjlJRh005Q6fx42gjAmED+xNlWHFg2eycC8k2BhxpDB1k9RuF3o
ZZA+SZXdPWmY0hSK71X/ttt+uDLOmMU/N8NjTBXRnSwstBQaPCo5c7wiJMv76evbN+GT9za7gG3t
h9ysobmueJ8dbtlXQ12Iqk9rrkw0ibfPJ/u01YjABI//WZkOnNbedjTAP2RyQGhfA1ZnuZGMdwmF
hpS59uMu2/NVLbggGADq8DwuiZ8/lmp45hDmPOi3B97jnGMtI/oEVkSp+1atBw2b4Q7vSvQxOAJz
FOE3PkODHLmBQcudQUoeO0M0g85dwXFDoE6TEqsXfnwvMVRCnNg19Mw07pgQo6Yk+W8T/ZsxB/hK
M6DvKI/bIp9pqapji8IoOGxgoENgSlt5jSxEbWNtu/bFo96mi0H0SmNn8pphXW/p/chzbWpSIOxZ
RkABvsV+re1mHqtJdKT8aQm674SKpkTg50QB+sLp/ESQ7hvHLI7xCPZH99nuY2PttETCK3GR4yHZ
nq5YAQpapr7tlfrSByUu8OLiQZj8mznnuuSAZzG6nRFojT28qCg6EpQpPYuh+xF9e4m4BZMeVFhL
EnIx9bT1dMSb90OykQ8hnczLArymS5m4w6HrgY+SoazdHrbg0qkAFJAQ97Q5y8rPqGZinUwCivWl
hbFe9JfLq86Krs2QpBaPN6I5P70uY7VTOPzbP8gVwQtCyZp9q57Nauxkx8i3KtJGQcBeCNicvK8l
U5NBYJ4WjHba16wscLD6wfeua512zyQ4AstspoJyXEoFf1gSX6HFTjBbiYX6rxN9ea1vxmkqPHlV
Wb5eqqKnknl6T3woVm32JUZbbPXwZEdqRWNXBKqgsmJd+Vu8bKAvnXKKoR6NRzLsd1qiEH+Da82z
DeJyNt5XxNNVzgbcvDrjqnWWJL3eJ70Aw3mAuQctmKuhU8WblxxJfFHJLIZDFHgLtBD8ye4w8yCo
N1ChnWDVmhedDWxY76plgobyOXjM40LROYPBJQoKaP4KTJjQ/PBobOoFwgQCYdZnAGWwsv8A9GmR
vWbSXixKw7CqGIqHmHMkYWmNW0sXsgPzctnPbLm8G+ypohWal2h4STnSPMfBhiMrAjpGcj3aWK/s
lREPpyp2sqoRo2y5aVO/Elw8irlLuhk4PdPZBk96+jrNcgn6rqLV6mHY497HQjnWfcLMXrvnobxY
w4es4R6kzsukZyC3detH/tG+6Qr3F3UQUzI7y/+1yO0zgQiPiguza+PKgwex0INWjbaXnZt4k6Wz
PZT1WJxMhLgx7hzfx3cwr2IuRZAYWZHrC0ZYTvbkJA0LWCRKYM50nLqeyPY65KzuVz7YZ8UnjWHP
SSFkiBTSq37+B1NKxuvZhFsNvnV2Iu8ErK5STsHo7TRSU7y1jXqHhFtYbm75NjigG7TebunkcsA9
G0QTUhNAAJ/3l9h7knaneObWUIoKJiKLXEBkGMafCTJOtl1uKKn/ZxmOUipuXCFbq4e0rNjNo4KJ
pyI8Bsyb2Wj2UVDbpDUs18gkBgBLnxvzw9/ubbQjSSRXimqovkgpqmoUylcpTc7Wg7Bd7S+3oEQk
GnR4/p/tUhV4LvEziyAN7Xg3OwZXB8YAzX4luWtvaUnSeCqBojhNEg50drWqlO8i03Mg7A38fG1y
b+O8KbN0rzfUL31gao83GHSR3nR6lQqNAAgqt13VjJMCOiuaeO2E4D+W4VBdj284fgx2gq4UZp6x
CMStp/EIp8huPjFEPlJsjYFNZBTBB/95QxFkpNX6+y3Ez/xypod64+z4QYBL+9LgJqRtAbQdghy9
6JAb1GJU+SuqbQiaWMqWP+Czgii2nRqWQFzS1GDSe3+h/EYsH1nnkqnON1XLPc5sMSDo6oOv0vCv
x510Jd9EnlLSmZUov/Qq/iqksGFm4TJlv0rSX2LEgQE7A7HgojnyqY8sEpuoyBu2W1E9/tcM0wVo
d+bBqUbAUXiOi0HyCH/5yk7TmJcSyFNnBfMZXgKs/D1uwKVlZmLFs+1NOF+4ixbi3AiSE7kXfDZw
R+rw1zWgePvrQEkVsHUt5+kq77An4pMS6eqbp2NgQYx2TD+xEV3uCrmP25xeT8fwV0alvdxmhfBB
zRBcxne40h01EqpgttYFtzJ2P1UF8RQ2Y2WLpejuJn5lwH5qRNvQtdhj/5zwyNd1Ma4qlPTGFbnc
SaDo62wW6FulcWCDcgeTPI/Fgmwur0w+IBnah+iLqN0uW/JDRIw7cfhWsWeSTVRYvYpCz9Ak2Tqg
EKEN00fMkhNyDoNOrHtGNzbSFIc7wTPF9D5fAbYaag6Xw5dFAkWF5BRtThFBm+I9HxfpGkS3dB0L
46xsiU0Js0EUfM7LjDvyTPaoJXbzcycE3UGh0DGYi26ow1/wjrvga9dqIW5GpZugGl0Q9zdA8z8d
oBOcDS+wLG28T/olacgsxE8zOa432N95KcNMxfVUUGslhWyfhFg71bXud43GMkrSj+1trmGNnRIR
3nKsCvFTDxcupq4tm4kSMfO1YTglJ1nFakJ+jMdOsr/8WSnBDCyNMnU3/Ut/dHtJUZwIePRVbmk1
Ga+VTC66FFO+Kw0kv+lmTytgkazbLP38pr27TvLhbPpCqFFY9zlmOFDE6/EDdmOKZq4pDZg2Nfzy
1GNTqc3GUt4FyYqzspUcluEafccIIMJYjJclRMASK+ew8SQNm+TWlr1eYKdYKj4q4M9qFR+mhkwO
RAm1i58TjBqjnUcjBdoKuzn+Klraio9mPCQp4eUUITwW+hldGgYJk/eTFIiF1WXQTHS+ZuZb3yAS
CVFnLaDa2Hc8YS7oxQ3W8m0NW6PqBfQ0osHSISHyrNHoS0joIGPTEjvZlWUzYvgq06xQ0YbpEVH4
Xg9+IWpT1B2RTX3xsB2X2E8NA+g4bLoTNTANrclGptGvRrDCI5HuA+WM5gE108SZMwgMlIAglipS
7GPjOXUP58XkVai4O6fZuaBcsVZtRvmZBOHUY06aCn8aR21FvRGLEnqvW4nN6UvOXNKSLG+vxJAT
YKy6HX9ammAGezLCy8HybO8IBfvhEX2baaO4rlZ2zt1xg3EoYRWCr3JziCETG2FqxJaTIQoz+oBj
iBvDKOBjSeelQAeK+Bv/+caSpn8l1wrcpFbGIdoFV/gAdWE9oH01KlfDZAwOJDPBsRFsVwA6daDD
yU5Fo50oKum0Y/VZicvT9Tz/NX29b/pZLQozjYNbbWt2Tad3kfVqQ/xNXeCbSlWRNUsrqi2hgwIe
SEs79xieRWWSU9KsIKivRsbe72fHpiXSo/Jywf+mn9w3fNzrVIMKDzV92B2wVettorKvBYZ4fi++
DxUNTa9dM1OBzVKQN7rpYALXLZCATO1adwjsQu/1drrRwiliOyojqbb0tulOG8/QuZELrtm8tirG
CWS8ZtKO1L/ToVE7ldD3kAptwOvjqDrtkh4as9vy0RdZyE9D4/FTaVAf2sN4NnGFI/2bo4ArgwXG
7mp4Fl8ihr1BZfS7hYox9kKkkXL45cr7Wio+PL0kCW1SZnHDgvyEzNklT3nThrCf/HkITbMFIyNy
BazkCG1p2JYNqMiknPSTusLN8+5rgBMpDA4kipKPJY8PxUnRU1kzzwdJS8KvcY4Wyhuu7oI6mI8L
+cDuDyEgwZ4od0xPc4B3LxyFGlglzrncpKxfiSmm7IaeNZCWONtrxfc0VD9MRFqAptqpsVSXTBbE
Ah7BRlp9MjQI2VgdKjn2MROoyVZzqdlslqxG4DcWr+gZ6nQBiWqByzYdmZQa1pWNkTgkfzDgmFnu
/aPS+xjBOJrtORKmIg6lLSlIuKQqFyPEzLunX3I91JYc7fnBT9Igty/DLrETerf3UQ/Y2gFwDN1P
x6wggpHyGD0PNS5wDqgCm/xDSVGONqboIOOM1jWVr+6Y9YLWkHv70rb6cMMwPntZ1b9zpW0mO6cf
JsAmwJMkfJBsquRQ6I30mLlpHFxyNR/aQR19pH+FaEFI20sAMSojq8W2AFGUI+Ssx9/5B4fPUUp7
5Wdwg7s3PZ/hR7xZhbFhFXNFuTmOQrCz1bMgCqxPbSgA6jnjzBFL559v3wC/idW9cGOfNRPre87D
P1AJGvubZvzk8I0lLfF4p8HcQeDOKRdRqxxk6UpmitD8Q0tQHJ4L6fkwNY6V5Jsn7X7wBhUGjfmD
0HSbEmQYQy/LRFni2DaEHZCOMlirGaF72cuWizr2kTs7kFEDw0sca0UzV7wHVDR+Kea8lHl1e7QP
ItPlWg5oPcqi1GCHFe4Yh/Z+6kSlfzc1sBPfTotZq2Ic2OrtjU+jZrSEYZS+yKMyY21CeD2zJKdZ
cZphpffL/dmE1XiTcctL4RBdZlQSwP4K38fQ64eIvh1dUwoy2ZHyK0yIyFrL+bxQsJDOEMOR4RLP
JTv4AYVXJyrZD4LbMfJeByns6d0kygvFKZ6xs46zu09TxC3j3K296NEdh7iG78anBA6ncclMH2MG
XTbEDU3svF5RWuBQycGweFFqfSVKLVpA/xq4XvOoU3fmD9Do6D5fCZ61vN4DwtzcK5SnpJelMg4S
wj6u27c92OVC9kD+l9YmebSEVqMcjYA6Ul5LsEGn8hLdkKYhV6WIz3ZyiIEQrZv6++wOZvR9pXrj
SsGE1cor5D5/Ln6VtdDU13dp986VBua6xvtFbmR7utrta7tL8IcxDgivma8LcfyljvVmwTna092n
jIXpsm29Zp41nNsgKm6e/dPSbeUIDuO7y6FLWRXxdOcXsSFCk6vy2MYuJfyGT0DP9qV+RVUjKKLo
S7Gnlvy9A5GIKrsZvWNeeemGZhTlktyP1+/bqPM3clHYzM+cDYWYB2OkT84tv9vUIhy+exJbNSIT
IeOCka8ZJthA9GSAYV0T8fqPkZbGZCcqXHGE/9A8ydaDjjpWNSC4dwsT1wNM58qYl6S8Bo99yX8Z
Z9ARFPabBT1mDd8rBUA5ApqLR0SuGTic/vsT4xIHQb2l1ojMEy69tPnTBHCqpkGfvlRCFx4bhYII
y/3ora3c+us1J81e/oZBv3SruVg8pLti9lxE6KGSZCvZlzVn+TU/FvbEJxQWQhnjNPhTqZ9fZSS/
X/dud2iWkVnqELUkw8Tppr67Iztm80RYM3YeboiMiQlZrMYpUHqeTnJLI3egRWJt+lDyQsk49lsr
Vs0E8YxN8Tc2ZTN+15DBjkIVrKHoy+7omhlXDuKqID+uSZxV/T68kaaFB2e56ZldPvPxS66d7E0O
J1LwDUS2sQWnHtv4/KEybD+IiQUxeOATRY+YDHmmhWRUqOGFwel66PjpdHK/iO26L4NAPpTJhEzx
LUDPSAYzYOs5x9DFycD1iP5rlz2dY0TJULAsn35tMASuBdHoelkUkWViyGKBWvY7REuibTHSuMyb
lA/2zKlQ6RDk/2vBXipuw7pbB3o9UT7w2PNjHCXhfumUK5HErm3qTzJ4C3CENjqUgCAIM6nbGEUc
eH4D9s6sJbYl45G1b6dXtLt4fU9y++/4JVWMzEz7wGjR+w284bczttWug5IjxJ6e90JraWm8IjWD
SxorkxOQq++UR0ikDNdURlCP274+ymeQQOpDNNNcX16ep+1rDgINk8wAlY/M7oV/PqxTmYxJV4Ln
VnW8mJWoX3/jtssP7N+EhWifSUcCa8QlVG3HdrlrtO6km2QsxqjiTYhZpFR/7RBS/skCGcy23Vwg
PSkag5NEaPmiS/DMTBa5PGzWJrcUXoXSPmD/Q8ouFQn5Cz2nzo5SUa8JbaD4e1J57YzzXmZQ0wAy
pBuX4MSNt8cp+PgpfSDuyK1LLReBNpwGE4Kf1s1Yr+FMhI56WKoNH9OObKyYkl39QtSbYr/02Qsj
To0sCtYC2K7EBVG6CT4FbR+xtplnh3ZKQ4TCn7vZedhj45XQEYoNp541y8gBHioTKiDZFJ9FYL55
TreAuhaDgbSfZpNSd65Agn7vGjef+/PJbeNWYuJtKyzqPkeLohLnsmK4BnhAPwyYvmex1hr6lp8G
j5Qj+49cQInOGK75hCP5BjmkFE97i9WxRJ+ZH8NdFdgEvkGH96wvIi22IcDwXyC9wZCLY9jmSUJu
5D6ywpdc6kucDKX3Eklka+kkeB5i2NjQSNVkYEG/N3vdJNzk7RzDVKZ4wqjKe0r6jTiEFYAeFgyQ
rXgUq8Nw5mG2bFonYFOrBqfrmOgLD+FBcnxLlQM7nFk0RiValGzwZNKCHn+xrUucXwwq4TqjnJnc
d6AiWj0lr5OQopFqOSFj6tcK/v1GehCIKFbf1nIngfst0Q3CsFuqY7JH85iz3gzIJ4W0+ZL5ZrDW
hRBPH8zjtO4r1zmiZYjN6HViZ/37DGmm5kITJ7Tx4Ffr4baydd+xmiGvjdfo5is0j++3rB/iOCFU
anKUyjhC9NWWpNPrl9qASrPnj/DhN5i0C+VuNdlB4qe1v8RAAj7tb9Is/0Xm+WNY+3cffPa3Z6KM
y/Ku/jEgwjNTzbul4b9Vam2X6YuDAh+Smu8lYk+hQfDEFbGMOmpSMqIE9cujvABynrOTaLaKAcNp
NHt8KwjRte3A718RNL1LzTArJdDpuH9nArXirqcKKYBPnWamjqi0d55tZXfHVaeDpU1RF0/3gSv+
f0JAs7kQbhTCOXwPmFqm8clXHW/HGnFpt4Zf/pyT40DlPpt6/gu7RRJOTRSwjxRhM839UcazhtIx
t+2FfAMX9QYBJp91ZXHMIlUCHskbzsP4TeQGu1p05DsUiMidIUlKPOpxAQQhGavAK4Tk6fJLTTmW
nav0eUxCexHu/vEchXXY5MdcYUaZZaq5MMOQ08yKjRtfIZBVWBchY82CrUB3LQXqQEXPhMRfQkkP
z8KAXeHaLWhNERlcBdSyQh8y0w1kr0P9DVLEWVQ7/pHwoWID9O8ZKg+jBz5dqMWJYUOP/i3Jjbax
C+Lhgyjt8bx0eYrW/XJgIqxfpGwRqoaSv7jTI3VQrR5pdHvOwaru5QV2LkCt1O+m3ms3RCrqya+q
DYonEapEJdhBAFOLWT5vAb3Kxd9GQCjeD6rPTdtpS9282oOejWE82E/ETU5hmF6wtl6k1VIjuTTA
/kKQbnkA28wqewAp09zK/mQjPPOQcs1mrmxo4folJkEDkIuRoy73IOy9hOwh6q1lGGITiRH7AKfz
dxsn7OVwZgR0jwyPLSmLv67jT+NgSg7Ut8z8AjjCqSRKnLt7LPJDUO5oaClTO2u6rIA3Av2N8+Ub
eQcJZI2kKWUq5dDRYFHb3UbSO1wkrefMq+0J6dFXCFnaun+kqtanWkj4C492mROlm3mYrfeOQ85z
nZpOgeDhtlbZlTTOzhqhJjvk3iOPh+1iX+LLhYVbhEVvBatQ64VS+8e9ReiqISzhTj7aeOP4WY81
zT0RMR0D1lNgRO3zIy0zkCYCijsJ96T0juni4+NcdND695Uq2C86Q/aZju/0d2r/RTN32GINeamk
Gcmh4l1jpA5Xut95RzFjaHtTXQn22hxTnkPIsPnHwMuq8QcS6+PpT0pjQ4mes1G8pCd5lNWE1AyM
eNiB4CWuhKmNZfvnmORD0VQovuvyzzTQbdW4lve0wprho4ZUOvGakqqwbg+YPzak9I12qJjgs1of
dvFSNDviucRhu61eMPKI5SUfGani7FtHhQyLl/+nwAwr7QmQn4voVOhF6GVtkYDw6y1mSgQplMiu
ScA+PymNlKnUzbEtsHHYE6HU//S81rAc0WNdDvrz+K3EdUgNL0ncqrogmROclP5EYIRP3b7wr+LC
e5edfPPQDpGIdwOxZNL0iOKMpZkZRHN02JrjbDFQkt2MR53VjVXmFzPwzabm8RRGTfQSHwMWQ5qd
/aGDCICUzdWBCNZ9aNSNVTMDWvUtXI1WRmX489/WJV6kqiHztr8a5REHt6Lea0RcEIi0luKFpqiO
cPBQ+vNv16Lib7BrTX8/+Vc+45Ggps997dmeLi9QAzLJeNiu0Cubu1UdU7bBrTRlQEQEk6YnqLNp
BjA1BTflfP9BS2VKzh817IGAXA+J0g5WrQLG+6Hez61xRlkRI1JBiHZ7Zcs0lm6sbXO9vYD5neU8
dD81ZZcA1+MFh3F4hgXW6K1zxbsftMj2ZVxayHh/6UbrBw9YIlQCtfRZgJTT9BSElMms621/j676
IiVw9+Uh5zeBtEU3nJSYF61uN4etWxUd9SUYOXIOz0Rks4n6mspnpDa4EW99sSOncBR6dFwSRGP6
rmMiJiyNL/uU2jmjFwjjM9GfroqoD53CkWqXnZRm+fFeoDO3/kpdswBSkueFEish8ZSO50uVLkWA
JIkov7DO47g9HDG4NtBXsPd6HmxUKyxJNZ2LxiSvc+puypw3vbM2Y5bFMuHWDAcnlfFZUKFqwsRV
3A3NR34JzMxu42IuU1dGkEioQGvJIgeR+Mw6k9RrZyrEY9duSF+AZLtXKA/Rp/vDn0VVA6Mx9D8N
1f4HcJp+xu3Ff7YLBw+QbCsjcBiVlLkQDdQVq54Fcccs2GIJzWPfznMy8Jb8UIgYKNJHOj5VVra3
0skIVeYkmUCgPYdV5YTByWQ9JDh1S5PVzRXKEy7inZlOzoKjKy3GG+2ihNyA7mXHxZJwoG06JaI2
/G/JzIPs2lSOynaLqtv7SQ95jK0/dWETG67HU9U1Pn0FM08VklMc+m62liJWERdCcs3s0wvR5ROE
6ukNgkRIB9fxxtghRxS/MxnrB8qXVUzoquW0JwKE5/7qDFDKlz+S9DRSRdbLAYauD9YVbt9aEruJ
KAz8a825HcW2xInPRHKyT2hwckBZbnG1y4+ZcWHLsf924+ey5SdYgxgFr3qyyAW6LLA6lo5NdqUv
ds+SsAbco21wNlQ9pb2C5XjNAQv2SKolCc/qUcjN3Ftkf4MDxalGgvQQ5XqYlr217NYF7uj7OMGG
1/oZ7eKgoSGTV+mr33u/dvwVtK0chTENRbH96sk4HULyrxc6IUVYQ4v3ptu6zIUuo2LGhHxsPBZ/
fmEk0w8IKhpUqCXfxAE52WDlgR8Ow/iQkIyGGhSlixF+0vingFVPmf/HjaO4jiadHaGAD3OuKiij
ebWWZ99wvuu0s/K6La+V2G3QlQ7g86lyar8ciVw3EEWx9z6ctpzdDeYbPOft6Sn3Y6QgNwdp5wDk
a0uQ300GRpBzkESijA29wuPUh/4C7GPbHuZ9u5yW3BLPn4GFV9BFyaRibdHdytvu8gpRrSLQ3V8L
5RWiFpaUAjEnqRNerYh/A2v+y98zU8A6s5RzR71jhLBAxDBo2I8Mep0U0dQ5c4Fy4j4HOo2EYe2r
K7p4HVlkSEKXc7otnHkwV9mCK3QW0uPwos7aRFz52omzvzG4V8tLaCfMYHxjKbj0iyhRx3sAAShm
GFVwCS8TZogTL2k7jzvfz9lzvsIhMl0UNUNWnOpP/Os/1749izYW6f0/RPTIKiXnHBdeOlvUGYHr
bZf0IFOYK2ynjLbSVV0mYf/kd9eJj4ytcb+y0YA7sjcTe8KyjJULzeGpYO/ctzuEX3BLXamlOdIQ
19s+lKqnVtkMSwqef905aMuOlS/9aFAAd1fDX9jqzeFKKiAkKjI8mU0F2fCBEpliLW/3VKnuGbgB
mXVDgpcWhjP9gPLdVBKVyI9+Zv345JShRE1FmiR1JlYhJ9RyEZN5pIMgZidUdLHdk1eFJkg/bO1D
Ku5D7RuPuSBS1QvftTDAgF8nJPkCE/ArqdHLf9GUK3DuZt/5amLDPCbaf8l6l/xKEODK9h4qLSsO
ME+oMx3Cb0ImwH+YAv42Yfn4jBpTJx+cZJTZwRZJvsSdbvzPM1Gfb43d55sva2LgBgaXZlpV5VT4
Z2mMxeDSigUVYf3ZOAVzbxU3k1B28M+ePO/pkEeHdz2AC9utZz08b7o0Lc7P25DisJZoNxez8XU/
dmhKyxMKuwapjuIUNU5Knw8XFglCx6wqEQxzQahQh0tufOPyeJk47+nwSDF2a7nIPTTONGo1Kqb9
O+a5OybE0wD3L5FEfdbMjwhok1ZfKMl8J9Q7XZ5mdORwXAGaqAku3v0rYc8jVj81ez0CgZId219l
dcUnQX6e2FOCMJlay+olYugaHPhDVQsH04xH7rU9udVH2+/V6CwAyDjxAYRDM1gd0COeVGEkWLFm
NjXc/fcVkpg5uCT6XZMOGl0BcT9XpaFPrOPFf18w7Xanv9h/bNNGUlLVoF6LC6dIc+T7Yu1pf4MS
QrO2a1VtzTM0mjmS7He+ulNrtsTdqcwWr0h/X6Zrb8OuUGiuGwrhhOkmR+EVsD1Ww+yDT4jYVMAe
zzIWbWOBmRXYeynd+u2KlKOScSz/ZZRxc2NeIAXVwIJEUWbssL8wcU4Ocg4PjFX1GodeoTF82Dth
tH9vymxUBG7fLMjFLbSFYRKjE7WAW2zHz7fNVlfZUrMPzQ794rbPCe/p2VxAqe7+YGim191J2CmF
QdxAG0vT+Uoqb0RnKM+ufdsHLNU+wn+npApPyKOk61eeLpFlmFkd3UNkxS8ZfrKXBWAefD07zSCD
TJa4f2Te4NEeWTNWXbjG4JL9oriGH7f1uc/MdWoadJDcZS02FhIhGk62rlKsd3OMxEYc6rHQhW8Z
8KKy2EGSFbsAR/KNMnqNo1ROG9qnjUPP38IWPweIVVzOAbFiserAkj+vVPqPpFD8X/i9/KHZ93/p
hVWbA0yovjWwjYpYi1QEBtmYjdk07VaSPJADyMnukt+2V6LXSrV5qeBwTksvk10FJWYgFZ5OhsF6
LMTBMZmQV8SJbYvbmN7/HcXDtNgHSdgSDN+H6RXw8TOX9Y2YKwHhh5zXppPNvIuMLOLSdeyo1lX0
/dsuQhYDcTADe904d/Mj3d/ECVWzjnJyRH46GZ22J85mLG7MarJBU8VslSC3CLqpwabO7C30nwdK
H3O/UiK9FjTm/yXHSe7/pYJSeHAzWPxd/KMdZcz+BmTXr//x4GrtHg4jh1XlyZhl1q2dPle83QZK
kmceodkQWoujPAKhP8EKf2KOXggC26+7vc77LwQrf6/VypcFMRgTFx9PsDos+TZchV+/2uEQpg/R
Ji2gzfHdPqdN/98gvKS9alHS2y9p4YdB2TtVt4SR5wWQoA58lyFyVSztyUMp+D6qRSx/M9NdZK5l
n5WglnKSayqVpd/45PnTAdcqXlxUj2JgKbPgHSYIE8Ed1RUUw7KuRcutKs6LHdoiR8+AUW28k+ch
rxEHDqWJGCoDdEanW3Z0hoso2mbDYxQdJjstL4xH1L/VFxBV89yrlpNiT3eyiBk6JIbaYYaW4opj
V75MBxRl7u+4IXqhBPuebD9AAo8Zn/YPvsLCeQKclaC9iVWlaubeJJBvjsdgaYu2jhNvbB201Ad8
PB7qoJZucg9JrdBrD2rVfrB8o5kzn95uTnd3vsGn8ysv+BPQFBefqxf043vzgGYWO2RH6+pqop3c
6XWFrUbGbEWMf0V5ifVQjnIuzyGGmWC3MWY1tra8YOD3i6evo1DnahTE3VoJDG1mEnM/0QwId/0w
92yWtysjY5g7piSxGJ4Uq9+XMslRyn64XJLL+ePVMO6YkSdjEiZt6ds7nxI51ElPYkRFTcA2furc
SaFmrqsipVoXt/K7coBsabiky6Jo8nOBwcaHUUAqcPA1oAjnfDeIXvuWN46OSMC/oAD/wbrfHtOi
wQWDJlWUnK1vjrrhLHFBEWDRGm3t0GHZGZh0/55zwNnovlAT5mt5t69nnn1uMHUKnOChSv0vPF4x
2u1UkWH4p4gSarHHxH0Q+1LK5AQnu0Pjw9Tm8YzmexN1wlkFlWBEixPwGqx/MLalG4pJpGwfmDXP
QDcl5Mtheph93/oQPK6A0S8iXZQt9aS/lec2QWnbM4ermdt0b8gQ+Otqu2t8+nm5BnD0wr9adwtw
kEG18ClkLGnvHZeC5P+MGMvOMkEo6jZJZ/qtFrYve6Y8p2SGZkOXWQTgqj3i5ALPIDYHO5IK+MHr
SH4xzRqKIN6tcUyf/HwKqXzsjSGZ7yRMsAR0PNoY66fZNTvPbnXRrAy43tgs9FcVj5O3gHJDR9ly
SaaT1yMzj/oDG2s2y+sjDc2e+h66Lyix2UsAlWqpFsvckJR/wq6OPZsq2i6mODqX8L4BM+AjKSAD
MOHfVJ6ef27i8T+tultR6NgLP7skX4yEH4ViztGGgX2+j5AAps1m39tPG/c3cjcMl3C9hct4uZzD
BrSIevGFB6kX3wGo4pKoCCi8XhggAFkALBl455HegL/HsR7yPPdDC5yaQWTW7VmPq8Zb5HnOZ/DL
sD2tXMKCPnGdeq1L/Ng+IPMfNEtazHBIIxoV4KSu5LjJ+pBcJAkeBMmVS5UUXTakTpfcDh9THQ8x
Py0HO6UFX5sBS/niZlJ3MzeS8loU617B1CzPOtvlVIiBRFh+hRNE4q1F9yBZQ06k2HzNdBkIl+ZV
xFm9ab/7+5ZaeF0XGs+W69h6DLoD6ULppLLXuacnlxXp1H5SNE7Oen/kVeN1M2Auq+zm/IffliXg
fU9RZ0WTgZ9c/njCyC8q2COgZbt37g/OGSUgmo+zpaOE0VRPAKPfB+e1lbyCqbSKrRXSDTbxFQks
2H33+RHH02dBEnH1k3qeGHBP1R6Z5D1c3rHiOXODTXtugd+pAgxesS1PXz5GdRF6Qh0X+qJviDVo
HUbcLJw1/jrCCKqgbXl0/Un56wWMslhRz+h8cZyTSI5TULWIwK6qZTWosApDyXb9fHuei8t9DtBw
Q2DwWXDDO0QlO0mBseUMOkIA9xQAgbiHJr4KlrJuHRTYrBmPmx3d2tZzMtwiawvQF/dopyuqQ8LB
7xstZlFxDUBJMPnFipq0QNtwqP4mUdYIFCDjpxKRfGiVtt5ySMHGJNltqI94dUls8I6IvjPjf1UB
qaLWUYZ1VaOIf/SL6QdRFn8vbWH6cBYW2KgHP0y/xBUvduuPmeHjtsuEQWGRncBL5mIKVeseep+P
DlUdrfiRSiXKY1pRpp9yWiOCgLCE7e48Q/F0ULbPMP8WcE8OcOJAtiSQeTs3HbXW4+A60FlnnbG0
u5qpoxOViRMh0uQ55l6esyAvZ4Js5oH50fXH5HwbcXrvMosOm7BlF247GVy4HzOVpiZPJjRQxXT3
oajaFIWCM8dWDpaP0+H0wa5eT6Df4IKOGSF/mVotWjZcRwf5Ayd0RbuLmZLwOhYN+3RSx9/yLbzc
NPIpf2M68gKEUlm30Wx60y5e1icyAUvm2a1gdHohSWbH6S0DZUfJpl6seTsycSvDpV6gPScKKoQh
j8Qo4MJYb9QGALQR1vgHXJSG46HA+WA+CUw8yU4GoyJBYvoS5jV09OKDkIbLFNdXKVmTpjVXyRPg
44cN+qahjNwWaG6pOLKqNfPTDF+8bs3QMYc3HKEgKHAFoyyLeOKSFwLPy+OF8ptzY9+uIlCyoslM
uGenKrnkbdI47qdgQPQ3U9Wisi0fwe84d1YdlfKpy/Wpvzv2MrBiTtPpkDTTJQOBRS0xRtyn+8LP
+oKToKXd+k8S1VYhh+8Z0R0jO6EKgDQTEmrocuVRwlRY+4KH/GlZV/Bj1VTbxdFYz4a+0im22V8R
R0m9KHQRp3FepgXvx2XRyn/+W/leCgtMz3UCDTpb18PQ8m4S2hTpRcsC0RVDl7aBWrc3GRC7wLAc
Uhwbu2zOEl+O2fT5h3HMM60vn/Tg3EUZ0DLjUCknW7eb0tPKXdy0YAAWU9m4hyqNzbzy/yZjNX3L
XBDJjOKud/hSUL4tQAwmqQJtPs9slXaPreSMOMSa+/3a6Dbzv3ArokH0sdouO+asrJYUlHzT8kc/
hEoWEgERHGZBlwysotz33dn1avRqjWKOL76Sy0xnUm6JqybHOM8bF8A00m8m+Mgk8pnBBmhS+xJc
Ahgn4/G1f8CgIuAMAyp25REwsJgXcq4CUiooc6l9tFJKaTqMx1x3+mujwz34snDb04Hfqe0JsKuM
Ng61wkUvA/TfyVEqJGYpWDgzJeiyz9LL3yR8VgopVqkU+JuEDRB58mPghKf9Xtou4yLi/bRQE/Qp
qWjLS1ArjqmNAqSKtrVgXRlJON0SpD8SEfwRre1IXzVcZ1U5fO2DMfIKsV6SfCD/JhbBoJGUx9Im
O21goeYlCcGNlXXo9fPXHzDZk8PGvEmQ8hXJ+0rmXoQ6Vx41SyBV/NX3MYoSIqJT2K8OIaiJ/L7F
DjU7LD8UdwVyWBaoEPsdLlMtihf6eWfusdPm+KSr342L3eCztzTh33LnfCblMPu6RxClqcMUgrfq
7Lz7dBjjm45N5KJoaKTBdnSx4Sz2h52QFsRoXUDXiMuAuxBbYZF0c35jboo5WvhgBmz16HOYujV4
EgsZM2NZuSDQWlsYBUhVqqCc/5DVjyqQzu27/4bsYDqVgrS0SpIqjtWq9v7SzT8cTfckRVLSDaQJ
j+2LChEY+P7OCdMqFxO+kwwXZFXFeTG1cW1sDy/X5zvkrxZrgjDdyz18O5oASewjQ1MXs97lLJQi
GhKiJwFGp5XIzt+4w7ENOsBJ9NNl5CmGmpJaOnyXrpgZnBacIU4KOOH0vBGtdCLIyHVAfZ9RlDCO
EncUupplbYydn/3spjPaT4Qtdh5RWk7LbDAIYL0h4GgJdwhX7Ox0t2I3Zoa63QePLT+js0cbxRYy
7F5gj8BH3Zip9oQIs/KBcFiyy3GXMvjqTcjQK8C5/EnsXKGkwM/d5GJR3Qgd9mhcCDQJkLog1jh4
iHLyEk6VBCZhd0ytlqb8PDlLPvKGp6o/OAgWwfzHZEhI1w9meRqtpWCf9PlCzojtZq3AMrqgcEIK
d9aRyZmoRJqQzsqnpR3yj6mJ497SXwwUNKqYj/9tU8c20w2sFEpC0vr4wHQfCsgbQpgi179ZPYO7
2EjMWVKssQJVm5OL4hCcn5n/4ltjqQXJaObeQWMqRfanbGU1aofZ2d2yybDUiyNITEx4yZc51xxE
OnD6L+3x0LuoioYU7sI8352jOjLnl9xa21gntbFTEqSeZNTdIO26xpa4AIlwfgK0o37VcVXYOVfs
KOpu5X62DJkqsNgr+7pWGHAt8gRuGVUTUkL/M/Csdn3QAUNEIg1ito6b1kTJ6eUDaaSGyZa3y6Gd
IFFwi+EAER9gp+SLRIMAaBR1crqH3RzFWE/lgpcmb4RFyP5w9Wjrd5ypT3XSHbJmXS764oODTUgs
7/ShGWZYOHUBcZcdo25IV1+DXWbmT7hrtrk2LLa/5ym5YOVHeG6eSTKypLQaMaHCfKDmHT9vNs7Z
KcqQLBviLhzjy8JtLbFi8cA8Znc/Fd45+PZP3o1yqGoqkNNmoPh1wSQX0Wycqgm2GZndCIi+5qMK
u9Fvgw+lrjKlQf664TYDvdo9p6RDyh7bS48g4uFMmunCjy3J0dXVn7Fgjabw4Yasdk6dxKmDMNU5
aAkNpI/GaYeSwcPfxQktIEh4crbcQ6s5Jv+hbNvNMl217/m5Qf4H8gig0EIVorP49aZNLdBRSyWr
hGxxyUOY/bQo2bQ/qH0gZmD+hybQe9UD3IwCTb0xYS2z8HLIc36hALyMEFPnLCkpPGeeq0KoZvAF
cYcqCvbSFchDtXLMSUUN7JvF9nb6WzCkJs/npfj05pXQOzWOgSQTkD/CP9/Xi0t30y+ebiW/MS0f
jAbpaPpmEOF8jzBy4CxYm5cfoKeT4K8pPm8L3EJ/zYp9xMUFHoRy7mqo5i0XLWsscGxme0bkM+7g
fAmNR22RNv77ryqztmoQ5PC8cgmbaVHD9yPo0+6CwkG2WQDbMnzXb0XpTZg0FgriJ5YoUwlUlBQE
RPMExI4wIekFeTouDzabxFQH+J9oLDvX2d3/XH89Zxi3yZCnHUJqP8JvuT0JlqoWL3kOg/1WiuN5
47z50ncjNKslENMf08UOvr+OBq0fEyjRLW3b0PDQhMsl21Oq2Q77wyyF2bf8kA7wBm7b8/tB8aHH
PezDKFg9DdR/QewSlM6pbxCJmlSMrOlALNuGB3ujd5/VRvMzRmhTx79VdbAGiBpxLraZLeoI6Eyj
M69tGIHeATjf7loiNBnai03qfIApWbhRs5bsat18tl++CiuB2lQlfb6xm2fXSegG8WWQI4Ym5CKM
d4aRrlyonGkn0ShYLI95f825R2vcTHRnLaMJytp1QvjG82ZI37x8mIsj8T9Z21Ic9Y/gaCGUtKvF
c7YHHhIsqipA8Jg09eh0etsEZ+4V+JytZmEENZvyjRmFfxaj1ketsZuLY073Q3qdH5EIJ6NTAFmd
5ZYOrvArf4+sxpP/3kHcJpQpBNBuvwAEK1MnxSC48zDV783R4eGZdmizOVb883XnOVnOz5qLqY8m
gx0GQ6cZihnWDcxgQhUMxe6p8ZfS34Sj7BaGvt/dpF4zozJAmO1iq0IiobsAxw6KkiLcz4dCURuz
E5/Ahi2Lo0BFeWtWPTcUf6SeegNFPRL052vsfLv+IseQcpbIHIKs7Y+B0U0izuDWIuVuvO97M2t1
W8VpXhZa00rXj/2lMpjK+aEWbQgXB81m2r3Jb0Xtkh2vrdNDVM9/J3g/9XwCu0Pc/ps+evTYsSD0
DJ56hgXSXqe93ufeeMfyWsHcKbocwOfzbSml4Ee3p84ypWbG1G1ViuEwOHTE9qKIxyoDy0RY2F1l
OTSi+w/GcXs2htvOc4jMC3J+axQRWvEjvqkLyiXogD3Tw8qhJ9eQ7pEsWcn9ov6p1S2drLzOiVIz
O6D+O2mh5tmwzqU1c4qyJoFhHh9Q28sVJgjW3ZSA4JZGBwTS83jnUiCX8Zou8mqGm0oo1OkZ4HFl
kqQpXiIiyBDyUiwSOJ0+XPfTVwdOJFe/48HRI+N7KX8D7CnjXFYG4RvjLjWatKk0viLtSxPyrniB
PVpnxa1PXSG/N4cs6l57Z61nTLkjQLrec4E8RAk6ABmOKjkI6n4asxbGedfhRmv9KFQL2EVE+Ny5
Sbx5fZYl5zhzkb76drCsHA1zmnH21tJeNLMu70aypBsTlsPdX9WgNKVQaAiN1cf30qbHbmIEf3jK
wNKzPh1upGqLDfBE2C6Ku8Wb0x7c2/RDpwjcBIJ2R1aH1CGxrRBQj1UO09+bjvYkzFv/nAlW2dTy
spTaVCVPrkiMtSuo9SneYxySY27XIOiOIcaVjICEwOkFl17RcV5HbnfLXCFpCzH0CHMimJb2UmMf
L+Qp6JdkQ3V1rA27ojrJYJghhsqwl/Uy1K3m1OLFoLu35M7JTfPlz9p9yTZOlK+J0QZWEA6Yh+Y4
ojqfmvu1AC0FSy5wbI1G537eN+r68l9WsAyygU5euEnxDrdGhZHO0uAhql9Dvze9E7+AhV7+JqeG
BAZYC1wJIB3ifWUbxYtEYQlxKkZ2d8H8Nnh+aniwgHoq1k8WFwSXycEW4pCcfgiGFaXH5ttgdPix
oaN30Y7bp5jSLwMbEgO14aJnXKPKC4HUQI9aJzTnIxCkKi01i+cmgE04l32km1HQirryhLudfH6j
g4lJQDpR0laXn87Mwfm1n3QX0spduoJNIXB5N/Tu+LAkt/kjL5EFLKqYBUYPwO8wISqMBk1o44Kb
TaJ1wiQ36ENEq/K7ERFjRNOS74LPhQZ0Z2pM7OCSIdN6D7u43wUtGVl87wPNglSSAul8exuZ0NEK
Rgn+FYZQQEgMkrjf/X1TH+rHu4RFvaYg6PeCdeVieMfSvijW9JqceN5bFXb/RY7JFxRHfGFzT4Ea
fWxvHu49+YokHw58zux2HdAcvnDPLdw+jo7L43C5oej1ZV8KYOrtWaWsuGDW7sWvW+CcrUUom5Uu
555M7v64HA8hPh5fDwuBRMcWwZ1/M08S9uhaJdsstVZA7Mu6v08gtxq/arOpdWArl4hz6+OhktgD
rS8EOyrdzhXSoqfORm7fzCTdSAdFiNK7mce5ncVgjcw0xyRZOjcyfrDgINKVcqlwL07vDYCW3BU4
2xJmNl2YoIm6h2JLk7ylmcDvnIlFMYlLkioh5Tht4j9AK7zCSQPFX27iWpD/5amNQUJw8jKvu2Lk
2lX/0By91IKnvKe4/MqJ5rQHUKwRJDZfWG8loPCjGmR2E2rYmnHXnVEqCPLddloTvlHT+o3E3yaR
YpM1joE06xbu6wVc1jdSr/bunAf2DSnFZHlP3BpH/DXzcOZr7VClrbUx0u56sNY372t50cHy/JA1
+woG+gpOiBue5N5GGsNNYBjLQ2RZAoMypZrab2MYCdVmOxmkTAtF45Kr+QWq0TYYZRUk+Qq5tV3j
WhkOVhXikqyVzwjy21f93hjEjWyadQDfLqjmkSx3SWWh/ljWXTRAZKnShssvstIHHllkctqLZ3vl
qc/klAjc4OPToUF6z3AfsJrrTqhEDe0De9IOCbl4KKrEzsY4FWdfrUFMYCjrQr5RN1tZKsJEVKFd
mWQGsluEGR8kmQvyCIGMaKLyBQ+S/IdYvCzQE86aA4m2Mkh0l00nsBwd7pUJuP9mwq23miqCP2Q2
p0izb9gWdpLrZ3D6rmr2d5Lbu4M7oBtc1vPxYafWjzNsaaFioXD83ED6pG3MAr1sp/1FhatWkcoL
yKmawiiiNJHzRlBGUCX4wGB2C2uSMGKP7L0FhzXNQVL63pvZoYlPJkABHB4q83Kw5SXpRl+UWGYT
x3infiOGTb+sL91R6NKfGSDY5qmmOJbVLyO8SPtSSWVfRm9xM3ggQc0XYeRmLhdHUtOGouKDQeUN
0GQu0CoeQXqTjREnjlaUGuZSvcQeR9g+/fQm+ogdjgAGLrAsS3dhpdjskF3JshgZJXf/p3PoyRfK
1OS9iBOxoe2z7uYcuCvNvuhhMDNFV3tCwg8macsTTkWMiYYA75rlKEHlC6TLOKimrDFOp1PMxtpE
3q03D8bNvxwUWuqKDIq5qzo57RU0wp4qpZHhKUrnUaCm35y7jeSngBeyvLI8UlFUYW945y3aeui1
OC1uIUNaVoJseASKG/QLPAcQKXSZtytXpBw1M74XvSOoOYOAaLu/0DPaxoUGPxbNERLzy5Ypl1Gx
7S+cLnR7MB9tWNcB+vmSmzMG/eI+msLuNkG0XexR83AdXsAdBEFODEFG76MIczghuJDPZAxrddHf
PxmObPrQfiQykyq82JmNf/ghEZ9PWDhhSlMOEJtPjua4/C033E5OHOK8M1wgMH2YRQpZ2agKkUeL
TgFf7QaUtp0sq9xxcbiy8GW71z8UcIzaLnOWz/n6g4F5z6QwFX1rruGr2NETQUFyeyDiP2SynZNF
/imnpu9tHtSQ2N4cVhd+C4jw2EFzTO+i295Po8/lxIDTprJZU6ZaUg65IfBvENP+lJj3lP/rENDS
XZhxU1UjRvSyh9GQIWRC3icUVIFEPLhZPobmRaZfoxkFP7Q1KGmrmt4kcmETj00UJqjI9wH66AbF
aAqphFBkdljkLvsit/86yIPesFcx84WqeVtjlD5ULdlv/Z1GShRxbpmIuDmNjboRWvKVkvI/dkGO
KffUuQf5LVOp7ZGh
`protect end_protected
