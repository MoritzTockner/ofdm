-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
URRjo4bTnFW/lrfsdGH35H1PJNOHj8E49s6Lin+5rfrBb2LTuQURu11setPi7UqTONu+iVywT/1I
Je+DjjSj82rKoksrz4DxhKaKGD5cbdq5XE81JLFk+s3KkB7FVCQe4wPkq9tZ5G5JDfvvCF060mNO
6I4XKWZlPPpNJc3A1CuydLoY97xO2qrARshJE8ZIUizsA66/drmF50Wwd5ciX/1xVbdr2yWhLcAx
Pkwel+SR8UYY/sn8r+afGYrF1XpNjE+EAcOzHueyS8/oOUaiI57V3u9oZhi2+o/LXtfGW6m5xPMt
4DWeAPdt9MQn6D0IPry6mZ/UUa5Cnx1Jshikjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1056)
`protect data_block
W+nfILIIosn0XzqcHKij9D89IBfwAXcJPfj/5zyZcZPYhX2Ovx3IJtBvKW5/Ti79TWuuYhsAFGfd
vcAD41MpIPa6NHSB8TLrZZLsyYIK9BtfxKXxRxUHpslKkeqCAvm5+YaQP87oxBKG9f5qeGHa1yNQ
YMB6wDV/sllhz4+Nkuh2bC7+2TMrseM9O6pYpuXemjRRwpc5s8thtfg1WQAqx89l6ckgmg0KlguC
KWWnBzoSf5gnNPIWN2+VSNGZVyHPIuRQAeg78pO06roUE3KlT8UhAuZ5kCkPcaSrxboUoGn6PdzA
fpAqv85bQoj7KMDfyM5okW04P5NEwjUP+DjBs667+oE98T5/Y7XwgTBBYrMvlahAYw0JHrbic12R
C4bv7yC4tqVPZhma45vBG3fkievVuQaZH3pvx1wNkGss8n2yQgJzbgcAaUEmMMLvzwCVRwGcNw09
gIEltDrP5LL6ENrwK8J3dSmboi0L0wfS0o+xiFf54e1F7SdqajvuZJf18Nfsp27qmWUv1rh2z3M4
tZjtFGigDy9UD+9Bfa1adLPycl4TTPiiOR3D35P1hn9z1kdlagP4srDvKRH9iBr1JtVuzAEfNTVc
nVki1R/csdmnKT95Nw1v7mlDnEStpXmILraOQt89HsNTBYi48VxxFn9XtSNhCLUn0iJ4b43NFAlr
kUD4f6ZoK24B7g/0nsfq+wu1Uin45BdIoKJhUZTUErN1H/+HSdqR7YT3ufiymTjT9OipxNnVcReB
3XnfRHQxLMJKue5TEf3Css2pgjfgualO20JevK766YqDdJgvKG2Cob/CaY41ibXs2GV0EuLmYxfQ
EgkD27SbePnILSezJYyhIxYgO7i3PjA/d6txJdiiQXz6zNJ9nv3IX/sbcKET+xn8bLsK/f+4TQCr
LNva6DMBOKGmtLkNyx8P1A36dntzG4OCpI3wot9xTPgX52yg0KE/bgmzoqAcLHRR8m6zhc53KQ5X
aklGtcUC4QL5uUeuvK/4LCm2OgGIuxowr6Uey69QdoInVh1DEnXMPB+jrj6jdv8/7F5uQ0f8aYRB
2STox0ELR9bQ32nsy4JJ5rNL94aJfDnCNIvCOJKAkWkJmR/GStZKzSu8PYGh7g263unLC5481ZEZ
J94WQI0gxBJmg5kaepGGHWlYZTHHj+9UGnz3M6ccGGjJm2eIEogq+o7DIlSvjzhCL9TD0o7es/Ym
YT//MQ0xr9XrX6XxmX45Qs1wvAcJv0d6hb6MA4KYk8QvHDGGLR2imRdXGXARVUamNlGILy8bft4n
9BXiM3vZjavP9pmDrQT2Ucw5YY2+WRaHLD2Li/+rmE2VXnLn78Az8tuZfvqLXWBq9IWkOMnxvKY1
oN/m8dKUBK3p3WYpCkhszg/LwUcjHEKOHZ1iEEh2
`protect end_protected
