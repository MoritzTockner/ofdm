-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pYQPa79FFCx956yqNXZ7hksyANeUo3o5f9hGSP18KLVxpWNMXjMrTgOAPJzUISn7/5zJB3Kpg75+
7oaDsn44T8TLwug1N4UL6SOKpqcnkunkuz7yYxrzhf3MKMZDCQSiN9SJ0R4Sat1qM71JEv3W00Ct
2Q4RgiNDu6E0Ic19T5mvWXjz6/HjC/eeftzkYTevrXpASohO2EacGYzMbFDWvkJU0kabKS6UTiXI
USciWDi8PrRUxjXNLgAneQmo3Mp07EXiHA2/XcO3ry7ecTghHIWPqK9KABhS4OU7vqc/1fzgfshG
vZDrJuQcffJvl1H6qx+HlbehOJcrnJnimnB2yw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
foYV+h/ZQBtHk+y2mDO66ZH8hKxsV2GXtZpkTqVUsVHpJ2fapSerEp07lyJuKa8DAH/kcOs52Kah
llO3aEgtRblpW2gO+6/aY1lPMjoV2/9l2MhkNpUBDoUy8cw7rZKqFfRLAJWT6NiSA/ClK3FB5J0L
7hc4VrUqzSTsa6vl0BLC8p2LZRIqlAbCkoo/vNlv8YGPl/yrMLOb1j5GHbmei9qI7GI+mY7w5Xzu
E8/Sx/isStf/DzsYKkaqhyO9R/gRd9UtLVdLTDqrJI8fVYBKpLh/7fvy/aWDMvUPahSqAEIMjl2J
RbE206ePelG/ytJPrNSo1pcmXp0sNfYNU9Dm/F3YY/oFMkKt2S8CWaOLLm8928az0Dwq6uPyfN7H
U4XfohZpt7WLKDtwe9di4blPrwTwcuObuqifMKh1e0AJjtOFjwZjBY0HVNlJrxMxcLsSTFU16QE3
OvGSKw7DCWweByOZE0dD+AmD3+Ne7SaMf48uBxRAteLr29+EzL7uO1dhpIH1XgjQTW/yAK75rJbS
TAMVPYlQTfdEpNc3ii94aMmI/SMKVwzwdnFdTK5FVLJH6saFrnm+Cqk1pns7XN35MAKs8JPk18tA
fg+qJdJH5K+JVC6nZKx4kVLg0KItuRsOBgbU5MvQVWPWk2k5fcM9/lKENFuyaJBbJDXd4waBgoCn
KaxYuL7Lq8i7VpghKpEczUbjSkkWj4Dg/eNgie5UAPYDg7onyn66MFIiFbTypiukZ+RgR1ng5tPK
MqMJWlClnGdlPE7arnlKiOgcpJt3lMn0M73wGj7hr0anK5Zjs8Xd9tXTZRz1c7x0qR1ZPOjLpGlF
XXLU9jxsUKeSzkTqJPQJIsmpwjYM47vFNl13kN8idkqWG2BuPWnDDEdg9UubXC+ly1EtU+xTpRsC
iTWGRfrmjRtOgjz3X/pNv7E0AhpghQMx2PX2+C3iEPiLDGnr0qXOYH/oBZd/V3jft/M2TQ0RG1Mp
Q+PTkVUW2Nb9qu7cVB7rbRi+gAm7lZ7iX3ZsU2NkZvry0Pcy6l8yvzh2a3NkE7jV6iojHq2sH4ge
7pYNNex3Xaz3TvovZ1ZdOwHCX+aM9g/z9eh315Ec+Yvg4eLFsfctpqYoVAoTgqQdl5pu5IfCEv92
KEHH46MzbXBgh6bK1E7M6OsN06Z6LiFGjqpjd73XTEjtdaFSfnbjDDq2DgTzHr+x+UFCBOSem4CM
HRlQQ3D7ZGfKOuDz2MEqGrMe+X6laGsOEW+ZGX/jw53zb63otwENr3tZ7EktPfEuDGAY7dl6fI+T
2qjTNmpY1F5IFPzyIyF5xFEmAF34PSeggtSTB6J4YKZFWYdmHVrXJN+gDTxGzXMp3zVBtw+tXlr3
41qI7GbmUTBhts9bSd/20xoNZNiSqOZA+dOXZwacgvM54oMR/CKUNOqDMw79vJz4Ra2VmtSKsWv+
IcRjEmSWTw6QIYTr3ho6GU6X97uavVVnMnuPCQfDvHOPJyEAw9R3insb/ilGCkAHAba38PvNFWfh
JAgZwoBau661sm2SA5U33tmcTPyxNOqJTUIakqf49+AoIuF3SdrH82F6lJh+XxRYCB3LfybGf3s4
1+FGN+hQ3sRK27mDcFKQkOetN1MeGkkBZue+7pStczvW642CKDaDbcmJYCqf64mGrfUrWCoD3XDs
L3ogI8eqUmSFZB5wU26CejVLRg4r9Rf00hmW3SimVeKhmMOOIG5ap+PE1Yv0K8AQKFf5KhiSuEZg
LLZ0jIcP5EVV647W2GQu6+JAG6/7Mc+SpDIAdQiyHCGhV8bphFI4NkeMtXoEHJYATd+JTtsIMkF3
uwerr5VhTFKEeWGKIJ+g6sQek++eNTcOj2IjYh2mFZj/0Q03bcrL8kchNtikgS5cDwXh6f5khzuf
hqplHGe12xrjtII5fC9WU+pVy+tdAH/RgoNEAcToF1FAd4TS6EAiRlDVvUo2ZXHUvFBOFMmiUzlp
NA5PMejQmrBHITzd8pPHJv86PRPJme0s9Vz31A0Dffx2F4A2chAqsKxsLcJBRxAc4iJ7Ks+dMRAU
G828i1WHyleorIt/fsA/PsvyzOAmXsGZbGN/LxUmCHj3rxSeszQJjKLn1vn4+8xkLVyiqZXZj2IJ
C/NJzTnxmRmrAtdX+F8izKjX2gzqXDGZW/D1358F310GIUctx/HQ4dPpMyx+qdt8M/ynChr9sHg7
zZZhqACPSCM50oBJVpX7LJSgpeeVF2S2wPGwqcw11jHgpdEDXqQ/EGz4PcPfGxehB/VCaWtUrP50
svTWp7xKZgdbTWxEiNmVZdVl2hwBrn+mAYWw6V/HGSjusbFxA5wISOrNxwSj8urV2mO9P6waES6G
2E4FbyYyJ3Cm236+jGE1l/mSzknnIfYNh1QLRvaraffN0AU48IFDAHALsJ+GKzx7XU1mszLYEz2S
6F6sQn9sN2LpCil2OWxDgq5z4wIbngCV/L9ExJxtWfqjjTRJOUU+GnK+USWyFumThqgWh4ClQMpx
BCZS/tXfNNhUpFnkT/XLGtFcQhBWVpl2BfeqI39QRB1zXNhMUUGLBTw1gIuRAMUWuX6TfEcsuDsj
iIdbqTxm5VjRsREbY1mvFLu/s9JG7Gwprgv0oKTrg64R+wG0TyxipeVdiPIzBd8cgAJDgq8Potkp
1tf1iouWEr7W3WZgdB9SwhNizAjMhNjlbjueMdQtbKC1elSiP3a1WxiI2ZOYsc6P/GC0MP4L3Z2s
esU9F6JjBSHCOmACtpREc3L6DC8n4SOsT5ZEnxUBliVAOkH7UvoTvj8Cg6gvFgth+O7r4MbxaTpw
QzHM4RfCXTuwBpTar3H3tN5SD0l7KpgKSjzCL0Id52T3Y+Ar5u/MF0lZT5zjc1nm9iC1vBDJ6Ryp
ERMhm8SeaTmKC8STWIPF/Txr5yMPUEfo2ACMG2bR6A4lTKH+5D5Usre1CUrYaiopHuLydVt1+JtX
JCJVgXgOVpkPBLVeiNNL1aizHkift+/0XWuGh4tQOkks7EiQgIYXGHAn+qjd72Bel/N+kN2X604T
Y5tj5bgOyu+inlWNuHGNRpu32lHc4uPOxGo5BxlgUvpooqS8peyFFjo7rHBTUg4p3Qi6eXxIIg5X
SfIvOZEFvxQYUIbwjhEainjHLNIg533nyhxXztVTmblUOXZBOwMv7WNO0nuN00mRRtkyFxseUAr3
hVTk8cbNtqGYGCTnVt0HYtSh0yx+LIFcjVxRU01shgioLb2lCXDnmkjw0F0NWdMYebWQ+8jb/T5s
mEG0F37V8I89uYHGOIfZQpnYrOO68YOBNJDSCK0g8qKt5WHbtyhDgaux7LH3edijSl3T4rYdAs/e
iLqIF5fAP0NSjOMuLupfhh5n2Idgq0gCa7X4HurjlMi48XEjZYRZCyrvHN6mWpzPnfZ7GKSBy8gf
gbsMandBknpIgoBmYBZOnxwQGezzw3Qn+9B5iq2hnpgep7Dz5r24/4qEVLiBQLZ1owlWczAmxV+0
mE138fNEIJNL/ZjpenyMuoglD0Ghr3M6JKr6USqnQYACgxEZTl/W9ZkUASTqGu3Ax8aMuJ8kInka
Xw+es8RoqrwrZkiw+b+6ee6Kd2xcnvwYLp+LJJ9eFnUMBRVGJvAGYmqhbHOu3odNfLqzHT7Aj4fV
gT0UPyJj0FxvzWc+drE3+Fd98/+av3jN6Q5JH4i5g0K6UuSUwgCKB8om7N4BwOzY2e0EhA4ChCrT
0XaLhyX7Ava1T89TMMtOYJ2vQBT7QvPiqAjKR01/dGUHWhRD0k2phZvrSQ7BGmfmdpg0sdjlaz/8
KWQWUfBxeetklkJsn/3bKLt1VeJtlTPi802TeE9MFebyYPwAtZyZslAr+CZabg9gzBcQc6QhxWqu
o/NuOe00eto2vQytRtGWO5UAledVX8lYRFWwUHq2LVauyApW9/9BRRR5YhM5v7A/NffzK5SHKtIi
rG/DC5MU6WOi+IsvP+QFDIStTy/o8VU/YJuBSyTCeL4X7y6+OXDYSg9bueyD5u/sXf+Feh0JhEjW
B6hULZX3Ko7BoKd+tTmJiCkL5lGiHdTcx9WXAb4dKTPpiqC9v5YbLwpJGWj5GW0uVt/37OAQD0Ho
2HafGl1be0uTVDedFeM3cSqjQRw0pxLBAFDkTmP2oRFcQbXb3rbvJXtSrE59QlveC6EF7yUhLLnf
wCCJlXPokRVVZhTiUtKHXBjXU3GSzqNk1/fqiBoWIlM0yAqGB8fYTndAhRaOG5txwcG4Q8E2vQbv
spPISEy9QpXP88CvzSITPS+KSsiQGSbePaZt9JfEzw+CGyDAfLnQYluogDajB4/oS/K7uyYCOT7I
TQt0QHjqze6fj/syamPPSymOitlrkrUl7d+ffnyssxinHeXIbSdOOX+ePtp3221ELdzBiKMWSxfn
8Irspusp6CPR4bvoZw/etPfzYgUXuQAeMCvl5EvWuuLmzezdXYTlnRnoivq0SQsqYhaFcrwMS3gD
XEs1EaGSv7SasYgixYuaa+DzG4OyxsCOJRgxGymbrSaqE5eFdpU/2MkYIwjwasfdxXidmujzrrbB
QcuM5U2+NNbPeLd8y0+bjFAUOXl1nXFirzR6UKcP6ntREfUvnQ+atUE+imJRy0HZ5kcsU6ea1CbL
hXlwFi+V+0POM53YfvlH9spFTRCU25YX1Jy0SdTlOnE4dPzbvowSr2O7aJF+VAqUy8fWPI1B9LEx
q+apF19FdfRgMpRwZiq0FXtBHS3NFymyq7046r0pwGlfs+z7O3rc+U20T3DexclljT+Ne9thJ0Gi
5AMTqD1Uh0Ghlc+3YRJr/v/d4HXBLyxKoPO+VtAFSRp6BLa7IAQEJxfqQQ4O2ftUY6KhG3SM/myf
pqH8fKI0dsF2vsGj6Ei0KS4m3qrrCZWVsvZ7qeLptsAYy939V7Lif0Sdr/7a/VFMuD73QXvyZVCK
Sx/9FMSI0CZl65in9W8fK+Z6NB80hQpQRZjvNWpsvCsXeMeyXyCeDFdgMN3UMebO45r+SNj80ICY
5a0sL6c2RW1Az+0AYPsMoq1p7iEn8fZYqenXoKES1T8RmVhaBSX//vIfxdKxP+x7eCMaI9wgZoLl
0etQOoKI6zbjHz3nQLUCR6Iy4NKR6CESLvhU6e+uCLiR10nVQZZQHJCcRn9+DWylYtzr7npImIXT
CLH0rQCPmIb9iBntH4IAdTmL5kx/pA0/0flR6OV6cerXAAefvZttUwlmRNwNjSQiNMl6+N15RqCR
fqK1YYgyN8XbYmJKQnlSUy4oHqAiwa0dSZHnAaCsYWQhtjt7BpF+DAuLHVRxZO0/4rB70EuEc23S
AFFqGnd18Z6D0Fqwsu/SQXudDHf6MmADVIWriCdsAHKYaboNK3VovQWitv/C77g2/XFXE+rNroR8
RPGnGHS+KAUFP1Gd9KMesTCeK8BvSHAhsT9hdPHrh+4uVVPLxsB6z3GQtFPSdJNrHFvTkCAa6rzJ
j6QQIZ7n+hMw0dsDrVMy9bNsracHSB+z9qvpBLNl/9T4H5efcwKj5zVs5XLhRLhOCxk11JSEHe5t
YQ04AtSq3OGXBldGcVQN2LEL1LOKKPz7UXgGXA9ZOpVjwlxd6oxpH2pv5SPbGgS1MH8JFfsX1WzL
tSG08HmY1nY9EN8+a8RJIdXXID/2q/XVC6LXpTkHQ5uYprXmEcYRoTFT1Tm1mli7H8RC2t6FMWMZ
Qy7y9/YfKaAkNqLkqqpgN4aT5WTQr8VfeDfe2fdDNxHedDdI/0Xtp4KhOHSUoBzYl5j7evcfYVhp
qjC8eb0CxSfYGCuVlciZWpe2+ongpZR815dde0x/8A8+msHpHWRiVYpiJsngnAKNWkFqxrJzICSb
GBGsTdS7bOuU8ZLQqlbrThH1bXLuGIfsFxaYB6DW+pNpUGMB4aKxNk27BwvGEZlFbrmfAsM7gGnA
cseNYSkKcEj1vIKexs6Y2I6eHXYctd3IYFuexc7Deb1Kd+UvvRoi9tlKl2Ahb/2Ey+B58kxIJxwT
XP7bevDLKzshl32qtZUoET3iez6M60zun0PI0yviUgvRTfe+T1EQfhUCjjneIOm1MMCQD3pqlVkH
Nx0J0rWuZxV7Gc1jhtgTlMuso5v5Ls2azI4la9pYj5i8GDnpJWM4l9+WOKO+IexUNg0d1g8AHLrz
TEdAFAe1takJ2wQWALtD6RVNGQ5/MblCY9tyHlOO/YVjpZYdrNv71MQ76x/zQD2uojIMSx5yCNO7
FKyPvgmhUHAhOZDh+JbzSkdelk7iLhVt31QuU8zdOw95Nn3hNAXnK1OfdDPCk5f9sOyY6C0XDJMQ
bkExW5T8f83Yf9N3ZA0tTJ5ihFWYZVvXgz4t+GWXo0fmxejj4WO6YU1LxUmFcZhKyjbg6ic9IzdL
m4Dldd0TEu1kdqRAHmkm1Xp448RLuu07Pmq7+4Vn+VyRopu4nFrnRxCGRMM+auFRVqheiQauPugp
jRY8tIlFIzithk7YKQ4pAlyPgiuPRfTexgG4gt+e2UzVSCzmCQnZN3iOL81N6h8CJkUJduNJavNt
WIxU/e5RZDvZJ8vPIszohnfUA4UFK6HdQfOm8IXmrlEbag2M4zA5FOxlv418kY6WCxeKD+X4jb40
FzTRH1M3vHRoIGHgxpqLiqVEKiI3yqFmkIYGSeSpKuTYb5bq4+Ea0+FeEsSPLb6VSb8Xt4VwYxYX
uRcKG8obn5Ds2v8rhRZqp7J0b0TVPevVe1TY2UlxRgyhYswBYihZXHnkYGML+1jpIuD8zoqyO7GH
q2oQS6PVpkhKoSDWbWzYJjaN9Q4tV9lJ+rIyOsnoEqLHNj1opeJTxNdrjhiOuSoWJtkVEk1Xcf29
o2XA1GwwgyOFwONmYLuqEdWxREkk77hRCai0X3eTFYmF/HvN3VvUfgjVH/BtnPTSYZlzFMmYuRmf
g/HftMGLwsLNIbt5xyiVZ6gVHIbJFC/mWL1/oVZ17Q/jOmbKj6/av1iTe5tP1437JQDeMjO8s+4Y
ZU0r/+nAewjZk07x6hCSVwkNK+zDhigLGoP+w7V0Nq7ICpuaSY0bofx5erwUrd+E15MK54FLsjdW
LVB85+/go8+x/kTyBDQfzxv77EsMwU82UKWqWF1iLgAFc2155sBoJfZkfA67R/owYrSuCQqaQN+M
b7wUGGskOdvTPoM+tYJ1DBDj3bsFQinVtyG/8vNKEY+68EaTG6qwsf1S3HYVcuqDSmqZOILic5u4
sHlIxwkUyoyl3KKQ84jvKMxTdzsKcUsD7aSADJms9RqZV3dACEYU+KdPAx0oN/9TZEfhQiXCwphF
y4R//wf9HDbPswQOoyzj48+ghbdBBiFmHvHlw9kuKxttLjV13vMWhBpp3qIR5T19qiUlm1/W7pAV
YMglIYrYTNkv5fYb/NVZittpRkJW5oatlZKv24deVi+s24tqpP9HTbkxhxIJYlULUtWAiCmXROvy
+Isg7ygXncqjiRpqhkKt/WwieYjkpank8jDjCMPnATZ+4DZ7tgXTYWZ6hSDpEWuId/WF9mGz5n1W
KzqsUMJdHOmCrAfzqxstH+eM4t9XO+zLweyxRmzHM2TX5RfLmM2cXaBQo+/uHv9y0kUgFAaM8RZh
sku61GLRs5IjeRyMPNHI8+NTvYaSp7Ez6GY2CNygdrv03d4tz3BWyR9usq04O894TFXP07e3xbZP
vXavF79GAW1HGeaTDTcI1aMzNUmZYj8FG1QTSwsXdbVrxiF6A8zqB0ZQLVt0fXcJFUliBneovzDT
GVm6BK3KWoPo7sGr7QCplOdo1bn8pZHXfLObRj54vqgECF2czv464kFlYd8MsGLHdlyUIbUjE36+
7+fYwVF/B7clzzloFRqXfOyUQHdhySG5dU0sydUsfzfxceV+FlUrj/QavvBVh+8rdXAsbn/fMLWu
TJL2FQzvG2WSuKZATn1yn2f0SedJ9x3+R+Unixm493vn565I7h8BGuEXyR1repXRhiGjxA0e/8Z/
Yx5ZGHn3UIj6b5ZxwYkwau6roeYvYNE5DlZ4OCSJ79FCq/P4U18/nQAYdDNGvprpFHjcO+QI5qtk
S+dkTk5LcADf9Ll/Jx0XfAjHL4AkAnJ/aPFGoEqvctWpJ6taydikYNRcgEYs0+ApEqqDFfiUK9si
SOY0CeMgWFi2BvYKSWn6gXMH35q6GWIpFO6UsqnIxiJ9PVdMofUi1AVQESF/QMn8glPyPJ1oeDgA
i/q0hYfJ1kmbeI9hBi61dD27bDU0qE8yoE7V0MYef6u7kcfPpdkUkAaxKHceSkkqGxk5Cv1E5CK2
XM4rZH0ye59Ab4r0xHDNvku6HpoZi0CKUJ8QjXIQRiVdwwWkp8gXbEK3ODGbOffvo/qMtzBGKb4c
IPzE1N1eszwN5acC4Y6jvQluRUF1hzGG0MM1ZrS5mCDq3fz7mYn8DdswUwMPKYOZDFtGLv9bqZ2q
G3WHfQZ0LCMkwc2NL1eWpC5KI453vqRHp0MUaccCBIHxCMcbC8OuO4afLleHX0JHMOJAepYnEp6Y
NU38bzaWej9rrnRPESTauDamS22vVvUum1g+KO68xp1gMHBctG0TMuZAU2Xf6St5MTM8VTKT3BTQ
3T/T+jDjwfnAubSskksC4yZcVBAPMvQzpYGtvNCpE2CIp+5W0BwT1JNSEuCIk4OGYavC1GrMsJ1L
5ZVsmTK+r4YYhDzdCBvsE2fKdUmfSYhdCymuuPvaqUYZNOvAYpBCSkXTB9xgZM712fDvBDXPEpnc
QSlwQI0LSal9cWU32qd5fFKvbf9DdPXzWis2CFdfhFqylp9WEqhV0x/NoYMgk/W73Lvd/XS9wn8J
FfJzI5Tn0AZCNKrHFfdLCbvSemN3pYWrWAzADF0bIPNe/I9Naniu8S8PVeLjYHYjjOgubizwsAlI
oMXUH6Vm5E6JZ2nrjs1IahtfmJn2/nfFuA1ZVPKTeBHFablFvMPwRYNX1JY4m1kNsmrf0P7n5ggi
wKK8TUMbC5v4lNsICUsVofr3Y1Twt6L0IJaFizWpwZUgR+P0GEoa58gSWSM+chpiUZ4tKHWCJsHM
QNkzKf4iIZ62ZDfynXVEoSARSu4s5Rk4NtDC6NpZ5Na+VV5KMNhuPq01f/fa+hkOnqmdoKhnJa+i
mp8eL3iH9BH8W38DvsjZLXvGraS1jWaNcfnti2Fh2+UGWeSusWtjMISeQndLQrmDK4QsZxiNXI4C
f9VlZoNucQjOfHnOOF00NU44qGXaTnfq6y5SjB6hefrLANmzkq8Xfdckw3tK7284reovGnMCnYI5
N9Uvzf9ndGBlMA/9BA87YLT9Xj4VM0CQ+184zPsj2N7lwJQ9JMANGMurjHj4/TwwgB8Biml0BugI
DHTrOGGOhfb0aUWZQcZfWDoUSI9bTUJpIZZ9c5TJ7PiSp7R0WTdQq/VCM5sY+ewKylnMFf/yb/Tj
QPbFiwZXSfj3taqcoVnWFV62TY2Lrq4M5CDTRgpLm5R8Brwt5F10e5jOhRhWOE3WYbZxIEqGCBKM
LGEYu8a/HkwGEc3cuPcKUiazy6ubVuRsz6V7Tx0HyO3bJb4FSnQbiWle1gjdvQeGk7viyv59G8gy
MDSylC7HjbIW1FSWpix2Ju3YpnoCvUsCSaxoh6bCjsx9BHZDax8MQct47U2nLcNjc9Acm3dLGY2Z
DKKkhftEgDbsjf81ZMzZhI97gfhwT7pmMEETtn8/C160XC2R52skDLh+pzu5slq4UpB8JvbZINSw
xbA8xdgNFCd0bTFzoc4nU8TVdjtSmFaZ4GS4HGG7bCpblah5/lLeA6prydGwQXC7LkDeFagX0dDF
UWxX0+d919Xd94aEppkam9kWSMcj6wPOO05V45wbAm9AbZt47yVzlFq82K5rj7/ZEAQ1ApNkjvR+
undqZaIriyaBJ24cbnI2vhQOMBqjVWYcKuS6QVz/tjatp0x0GSGuWpWTiUK5P+5z1Mxn/aUCIkA5
2uV237pqStNCfcI5ReE68/rHc6nYPJzhFFnk86I5Azs/3jzdquolGaBSDFkNk7hRgcIPfBc55/h0
a1eCqk+iKy/Y4Kt4qRRBHKj+uVtGbl+nlJPcMVW2OQoIqMwVTjIqwVRL9fVDmdXypUCpCJCQBnKl
Qf6GPvU73w1geaCE9WYG/I2xSc4KDMjU6upxt/VKs4tYl15573O909TSjY9CJe+ailkD9+DPufeP
2MSQjeH3unamvZSo6/6wtBSvvV+YqfT4alr3ZQMG5JD4LZ2xzmf/Zb7LVuFKgWabahdTU1lUB6OJ
TA1Ng/GAi8HUzcpefQmrmFFOrZkJM4HhCbR2CtS/IgV5pSQQm6dcQEuKi/7zeSgZrEA9c6U6Zk6F
nlQmPm3RCO6KjMkHayBa5xIhC+Iat8WeeI3wrxqmnTscetYljOfgdhFn+RD+gwwgWJujse2gg2z5
wE9n6X+ZgB3SHOlESBHuc2hELcijBr3hHtKIHvUgYIPa/gQESXQXVf24DINCxGtHiVXd1wDHFEmy
MGM+Y75sB7vaZ4IZnBIeZnWBiF8AuuWQKedjRbmLd2HAn7az6jK5AVOCmga4qRbfD8I1IQcIAntG
pJO6QMxDfEsDjVXKrnbIZnpYJBaLAxB1jnzbQ1b9LtSn7RQBI0ERGIxElghCen6xjbndyhD7jXIB
T0SigrdzRhWUbrt4kogXIOLnF7WqFSuH1g8pckoqAh6NJ3ZnEW/+Cbrm9m+rTmN4tW4Z0mTG8Au1
2iOxIvpIquhleq14f/5Drm+zlfAVGyxRCnABuV8loUXJ41jGtgl/stqzUYeWB8ndk0a85gr0lTDW
e0fRhevkdHglUdktaKsyhAU1db2v/gHjfMoq0L75gXiEwfK2ko1CspQsPWS3D62RaMAato3hGAJl
SUZddPZE+B3Kj1bZQuavYdpKdjTFxIpBQ6WqL1CXZ86ho/tfqebZHRhv6cwoziwCur4CuOq5WjfL
2QmwSM08YZhbVM0K9ZU3+TecBR+3FGRcPnk9xEyBs6O5XXpmnADZcnkyeNSwutVPw0XfSrq5jZDf
s5P2+DBZogiZiN7hX+1AX1QQBrS5MgJZJRpG5JmkJ3W9X7g+kcB/kGipoN4/ovxLE7KEWUYvt40e
zbx+Gu4hnuE9IdUVhuj27i1Xy/ab5I0rQdnE9V7z8+r7Sn1QqRjAeIrDRF20azD1l3fA5Pt+wsBU
h01mYySHg3dHxpaPjNhISZLboP3yjAsGVDKXTFL1unJHPxNUKl5OlTGhYxSVJpvqmSlB1FzI9FEz
HTZcETX0PygCxwroF13iZWAVEplkz6jqKPvZfSzHN7MFGDgOkTOEh4xwO3uLHmU9v7D1GKt+DX/z
1ss/my1b7jc7WS0KzXfI4FbNOavdo8fO/KrUN4uO9O9Nwm0SS1cjtm56pHdiykwt3w0KLaLA9Jkp
rY9yfUnSdiUvCaEnE3mfK+rs7jIJI6A6x45uY64DRIQKuKpr0INg8i5SzAVRei2OwbSeI2SQZ8Rh
0E3+vZ3swpiTK/oTywTtGel+zE780d0k+S6Nq1c9k/RNoW4HcbgBD6uqs31SWdD2/hjY9fPywtu0
mDMiPn+ZQLbHwHkKCDFwomDSrLtrg+/XrIsdU7wREjmPWd3lFqeBv3QCbCnNCwBPMelHlOc5slwF
rdNCPa3M5DBZGJ5wuhBc6elvsN+FKf/umdFK+kb/Hzljn5Kv7FaTRbcuzBqAHEJVVPYX3kCaoNJN
L4osupz4Gxh5xLq8RkOk5CyMwvtJbognlYN4NYHIoJ29swXGEg4E9sGqsYExoIr3Vvj+yTzigzmo
OTr3Sf+GoxH2OJAwHkz6Dmge5h4B8u/s6d39hHDAGEqd6nFF94G/ES/Xt1y0
`protect end_protected
