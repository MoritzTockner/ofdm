-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
J1Zm3HX+GU4Qzw/wvaPSf74xxkcSCvIh8UksF+u9gJ+grrdfGDy2xXy9i0eiL5taxLREFQYLF4zb
xw8d0Ib2WlMTCwUsl11OZibWyL0xjVD0is8FDgImavSosiBFSgr5Oz7DVOdoXBMJbDzLqBkS0ZmZ
rNg9K0enhMoFRj1Hu+QGT9kvtGo4+Ubqr9lh6bk39WuOB5TUZHBT5msqtir0f5x4sClU6gDnJlER
U0otb9IbmvPJxitt1OpgyrRvX2mGGFYZOCind7vYzsEm96/UyGFSdfngcDSNTpymcmCIw8eUWS49
8qQrXqfiK5YsRm9lg/8TNYhKfw6KsFYUh/f4QA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
vh4Ckr4FkMz+AaDNqgujh4M8xnIuDBeIyDm+a8DdrgMgqQxwujY0IdJNjgIir7d0clwSRGgkQyXD
FxVeJJL7vz+gGtBJcsNYP/tUVK4xEBEhsfZXtPoSzrXjVPmVu0TDdveuda+v9567bdJqEnU3vYLz
fC8vCR1/fGEV5u/BWb5YO9pVOI5uzqxi3TcSyHx6L70Juf2kBCsI0klIyqd7u3/wFp1LFNm+Kizh
eTzQQActT6SIoVxpwD2yQTi4e4P+PZuMPxOOcWzytm1q+9eS1aye8mfhuZ7nDEM2IZ99JtHpm7vG
nvMDbdyNeHquea//oRIi2Un7Q84gRpiISOoiQm9SMolmdRAqQ65kc+xQyCeeXrpQ/6ia8zgmYTLy
Orfln12gDe8Xs30GcWJPlgytWmmYa2I8S3gRlJ44kZ5HQXttsjNSqZbC56/irYPNgQv6lXnQP4AI
0F3KsAICFP1g1aROHTt4HKp0EJNrGKWBsHLxJu/Ls6b6LHGhUUpmvv8y4jwxSIGocsD2UleUfj7A
Eg/4zgZycnB0lGr3YN40SK/507SL6lM8bD1sAle+wxqtKb2PhihKMXKlO6rpS2Fr6CgydCX3poGw
Hz7CAuIW13xFYPZP1hF8vCLEktQl7UFkQtX2HIlgt+W1lHFyhvM7SP2jcdIunYxijkPcQtVcMoSE
XxghVETmr1+TAGszpO29PR+8FWGqaK/Tfagq2sCoFTjdbD3Z4bIVKtJUI3Cvuviqoh6+K84GTWB5
nE1oZyxXVb3+LrUkkvtELv+3ck3r5XVIBdW7AqwXAzgqXMAnn+0XsM/PdTVmpmBy4w1FWHwQAqXk
aMt2zNVFWNBafu9FPqGnAv9zpnhd2ZiJbzbb0+jVbvsK3n76altDKYj/mFr7DOdSJaYG0lBrV0eO
uKAzySkddzrPSvaLli43NjniFKOcvQA4LtlTk6c0MuSuSz9b2Uqz+ljjXgSMqMDztvj9ZTrrAGP1
dQT8SeYevYEhZm4LIiZJsJDfdW5DuaNr+6jKZsRYHBo10gcZ+bgo5/SaJzLu/hUoed9pxgHMfabk
SAc6PuN7H1+opnM8BWAuOWCPkCpnX5hYnYxNgTQUrXj9fxFELwpmG9Z4y1lfFjk/NHHhUxqc/0lG
7eHzyhvvk8F34pr90EJPJeRai/EGy/d1TjYe8aLMSdEUN468v1kAmySkx/tGxGO5T5+cTomkIJDz
h5v6PC4/GTxbqUkaGNAV0wHHWGdXK4k2E5RpBRj8tFWKDe+34qJt8n++quGkSThCQQKLdX2r07cG
oY68DkNkHOoXMsbN6M+VTujb0OtDfr2yYOKnUjiwKn0EujZjrhtERRRBrZCLJXF7D3ZDrreDYetY
GuNWNfVzuPY5MZGrAfNIus1Arzt2sjAdY16upl7czzsePdiG6RmBbd9X1idKlxQavq6iptAeJE5F
8CTBBFagq97FoGA2maiLQxVYV+S5Q0J9H3SQQRaVajoV3CvxXzkozx2JPyKW7mJ53RTGlRoR4PVw
OQHI3OerfjISvhaZ01lQAEdOlziyEM7YxGkOrlpbAf4BBdTAy1xu8xdqnn5hM5zoeBN1WC3PeXIo
YwMtVsyrrTYAIVR3B3c8o1q+MhTHJIF+rh9Ypc8DDuErck8UYux6BT6382xUmxBadSDZfFXZiZfB
w8cTew6HIeSsOpzaQFv/Ah0qWgO6/SfuZM2pIHMX3c2oM3kTSOS5oW6sTqcMOBZD9zpUHWNw5Gvg
Q/8CkjfC/mRUNFurDHj8XCuymjWeAdH+wdxH9S7rAcA/BAI2w/sl2r8aA/JRWQQCTtlbDrzHz08X
r4DAJjn/97sqIQYobkhmUgmIzjMSyxVNmo4UMNV0UzbftmKyEFQmhFpp5JoH218xnMSAJDUZQoH3
Hz0T96svwwhA/tAXIXV4ddpWvx+V0E6oWv7YwqC1tmhZvAdjfAd9G+LW7xiP5NPWEAevYV00oeA4
DeOppaLyoC7S/k3vHpInc+WerAlQ43ZVymXEShl6rytk4I/nHmU6EHgk7KV5bMZlopADttdVrC6/
8MZl1EJ0Axeu93pHcVVxrnfeJGaNX7Y4G3B0MkNzlRor0y1aFj1nobYYKQFYmVlZPxDtgZ+o6gDW
GtsAEpgVejOF1eiAoF75QOIXBGquf7ECN21dWTmT7MzH2nXbkviHubRNcHISrr+/TPWOHErTSYO1
ybEWyFPMVvo9dPALPClYKwd0mn0LL9/k0D3KyvVLWXwtc4YxFTbnryQT4LKAehi2g1bWQr7P2A3l
uy52tPTVBLeu50JaySHR6NKf6IJzRGY4wPfD1hpoLVkMZ8Vyor8LirGFD0F8L2DynuGI8PQzklPr
oKmXz1FP8Z1PJhPq+aUSRQsuWMN4iHkD2qgXVCvOO3d2Zl65N/9D0d98Pv+9PxyhmnsxKMSQ8+Jp
VXuHFJAjlyg2KNB44LTbBev/muInuROR+sYhM8rkFgZ2J4AqIdl6+GVAh3tMpP4c0UYuWCBm1DWb
OGWxRnK1vWJO2fZjk20dSW/RyoGHXNdagI7ALG8wbx+TI8UQFc5AJg37LUUT/MXBwzB6AuuC04Oz
JFzu3MYJyFewaUz6AM1sk9XIQLSBGn/SjGLoXImL+SI8S2voNyd3ioA4KDP4hBxb9hJbIIOf7LVf
IyUNorcGex9ZsSmrxfYhvIWPyfeXFfQJh8oebL2klbeWesGsnH9L/7eKKjzu/U5Am1R34tDecL4q
VXe238GO0SOt1YkEwdRrKCzrE2t6+3hYGb4Xr720ZibIVbQoAeikx7wPOyCr4Bw21hrHNEPxHQ3C
hAH1n0Q64oAa4ANVz8XQ3+kYdmtyewtXyT+8zNof+SeU7tdj0lBM1eJW801gKopcD0w8bMuFGDlX
vc89KGcDNuUbkxa1neWS0QEL78HOuUt7k6DFz66L5qz9QpQLeIdqoBpYxpBideDSmkE1oWv1+zYK
IwdClQ4QdfdtpwmyS2deUH/e7FnYsA+0Lsoicx7cfpa6K9WK59PyWi6719P04XPdAnZkV2KIuPLg
UC2peIyk91wPRZQelUPUZSGetBoh+AvguIkGJd+crUeK4t8v5CKKvEKA0BSnUd0EUQbzLD9hAMom
ebI97ot1dDSjwFQystW/YbfKMkmWG9fBQRMpog/KEO9wENvyA25jyxBfcln6ehzit3WOYF+w9Y/l
xGAoYGKZPT1zpUIos2WmjeYUqAtbjO5Oow1j8JnboTpNGCLr56xSKQF6zuHFTjx8NA3Db9QamqnU
0Bdhf1elZXg8i3pLpm+Fo/YCwlXnVKnP6CZGbSET9N/U2yg5EavRG5T5uyXW3EcMC1Lqogu/Kxnw
TAf0JSjmBSrb4he6i67vvcTSXdmuKeA2BBWfYP3DqUrnaqkXriJd2F6EBEH4XkFIpyD70Nhe5ypW
hebNzIY/J7vFScuxOhWyUID52yQzVpMj5VpTHmbiFJCnaEfJ2NMZY4KiP6Ulu4R2BtjvpXOiQTUc
u41AcrmX4G416lv22z1UU86Qo9t9qf+WK6wj/kvUJC00XvjkGG0GsNV+43ormiT2EFoluNBo7Pyr
Qsnw71fMgpurymkJBRCJlJjTYxvp4Np1O6Jrs1H/7j4yAAdNpdWx43gVS8UQD4s39QSjsb2fPCGt
Qi5tfd1xkTBHVFE2UQVIqkTemuBNyc4vPlLReMzdj0E+LF/m447///9JklaT1+Dc93voAt3Bng3T
i5FX+8KhVx+/VX6oNcaal03a/5ksx9gI7PFbHLElMsjg8iSqU7qS4m1ncnlaDMeQRvh6L+a99hif
ORAAmhNZKAgZ/XVUUJ3qmzBtwCBs2Dm82tyzkzl3SvbDW8UYDgrspkzUvreU5NeXWOtSd/70Ghdc
KW3g03YPtNruu+kT5z0l799Qeg3MUS6/J/hF8We+N0dQFoZ8kzlGTaMLUzcABd4UzgvP3nw8G/g5
nNAwYqoxIdRfj/u2RtoBDGfno1ahNNJjJnp6h482eFWuabVCHmQPXvH0V9aMtUDoycQy2wP62Ol2
5Nip45FopXsome7/xHHBZpQJoD/+sE7tExxX2sPslkuweixNybZAEPzQlT9F2sp+f6hrI3SndNiH
nWEAU4jNlxxpsmV4fKqrk9AQ/6Wo4+BrizBmmrPWpBb9mEKmn6eqXXHvGkW/pDlEihVd51CkAfmb
iklw82iy6pLJF6kAcekRb8ZV0kSfw+uu6110TcfpWPSj8nm5YiRaQ/bs4FvXWP9L0jIp2gd2+2Jh
x4UY00sADV8LxQaNd74ZwXp67+TsAUKPnFqlEbISFAJCgFsHqDG1ksu2NW+NiN6fuvpdcD63bIAS
+V8Oi6tb8rdTVj/P3MyZWIw1+VVWybvRL9F/PJihXjOEag8L2jeBUIezfzY4RUFZR4w5ib09U6lI
QUJHegNb8dHmEBMMF/HRptB1jFywlks/6pPG/6ScJMjPe2lWPeyeY418mhtrMPHPUXzcBmHl3IA3
yiClWL369NCObEqagNMhd/PMo9cfdGhCKcnQvLNm9BtbZARMv1kzAdZZBr28UG6M54M7UlhEa3a2
qzc1/HfVvlxyIcP1fnnEuX8hK6gTyCxxCLdMl8BK3CdAKxIdOSNXeoCfWSF9PASI4HvsOvE6T8Jt
aA/S7R69PR08fUyuXw2naudwpywBndt2Z7gwAPGsAbe1McrrbEkBJ2fJELTrLh5Uimy5wo/H844j
VFEX/pn23zuFSdF/Mp99ldCqvR/7lwRSjn55k3qJ1iHIhn8DCHKGJFSo0FOJJoBJ6igz319ar0Bx
vVykIRezn33dhC44rtC31u/OIWme/c7oDjYUppG6VULVj89IWhhwhA8ATzLuCau4KrZu0CikcLWb
WFW4td/YXRlLXJ9+AXSuehBXWEqKHrGoLo2oM+Cwl3uXxL6jAHDY9EjoMOYnfnm8PhGMwL4bntrp
wqYDmOq7RsRbi/dUGUIT4Hm6lT8CiuFnGdNGJnFibITjcayXOW9xsbRAThGWwU0Y3giU4tnX0j41
bGjrvJ9qIzfJ8yhVAr5FVsQaKAYqgKDhMrq4Q1YxAw0XBRCBBTDqzOvvdK6umYvFfOJg+YSy4tBg
K1nGl01NBfEByNI7+/eTGm3z7j/0U/uBXMK2blwk2J8RLZuziNVHUk3fE454KUs0BqtjD5iRaRV8
dzTRnrFxDVwFl/axTRMeThbgttZnMU+6WSqs8QH+yF2ApgXBqkDAkWDI3LQe1rO3QUQri/WGqovi
xWPEVzA9+XTdWa9aavzkLEsxoIrLEaCmUxlr+E8KNYXGYcLouq9LpOT0QzAYMvfaijAAD6NnEkaA
73ikV+tDicwgTNJcFXGUegF+P/EPFoa4UFITmNDDTe7bjTD91BgOqPZrEVLGfWHs4kDD5sj01m5s
s0e5dBoXqajH31A2qi9BrsL/Gd58hTFYsTEjzDhR2wJEwRHg95Wju9cxiq9tnyB0AcDMb8U6yozn
960vOlP/fY5NecQnk66SOEqE9u03nuLYCK89YelXMm5jgbE5fB3UMN6IzGYDvQyOv5YT0LhbtJJZ
Bk93mYAUsmmJcBsNJ+JDC2MKSEdKiEhuHH8Gi7zI+aEQt9U/THl8+gTmiYirwmeGvc77nHKkhT3J
icwAq12NiufLPZGmvZ+Fpue6+s8g4tSrNcKpyzdFV8VkYLSWB+R2nB+wK2PoWztr7IyY7TJQ+zv3
ya1mfKLzRuQFHkNds1S0SeSiheLHyGHP99i7BZXkfeCZ4AhemqrMc6IAkx0ts0irv/RWQ2gA8FKI
QSona6IVS0o2BKjl6cSIduL0e9w2TpJUKQSupRSgsiIUJITA53p+Q52DU8e+MMNzBt4z8N1YnnKh
TYS6HEplxU1WTE4cYjG30zdveajFwhlDGNsCR5RGcKWqXyKzXSkOuWBuVKWIYaiGgvpGa6vO1Ys3
NAsVvFPLAWIpSiS3lK8dn194l7O43Rmn5jcRj2v9YyXHFvqCezSbyGoYp8cbvHqDgVzRT3OsqH47
ue3yx4AJVFovfTndi2iAarkw7lXxUxpDPw9rYez0G4nGxlgVQEc2/SOU5ZDwW9bj5+FuqFcC4+Xe
6nPXEXbpbo7mfHEIbZSfbYRcDT9rfU1vfBYsrERS9VkHRweY6mwfZbQHA37Cix2EczsjDwwvYyIT
tIuJBRYdS9oTUlR3Jiq5Nux+7IAr+Fy4XF6ZYO1fKkMXtAJl4ZRJ9t/vkLOAxUSkex6eE+Jw3alB
5a3GHdj2e87w/3ws+dKlNRp/pwr/3sQQJ9hEqsF7PqHDby5ccItYN3tktDZS1vbKtToiCQpKb2vJ
yrkytv5sXeHYem8nDQ4qI4V1xAZsUXEHsNkCbgkbZs7yUNhRKxDQkTfBRf1cBmo96Z8qY/fX6red
+3TmFtyZ9F89vm4pxKfrrGywr5h4XTZU3rEM9vEYkyYJKZnc0l7VfH4+Xbk621IrHmBhOk8OE+9l
SoWbICdQ8dBCTr4lmJoXMSOk9SPhR7gq+rEJo8hKgB0dyDyrcaWPOvA72Jdz3IG+0gxFQ9yxXW2j
rDGXr/6F6r1Tr39/2SXdkPqErbAkUiY0B5QF0PeH1sBBUMdWQJQh5y6oawk/OzQf3tLQaoT+6Hez
raK9cUMDBg184xHm4gB5cipQh7wGlRhPRFpq4467hJrA+35GVgDlgjmqdPZrFoZmw7lPwbvMsETo
sDY3pTa5XJ7QJ2X9nSO82bE6J7jTSac/moKAShYV1QDrY2nC7v1JrvUNmo5GFB8P75xJEHrotOzk
zxS8BSRZLNyV40MFxYBiN79gEUkcC6Oq+Ds09d+ZO19iePyFO2ATEAHCeDNGNgJXf0sWKCtp4xfO
surm9UuiYY3A4bHzI2bqP4HaYjvjZwaiC7UUEtC5vilpmYkC6od8pQGQ3ZmQb2OgqLAJ3H7BfwGd
cS3uMcPEJy0s2xApJiFfM/3QU/ivutgyi3Q+2+pF5s5AZD1Lh0MWEd79/lfkLRFDKFu3aDG9oFH3
VCmbWFvgKk1/dUskNJgc0w0CLjJuSd1WgKb9oNnRgaD5LbyHERWb4J5KtDR6xg99Q207FhfUJ1AO
E4Z8x83PDttvehjd6rh/SeSWH/LyD+NLQ2nvnFFL0FWNpfhrIQ0slCb/ipVrQi2zJkA1eAVdllHl
8pbPUf7j6jVsAxYt92nH1ysZQD/tZE5tVC1GpbftkoWYCh7KV3sqBgJ9Rz3NNAMTIaiAVF2T0brL
Fo2imE/w04jRjJipx9xUKw2ZZP5PE4SE7QxP19vpBd2l3TurG8FCImZ3y7H5I6DUqbHb2X4jrUoT
Ec9TZx3Jws/E1lb6CUFli9SIi6jFEGs7XTOpAdV1Grrn8cLabWY2fBFOoaPcarTLHr4eoljM8bbe
Jjy89wmcZdpFaPiXFm5DmQAe6VAHr4YOw3aATM+v983dRk7DcrvW+KrHc8VhWKiGo5MFtQPoXniU
08B69ONZi9M+QKtqW+i/zyNTX4kiPEdt8vzoMmVdzbAIVvyKMFqdXw/Yr1XOm3WrVIzr9MfcnDUU
aiXAs9yfAnibCl+MytdAl9uSNyfrr2xB0QroLVUDj4m6km+yZcV/iaBDVjiDFdY8ibekItkI7KN7
RFqqmIMQUM92eknVEw+UcEmUaMadHWq+SKqJ5cdx2RJJX4h+mwjlOxcyQz8mi87JCpDudHRi+EKf
Cez1GssZxQ8MwXGVsva6eHyG1zcmV4ulSMLBe1Twun47PY58Rz9hZE8Ld9Z1WQUNlJ8q3KLABTeQ
4uPh16LrDgUKwDXKBgMp8QUXayGl219WkW7yw8ErijFdEucf92M3svGQHZreUPbe0+tb/ivPrFPg
XpYcbG325rGKKmDbsTTLObA1FzNH5gnq0QhuD6hqOwgZISMlV++gNjI0S/IzbMmuRO3F+Znj7Bmu
U8AOBGPi3bCZFxXwmzwk4Xls/mf0nq9ed4CEkI9RnnjKfumxXPpeQalikVYBmhp8dpKUK3h3morY
VHJuRwcNRkgIHDq/vBAlAstYv3ZOdIFmcHNo7c84XjKPkGDZgWvrQ/d4kDteyYWypHFp58IvmCKu
gAeNXsXj3Hzb2Zodeb+esgXOzkC3c3IlyKXo9DyeMCy1+NHqxWvmf1+4o5ybYzU2pPHPWg44VQZd
N+51IDjVAYFskkA19E0Ceu6OUQJBdTgYaL+BPFgeNeYA0fkwfovaDX2HKk5ePFVTXonY94erNhaz
TO9U7mdAFRerA6jeIAMWIHuZCFr9yysWYAjkSluJBJUuaRk2yVcvCN/CYr5nZpJdzzOTmCGeUIW2
cZ2O/9jagohvTsoNQup+DFCvsDCXc5g0OMJ6FvCi36g5yLZ0CBBoHEuz4baR1Wg35U7W4sHsleBx
6mOHntONnuzLAF6ZXo5baE2OSapQ+7WYTwYRcXoNFTgur025BlCKm+eNpOgR87fmlKlV+WgG9hwb
TTZFa3iWIF+xdVexKsXFcM4fdCvAJ4sdfwRr03l7u1P3gLah50tjhUHTz/QA8lHeY1QuNctFSfVW
rlFVX/ZeJQP5wQbSZhOeE4o728WsoOug8QroKc76waBYJEhf5BMPvIHjJevbq8K6QT32BAtK/ceD
+gExqMHy+BztJ6GQ/j/QU99bbulcLDTQfei+dxEOi04VTjGrzlV3QZmXd8Boiu/zSO4dGyMAyog4
GSHMskL1Oid8ZFwj2lLliVjkjSh8jY19Cajz2XDbPAJAKbvZ7tzHtegir15O2cNugTb/BXGUH6c1
J0S/Pl+FbsYmUF7MpUls8muIyISIrRWw6PZpxVSpVEJd/rWQOHJftE/es4aF3wjkggSAkb/DMO8Q
je2hJzE+PE4By5JRx5HXMk3hK5pdjNnNZ6G0ddt7oGfHHaVLoeQI2bKVSIv9XokA05+bea0xC48G
3SidGztAGnbR/yv9Ak3VVFk5mmtuMfC/MzUlbga1Z43ZtTw8vLN/x16OpXxzCpB+M7QqHfBi8rXQ
2vw4K4jbAzSbrscv7hq+A8ggjvra1Yqi0GTNMs8FCTxFn8AhsWhq4mey0u53XGOl0qnnpmTEqVvr
gj3pqvTaa9DvXvjG9sQTfExGmIFr43qBoaMZyPvgHleL9W/KzOh/E27REnyEi3D33hRZUSR5cEJV
XfZUpe/Gi/WGb0mk5jTAfySGm0NZ6uI6VX4FCCgG6cmZzS3PqR0c3mqG/gMe21PkKDFhOE8agphp
Ws8dp2S9T/WBe4+V4wLjqUC9kKXtv0OicM+CyGuH1kNQ7FGD8kzqDMj7AXUPNgBJ/60DMFuFFKlq
YTswsk2zHFa0hqnYkCAbwMCCuiS7x9/axQl+B2oYd8uFYjXvqrkpW9lYZSWEKURYtxhLnhDj0quq
Ornw0ZTU6df5jNSNHyVbativaypmWR3SpUwVbG5Q/Rf5XEZvEKSPsn0NQjXH6bGWgYhELY3em3pi
qYVroLiRyt+qmWjE0/tQxxGjEk5EBr6rB2jpUPrl1+IKHinO2X467nH1J11debJvG49Da1oZOIQS
rOEH6Wfo3hGDqxESJzKa63oHC+87F1UB4jFa5eHZ8AqK1rIY/mq77I9+k+W0tAEldmx3aYirW0U/
rpBjOMeQFBBl22i3SUnc5sD+yVa4wPIt4ky/YF14O9wUyNDi0eYXGryTdtoTYodXQlUg4aF2C3Ze
3Yu14D55rrSvCMr+nOcfOAbvMXgJCbZJ6F6f7+0S0AJgTsRBdlFdhB6Ihp6qX2h+26m2YSozCeT+
gP1pm6uYJPbicS2YXXScEb+reVZsILzFcDgtN2Np3E2PK00osHd7ebb+m2kUEBhSLvR1SSEd11FE
2yBpfFkUSWc0HQBQyfVNicBz9RJLNmMk410yFUN14zunAncL2k6b1mO4c6IG7aIJLvCoG+5e6GDV
jkizhtRTk2o6XqMY7XaEMVjxCaNqUUaeTWMRy9Yk5hdnfq6c7eRcf1QlWaDwvaat+U+h/0egn4GN
F3U+dSCT4HAFWi1SJDppHJi1/2UZMrCcTePcBfqP+OszhMKGsTxNaZS5dpkvWw7SZqZLv41vOoqk
qnWzOhwIUVf07EbOOzhzzFjSRMW5vXU7i81YKY1l7HpEKUzkU1J8kHTNVdpKdycYX/OL5gUnikkx
Cps5lORzlNIwNnaxCRwPBMasnQPtn8z7gEnW5DI1huHJy6urx625vabAcBenzbOMNTp/HNWsom2J
Kscml0cKbRhHUCt2yEwLD3AItk6GRdYdbfLEc5c5Z/zg6ac9XJ/D9LEOL7H/LY8B3qmeRkkFp5SD
fTt/4+oAuZob1NYxB520A4kYaaaPRrkF90vWEp84UlQwUFlal6KucFZyO/jQWJTT+nJh3XIp3VK+
KkeIf445/uc9xNoL1hqq2Cjcg8Pp7fv8XtnK9tonq8nC1beRGpmPc0qZHh7pvzbgIdFyzHqC2SsC
6fZ3HRojSdNs8FQ3fcnlsbVqCh23l7hOc/idk4EgxcpT4wwH2jz+5hRMJNEwjAYrZ43aqA0jGfXp
BWooUlMPjdP3cfLlVJo/q1ZiAsedsy7siI7vBq7sz00KDFvfNYwm1gxDO9NiBpUrpOaeG39IEnch
k0xPPi03PeE4R2wf4OAKrTh1OIM7qlaMOey09z4Jn6LnrKFadU5WScEMOh1588Guju/xPI9Bfv+q
OaI3lC2o1zwyhuwaVJGmUyVX2iev83e8YIFj20lpdlTtf3M7gWFZtfbrN71eO2i6SNIK4feHZF/1
S1C/+xIPONXSKC0hPJyiBUvIVCfa209xRpo4o5JM1xpu7ycrvOEZhtmXCiQk7IJnNd8TmAPx55UN
wFjWzITjknf6hyl8PU8iRFFTFnRTiw1BKBJjSDSVzibKqrcaKM0QzBsCK6KHPj+JhUSNGxXtZU2d
oS5D8hSD9+S4DYGVSCDMX98CgDUjutJyY6xu2EeVOmx8QoPkqUTF3/rASUi30zAm6PkGVJ8Lj4cG
CznSfnGQxTocin87JCfyImV5QmN6lOpeMVAtt9oGlGx46DAo4POt3ukzmz5+aRNLdhTXezOgX2dl
S9/MMfTRCfq/Eux3uJPgK/lowqehc5y4TdJLDgk2YaDH9nK1w06IlkJAhL85qOdDTeh9GVXWRKer
RNSsIGJ8ZFuA8EegcsoayhIXShXXPMKpjiMbExHdtnOZ8n9/wK6IE93KLO9TEqz4d1IQmaQ8OaIL
UwpWe9lkTRc2wAv3vype77xegnI+YeEvTdlM8zzmW3YX0xQq4Fy19IGecuVNWgo8X+fDwVoL9bN8
bYwll9svIEN0/wsu1uffe5TSsYgME+hMjRnor03TUYcANjQ/HbDq+ALg9oNF+tTKXdpSxE6QUKN9
sLWV7+cNys9wMy84Oc67cr/aI8zz3jqfhF1PJi65EFc/CFA6B/7IKrposGK1HDHMVx+AK+1/qKza
lPI9rEyL72gLqGmxls2sBdAEMnVwSAYdj2Ymf6dpJcnxNPT14WjXpg8tTA1A9+jgL8UXHPn4fqc6
KrXdvWxRyOX5KKhB2F/bR2vVFncYVsIj/70wOsAgJiD5jXBiweLzMNZeFJPX1XFeb5Dp+GSi2PcB
Pbi05Rd4M9oLW821XJ8a7C/PDGo0GT6aKA16Gz2KXnhLtL+sUND/iK8rFGdG/y3vYe04y4e6TYVq
RiPXH45PDr8RU4iVyk0GgW6foKUDoqntKMRr3QLpDlEsRE5YmK3gLV/o0w2jsri5Ps9XBmChJ6RP
0mBTp+v7rpE6/8UZRW4hiI+7Whufl22pRcHBaWOKQOmXg9Jf+tjK/H86m5a8V6L0uzk+ECcOi5aD
vAcVvNVt8S3oP7RriLZtpiwTopl0dazQyHzj2TNXePCyZ9OdlslRDQKDYTMQCXAzNi/I0g1nldaY
BhCMhXRGTofV8TgCqbHTlZNJ0alHzA10JYagAJdg0toXYpsY8jgIttNUKCQ5Oj2niXIyDPs9us8n
ezFaJvZvRxlwOGEhU4ZnKgQVBQIrgBLSu0jttqZP3xZrXYFkzY3n1esvPpYfVqHJhNMHcdmbDIuP
ieSdjuTWtloeiJ0GXWdmV8VVLckpSIn70b4HZUfyR2qIz0wyqWFKPyVNVHk7rk2H2s8sd+67c9p6
fa9i2C0MtL1gnQoW3lyUh6QdT0kWrgFs/gKSQfaZqq65Op0Ax+xQcuD4D3gZ2zgxK6OO+qqrz7Ep
GCNgrZF+knhVUrBCwNqTuxHkH5QVJ2BA4Y3BuhAvFXmN4KMM+F4UyuyO9/BFm6NEGrVLr44BmseH
qtVvJN03LH/wgewMQfWzEpyi72xuKkEnF9D0nRw4CuOoMXBrhfpBy0s8SK/3102B9dWaNFMf/DYF
NRSmqk5ikVh+gycaL2V1SpVXcKXg6Jzetn0ds4FuwIkxgdwHlkL/1idELMsacS3zSgdQaPzgp8yb
ipsV6mtBMcsdWvVxUk5cgBfCmhsUrPEO8Uclqbo9qrYsnSAY07l2Cj9ggc+aEhnC6/PM1xJtUG00
U/iP+sKJPXfq+MeqSqyEkzTbWkQAld+lyRtlegxgzu7S0zX9c9wOrrIDn5F08dZ1GoKLDCKz62e6
B092ZTxB8hpAUkfnGY3R4m4cL/KZv78OGB0tW8b8MAexmk/TDWiPFx/3807mXfGpM5a0+0cOM7/f
IJJjoJ/OuCbIy++b6ftuDISDVW8THumIwvZdNYip8UNzE1e0BzpdTS4YOLGZnMb1Zb0m7Gc2YSKs
gj5MJ2nbW20CFQJglgrbVxkWKkBoyMSRj9i0GhbPyVVh+qo+tfEdImm/oMsOtcJ0CBQV/OkmiJ7C
TU2dCiF1sURWarJ3ewTv/u2NlsqeCmKl7VkvMNofziqpyKchVdnDhWN2plVs6x4iF4tsmIiB1T3T
KN/t//UFmBFbxRmLT3uArCdM7DI8eQj3SQ2KfxvH6MddS2GpfCM1yh6YHYNQXj1YVBPat3Rfz/mO
krluyVYPJL3IJcOynzdr0MDoEeTlGzXsgCV0yQ7bBs7yl3aWSWb48rhDfVfCAsOqOlg5uMwpRyl1
R24DEMyhr/fYiACm6TOnX3bjNKFRByPxki628bYoXuN3qCMFxLlp+5hceTmrCtWiEmFb/CmqrbEz
lIvQbztQT+/IMCyBhUUK187azwMtkyGX8AmbA8L6y7RhtpGgR8kPtlNZ371MKNRlpoJPoCSeA6k4
p1heC57Fh0/Q2VvxcUq5ePNDPPRDt8A1OBLg5t14QFsszY596BGH2lHn56i6GADamIwFGumDiBjb
l2BCrfWlVW4ChdtUCkRFHMU/Qyft++ijgegyZiGKn2Z/x1++izEcPeAIGFZEJI9knZ9CM8k/1pjR
TFPuEF3ZCYMcHdfLEnmiEwW6rpjgtzt8+S1BA7XXaKjTT1aGHeSCU3wnvR0qaPRwBmnwY1ifCp9v
+BcmsGQxpdUyOT4ngLs8W1sM8ngPHJbBu4zNDIp9e/O787/dPXyl7KMEkD87o8eYT1eq3zj8n/X+
An4GVoJLaTy/9yQMgxf4FgD4T/JbDVYaMC/EqQWK5uIYsvD9ukZwYizGQ5dL0513MDF9sAhCWHnX
QwZQi5GqEV0WRNhh4Nt6wi2w/RzYk6DWOLy5bJV2/7yJYP4KHIc6wXREERfHQe4xLK+DlxGu/Yq1
8YxxHaZJCR3qswSMMjJUwo58wH1EtID5RVbAlFegGfQ+BzlpPlrHtncNglESvUT2CGsMfIZ5Nq+v
tx3TjWcpzaRH+8uEUMqlK2cMcgmiHEMfU9rhhhoahSjgsGSywKfFyrn/7W5QLTeaYzBnC35RmcBb
j+ZELnj9AGAdrKZj+EnDXw4Vuw3Xn7AMVq0dZSTSTYGHuKX0A3K9z5222gq5BmxxOTJRlFYwcXsS
B+JVaI0ehgEJkQrv8XnYIzUwyeOLh2O99L4nBUgi378EiCzpUKkXLPjuhrZPRN3xvdKKU19I+ft9
qEDj5uTbwcLhcbnIvTGj0RyrczZ02nQehfZzvpTkQNQmgTVIaBjPsRClDBdeW0NEZlznIt1Atb6z
2d6f1dt5t+LnP3f0kmg2QsvYOPU+aglR3XI/jtlYQRdg2Wflhjmgf7B8jZ8iYuQjLoJigBfFNWVq
xpgq8Rniu9S5hX2Kg9XhsbG+tK3dzzW4RHCrM01wbFn2BNTdGEV5+2ztxtZx+GG8N1xeslDZdKR+
PLk3P2tLFMIXqyyWMnjDgXa74SkUFUaKbUaGvzeQsEDcR4C2NjLmGRfwLgLsYjyjAYoF2yYNTk3f
ALPG7WpNzIL7cL0k21Zj2tJp0nmzXuXjcB5Kycu+/GvtNsZA0qNiwWob3zq0vYcn/dce6RM+VMAL
bRUC8iS7xBj3X07W0otNghfNh2y0f9J9+rWJVHELKDMYmhwFJptV2PLqCbumP5jj2in5AVafs+mX
jjMM2Z1cnL1Jc87u0XLSoaC08bmAWzfNQBwBmc3YZTfnb2XN+5qAcZtDZGelfr20xB2QSZ0PfTaz
AbC6OZRa5ZbZVmmYwTjCv2xE3bcHQFO6NrK/b+NEJDntogstaIAGEHlz7Zh0QZR1Kh8Cyio/tgmt
rxumle8oTe2bnb+s+G9yIh3ljwaqMSCEC5HpNhhmBRrqhHIX+R67RSYQcMr2QaHDPr2H6KL41euq
aW9m/FCP12DKgnHZX1HoHYuYZ9qQhQ4AqraIpPY3FtlpIDTQlZXvYeXJol4MUag1kqzEYUw45A2M
ymaYj+G1s02Om37i6ZZYtOTu87gxnep0f/ucuZNO6oM5IzldmhqLcejzavU6FaU5vgIDZgX4acpW
H6P4y3c/zu7F2G/azrc6qw/wSao883oUFYZnB6G0XXq71Z9PAJQ8CCHxMQ1A36adDlgsEfOegI5L
NuHGL52d3GDJN2zD1mWRhJIE4RS9bT7NSE/Es6Hlxugdmo8eOwLr7kTS84yTzBnpP4PZ82ZltsYA
nwtbiHJJVJuQX4GuwZrkaeMSDrGzqpL6n/MqH8pjpVRx73YuSWuIRJCGxS4kb+6m1kGgOajWjPyL
lLlB1QoC6vFF5fUSz/dNbXaEUA/Gpv9iJlhahmWyC1AEqipu/W1x1rdhviwmF+KnG0zw8Eu6T/a9
bY1pr9SBXS4MVvRtm7EBM6z/6V56CPTHGg2omzbB3za564sfFnWE/Hfu0iwaJBhLGhhn6lmza+fy
ESThravbGt4ecKDQ77K4J1PihGmNwucxRGwvBelkfOOly/8o+JZm+OxR7JUtPkPZ+MgEqBjak6ke
6/Iq+S1ImnEvgkmkikXcp9wqQ/MboD+JLPnx+/lpE8V7Su8HNs3o8lWubkT6v3tUmc4IQsmxIAj3
a8O65YVhKPwfnpcq6wpioZWSDgGqHolMrmBj0V2DEk1HacoFx+tSJrT4huCoj+3rhtRx7JurjH9f
O865N9zgdbyHrfIsMrtK0D4YTGScpZLDSqLmxbMrXzR6Kdz/+Vak8IQ/crRRQgM0liLjrEi8tHdr
Ix5LiI3iix5FWwHOvej+v8XL15RfDvzQkWkrNBWoM9snFvmnVOp8rNZ/eNOiy+PjfvWQWEEGCBBc
JrRxaVdG5vDfj2UAGsPQpNf0bh9OPfH7NmYhAok79JrnSWhSGVkOb17XWjEwXJoNiy/Rr5/uRJof
DcHL8u/os55wMvweqcGmdaMklQrLrDMbIWfbwfir4NhxXhcTAhKsTuWyLkdKkiFpQ5zLPnazV03i
Lryl00pLtMxeExMwnVXtEV9gnFxTP1yPXfFqjTc9y3kkhf6buIHJE5ms2owthXx/j9CMxjFyl1R6
Gaz6ZhWX/k2AiMQt9aVeR4CY3xj2cSgoFJLuv51kYMTzKbSbXZsBlithTjGR3Xi0HsGzSUZdeAcw
8WkrescN72eq9zLKsExlnuiF7gd8LH9XJtPRzEfAsDjXbYrQw+djzEvK2bA7wp6K59lMTcNnZmvE
KpEb19sdBHyJYW/mXdMnNPU6oAc49MY/sRc7miwhROjpNWBAOyi/yf/sRVtySCbnUfAXRsZvHbug
RjRR3B21CBLJGkEDhWJs4Nc9Je4U/VhadLfqfeNzWCKOJ9krTx01/ra8OMDAy1m74bT3ws/9o9+1
dJVf0MCsaTJ1L6gwlBOlg7bceLPgnWYyuoGTxX57V/pD9mCol7Zu60e+dGuZ9nTM3dHl8oRoAk/8
Xb5MX58C69xvWX33hzhXLKyl6XyXRCfR6yy2tX+oLJZ06b78SV6Zu3tRFKAMZv6g6bOxi3JQDlKS
niryOMbGXJIkBK99Tvv16C89qvJJYbtAEzWpiHYbM+OG7qqW5gt3+cltEPxWEsCQLgEZr7yI5+zT
1RCe06XSx5ybYoUaMNGDahfan78G7KiiS1AOT51P/AHgTOUbjqaJPRekqDrgkAk6n3a/Tr/kFSog
Ql9kVaq4aUdvn0kAlmtr9MgcDMp9iewOTjK1xbPMwih9hZIlP5RERA+bTFUCpp2bwvyKbieNZa9y
OYI6GcGrkrr4yX5V5nYdsbm30WBHBPcO7IaQo5QdCF1p8o8d20/qJeNgq0zlk4vXn9vRsZ+NPApX
Hj9xGpd8da2xONW/gwC9tw7XG0/cWKa6fUVUGZeOirDecJ7ywdfB2A5szX0eDD850lgTShikwQHG
08Qm4zrwpnQIvek1HoIitICpUCaulkV41IbwlZvIYBPGpyc8F5Mg3I86O5DhoFIAxAVRj6FeRyTD
UffhEUdXa1ewMUATBSJ8aYrbAdg0hj4w7z2ifCK91i20ORKPvvxgwZKTWkzMWKaTmZvs163Xjn38
F8BgQe9TkJRemGvRZJvCrk1BLiJ0lIfl5OgCrBb6WAw7jdGicHUoPkCIoeThclorv2IHLhvYibDI
1JNUU8DJnp0L+WqiMZ4KWI6Tv0CS8oudjNmiYRgNSOpqCggw0usp0LgLpsqVs1zsi0xFaKvIOhcB
sawck6oqb86QQCwWcbFfQvX0BYm7xJyohW4J3ExzbnSjYsVk1jBvEOqJBtfS7pbwXItYfoELBte6
tjGgmInT9ot1UDTUjaRLymMaNWsZn+CYdFirlVbs5exCQe4IDh/PQGvVeDt9p36J3AcjRzfGZlGF
VMdNYibS+sTm2CEN57LFBoiaWZqNEySiQsflM5naMK9TBq7wJ3D2fPkNfbxXyVo5ebeIrN03kiXt
8dJ45AA3mTGXeZ+81awKV0C+hl1E4pExvNYmMeat5W5ijjBSdNMUJc4/HiC9JU6czfqfShb9cNTj
sKB/q8/lqw6biuKKRAC6vLHcbPcHlnKLbSnC/AZiiRvlO3qG/0yvpArLbnJIZKn0Fx0xG6PGHKT5
U1VdE8RGQZDoIkQYL8o0p15HyVIlHaZPFu6vNQ75A36gtooBp07XtpVwJ6k10fgAquLq0JzRFpKk
+Hx2S/hou5f8xnUK4IrUs2Oy6sEvDXi4BLIwWD2QQyzcF6LeymvCGyoGqOQ5UI4Kfo8RLOJmpG0r
hfOWq4vxOsGh+aOD8yhBVBx/5itxSEY2uTBQptLDq1bcVhpOJw7vS6Bp31Ha2rwpWsl2sSBGDAue
tLLYBr4EKHYXl/0RpAp5VeKaHW3e5AJ68MfQwI0vxjpSVgfLFusH4Y7HMbB7dHiNmWLRovb2RQU1
J22EDlXVmWR+jgcYC+I9wG89PcyJQFOAiqkWyBmm+5RIyEB77n7523PXv+lC7pRpGRSPi5VBhelh
oKraCK9TSvql6KfPNc7ZTgPqb1277NSyYjd2p+q6GFh/4u5XDsKNgMphRYR4tcmr8qLQXZ3mMjgt
JrEIwTZiSoG79399kOXFy+gsAQ6oCY9kZA9pOzVFRD8MLFjsm4OZDDowHrFXyzyNRkYUnkVj80F2
WpZSErXIlvrri6WNnM4XWI7CebOwbXBEY/XXmucwxvHclbps5ltWp5Ljlwcnaqa8WMJPGgyI1Gcv
w3F0JdLJpUyBHk2zgyEszRA2hicp2V3arYUMMOPYNyOE3q/WAZ9Cy+71S+MaGXeJJqnXNt8qctcq
X1cJl5f6L3zHDuZO+G5vHa2wY+21NK6jpbe8FQtfrz3d4TmawmLI8asHA9HzrCLPt7tQHkwb040j
A/zCJ3dHu6hwmt8DxIbbdF0HIGqftihJ528iQwYIAagk1nf936WTFXhW4aNXMdw5lWEthWIbqhmW
nYe/w6pvIV+waTjCD3i1sPNWAbv81LjuUCwRBSt5kk6W13he3sOdykyErJrNRXJklYofbKPPHXE6
pSVOs9mBFIhBKDNrdrboYWfwMccpF6IVRUMuDYk1OmE8aqAu12VKe+LskGCXEiF9Ksc+ERyeKZYh
agy8/Lpp+s0ZbSIcUnKZNeUtIwWqneapR5/oTxV7o/yYSJkk5lORB9TaelBuqNi1AG42OOrrfS40
/VjA/ab2PdkRqWOy+iWy9aTfwokEi1bPOPSjaov4rNjzBXRlZQJMhUAIo4zBb20Qr6SE2Nl0SUNl
P6/fUAgxu0mEaq/koyg6LpXmKW1rEM/19v54avkiGSPNHDFmJeqXOpnQ0FNoSSdH8Yg6K9SKqVf2
WajvdG7JdHQQqUq+tEWo8T1xuqz+FWxBmqJ9G1jqL4PHRPdtqQRCzCw6irYGtBdAz3ByHJlDDfhf
u+HeCicTgZ9tzuGMAjMX8jyN6eNeD+1fdnULZBQTbcgF4aS22DLccivcf/rGLHr4qrjZg6lYxvyA
HYTTTVhRpU960PJLESq2vI57QqRghP2fAsWOjovo5FEgxnuJ7Lm1OsRYYzX4gGSsokArqbPG08jz
nOlKGxGM7WkC+NxOT2Eyl2YuO7YD6XJGRLu6T+63RMwjq9P3Cz9xPKGvLJvjVBNv0zL2PFbXWSvk
LocdBCbCTtJvEe6cl82Sjb7fKepO0TVE+beAF6N7VUQjyl+QbAoL9lG23VVVANSxzo7utTlJe3Eq
HWU5vCTLTCUUAbsE3a4UyALwUrdHQTHA22T3VDFRc7QP/Nv6dfgrIkT2COkHGDo4cQrDGRaddWX5
PpAPpaPXx2fzw+WKh2Nl2haMCDRtSI3nE/zXLY218+4oW0ZKy5uVnCYnmMsh3gmdQP9nDsOblJr1
iW1LYejfmDz+YsJJmPdloGuXMSkqD3JMOjbsxAm6A9wDRk30OLytFOvYJ1uii9Ue1LuVLLYk+K6P
kj4Va6egZRAnd0WnDfpd3YB7XjN6HiqdoqiQFN5MmNG2+YG3P5EUlay8YymUcatLkdwwl3wbyzSa
HYVFlmhdDY6lIK0WIDJaYRLUxXBY3/PKedSsj/2LLrYvoc8D+0HnOtylJV3lRmV8EC0kEo2BC57p
7tu41uZYUUZrkXKnNNbb1m248/l5eIHBIE7uIXXC3z07UrafqGRzyQ6pJLMNeSKkL690LZ2hmAmk
EXMxnhbxg8hRTEll0koFaPOQeUM6ghbhelDjwc1vlDtfnpaBbBtVvV9qrSiL8bhDqaZhUU84DLFS
zQasaH87zZoqvQfgSiSw7ufACQ6/Nr7dMl64jiWJXz64IhBVubKYSzNirleX+9U4AHz2416zAySM
szkEwnLt5b0TztxHJcnRSIJnXbci9E3fHs1HFqu2JOV6OPkPK3Q7tpQEIqjBjwhtqEK/L2g/Nlla
Z1R65vFAGXJNGCihBKeoi9KfSMPQxjxtysJu/kE58yrDWA1zELB+rXB3CdmBzwcaAwhgt0rmQUAC
PxLRGDhyFL7EEoxc4O5gdEMwJUjj18gDSbAH7hmlD9v84RMD3HSGdm1ZYqcMivd6btrmahAyDzgc
nbra63hfFPdjH4AXb8EeU1SRrvItsglTdA21oIP/aG27H1EN2q2RxSMsRKjMXHFTrRm0S7Wlf8iq
MpPANK4y/nLwPNejP39xkcllmT/L3NXfUa22vReepi4xo2jzwfRu990bkaznVbabKozm8HSK3IsZ
Ui4RObnKY1Pw/GUxxz0INo8qYYKoR7VyjJLGM7GDpSzKR7oQLVasj97o9MfzIHWl1O9+whJrJzrl
3qfR/MCSja6xSzAbbIsxRFso3d2aEKLUoAmEU71G5AF2iEoYStaOhxif8iz0pjR/gxUXw0NV9iTi
7tpSOYc0C0Adk2etsh8lBbQAV53Mi5UQSVAVjDuXzROQ+IgQ3c9+Q05inRi4kUYXJgsytMQPi7Mq
/KooAsL7H0kj4OpCPi25iBus5Y3XQ6O/7zikM/+AvaZrWecUW39jF5Y311DNusni/1oOKZznImn+
R6OxCERiL3X/idlbLJ0pASL9NmqRZYX4BS38z8Guo9ITSK9KqtlbKrid52In/O2GLD3FRUkGHBSH
x4jmmBMMtgOzw91DeutBUGH3ZCk6YlQqgS31mLP30KD7EXhL5EhlpzutvDWdMDAg1jORNvdtfeHr
O+JnudQaVOu9Df7yT4Yu1+SFrVkL28bmHZIn4VOkxP56Z3S7PO690HB7rpy/T6BArY+hKP2AWz1L
qMul05tMlcCbDhg2fUM/1/3nnksQbE0b1qT1fuPHBJCWhj5fEoffhLMYTOCgiXfiQ4l+I3In+WBd
K1LOuxTQ9yXVWNbp/kzui/CufG8xu/D+UnkEJSBkjwFGNEE7CFEiQbN1gsd75gTMi+oYwYZra/1Q
c4kRrDZYhqkxBwDPXQHtA9m0uBS+Gyd47mzdwC5UKppjKJXU92WHycsxMGZREkThCrIXfX3vpaG8
quVqaO1RkuxOh5Mm0G/iwWmj76/u63CLuOrR6VTYDwLWmZsgQUGJvLjL984fzjhnk9kfH1hVei9L
TOwsrM6AU5MYQqPeOKiBa09RF69wOj6aEzLBI9xgr8YVAfdpyCpjwVrXT3oHHpziAUEnSlry2Wbt
M42XFim5DfboJDHa+ZiXceG64w7R3iBHcIgkRxaNzufGN0knmRf6VIsbxYJiRyS9PG9oNSTMm6Er
pxB9DBit2QhOJ0K8Ggd+5JrY3DrPr3/FacnCSz32L8dA0FpAXsyM/Ci6lbUgTe9Ns6lpPd2C/5am
mgtgqvAlzQHWvS+OwXQb+5fDm7nRV+Hb4G5NoQ0+8dFhfb0+/NB/m5hoIuMM/UMrnRy2woW3KVln
7BRL15aef6l8IKfDQ4vjvT8zsu/6VbThiP5Ocoj3YGWa7fASnaa0++WFdGsGBozd4H60cC+UgTDA
BDoeZVTaINCEd0Isjw4WMZzV5vdUCOJhF3uYxQb5Z1PMlIXiumbGF/7EEIWxrhG1Vo5BLP4NaTju
3I6vQwqkxCl7sCBqv+yVOMynRk6ZnM/htX8T79X/z9cOgt4VIazWSEZ7L10WKAuogFbcCEwSLIKR
4718gK+extLqct6/rZsZX/LDbAu07c3RpSkp8yDZNzsBQREBVapvD09QftjDLKc141bP2BEueWA8
AhVuvi77k8/jR0SEfpOnFHPyBJ69gzdmycv65D0koUCiR0+vrU2ANOaU0YGjisEF38lfX36d6zsQ
fEJLpWwGSm2QsfQgLz7GF3tCBS5JqIzuqx+/0XwQkTGRisPcDLS0ZdI2B3gsXv+YAALekEH2dufZ
S8hQ7seJeNwa9Xsw4PDNRRYvCVoIAfWt80Sfrx6M92gfyzBYPQoBkPP84OxUAzk2jQCofG2hH5O5
ryKQ2Wcwx3WaG1MBjgYUFv/VIprYmyp0SumsJ+IhgD2ombB/qyI41XY1NrFZZkbzVPG7A5/2aSOu
L/HT7JrH6kMnqqeWXHtwhbxDdIjscSTl2Q3Ae8EUxvXtHh/l0dQifHKBQBuOilx4Z+IpOruWvUjn
x4Tc8G1cqnz7T2cc6TEzsnYX7ihveNVyf5eZ13CYgFsxOY7KakTamJojp6sXqFaqzMstyu7E7cqo
NnXNEw+dqMSjvtxPkTb0yHoLRZHkYfdRNoyEWTT3tHWON9Pdd1IPxL3ulIbkMUXq8/3AqTwfaFLl
Is003/8pOHNzd99Mi5VEe7oXQ5EYkPsBStXOjHrsyd2YcK4vX8CRGA7m4a1JSVTMjKrI0Zz8d8cz
k6Ve/ozwomRaTyQCd8oP0RZpP2c1E3Z7Otx3aaGXJJAYvJbAeCrTUEC1+6Q/qlR2czjcPJOn7igh
FcJ+m+PyZx0l6GHYNaHA1cNTbl3hX9MkknUxkQxKhYbuY8+pBdQAdGgSzkPTZ63EY7K19BdFnvqA
xiFm6/vTpC1U1RlPm1bdn323goq3TQY+dlvdG0sucxcUd1DyZ/GzV4RJMENtwEadvB0C8meRdiiU
e7FzQzaSK25rVavzVJZEQefgQfyHpc94B7plXLEzi7aETAsHpmd5jBriFEpxtxr9EfbmfhptPxnU
PQamThl6cQvqkveXQjLgCalCtsim+SIidKLVZRCO4X4pUJ16rG7aanKUsRL34qyqYFyFwqcYZwzL
UvHUEYYAtDzo5n7nTelzh8konAx8gUWDjbYBCcolx58zNGuzJ7Z8uavnjFbWzFVHCtJXzounHtqm
mLnmmpxRwwGyLKwqoV6SqpLraxNwp4CZP3ZakW8PjvynbbnYm3KQABT48I2SxjqwNxoS3USgQHL+
pVoK6ebXczjlWMGWMHdB2dlaxxdyB4hjZBjxb6bWZKqf1VbR4NhsqixAREMgwK5oMj6DaG1VwsDo
XtfoqdD2zpmOfQ/EtNT70DnvnKoV1z0+uHT6J1+6b2wdAqsMgut+zdDHd5CJ9r7UGfnv6BDDAQuY
GrsduS+zQX6k6JVPevJUGaGPmTxBI4yUOsdwkbPJW2GJaR6rEcB6wwRuX0dFT0iQW2u7srjmNKt1
7+y4rTd9SBu2HPFwlD740CFVKZn/p/e5iR156NGPur1w7031jnO2wz8dhoiRhG4FJUIJHoNbZ9rn
mYHrxYvkL54H86GiiTE+MjWuKJnvLWCdCaDGOECcvi1YwvW9mihmTWHsRXQ5ZygLylOshztFQMi/
gToZoyJwS9WH7mJRBCSndGYixXrv4KQ0SkGbBB0FnZltjTKwWeSibdSVObcvApKmQymKEiU0ToeZ
MjAxsCSKDNq7b5Rav312+6seJLxzItapkqZuE2wL6Rlt4PZo/e90WbHcjVZepSkyfA3LpNMxPqj7
N2VJ6LdXPKYGrnSNfQ4jZrIISc5XyEjTUkiM3Vr1HCoyz/AUTYTEeLvrewmqyfKpreJNuievNGZz
vnnSepWC1/R0PGRKcPp92JhrXViZD2OyymgnmcC2OG0sL6Ob1XFy6g8m7u4ebe9YStvygqn64yy4
OvT4zBAUsLONg+sL+R2g2MEaniGvafahYG4nPrfSAxi2Nu1Fv6ZHIOQkdn4J10Jq0hZ5XaVV+dG4
K4myheBGJS9U+PmO6djOouKC9dr2us0s8T8K7ppSHWYT+1N7lQd371F0zMjNdgnU5vQftkzZwbq7
wWw70/HNgSLE1FWXOV7ISstw7Lc4qbRZoBgwsMxECIqTY58O/WZ+PA2uEQvG0X81fdJYr9jPugf8
hgblgNt5f7TlPqzMWTvBkwynxMq2w5uTvsMFo/YQFgmWPUWb82ke92EEORBv+uXm7Q42i9M50IYU
C0IpTqV9ZY4WTCW89gYs/C0Og92MUGcZc5ZF8MEQkhLTrIiSi2dCIpLSOXa9gHO8bNzDjvHl3WnX
TvNN93yMhJrx7PSWd0ZC/MlHvfisjI0Ybv1kol6E7KsBoNOyBu9cQ2Os2N9e7w9gz4ee6mwrifDA
TGgkx0CoT1wBaNTcq7/nt4t3XEZ27YWRfvgYq9NleW38uV9sP0uIIkdo54K6hHTXPv6L+k8JPkyA
CSiMrTRQ7/ZFlPvaCtkZLqnMSRd2WKpBSLbxjLICR37PK/cwU4TxJDD1q6dgb+YQ1EYMaUQ13+4x
hxLeoOYoIOeJl2B8uDBzkWvvMU0/ROAEEsbCiZM/RFFZzxvIMwEfaJP2m+JHt3icowe83z2rM2s9
Wzzp3JwsPRzu8Uz8bBXzCYcJXMraqy5H9Aw8it/+QzfdvTodQYPLdAUjphNqhNcbV7IsCsLOBe3f
HQomS6UTlB54ba/dPk3+LdCm0ynyOZY0onj1TiBBtHlqIAZKlavrSF9mQ/QdNkwv2n5Cg+PzgwJD
oe/12PwnlQwV82g2s821RonuB4USXrsX1qswzZ1SD+UjOQsQyvDuwbjbjWGl5tIDVCHOhaxZdTIj
vLo+Xrbs6i85T/kgO0eTYAfpHgvdlMy2Q+E1lAv08zdmZ5sz/ZFkiH255F9i7hPSj/JDejw6qjpT
T/kxRQCfp9NuPUY5Tb83vrYW78eDYYNRewLpjYOCzCtO3W6LW561Zi8iTJtH6nx0UNLOlsluqj/u
2ndavh5qH5PQE8v+DnxHipvvy+Rd417klqAjv8Hb5ujzu0Tj8RoUrC2+VFc7VaCbAsmCcCm1y2Q7
pzuer5m1ubGBU8accNfiOr3d2ngrZkZJtHbRi8X7Tq/2IN4KPIZXzSv3CWUxnB29kjf4Rfq9zKOU
NHVsZxpKTaUmyvOuG5F634xlXHXay2kJMGSwTsVqd+SIK26QDujX2kaqDzZS/XVP8EwuPqgH2A9I
DyhaDzV0RIJ7K0T0ajCEkMidDkBW4efHu+cmGw8CkEGhnaS9uAgkTzaLDYBAX08DGj97v5UM95ag
WViDlDoY+OjUX3cgv9vCQRByS97/ITJjTE53QW46n6gkd77s1SkUXNrliv5lfK/GcC7RGNjgGA2F
la4qUcZtmMvVQnmNgit9BSkE8RKUT0FyWYcOTaORu5kSaTxkvehvpcg6bx2ryK+4b+zhB5oVoejW
BHGlZXtzim4az5yEuHwapJZ769C9v4eMbew1rN9VPZy6UAO6mpf1NBY/x7dh/jVn1okhynQ4zZmn
GAYv5yQ/5/AmkxcAt1u066TKAp7YfoK+YicW/q83PLFODgoH9a3d1jFuT+9/rio+alzrI6kCtmyO
a0Mn/y3wOZjUHkJ3tuXSb29dt6bvS7ZJaBBr+ls19XbFw2WBbuIAoFXhDn1/pHJQYgmGMyQkWqZq
6I2vY/dkLw3jxe6WSb7PThHFTNlIt6uS5/nQsjZbmm4QYFgywrVgN4AFiNPzItHX1Ym///fetxMY
ToxZSMtRNdNqCDxQVhtPOi484anlR8Licq0korJOaynJEExB4AWXmJGTHxfoaC3My4e8mXrcQ+hW
dXjIwlLWgsL6phHCb8sUYiK16W5NaxOnH+fMpx2QB7Si4mk+CyIlMMxC7znlmPrPY7esbwFYZk4T
o8PG5DT6A9ubtZ+GiM9fu1w6FpOs9y8eskSJQiRRy3GXPqc8D99smsp2hL21UDGQZqUSbVB+Hdv2
cUrL9vi23wvHg8k5AeBmyqRuZbGe8tEMdCUmIm9xxYgq98l4z6zt30nqS/+aukubYhUGVBJ05r0m
XkWQBY6sTfRvSTJS7Gk4sqVEz6crA2Xbff61XTdrgR0G/dDm9XIKIxAuMHooxMoZwqKlErG9V9+z
nu4N3x4znlViCgX/PM37wuz3jP7rpnCWbLnGBUw04JyJyJkrO9g0VRGyIwMl8fH8ZqUfzLvYrn+1
f6HLBOipJ/wYrilJun9j8FlhkwAFq0OzQ9/3OuGZaQKplBkD++YLcttkPiG/O51N4xNoO8HyLukE
HtPridqlH2KknS1HMhvw1cy4ub2DJ3bqA0MZ6Z0G1UqnDhVH9wco9SLgWfkeVP3jcXtgDd1ifF7S
fvlaI9Nvlrapr6Frn+DZIydRojJ78jIuYVGKSZqzNlMTweKshchKwJgauO01ow+A91Obdug9cSEd
UYjhbeJ/mexy4a+8hy57vJYvjdTucGvboaMHhGfJuOBt24JPN26o38/z7TzKZdEYeGk7fPl0V+kf
iqkNuS94OLdmpBy8D/8SJYkkZ3nmVdVwiRqjtW8HWBb/lvKeo8ThSTWLzzKbKQFfxIbonavlUuGx
u20C2QP20EAjyDH4IPrifvvLIMKQmfdLpRPOYq3tLQaLx+Iv+kluuO2IwF7xQC1Ouhbjly9wwyww
IL7axDt2f+q5tkLfcn9DoKowQ5F+jTMRNtu+0faaHdVMMcTguQ7dP2PALQgDWiYzPZQf1FdIs4g0
PZn/uYo9H7tWL0LepMr6lpvqYksuBMJnAsr2f8xhDF/cjCOPRtF2F8TtW8Z2wx4c2oPs2H/4IUCF
cI+cuvVGH87f2AYgfh71w0g9Rn20RT6A+r+CATYu6vHcK/kdEUsVLGl7JY8X26sqAzuPJQHsDGXS
pLXYglOnUMlJz+lp5Dn5uRDRR3PXAFmj6LOMY/fWeFMr+A+5uVZmDQiDDopGalEJ2Qo5WTPsgvxI
rVN2Lom2RMrIHtE0fXMWN6eTpU1GlGvtfQYZh+zBYMDaNeTZD9zd/3HHCsiaFh40fZE8Y2u59Jun
CSvbuB/E15vnHcCAVxwcJJUYYOyoihZy8IuyXPPB2yQmGFN+W1J+RXTjQe7cHHm5xsEDAdPc5wIo
krTfLCwFJBcxH6RpRr7FtNxXTTQj5bDn1NLZFFbnj12hHMSzcZU38agGlv+uNCpN6KB8vmBmCB0X
XqmuT5O0MMaDH3BS++CWjUmUY+kM7WEwWa0GGhBYjdxjeVaW1N5mYOtuQi98wLaqv5NjgsaH3vEH
LxLDNFjEDqt4/vDMuJM6ta26yM7LnkxdgSS2Ecx/uwjnzn0YBsBjpKwLytdqkPLirsMvJe0iSLGq
uTAW+fMOOyZV8Nwigon03q29QTxE0UE3LX0L3bL3EymHKPJgox4SxMOuq8ghgnKwVG2eidw45lwB
8mVuCqk+nFmAroVtQi4dtgKocQOHRV+AklxXYuEHUiHB3lbEyWJyKAMRVUVMdozdB6PKXuvja8pF
ybPjSKnrSsqyv9eDaqrrhXeOydJZOELCBeN9UFcPxVR4HkR+1yBixYkNne7tlsUUa+Cg4WRpdTlF
B2HdHWRG/9siM4uk3jPRYcU4Gfnai6zVbShb7sY8B9PH9sy8eIyucvhHt9W2d9vElB1PtiUBqJ+T
NxPfaxZY82GzcNYAh3+jzjGnwSEfpuOZnEOm7DjHBYfEbmNMZq65rQI5jQmBDDRtu76Wz3HsAD0I
BoG4ckSHIggKjXhEcapIKrQxTj+h5nrkYOeAee/ZxNwVUJZr9OUbj3XiYuPi4XqoVltdAfcg4ei/
bW+ZauHITytW1GlMCHFE64TRp7JgDVFHPrcIv21NTD2qnLre5dF2Yzki3Vp3LWepz/rzuhafHtVz
5EbKV69cLoODrKXaKJZ68Qzu+myWrm2+rD6i1wRwu2OcHBcxPatwJbT1lCBoF7/Uf+6un5Z2BRFI
K4Z7RSyxkhie0dXCXgXpRCz8VePYfl2Phya+uvsZvrAA0USBMCuz6cHrO/mn9ZUIKcTuPjRM+0Rc
Uaf08eFY2hF7AmD2IluVwFpcFZqAPu8BycZTZtgc3wmpFpu6ez0lX3XBQaxZ0t/t10+RDMBi7aYr
0eegK/4zazFGM/QDEhoAeucQwGQld+riw8yZQmjQFAxlKVBYyIMKaYEG+n67lU75xbAceSYdgqQI
qxFqY+5qhvUlSXOiaHr+HCAp9nEKyuk63fLgrZkf/x8vrT+KPCV4f0Sc6aTyssi5qJxvPwSMMV9c
rpvmEQYbRhdZRBa6DB1Asfbw2NG1tqbtF4Uy6Nzd+a761j3NhC61MsBdqMQPX+AA6aJWfP2v4Gph
uoRw+40E8KQMDe2cLh0VccBq2Fpm9QrCZaZivx5y3hiMm/ksZFaVzQyF//OKYoNwEmvhGNRyvOUu
zs0q8DJctL8fhmQ3/Bkyq+DkijltWWp8BtmTInhFd6Kx93ZlFoydy4Axeu/g08IOEjflxfOaaugM
P9sIOEEco9Yg7iuJyQHufBlYgj1QeQSsTBiMn3u9FusSh4crPHnTHbkv4BmG4BhOFA7DHU7H55ng
HCGoXjgX0Rl1WdYO+OjOJuK7Uqaz7Id97lQRdBYztQ8XTvOlVt5zsldhjVRqtmfW3ZQkRonVY5U7
GnlzvdqWdTmUUYi+pF7D1ga9K/XvSYAaC5FCVy3gaOxcuUcaocCI1RAFi5u6JBjrJxWJQ6oIqh3K
lU1z2Hq75YlJi+H9VRbwA4HDsDSKD4z58U6EXbQr5CuPN0txkJ61IDBgc65kvFepb/su7pprQQI9
XsjZJarJD1m6TZnqJSF5ghER2A5rbNgv7GUPy6b7U0ZUU0ajCZHbiUyFuuS56uow4elDc/n9A2lL
O+2KlcPz70pd8Azm2i3kabSObusYQSiXbAx5OYV0K7ZclbAERmrmsFgkxGQhJnh/UljD06PiN5QP
ZXn6FSfRnqRZcZU7VuL8RiFht0RPW954tDEsdHlCqF/xNZXNlNLRJN8iSBdbzpfUuOdZdqJEnrnm
hjzrorZVz8677FydJ/76kmvLL/OyjYOLrzoy+I2CUdz729hsITxE7mEoJpYl7jpejYIkyh+niT/K
JopTtpjWsWX1infeCPNskqwPC02ThQqPMWQWek6JmOtBaUXIUyRwPitFjTrzznlCDCc4F17BlZ9L
49hYOd1W1LM2AJtu/WgWPWkUfUxTw16uCPmWcnDy9x01BECswIWUuQhBl9wbmf5+VRoRtshc8GXj
wMYQ//P5f3gAI0q/fkBdCQ89MU/EMH95LM4l3u1h3Az9/JsuuJ+MbWUSM+AiW2/xLVlg84T7zVZc
Q8i1xZEh1Qj3VHSjyKXrolmwtDGmdVrCThZcEVQ/AMr9nSJ6Hw9sc1pnuxxG8UgbFy2UfncArttB
xDTqjc2RXhb2m9CjMrquqyyViPOzksLVbRyf+uK99PZ0xCSG/dVgk/ylpy44rpbNCq1tpDEmjudf
5SMxH0Mbu3xeG7SkuIqZpyWW8TK/E5NF3UjJ8psvVNNiZWZw4BedJR1xuNZhXBxoxTsUKDVdl2hn
FQbX7dRBBrJJmkZWm1U8M/7dMUcx1LQQ6Zt6HXrnMfGII9NjUQo3FgItxwzuX9jztIPlgCxZcqeG
1WRVYLIWV9pM7COqfZer6cHpLRg/xylJMYsgcB2VH3TEpQ4oclVlJAyE9a7Of58lmXTUAfzwM8Q5
N4Ay+W/4UUz83HH4F+OFFzPoAmGK7nqlAvXCePHIxVg1rV3fUddh870+9nCLp4TAuui871x6meD2
TFnav0DXMKOSOykANG7Evt8RLnI1/O50tZo6XZj8rL9CCEunVI2WQUK+Jtcf5AFb72eUCIslllbA
G9jM6gxNXz5QKocTIac+dQB0pDWC/xOsQjDdRwtmrhU+Lv1upxTrBP2lBYw9rQ4Bl1d/thHfirJ5
zxjPWGFwMH7bdBj48p4kx9GnG8azwPnqQ8U5etXLBHHMbYgyOHmk1c5ozkFK2ww/wDHXJD8TO0wp
1KsmFNCkRJ6U+rhrnd9PEUPJnwc+1/l/woHluzUpXWvXPlqZlIEw3AJVzNgsdNSOB2+rdxG21pM3
6vn8e3NCk9JfOV0rwTZELOcCJDj0rdTilo9NIBoEBiQIQ3ZKxeoKtqiV7aAGFthSQ0Y8v/OL3TRm
QqB5Ds2e6pb0bHToGYsey/+HKGrgmtioy0ZA2hktH80poDQyB19gP6oJIfgDux0bJVO5n7kabgOg
kSGofXDgkOCOujzjXxcncoJQZEOAfaBL4rA1JcSW7u/8fLAn8l9NYKdBpjGgn3E1ipmSJPFA9YZB
bt3oT61yUkngcWXCVX989f0x8P4LoIj9oGS9D4kvp9MdBNWDKtdsnS8Vx/aTEqK4dLYmd0EdWGfW
WqqPKo7/8affDIMWct0InqHgv8BMQNxtHrIO6wiSFXbmzXJ4QdVCyPj/LOZ0WZyK7N/RTH0KCFZ7
DtHt9r4VKyCK334pZF5Xaernv3N2d8a8F1Qx8FRyf7lFV/rrNNruSf7nSVmnVNV3dUcHF6AG9o09
A/dK5u30CJ2/ve6qkBY2jbYpw9Ilx/5vuc5YYalpUUtyyNhqZUNql2kQmysV3SRd0y1Cl1aq4es/
j6qC39AeAf74YnEyxJ4aHIsrfFK+ZZPszAF5Bv1SSWJekUuNFqRsMSrvQ1SrpifQhKP/HHZ5zSaM
JnL8oOR0oufyCyGH82nQIq6FQ5OQ3kR9x4UdoaTONlmMVsVav6kvJ6altv2CbxueWsMKiLh5gcGe
ZcJOtssrfJBAxstCesB1kdrUKIUoUgXr9a03iMDZdpkatwiLOLrXPhH2e5n0K0VZAr4LgSa/llAg
x+qaNcOMfeBrHLBw/Mp2RNGrqxKU88+R8r6yEsS3kZiZ3/tQK8+uz++ip8VvlPrKujDTo52iDq2p
f0sTK8EmEMS+m7g7561eVM241zMIM1P3JkqFfF76ycT3Ro/mKOi12tnXrtIzLFNbTa6U3OWjOEiO
uH3ntj5N3fJry4w0YSrHJGXX13/7EsuPWkDHWkN8ZO8Goojzzn/8UTKKs15Nb/d6WOjswAm67ESu
OPS/K9w8gZl7M2aanNFd9Oqu/CATT2gqlpOOc+mVU3Syuvtr0ys0JgzpsvFbwZmw4buk+NUwaJ+I
M9g0PMbvv4TrAScno7m/UDDwIpvMyGz4zV1o+sYrOee2MEEzZbMR1Aj3KqRvbGGP/VSZBvz09YnF
ZuuDgGf0NiRXW6rKs/VPr5Gn7U3aQQxcRq0Iukck2dn+CDjEaj1bYb+6Pk4xa7zRuWB/092W+NQ9
FcvCoXE1EA2O2O97vOl7h5XadlT+/PHjV72UueIOskZsYSIVYr1kveE3HPEPR5WVIqIaFwtqJRCA
esxEftHCX2EPentGw+HODtb8NO3DyjEo0syF5p+tExZ2MgOGUbr0kK21s/NQ26P9+xzdPK4e8bQD
NSX6tc9+4TqDnMl8cpZ79J2lgiWmT9gvGMyBoBycsz33T7fuPCHJ+tlSZBcHgcbl/XA3/MEY77Mi
OrntSkwrUuoAwVizi3uCtU0bOyivaEULKIJ+Uxsb7/gBfO9BvxsbukFYd6q6ZIfWcBhdVerW9ivF
3OWIlUheSTw9BMSYL3rg1zku3gtFxYuowUK4Nklr1sex6PpCJHQnNvSvqOlVpDyGchfCouhcb8k9
B1H229Cw9cZyQqbpZjEx3FD1f5yqOeyk74Lf2xNFtjmtstuHiAiIRu4247IYqnswa+LAM3+dHBNH
Q6bR/gVCQn7X+bKt4432uut8kbCie1XHvWPWvbV3xx+9gzOsi8oV0VvfQ2hmIzaVqnDdBq1hAwba
fR9pkUSW6sV1SL+ejxqm2/lpqJWfLfYkA5hXJlS1GK9E/ZhrILcfgRuhtl907YLbwrML2a3IskRP
ryLhchAj2zgsSqNzFHlcjjg8H87xjysUwpGc8yp3dEjqX76wHj2C4Q3chjWjRV/JTFr2phOUtBE/
2MgL8Be+4bI0vW77BQFdlZIPfH/Ac9Jy7PCQp6EgjDj6CR/zGP8idKjA0W8o9FHENMVSsFawI8cQ
HD46WbUXHS0VURmIj8RWtDHD/xxVYJ9skwvRNcQy8CIFDKE3pAJqoyUffn7NG8ijrzGWBGTRCLGO
c3+u2/DN/2XPwsMEThUhjAXMv4+eP0Y5Z8MF+ml6SYzgymlZxLvuCRh3nADURVD3AymrFrWE+jjJ
eboE+E1ja/l9ErtYuhWzR3+kXptAm5N18qMDikLz2Gjiu0nfAqRT8aW371GqWC+NmwgKM2MvllZA
A+xJcTVP/Gjej5R/7tGBvSlOYzMrsPLUSGWrMeaMKOz3CudDdGdIoy4l8eEMkmUPnCERlJkgg6ov
pm2miAks68lGoZjfjt3xIjKU2yht0BeAQIbuOGLij0KhdCadNTYWRg8gf78/ftj46nzV0pG/uW2b
8zHWaZ42itExxJUEcCMfvkwE3l7aDOit0pfhLG2G7wvqLpj7FasFoQgwTiV7RElKx9Ug8FqAzFUJ
mDBe2VsQ7BD1JknmVV572N4dlKuCUbAZFpRubBcgfT3pn/rdFo/5+4uL0KWhnNzKH4JkYFJTW0BH
O2jDphmCAd+jZhukM3DC5jtJpd0le0nSTetLLCEOnwCO+hbKBzpS7iJZOVKGzheiKxbdH9bYrC6E
oXQEY+CnNDW3ZsGztt86gES30DkO+I8PwRI7bBxvg8uo5GTVqoi6RmrGiqA9RfttmGzqjKY/ZuR3
T+I9lLAOqmGyTtXGaQotjkHh/bOOjlCiTMfTEcOrKG2SOTVDqaDKzf9AZoLAY4CjULZ18wtnpf/f
3BSuUSpd64tg3g1m9WZeBtwF01Bn0HgEFUj0lkP2FRw2ds3taO+WThSRJtY53pIxO8WSvjUXIc9z
yU1rnsW2qd+JGQYfkVdNzhVBjB83SXGB8vbhbWL/AhBBzFkd6sSSgTU0nqlzSFp/v7VHX17KmFeF
Unf+t0kur8FvAkq4QtfQ2y94G7DBeQq+TjKLAo8ZAIyFIYMLhxauG92/P6PgjADH42LCzrPu6YDG
+IR8zbIXoty28IFUzhrprYgt9qw/wKHgHODAwt1sqgTISr4HnmbL9PKnEO6pfuB0dE212zs05Ni1
r/3blNIZe+/dqBw2UQjQ3X0Gu1V1ZpNbRxPQ6sqrKIRHAtxMxqgMx4ckIXS+9CyftCntBnk80sTZ
J3WjPWbTE+pJNr2bvAioKeQgD+ABaEsJg8Tx91nOfZF7zwpyeQ3I/gf2nw1js2mDAgI+nkh3yHNu
qQ4wexIPV58Mxvhg+OLMo6E3DjdwnyqdQZLTZ3o5c0lPp3agV7Dj7JBCQnPSt6P/8WEmFObHWiwi
EVWz5rmb7jyF2EqDxorgDmEWdukjRJkvlrMtYehDo0JP6mPNCYew88LQDzQj6er9QKMbsfUxUv0x
9XPyjC8LRFJ+hy8hzhqu0xQXsP5EsQPfrAxpGkrXb3zxa4G1MThcH5zRZRQa+J9BgkW1+lg+m+QL
ovU0NVinHwuEo6HFoHIY8GdTaLnjnA2ali/+N9gdK6FXYw9Yu3GYcnYwu0IirwQWHjY7eIjGj9L0
JG5R1z1ur2GgL3/ycCT200+323j3ekKVJW2ye2c91cckJxQtfDChpnXcQTvFcX8UVv1S7SdAQEvO
D9qW4zRjNvgEKoKUWRbBV9cAqciWrr4LfD68Ycr7moCEhpwZt5MHOXJ/3QALcJ7kA6WKntM2gqnL
PrYlsi42iRUiJbo4NvuW7MkvnBAgH/RKwOiOi9qAsgnRl7RTrpxk1AWssyOKNI4fwLW+8+4Q4vtD
yzSqHtANHCvLrwQYJ0WTaJij6Y96g+uHClV/QvMeUq1SpJEOyb5ZagAwqfhRn4vGk5uE//bOLU2W
+QZiCFXJejXw7GFRVN3bzmm0cstXjyQZK0B8y0RqxhE8eETuTFvpsd12ATDslm6jH36BdtlevkAf
uRaxEVTZ6dgwBkKHCl0zW/VmyMkvRl6i6uvb0QhORJ8J+p+kQwPzoiUMoh+8dYPQqrGJINVfeF+E
sTwap84AmfIM5ubiRsDRrVrwXEYpTavb9Wk3btl5YPp+9QJ7EyswCgl2ma0V6AC7KwU+Jis+FTJn
+F345kWPdw5021lyCZjRgKChaK1GMeCv11LkW/R4ga7ubBOKtMLY2vvNChjKXTj0DQzXDzL2VjVg
PB74K3xeKvP/bz14njKgytUWiHBBwnI54CPKjvBdzwRqQAENq511MV/EhmyX86djBx/LCLv05hMI
WynB7et4SyGYRKHtXgcT9aWZpfM0iK5BrnuvzGgkS3MYMqGtjOZXV9CQUrcxFzmiTzeWuSEfAgbT
m96e3PlRoYIdnB7XNv6Wp9GzRA5xJ9SQSggZ+59/1pBXJPis2SE+EddUPXrfOedqEP1x5tdY1uol
N+SmA9fX3PkMTYoEoMqRUg/MvU2cm6Gi03c/1HCXowy/a2zVPa9DUSJl3b8oRapO6mlmkQH3eibv
fN1Z6GFTpUgkA6syxRlaSMQrxxaxltDBVuyMbNGVZp6luG+cZUL0y7djucQ3hNsEJofTYIkeE05E
HTH65tGt+yPrcRdlCciRWkknBNBeQx1b54o2lALeu0YFAa7kOQK/+GkaGMBQx5PHbq+H9dN7oKom
/tJSHnJyfTxi+SZTNXCazDULCHG75/yB19Sj0/pq1LiloXqwaLEw8dvr/RAGgeNaKPk5KadBnNKb
J1L32dzmK7n05yTW3DiQ67BGFX2wydDi4hyOrjkXShP5cY/mwqiCuY0dnACtikTH24gDvoGdiXjd
asezULnYAsZqny/Y3zhyzkxRfKD0gheOxTLeblT/sp/n7rY4j1M86bEVMX4uG14OSt4ZofOoJ0E5
PBpU55tKWZOH1GAOSHqdHuDYr0R1Nwrd71JEAYNlnUjYnXpy9nR+ySX0Xe+Gd6XuqOmArpfEiz9w
Mspgb5RCkzzq5I6fUnw5sAqLvKQ+2Unvdm4CWvOV7GAc4DM++sAITXrVTYY0F9dJcF4XD6CqlZdb
h2toEL6BXu5LXLGfLHnPfGGAaKPvSRz63OQWLMRegRAItGHSHMkasll7w4uNCYLNPfuTD15/5dnm
6d8HbXQLM4VBWC7yy14UNIUlpcfgn1fO5Wkek1TwUxz9mu5WVmefcNv295aAhyKxavWOPSb+5H8H
zVuGZuI7vg/bY8c9k639HrhPpaAi6S7cJnwILR9N/O4bQbzBJY4xuwMXokLXg8NuYgvNqxHx8aCY
atGXxRtoGS/iDsz+nYch3ZRc0ZX29HxmO5PXN8ZJMVBBmsZzqj2u2hlvC/qCBok6/e8c/xBdF8Kc
ojXISwkSkm25BTVwfckbHPLf9tF9XSkqEUjggKUc7Qf9xZYX/K6NDsCJVxB0prUgg9zdk4GKqXqK
i7cqze4FSrXY3YOtShPkenChkJJsYG6niLpnkU1eJZAlDDvaLuKTJkFvkQKkMF1orDeHI6EVZlnm
EDSvMiMyta5+RnhduIvrkj4l8mV1GAWzzezKvZeiQxRPGROl6RB84w8UkeIEx5qX9CMy/FR3go/G
8LqF6nMI7FCaHuUdBWPRwXzwdmmBo4BW947Bk9chjghhkLgEsfkUbImQ+tO0kYnlgV8YlVxhYalE
TQDbyPCwDy5fGBxHVeRR4U9Xu5/pBtUS/j5ouEEP3QUatw5boQwG1u/6EK1fowcRnesAope6H/It
qyPqfX67kvxO0niUlVqBcqkcaJF7UMhnleU3T/CeywDX3dd2ei4+Lv9md4UWPiRC5roiCXkPbL7h
xZHNL6NcXw63tD8jRPORT782epyo3xndb2u8AEmdSEk21cWYaW5rfgnzfK8MOlA/2SVmmjLVFFZd
gDEMZeWrSNk+Y9X4WxSG1Y9lAz0DpDxXiJS1EsKqqg9UaRl1n2vI2iOXiCmbhlAc0Chef3yAq9WD
DppfE6NgdSauhjwSooJga+sRkyjvPmOe4vyKyxY8hviahxWHfyUNqVwBiE096JMAgYAeEqMD6nwm
gXY0cM6rcts7QQupx/k+izROdUSEUMCWoqYQMy5jKbEdcwOaEjs2uzE6OJ122jHROlaDvopQYgdS
kAeKfFLDvfLXeUsCjIj0EhGtk2AbU9syPCJb8+VXrx5cJjGXu6fntjymh+mxmvW3ZsNy8VVyZbTu
n6+KySHGuZZ1YJtLGT2KuUbU6trqGUO7bU/wkFy4DONJDWWLBCUfyilS9MSBEWLALcmKO1qnRrEj
elBFJb0xvosh62srTEdNHUvNd0pjymR6MFlAYAzR5MMGEHvffD4g7V6e5+yAYIISi0Jkmt/Sjkpm
y51Ih3p5rWuahNE0AyYPKY1oycAjh2FID2lIwZ+5kBJg+eDZKoWQQPEqBDBzol8Xq2DLRoPMWQ3g
xfi/9v/NJw4M2zK/JPN8vTJaz/rkzXwrJ5bHeZZJB5j3ekv57MkvbJQODBXpeGvHlrbvkCt/sdqE
jmKldNPIRGCdCROrdWFCV+JnjOY0VK2lUPqB80/awzIgOvP+dBgmMRaGsjz73rxY1+QmvReOAYux
1LbldL0Et33xGLHXvFbRyx/L9iZ/DmcDBJANdDTKGCrrwtxc/sK7+4y/HgM2nsZ/BGIDRrHaES6u
Tb8wLWztBizCKEtSn92u3bmzVBCiu3xWJQsEblq9ZAZ7m7rKB00PrzqwL3SIYiIwv1YzZysPaQxY
acLbMbelnqVdPZOmch9bmVEGINeCgUlRuLCHVMYIl36NKPM1MfYytugoHneOU2xxrRO3iBfkjHDk
XjbxDuuhQLnif4LgLSHWm1RwPiVrChHTtG/d2IcWQwKde3uSpwQ92/j8T5yb0fotoO9WirJKrv9o
dVKJEefeCoSqN8YphzyKgGsS/soF6bLlefcNVZ8/qT+Vmariev5waPbEtpAeuKCQCgSTga+sEOHO
YTmOFP+AFbNDfTswkFHNcriCUyxf6AZ5Yj0jH0/kJRotiTN+3eFvswLdMdj+9T94wBKa00ljMdEN
hXXo4mfYiF8SoBwFGVXSZ2sAKjMcSEa1jkUepd3iCXfjKfxmURlLfGG1848//2VgQeMF20CSxqJw
Rz3RRom+feihVCVgb90gVTlkmnW3i5arVzF+PR3YGMVogPWwjqwDWFeBjb67TYEktSpThY6h94T8
cwdQDR/EFNYzGWuwVJoZg17+MyyQ/Y49RK/pV1Nodjz+tMMTxs6KJdYyKzXhPo7VF0GK0fF35bZm
cj9pmK7LsrmEPEhhvYTFbSsIGrrzETmQSfkeXFEgnRQg3xxpvDPO4QgOlwQ5JCEvfjo7XxvIH1Q4
te0F9hdBXH939c+BL3z7f1shfYKUwJyw82EJKqTvypVebwBVaAzsiP0i0koiPYkwXg1HO6szdRc2
Lvzc5C2g+4bX0oJgCvbrDLXuj/+tmlmFtrDszsRcaurGcKc0cv3iecoyqqIgFmxAJgSF8G8iGFKJ
4csm1xZpB40AWh6JNGHBZ/1lt89dq+u06jL2SwFoPMjMHFOxiO+OiQT3I9HhYEaXJZZjFwD39H4L
bMHh0vvM1yMJ/Rsg/z04wCTwAV4771XUW5RGt+55pq+Gs99n10F8n1Tqtv1+0LmyK94qR3zwnF0o
2QF2oZeHosWq70RQpgMaMFDPm84dLZGPQVYinIc+96QQlfRYrE6sSzAb4z82L4YvSCDT1er+VBTu
FYMzdiKnRr/V/JdQIPzdLyog8kT0Fttop6bx+ZTe/0ihX3L+JX5CoRqTv1qXMFIhuZuz56goRe7h
A4j+t2PXcD/N2BfC6iuQ5kGyJ6KADVtf8Qa2cS21oH/NhbBLMg4jY9ZwH+5pjZfZU53y20TyAOF/
pBLtCmlevPWvpGUYMSd4QEMphqsKOH0cJvxi1z9LnH7clAUuPcThxb/QdEbAxdFpr3jaQN+TtGnH
71oZaIL6zDZKw6NIVibIdAKOpPtESUVl14CgTV+EsKg3SMIuo4e4hgQSpVIk8TGXULMTSPIm+yuF
w/yNWVVxzgk3XKpPFpG1QUsbVcpsCqsEA1jZfVsw/7Ze8iBbQkg9TwcQwuRYdDbpWhkvyCLF4mQC
I5O8c5/ZYMMWesfXNrzZEsVBF2ofDehJsBj47VGymuT4teMamTN1prX5x/tU3yHKhTVDpiYQQfUz
qhRqWiMMW81GNkvUXz5bZV5bDf2b8kkyAA9SyMGzf/u5tZiockBxKpjNxKW9zgVZE4wcwNHFeIiq
CvID/r6S3KgXLu/5xs2D+POR6HTreZyUmAGIZRHCrfPbvmGtZOOi5324zLq/6qqz5tRiWubkl0yb
lib5VQX6SXPjT1d/iRqr6EVBICmhnQ/iO4qo9QDfLuwMbcCflD6jnKGAqjmLRRadiWTk18EuMalh
0nsHcZqg5dJ6tNZxPD7IwafknAX/nUxR4ZmevC9+5ToDPbHC/usdcxDA+pXtqz4UYM0DkgAyH5K6
QXqNI7NZBQ+CEYAvUbzb7HmaErXS3Ylt4ZoHdSpBFBpqRxmPityb+kJBi4MFVBCNMLATXHoHgbpZ
5PCCk5mQIjMbVg5esKcaocDKV94NQFv0VUud/jVKcQi4AGD89fhJQ87M5QhsIsORlLqp9UldF9wg
GUPohN2i2f5WO/K6ZDFih4FffsMh3kum6oc/5CP90NqNc2u7EYWq9aQJbBDpVyVUMYN4lzwD5hpF
dIyp98Ll+7XKhWM4qeX+d5K8gYidZqhMf0IpcqnsojjVioRtju74iRvrGVRgyYO7yNyFkb5FIbXx
B3NNg1SKDgt3kYG5d+/2YnDeCLOvp/twbpRB1q5DFfYgDTGg10nlNkCm+jEezOv2wM0Sp0H9OOW5
t8NjxBVHx7pCn8dNFi0xP7SFN2Ur40/wlvQIvLR0wztPWO3BvpvMASLNM16ivre6rXMwJxHzyj1G
5Dh1mhBLX291sxZo95h4+c9IHCMI088eIxndrziWNVU8YDIaA7MhVgJbi85L/NWQtuXYSg0Cz6Dp
CrPqEwXED/t8O0PT+szqcZBe/0PE+QOp5XGieGRDbff2kJ4y+Ytl0bH11NcUe2BaRCKjIDF9NLhO
5pHX6X8GioH6rPigQD4maFNRKrsRIUM4NmjOPzMaRPUnN19dmAhBJW7xGiNwg8Is8KfbmXC71Wjq
2j02kg1D5F0Dru4Tzs9HIRFpH0ZKCna2uhN+iQGUW8WWljSq/CKcgp/0em1UjuUvybUz0FDmmT8D
8zI2S7i2UaPYyog7E/0e9G1d/d4RyX7uvja1r2G316JJivb8yHN++lTgTRaw/RIcI59sWX22ote8
fGjUu7LM4/tDWIupR8/xCTaXSpM8Ih0MfD61Pj49PMU8UMx7QK6tlQLbWHVsdwkUmg7G1jGCIXHo
IZ+wQzhWwKM8JBaNTCmJTDzJxwcNVNjJHNadrO4oX2xbi2C/M4SNGNg5wwXfrMUY+XiCUqHUJove
q65R7+VSh/l30h+0VWuPCIpzlJ3WGdBwFv8A1pmXP7T+toww5ApC5JswWUf13t8cLK+Y7JUQKHXN
jXpt7bgLS3smVCiffLo6Jg1du+yG39vh+djtnVYa3UA0+oLwnnx9oeMx0zh4sI2BoNjrkil+nudp
hxYItARAIzscp3iZ+oijn0Y4hM81RZD508PIczOGSzgFTK0gCpFxdkVE50lS9F0ApkwJD22d4FIP
mVP9q+qZWI8auH/YtgRU0Y1AgAyF821PFoS+K2ThWXQFGFB8V9FKrStIpMC77H8rXoT0H77uusu9
Qe2Da7hNQynBrQXeEcuk2FG48VSGBK7LgizlxVL2YcMyMyuvYhseRaBkuscy52NKsrXhJ5VwQmSX
A/26UakqJW/3mRrEMEm1G1AlZIhkcneEOcaLYzGaQYe8YvYqdh+o0zSNRAmYNnPfDzPY04xcZxHn
4kkh2ujSzMx85u/44x+MprTADak4uvX7XFZkAvXIma3eOyZ/dyekkR1hJcBboZgcfELN5D57x8q3
i5FnI08PY2RQHdpcBv86EKzZIrVBvAetbBdlf9xaLllaZT9wPshwRMGb7RPXEEQ9f/PYy1ORwtD4
vTR/aR2opdq6rpKue/sFJFuXaGExEiXaLgPUsRVmxfJZvwwoHzPRss79tGVLTfxdRpHENm/rQeKr
/T12YiFj32mS51hRTli+z42aUxe53sEUezSWN5neXPa9HoAJ1Eqj1J6jf8AqXUTbqU8Iv6KqIjBS
SIiI9wX0/xuBQqKnQ5o1/JJq8XMzj4iP8yfvNJ5/DhzsecYU7eDTwd0YycxTkgXrERXHlINumZkO
AELoRMJWu3iY7Py3M3PThIst8bnu45FQ+ywrq/Bw78rwH2TEXvcOAEKtQ711xAijFSzF8b6hOSGF
u7wkp8NnmdhKXfVBFRTPrRQfPg34UthbF1p2+fxhph22TKPIFSibWxwz4kDHtCAZzZPVbXx7bjLD
Xompa24KSAMCOZknLcjnjHWVvhB/hgQUmg6Lucs5mLdnwF8SaHGWHJxIbnuP8XOxRn6l8GdfSr4r
xp5e73RWwr9S6LVo42U4cz0z0DIxlhP6EL7hHOv/4A+j6P9AKb9ruZxze/J9KTlVohxvTJ6EJo1f
5Hc2XqWxwSpR78zmw55qwMHHQhiucTUCF4B6ie65SOop8rILoShb1S+2ND0RVaW/0ebIxfiULQxv
6oF5GEbczR2p0SuotTRg29Hh071zVV0G2Jq63IFDGU6QMVjCdei4CmXqef4AODAytOPkzUBiUW/b
TyaCCGbrASOFKtYG3tRglYyVrJijKabPaHx9tKX+C5/b4ijA0jiKBJ6Px4AqeFYxnD2HW6ORNOjx
cAMvZR0U0jPpzcPtTnaikk5LHZiBgkJp7yMxqp2NNW6oD1yvl4EPVfsb61biYYEFf4GNGmVAKl5a
IbEZTDAZErezJ8X8yFkgNdxOCtoNfb1aClTLNCE//ztfQXNE6htA3wV7kGTH2J6AHqG6TI7Oq8pV
O8QR5NbdMU9+KLlcRdOgPi0xRtYACasJf9LUOQ5TOyj3zABlXEOocpaGewZ8/qou9CAmF7+8sZ1y
WhLZGHakIJWO0xod1sWytPGIabE7yX9utx9mybqiRmROrlP47VqtGSWewbONy9JpAoW22EWXHd6c
uFuiSIUfip6SgfhV8uq2FC4xna54QfP2OwguuXDSV5pcx3mNqWns6r7MD8XogOFikzyaBDyicryK
HdyJcLgbgZ6HtYtUhzd/DUdU6U/y+OiyhKczZX8RzjMgtCNu2v4IU83ljRd9vQU61jAn083FHDAe
SkWaYnREZvqCl+V7Wa1qDH99MywXj3WmRGytFv1bd312/Ok1JYL+K1ngcZmEMn07uUFmBNUW25/b
MrCuRjefWp0tv2gtadvVrH5RQdsa7NiWWgQAuaY0Vg4KSeyedJcJAW7BSaX1fj1WJEOTgVYIA/h+
a042FeTj2eGVvJjZXGHeqn/YY5kyuR7JnfKB1l6W2HHslDHRc2nrKv5EKJhcZLDY5wYFOSpjatzs
ZoycNhqLSy/rWRr+9qzdWcritt4rZ3V1SagWpzYu154t1F8yLA9abw1tdmS6PsGmuuC+eAHyNJNS
6urITvHC5hCxSIoN4bO3U8dPrX9icaU4alHxCjt08LYWTXfiB4X4gGiybrAeJgRXb/muul25G49w
rENbXfM1jUYrKRwLvJK45aId1U7Q4kadrpx2K2njbgfpbso6qJmmn7LXIyBo3aZvlY78gizuXFsp
CWokeDtrcY4qJ8tNKsHztxY16R3aS2HAEvolqmlugSkf05X3LAtsw6TnIp43hHOmOSF0v8QL3172
6U9ZP7ru+npoL3EyOlUF3oLLbZAdfuj/O+UXN74GaeJzokxTRLtrA4Z/zt5fEmcjQKGYQtgm+xGS
B40Qy/ZXdi3N8djWrQ2jdBaMelBauKIE6tt1p0K3wJDmUUxItkmfAxwShcbS416LUq6AiVjNCcVv
a8ba3zUMWcVhL+1Y3czrp2zZrh3MLJC+5sYIsj2M3BpY3I5k4IqAkqA7+rbR2cKKbxsAjKOvTU1P
RkMqDxVVK3HjZq5zVfWYGruaZrzApMal75SgxqdZTSBwey+lO8YHC/WrP4S9zqVTNPz2eSohIQZg
vFDJ5ogaZQ+mMSuubFFNptp0qRigi6CIhtSST+xDrTYV3REx3MsHNI4IGTg8iow0RNrgj9Yr/yu8
qTgu7bowTTPJyALhi4DP5UhRxUKdvki9tZBIX0D3wKRHPaBl1VwgLXOh178urxNmnYLOigxVbLxV
eFlzwzawwVoo5VRnT6AIsbzz6caSrv5sgLDmArv7mOS1pYjfYkGXCQxkrqyRGGtDU7KIuNxw6ev4
85OC65S74+i2GdtyqpwL4+Zv2/pDrQlTuPjKRf8fquYbTSmpK3CuFCxjJSMDXIA1bEK45pSpsgu/
2hlpRjpMWw+qxRDBcefexZ0m4lhuhn+nKaFSeqoE2vUuQlD0udoAyOqdmKjEy1Qq4rbMNZDOapVi
cUoTcOeMmXdB8ChoQKuDwW8J3PbhngvqIcmHdM8EPSM1eJPbPWhCsvobG7xS119mS8AOhX1ijHXt
KBVyXDwTfIoruH4R72oSuTiDQ28+tcmmrey/6lUmBoEB33A30U7VwOl22BVygWAmLJWAFQRoMg7M
0O6lQ8dxOXB2oOz0liIYNVyFJtB6ZL+4y7nzjwzQNKv9hMI4YfKPCop1eY1NxsGiIquhg4gLmQk1
V+0EsYRgQLEWnwKrBMqRVEe5NLst8O8XEFgf2cX4Q6eGGaD1DH0al0f98q+BEEyVdMbpbBKn07KF
kmtDScWCqzEwk6K6pejvUM2LPM4Z7BF4TQc5YgbOc9FyzEi7iFCWfXsLO/RVAimhaT33uKA6hr1b
iQgWVVZx1+3XSzTKZK8FusFZu8n/im5Msg8xX2wafEMTgqEwkP8nLk/UXB2BVbEp5sheSK5umoOV
Ej53PhU10I28khOic9x6IHy7miRMxM1p+YM4Pe+ARuJeP7bnnk2ElUmrmeouYoySFtO+wVXyW2yE
vc0mE9RIIWbUNpj3XL2jimgonugn13ddOc4lRMvJKLf+nMYQFT+KCJUP3tOnBt896wi4k7lKJijp
TJi6KNuOScTqcH0to/jLd/1pdzunETNxAOWMFOsqgImlBIrDCvKfEyQnmmfItHrtEa+8mA6fXgru
/PbkN5CAqjyfB4C86X1jLzmEIlMxOdSGEBHQRaUi6Zwp0xmWU8tX6nB2mW5ybvOvbuDuINjK7IfL
dFQtyGnLa3iAisA7MGBQqnL+8psa2GpzRs5IEkc3WFeQuLsWr3svS1r7HaeOV36oFVcJ3Bwx/XcY
+0jFG0RKUjgBjXB3o/D02WN0AWMlvHmvqo5D5lREx8kxauD96ypt7BKjB1bkKf2Yzk04ZtuEg8x7
3MiAFmT6C99Zhn+/oU2zH4j2dtb3q+NFy5t1qV+yrKX8Ct9wk0tyUgBBNYu7CxPdTWwGs5qvb+Bl
cN8ppa97//7Zt+FDIRWewGxRb+wJJSRoVqvP1KvG1hISFI3DVXASi+bxSOxzjgggrUoADQ0MxCDW
GyYxIvO6XbR+YVJi0fjB6g1tIi7pMs8Zq2cXE1vCL633rNmTkvLi9LAh2T/FYLKOycxw9uKX2T8J
t0JHnpiR7zIenqBwU+gcB+h61KjBQHl4/ZpOnqx0F4q4xKsJ9a3EGW7FW1Uaim6eMSSqNsMzT0/I
jXtIu8oNyWmrQhvZjE7eC1R5gsxnJWidZilnShgaVBPT6CgvUi0Qq4iY22mCA+U6Z1bHUMY+d/RF
XLfBX4ZulwKvQh9PUTxYZdzZTPf6ew+v9OX3BNFkeebGfbHD3LVJviD6ORj5OTn3u2amgi7djpvK
uzf4XTvP3Uq2dz6SiK0OwhWDZPOr0deiFYjY8tu+q9ejQEKIAYATMipErbt5FzpywUjPmoeQSlfv
kadRliIny7J4jEpohhRWuEYoTH5pE3jCz16qgM2WIHaW7vZAC+Hxyo4d4qkLhUIUorPVGvu9Itg7
HWGZ2XWu9f6kBmhIamW70+rfGwdOckAvuy2AyD75iQyE9Lq7HjHYO1VAnMgE+sYNVl+ud3MktWz5
TLNlSWifnQbc4LTB4ek7AJDcIs3Dull/xJ4DQMzSJfoCXofnqEsFFAxuh2M30AeZ4gj90nJMz0S0
kG/RAZ9/w44Qu0IjBpSwFPCxdf8S1p8cemXvgnNvpbXj7UyaAHrayr2tzLEMydms7nUROqEWW3au
Dhc3cyiEYEFFXSClTwlhMPVWUj/CgI/GyiyTpGKU6IawXS856YgR88gc/pHyaTeBPNdr3vcV76eV
ylebTx1GXWkrfUGYV72W30UsbwH1ulB92lhxZPAR+FAJv+eoyrS9sMjtVAtfsJCVtYoAdL3YuPHv
oT+2CePmhT3aBcvJI8+/kiDdUXuRMtqCnxsNXZJ7nb0Hej+lFfCV+ybPm2bECN92hLgh/IqJwwc4
uVrRghKGSTD6hJof2iYuC1wVTE2zeuTZ1sQl2znPMEcDVxKlG5flYo/6opET0ghpx6G7bkzYNz/s
xl6HsEFLlTuc3qpyHZFIrw9czsf2GDvwgH/RyCs0u46/5c3/yau1oqt32SPoAuxM7CVO+Wph1+ql
dqGe9HEir/qvUhOqJ8FhWYpUcSCBDTBcBCgtSWNRdBlqbMTxrK558fuBZLs35dpiJe/ww4DN4iGh
DGsIdIfGBqcjAPsGgC3BikKjjB4vbR8CE7QxKyeiAm5RO4IedAgu8ZWDusXK9dQ8B4uzS8Y9/egZ
vh063c8CPKYihnRXE4HV0Gw0QbePzl7GVGYIdkO2QIpmb7WybrQpTQNYrQfQ3QDZKrFMmR+NiTai
PGZgGuky9PdzlW3NQaV9SidERgHhLOVFFT+h+hFhaygDsio4DlVWwFrGlsxeXD5BweNHTCd/XDyL
GXWuu1m9Ku9gjhlAmIszrJw9zD96/lycEgALL1OnN3mbFkzfK6KZ0HI6UYb9uDr1IqBGut69iG3r
tFw8l4lUJtLiYesxRzWpZeuKvHUmM+/PEDjnxHtz01/xAjfClZ2ebsIbvapmeAHaqw616UYA2YrC
+sJmIyKeTixaY0PA1/MpDm4js9+PQj/WS0Pi1DFTDrc++AOipb59nAh6G4Tupbafrco6gLLbOV23
yoBKc0ZagBb//4uH1tufbcnn+KBxhqTPt98go8wMHJ5Kn/v4DoN1jIAe13Rx2VObphkDFhb4js47
i7nknQsLiwHv1+LsHSKgFaBSNbCe/eCZrDgBnMYLHZ29F9LlQCFsFQMpY5/ksf4yhXuQbKOw0tcc
XA98rTdi6oAbixBGqjXWL8ASkQ3YV3gTMyMXk/+WkPq+VXBj5GC/ovbstzMD00BuZwAGObfFnmR/
1oYmoZR0Lj2LM/alLdvEjE2A6FJNFAqT6Xcq8DItoyhvtcGPklT3Kq5XnAkNJo3U00Ahdmx4I3uj
T9iZjudGkmLXiGVYjD08JnVPjdyHJFVrwajDABYd0xnbEweale37ugh5fp62e7pWY073vebsuenI
72wnbYJO+x+RoJdYucMweevXLfDJg/SMpwtGPWEjO/r2sJIvdo2xTTSvsD45DJ0fSc4D4x1O0aZQ
KF4p73ZyeOVhcndrhZHxyBvJbKF/yTZUk3wz5ZAm1qvi3AOSybRJjeZqLlgmk6RZOTyKE1CJego9
qeFQmmPbR7nYzOwYCfGpBbOxEUSqoRBCXZLCUrAJaGzVoUNLEqla6XQUQX/Pq+RMp2ceQ7onpVcw
3jIM98eTUOI47Rp7Yuwqy1vwNJ3xSMCQRbApUMl5mdx6unzQXRgM+smzWgrkIuGTbHrYd85Q/09w
UF4GyrmAfRmpaGyH74dj6jCt5LjxDGlDER38aX96zmo7/hLFhgreDJQHB0QEtfQPzr2+4YVRRKqP
MDDKn63e2Xsh8O3qd23+drxCdGa705VIUDuucQw5+0MGO+cNh8KJlCAjiI6XTmdiPViC3yQME2x8
IQwsRt7uQWU/lTgNpyfO1F2xm6mFcWfwG+tHC4CqBBgTx5zQShn21dP09C1zTj1s6P/KECVYF5pa
nmoEi4WKJD6y9QzWlR0JFBH0MtSIJygHhpBCb9CfMZoiBGfIe7Ya+PfijDii5dBWqxdoqbcca1J6
gbHmThSsRP1Dnm0RMLqBLdRSHL/9WmNc9QQVo5UUg4sUwZF5RZb+3/yKxMmO4eMXJC5BCaWjp6yQ
IHpO5ZfdbXe+L9Wgcv53FnHjUXXZDRTkpmtvzxwWz1EG3KiHe1lUhKBoCZtQPM8mIlKw7nmjjTLJ
hRuLkIuhC9MBlxOI86MsZP77h7N8nCdPUJq48DDR9ovpMAdsPs80Jrv2uDpNaVqafK7/RxQMfIYJ
qP1+Y+1J94xpDtvqDQfBZ5UsHlTMxbQJvynsUrY961lKjRCOghBwBlz2TqDylJX8gB2x3H8RONqn
n773W7SOJOiyfwToqxbaRWmpl/kI5ObdU3GZC2oaCaRNkgYEkrsCXTgu7k3zhaggpx7DNSwSDP0G
CtFr6GO1SGuG+cx1FPtzIgecpyjTAEKKgeGCpIqTrtDIWoOw5EHPo9P9PTWpnNBPdqz24JA2B26d
weNQPMy3MBLI3VReB0zA3c4D6vwaSSm7mjJI1CK7oQ2bOQQ/lb6Ture8Kado18IovyD5IrgD/j+c
PhaupCj4ocplOWLU0GdvF8KAt7/iYkdzbpIm7HMCeJFwMjO7vzyz/NtDn79yJv7ERJuRjP0TU6o9
Eku7FEW/gAofoGKvG6qLoNd1o0bVStcsYCZJyHx/X3ch/c7+jkaCBF+DLLi+2cLQyQ22KP6BtVOt
sm4/1zfKzyD/WptpSjg8VUPkqSIiiWB9CnWUEhIXmmyCP0dXN7sl+2o9BzyD06J2UbJocg3CVa3O
HsFaQe3o9oB+xBQb/zWGaOQrUBfvxey6T26RvriqVPRrea/I4pIFudtqx5s+ldm238Mthg6zOAKb
8vsT4b2mc562zm5rmL3OpNff3yKTSLSF1PuE4bHZNxVitY9KpL3RT7TLfMzTPkCjodP+NqCxv6VG
On1D/e53BMztsELKLQw8M8DXFxLcblmAu8dg6HCEu6NlDuYlD//te26fUTP6BPn1dvicvhPnbEhV
+9g8IJtCjJ8yh6RjjN1YL6NxyrpC6x5YBPnftTdrhjdY1sTwQDWwwMUKuu9zx77bPPs4eP5o4mXq
bav+a0b24b9OvJXkYunyuSuM2hOiia0YELTet96u8IRUCH1ojLcMimAzQ8ZurJQ2MbPQrzXjenMO
NHF33gN61IoK3rfYgR3K4lSF+kcvULqcZQSAWeIsPjNcPtkaVvrOUDodiraX49htooRVg/703JXu
ADAXUH8zDP30Yk2KeM51jwp23yrHGmFChQdsGbVIvpKCem/qCMw1muc9tJd2mvw4zXwUPcuk3q4E
XEWFaf5BTQILX+JXHlF7SNDgEARVmmTNoHGBSuGUb7+KgoGYTEeQhrqyTUYyK2fZv5qaEHsFEvRO
hkgwHDBKvTlxwz3ksTGHMsdKL1aiPPJdBc9NfSPDXzEAlAFdB3kzWIoEzHsYLE8cMWBGuGDMs7O/
erNXr+jDigsTByN5WHklz/J5VkDC592eJAJduO3OH2kuezbst4Gbn7TIt9Yg3CbfnJZTAovK3IjR
Y3RQyuwzw9JoZknD1BbR7Yaz1ziv8cplaXRaZP3h3yHH4td4FRLaUXw7cgFXTCh0ps+jMng3jtY6
TRdAf1Jo8neDZ2Ow1GrpErsRuBT3z/CX+CxCzhv7bShAqgbpUw7YoG8noZzh3mOkBttD79/00eOr
jN0Yvnk1EhkZb7Li9mMQtRqBIJYu+VX9G+eShfKph+9xbtDtTwieXXWbbuAPxeMUe4bRxpJMIPM5
LmCwzkw4mxak3xBdP1mnoxjKcirAtKZbfMkpIE4cd0ka4sxytKhCPX+xI8o+pa7rFws92CnjerYJ
BRgAzTUjm+QhLjcJ6P1APqhAxBot/rt9/eJuAbvYzopK1lpyoqqynwawL66dYoFVNhdnESg6K5mf
M2eiomQrwqoSeOFoYCmJBo5N6MBZbv9iRP5QcYnC9vu67wxIZm3bNZ8Wc+UE0o8EYsR/WmVX87ok
4kkGUZTLh/hlbcNjqPfa5gAtn72HNhwr9JjM84ahsW8vIX8tQViPZekNe2reuEPIAsrouBiD889p
zgs35v2CXN70WxuY3/myBscVcOMIOTGEKzE/wc1nNwCvTd2Ihk+MADzj2W0/ZSWsXCiagzhIII9q
hrTr3iZXFB9bcv5Fb39f63faaOVT1w10MzBLNOF7mz8Ks6Yi9nqu8PGSn3nF5grI2W8INYc4q+hA
cx2gnx5QkxbMXYOgszHtUN+FN6TyNUzj/9MM9hgJjliXi5rfSC8vxmXJrl/lDl8BEoEBAX+lVhZa
eXoqBedsghak6pj9PfvVWYMM1Xngh8RHkRzMYhWsnlD6PPo/CS3m0V3MpKYzQ0a/YpQTuuGch5X4
N08FV1OxkA84C/iW/eO+CjMuB5HkFsAZ2nR6bjw51CWZutvvbk6v62lppResbwkMUNUQ7LeAKFCm
fSyicSCZIbZ9msuWFec9Ik33I3DMDe7WahCpGtURm6fT+XIuvSEpsOAP7MC4eq+cMV8JrR/4y4wH
n6j0kT5wyk9vEwbrPh84LOkFg1zzv81y4OvN1twjMSNFcEB4AbffPO0eo0PYjWNDeV3EP60C1tH+
tl6Nc4ptptfRqXVlOTXZsdyNUUNU8kvuNgzENz12ZAEoz5BNE5P6Jsz0vNOEyHeG+lRwiUqhXUhm
s0JrDNp4/V6SDW+lIlezKmFwuEDtjvXRTpnTlYVEmPQrhUEJ/LsarOJvtXm4TyLUfcu3joyL+E4G
DbZPEll7f4PChe8l3WcCkhIZyZN+pLvSLeeo9pJKH8Vo8tjBU6saO6VRKnGrInX0lvTefCQ+ewXf
k3El075cVsCABSbMSyn0Ceth9y46Cn/jwOMMBN811Bi5VwqvBkPaOxfxyY5YrvMeKguKGPD6X/9d
L6vED7TeMKN/ELEdKGYtEvgy4jTUUPdr9BBmBjebc1rrn7P106pjJos63FMp6zHpat4McoW8OOwu
4mfM8HcNTwQv+ps5B5ScoYqDWScjroF9S/7cFeF97GHSMgHUYAjY1bzDyLSeYKfoFZ8KLtNCE+kA
orK7oDAxhA8e4QFbX8CkAV8nSzIZGrIHgqx7nfhkM9n/ABg4NiywRdk23TiMFCzIZ6Z1rb5sLtul
xOqwoxqe6+YveuCAXLpMYTYvLFKstXtwrCPx20kdvT8N/5cF8S1xtI7hGR7qnjwSM/D30J5HLLyc
mahcwfJS71epMbG9Q73wtGvR/Hi4+weQNGbJW4r8c98l9zGw5won51rxMjvVP1l4HEFLhdCGBj78
q0VLcCj81xHyyG02Bewx4k44IHmudKx2iLvebB2GW8VjSPO1VgU8CE70roZSGeOU8Nw09ahjdFFE
nhLreHi3UMNXBntU2cflDkLu7hng/m1jPgqLLT7Xa7Q1Z1tBtTJJeHjWRIeKbMCCySN/vV5ahlai
GOxKCeQuokNjMaauCUx4zHsQrTIKO5bJDLZdCjJ1hNo0MOOAgqbHh872JdY0kCabPq5+Ch6iEbZI
3QI5Aya2fhqX4OxqJZm0Vi4BhOylj0nAW+0YKMTPs1+gpEZBMsOf39knm+YiYU9JSe7EwZoUIoHe
7Vh5GR2TkbMAd0581WpBy4qgVBgkowFjaXhnM19KA3Jx4oWFuPTi5ERCzvsZWHnKcANeh1yFtmG9
qBh/ZxOvEMnJ4F/et6pe6OyNtmTiXPLOxjyctoTBetzthwHClfpvbEprldPlazjbacktxumq/hF0
kQK8OECdMTJekQ2s9Wlw9c0alaLjup8O0ttPFyz4beoKFTgIgvcOVvqY7TRpuy6ZEWLrIVrfpnqq
EwRrPX81DXfXeR63ds8YX7seAGpKtRJOcseMz/ntyyxYO34fNgPTxwVt0Fx+aaaoV/kJN1M2z/Af
freTl6jJqISnM19byFimKTjZEO6LSDhvRLVU/XKYs0D2i3ActEeKvKZsKAvKRlW+XmFZqIEP3/WR
bNCh2Nl3OAGT+rr5p9BtQ62wCxYpsnf0zWoGUs9bAdHTiUVDcq7YmQ3RU6m4xXhZuunx+xP0mNcW
dW5x4bUPo3WX3sr1vt52YRINm6uH0hGUcGsoMIO5Ioqc58VDgNKjnmwQ11ZmXDqhW/uQAvWPG/7C
azj0m1o5e7ZpGuzaFeuOSClG5VjhAIoy/TO5TjGJHs41X9cDewLslI2JXKoOLhOY3v2jMrAhnv8G
kI93A81k4HyD3gEG85mAYrw+mk0nAjftR45aGAY96CFEdFccpP9kzRCJN+C/kSaoU+c3dzIu7Il3
dgyMJEQcKQYetv9Hq9AG9kCULehlZNlW39Qhe57qukkuqXyz7qsbo/dh4669L7/1nYK8rgd5W+rn
HgI93CT/QtfSmkXAWYIuF2+VNuolnIzKBQu9iSI0Qi1ldfcxD0Z2pnwEu5kZlFj6YppbYfQOrV01
H+A2E+MoT1w9lbop28DErzTWEnwAlaLhsjS83c76Fszs+YXAxt7qzaUNGl0fatJGkCnKBkEX92kG
kLBXrPVNU/+rkpS/aSdl9r6YiPLxsZcuNPtmSlGGmP5Hw2sDFiRjr02KW94pM6TOhGdTbSB5SCWn
8YXoGlrL72pil2N7pDVON/p3ukpJYdvQ3u+SQnj5akT9XGBZT84vcMJFUkl/EN/H/Xn2LCOulfgt
KOV3CVMywpoOMAl5mveWF2tXD7ca7kuA/OiVEOzn7oW+zB9w+43obAFquI2v5wVruLSAbm6b+XGO
JUKlU9uh/2d3BJBBDeWO646+cnb3kZn/peGpBpJDjR/LRQVHpcAWHVg+osHABTS1xwGK1v6teRIw
ke5ds+7paCVQ9c9oNzq1KC+3c4Epzkwu/KDQUokDRcCDpNvDfRvwwmi6Eg7jEfzMtcr3p3pibW+T
Cv+32Z+VHZg2Jaki3QPK6X6q9WCdCH7CX4zRodBxxJ8yOTowxqGiHNNn2jL8EE3srALrgHNXzhW7
OW6nLZxshl9CTNEptHgVxeWSkk1SGAF6EVUIHyHHqjG+zvhPWIMmP4HQBszsq+r9L7js/+9OeAyW
cTjOPgm9OFPV0XXLarypbAvP9tDdF8OyM6lV9EorogBmNjHWzhFIycHbp64flNhIoDdzKWBTfuAy
gSce077Ww7ZAQjM41xwU0DtQYBbv15AisHrooM/3t59WaBBwcCSlRrVyBHQKASSm25KMPVfOWrUf
pJ5DmnJ0pOyfR7NvYFdVoRzc6wYGzXjG06jntC3BvaFn0MjZEECaguDqjLGIqr0MT2rocZ9jC4Vn
kA2OXLqzBTp6UTV5uSFLj0MwKO5yP3orpmhkjNik4oZTggOS0q3v2lADjh4Ygw8uWgoPkp7J5D3B
Q4xpMEtx5PPYnVxiBmf6E/J8IT/28mUmjYriXFX/FhFe7OqkRYfmh7qCDqNX5f9JYzmF4Yp74Vyk
zdJj3g8s/gflYcb2Q4hYriLhZGDzLO/toEIzWC5u6aThdT+GG/3+qlgNnqhOVS8DXYAlDBjYpppN
gi0D5CQJ8IxB/FbZ9yCD7d7PHoGaWx3D+eRVZc3YLcpFmoOaZtK1IAHlipJ7dHc2+KA2OxXqWCTI
0/aZil9lefwbqA1t6v+PW3V5/MpP7iqqX97FmCBZFcHQ1Ldi+6X4T6wwNVwTJofRRaU7Pf1mDNDD
Q1aMKadJJlAbxwdu+ldRv9sHdUqfgN751om4l4bp7muq8J+1XGN/zQMYNqFDLeuWox2QQPSxBZA5
ja3BqAJjvZl1P3gXucu4zOntOSH6XNx4cf7bPcvvbir4kCZepli/yMwgASdqjbfE+9JYTOAmpnF2
ojMDgFthfJDlcIQrm+Sd0VIYsQuOaW9Wrd1LbSYAxlF+pcmaXXgdzrSJJHrUCpoIy0+5pm/K1rZ5
6B/dGhhUEEp8cIiflTfw9aDlp/4fSvlgHPdkUJGwZ/ZdjjyFeDmd9JCpB7Ii2jKHR5ReyyFeXzhY
X/YtgxfsfKc74eu1Ada0sDO+zYGJXnrBmmptOfNgENC9/V9s5pCBpwyAst0E0WP8TlxvUGXTE63q
hjPRWk3bwXqUSbGmQ/wH8yZEDcvrXCJo9IDzRJLUcK1CtJ8wvxJd4zZqI7CoRPUd0Tgrh2neNu+w
tXI5ViqnmnhUMKXCxBAmM/pdLYQz+KKk1ByMxOUulT1kn/EhniBvDeQpnEW9YKzynaB+3CQJj8vx
bU6Si+mcEQiDRiQdDse25WLp9gejBWxoKaYWURah2YX+YgaFTPvQw/a7EqN4Ne2b5C+8co7oys/M
OgVg4mO1y0WXc3EUGsAsl/SIsDxf80rTZnm/A/LvvUYO1dNnInDeUo3WulAu5RQXfi0dhh0ANuLv
dEO8rh0UAdAYtf8NVwikpE9dUuegT/Yi2FgS6c5q1eov5M7t7DxSwHTEwxfsPyGqQfwUgys85ms4
d8j5dEM6a2xGAMER4NSiHrs9oC4ecUUwp6Wd3AJxTLGCHvBo5r4fX85C+XNkPAUnjS1CNlZSWU/9
+2dci4YcJ1/C6M0rzBaECmcSIl0cArMLG9YZUcGcn75a/67qc7V7H/gm001iQQOty3lNJlakcyPO
iJ1gQqPu5rDyTLz5pRcb+2QdJ2Jx32BvdLSWYV92n1or4JT+H6FsNL5cxSTgVgeZIIbADge8vafo
QOlqH7Xp00HVzj/YV2G3yG2/sjMsF18d78GMmsm568CaRmqvsz8mHvE6TN8DiebAGxxWr0U3i1rJ
acTQCZ+YhQdH9jg43QUxC7xidAjBifT+PL5qNOqpoa1dXQ4rpCsJRLBVabX8B68W6hyEVKcyBGYW
e6daLiBtqse615rueIGMjGGddGvnFGMRVfZNOS+ZRwgiVLZ0LyX4SER+EVbxExPsPCSrDci//9kR
vGWK2iY9qpHcrnwLuQOP3+k+Iw3+EPjJWApkdQNzZPZFzYsOeGdJgq4YruujC3XEgq/GWuYvyLBL
2xLslcVlQBLHuNIKVuyirtfC/EX2bYPXRgn6CkXJidCos4JFqJWshH118Ql5KoUqAzlhSfdvtHkW
OVjGDAVQYJGvHzhIZ4AdTRdXq6C4Lk6xJTLpVOCXoU6f29TRb3kaHF237ubu87qJuog17xfWSX+X
0R3AHl9j9ZLDPY1P/MUYTTm+pv8jNvYmdY3pxZLeY6MpRaz03Z0JFu+VppCKhe8nQ9IbC8mHIANf
RjHcnkfwRIBueP/FIhfqgCBV8s96nfnqWRX2MnvoiMQdBrmLRwcIHLwRgj8pGiwIku443blz54Em
GrS9mBMpOB2zhbOTwiDRTkJBx96L6cplDcEwi3szamhitM+R7w1a7WKSXoLW92CadJXOKJSFAwmF
vUMeGOmBf8l9zgpPwxMvxO5RyHnQSzihJk640yPqbqW2/PKcVCn/O3NuG2FpX7GHA0c/GNFW+eie
duAqQslkRBZ44aTG0LkIAe9vLNfATvJp6+FcpHTdNj2eIHOUimesKG6O22Fg+KsxJAVEaeO5t2Ri
4kgq5lZjXB/7Fm8bGYXAJj1e+nA1DNcFPsxdYN2Iw+YFSMcyP6TOMlGjJVAWnC9U7u9O/NzQ1kfq
95i5Cojhy3rselNvi1PaopPBfsXBg+XH6zyzsivF9FPHLQxGyxAHKMI+b/kk5pczZ2YNO2/pAa8E
SU0mwT1j9+HA+bXBQb+YACvo+MwUJKKXkkByVbWpzVtaw3s7J4jN+0q9r4S3tLKPNNkj/4GafyHl
EHI+7w6WimENzZUgCTH49W/pbkQe+KfAMyOuEoDcGDcCWdKKXjzsBM6U+t9RGVunABe785ZZakw2
lTtirHIxaKZT88rWQy27HMIhljDSNi5xyf7wyBoF3yD7PLwVsoePONDI5aUWlUR+JGukDFW4NEtG
NSwmZzPn5CEmx93YEZG45pZyb156dJlVV7YtXOr+zgEdkhCrkhl9bXdMfroqwvqQ+CHS0LEulcLB
oaw7nqWtVi8EsETt4GKdxTpllvBFmky+Cca/aymx/WfaSYlTzzwN6AmvTl7M1s9Txcf4zr6Fd7Bq
vAhwRES9O8s2pSUYhoj6t53VynpU6I3tjhAP3D4P5ug7ZeuEf6iNYi4M8XQBPGPfA2ucTKzyxlkB
LfY0Y63oD/ITgvd13w6sL0fEnOK0dig8HO6ijX6vppL2lv9rnFN3MGHR75UBDqzEAAO32p7Q5NPP
2Y7rTSQFpSyKkLfMn5cUpzMjE02bYAcGWMCkMXQRk6pWzejxoXjNbh2rUCXpGsewRMmhAKSF91Yp
PcTxOnLJ+yeCSu1+6SyEhip6nJHSkMY0U/QpolJnn/zdQ7s9I1Mz/jawcGcJv3cMJFXic3kIr34W
oW2L8p4P0MjIJzbNK87sSVlph5whHoDu+UG42a6Imdg2DTXaFInUGLepWH/ZqqpMIlqS8vELK4Cf
SvJsEjO1bonse0Y44czd4Lbt/05SVD5VM67fn2I8StRB+MaAwU5UIy2oNYWNZEk+o9A6lv86TXOz
9QBG77aclgKTKhx3JRpRj8I+HxEtbO2CsHDzR5+XQC9VVsfXvWQLMmF15yxpCxZC964PHMPtowfk
hfKHfdBx32RqcxK8MB0zvS6ZrI2Xm2V8EwONBvI1wCVd8Jp29MyyJeDTQokDF1z413sJft4d2uWX
doyNxZQFZf3BHCGWc0gppSxTutuGXkGcQ1ijQ8XtLAIvsWVbyfctDGdj2AJ3phKpZmX/BqPzh3R2
VmIKxx1LgU/3YOtoVLEs5qVK8lYkDo534N6WTtARgG2+yHlNrKrtMEM6dHCiKgJcsSazw5FiPmxk
rd9M9j/rmClxD0VtIcWUD7F0Lt/WmZRlf5n/K4cdy0GKFsm973KWIKpERSlqmb8l9AlLxiU0RM/L
a+XJ11HF8ly6O6n0MHBlYn8YNx/t91WO4PnqPiHTktu+2YKbg4wt4cM4W0T6a5mvIWYoc7tzNJ3W
2OYHlhhuSaiGkEuMA/zbAzJ7P9VxZgZx83AUwSqbpT4ZU0TMhEPlUW3N5FEiGb//M81vFAMVXYYj
xXJMU/dGVsv8IBpUa4h9N0g1xSMAXELOTvoAMh2JWa488PrGZoHr3LU1gQZSaLVw0J0yGFbMURIk
XktWpPB6K4zAytri81l3lP6e0LiJoen8io88SKwyHWNEod5Mzc+j+B/N4yaP77YngpdFY7d8/MNw
XqSddBANObSqSmCT+HwTOgUZRJtqdvRAe91JsT75L5sPY4ps5qJinFqaL8a6L5IMpXCs6yINZ/Pq
9OZDvKpohMeBxRJT8sv4kcalxA8Y39i+VHyZo0aN+mZMpK0PBM3jF6w5n9NMGiAxN6LV9JC/7OJJ
5+IWJ/NkROzzoU3kDoO8qFdhsODH6frfuLUZZ8R+GGOB4Pz60ECHNdax4fxCgtUbcZ+G6x/z5V8n
kIMt+5d4w37gGkJouv8A5Su/I7mKJc2/ZzFEGHdlh6vgMNruyUea00No6/LDYwbihry0oz/9lRXp
peibb6n7gMnYV3lkyMYBPpTZvGaLk/8nxTyEXmE8WECsedVkJXU0HLMHMUpe4VaEESVrnmfug+cj
DNaDNmBiqiiMTrBcPHYpgXPtB+Wn/Y5nM/IOi7Lg1tBUEzK5KqwXPh5BDHBNSS8A6IH+RSwyDMdU
l0KGRmqsjf70FCBMoueqQKpSTmqjmTYdTrmfPKVi5UUi7k8/GvlssU5Ztcf1BdsSNXvPVYh7HTsA
IlOf/m7iQ3Igce0DPJyszot+Z68ZaPISFWRsBMTt3ZNPOMB0MRvCEZVCclfaji5JPsEc4vKSpLvY
12IaH+suKKtQfP9Vb3ClQYhl1vTJuZQdZvLPHVRcy/T/S2/gRDaY/ntApmhdFNfFXT50J9oIqwVx
/ORhPwE4RGlq06g12V9I5hJ/IkRuFKx+Py5w7xr+yxKe7PCN/hF04F4unMS+cC4tfhKZxCXzbQ1d
FbCzRzol7GSoaWTVsgBBdE0QntkmLzqh54TUe6fZOrRwARrNpu05rthXJWxPP7Fcyq9D2roRD5qe
+oaQrS4jFwDyPM3B7N49+EpDPZcHpOBR6odWwqRryBl+BIMjjoWYG2DTfQrLOXv3MTF/DAHTeAZb
KzijTLqPmcv69p3Qj0wUcGX+faGLiiYdSf27hqsRZJd2DbKgbwlW0IjZfAlz35gRGdx2UIxpmR4g
8tcsQ5a/SxB10WuKC/KfBbczPBWhELW9NdVOsFJQVBysAWCo5SaK3NFjV7i46jhO4vDCslFLZyyf
Mljgujxo8GYUwBGBctcOEkgwZZQ949gH7XXUr2VQYPcXCkYzvt4Z+JaW4oVKtniaxVObSgL6Ix0g
eM+crhuJEF5KgKvzNt42b5uH13dIqV3b/4Vfkcd865r8eC+uwlUiWJe6qm59sRd2HQ/JXkUdl/u3
EfduWOYYXgddm/ekmweJKf2ScVJiXaXHCUAb4L/U7oULMuNyALnveY2nNBV/Hku+9Bv/2gzHRLJH
YJ3MJEyjwC4m9Jol9EVaNmpGIkV9wwY96Q2uHoqcYmkpwcLkvlRt8NjPpuOSYRlieruf5SBOpZBD
rya5Tz4KqZvjqC214B1zPDpHpmlUmkwiMxZPsLx58HdweX6iDZgEBPhdEBkS7el9Jb8Q3KrfL0nx
3ghaqAkcRVDV2Q4z3fE1pC40JrMDCpZ/0AeioxK1Dq3So+qdK3ACnZXUIp1aAL/etueGJerRsbId
mzFSSu+URD6JRjLaaJsbLjBJZkG5xPC0VsW5x2fp0yB1tCmcDcqxDq9zCTa+kN2UNQ9Wh3gVT8Zb
8d6zOA5L+EILtcAI42gA+40TvHn13GEBgZTwHczR3h6QRIYmHbf1JhenDcigHIVHci2TKZ59jkLQ
Nwkm6QSuo51iddwuTRDZufDZn9xW/omqPXdftPg2rPuZoYMv/pMsA6dsCmN4A6uWSGXWjhNNAr9N
uojZvnnf6oW7jn5Xoc2ikwfSjLFGRGVYLV6CI34Dy9H8EXengLciKSRvag1sHJJiZ5DxDuWpxy4Y
5Hgq51uA7NODVzQSPNpHJQKBKBEELeZLCtLEowGJJ8AYIGZ5u7UoVCDibVYj+NhsHz5Mx6kBcg+D
vBfgvZ+YnIMV+fbDYtMUbbYyPi6x2gTqvy3tzNij2bl6dlZ+URQYN4ug5yfiCV1bBmd6Mlcu2Qej
4E/JM6ShvR7npHh9gkgbFcu7E/K9UTij26RsxxJPcRASE9IzlIi8YV8IovEI3JXOhwgSzsx9Cwr4
c6UaAP/KwXMgD8xu78Zw+ECfO/Qi2FnYemm5onjX5Qn8zfcVGowZQvpp0Qyn+BY/+Ak4ifVEhh7X
lBcqDV3L9GrpCA4+OYeQHv7cjFfxKHfTPlO3E2I0pe/vLlJ2j+7vJKOvzvhKLwqsHMzraZ4+Hqvb
n1oCxTT4mswLnVYSTV87LZtfA3ze6nNa+WO8QMwG5aHmn70fjHIo0W7NqQuYeCEQKWjyry8Rr6zA
0OFct6sO9h6VPcn52z6nMfVp6tuHhyEQxytnSCqzObydGvj03G7QpTK5m5aTjR3QdYWQ2k6V1JNb
Q4PbwZjzwJKZ8rOGJ+6/sPUJuXWFweWkw5mrgitq9DOuam5piQte2O4L9DfjPhZfH8M8XyK3boBJ
IiJYSHsIFBOtN7qEG3/IH3ArHPOU/AIi2JSxGZAb5Ic7ruWXfeolxpnZbsjWvhRQD7wsTU5kFWAD
l1Y2TZjx0HV5kCQszW8YdV+UjwWkFqfZWyVypxB3/884pmg469hJfn74+8XGoS7ZvK4nyoNQso+4
JvDsa2dr6gNNdBofkiYJ6beKNmT1NOToX2xSIBUZluG4e36VC1BiccY8j3cPzAl4VfQXqB6G0hVG
xCHsJBcFfby/7LiLyLrUAnLaZWjUcL3LzF3oSiuEgsqFUd3sqeT31LLgQ8drPKNewQT1o/58MFcj
NbhgGSfUkFWqWBTjy3KTwceKUgV1sA2/fFqfJOQ8Jd6sSkzcyqWKAnfxNUrOkhX/XV4BUCbh9Z0W
O3MixJTr59+xX5tYW4g92m/Ppj9n8GWUg3IxiM29MXLOMwHavsLBbkPAI50ZpZzJg0xDpkg9tcsj
xKkRi8wND+eqjzAf8sPrVxaKUEE1FCSzNaOm+uulgXVSU5ebA0ow8JQxALTGPOFpzgnn7/BpjtfX
M5HMsb7fdWjwKPZ7tKLwjXrPtwRvm//eVLPAsaUwXjFUwi1CZNDwtuPGE3/MKTc91Ox1g+cYodqO
qri2NXX4REu/UTcW2hDaPYaOHlFz3XiTQHZULUl4UPg7TpSsHz9Ch+2W1wQfSusH0wIuz4p6BHsW
vrPYaX4INUYErBlRtmc8JohSA4teniX0STivEYWM0L7vajmmU42CzSa4p5L4UJwEhsAELjYtDFQB
tBfxAyjNcrwMYu3FGmbpt75anfnYDRQM/NkYiKXRFuqBC1xZuwvW1zz7OPDsvHGoHCx3kfNA4O7i
b5Eq+QBcPzOHevk01HNdvgS2M009grz8MyY1vbl9vIUiYVDwEESvqU/jaGpj7f5jWVeQWuwPE2I2
dg1GrfneN9Yrnr/uc9W6aRtu604SAGim4xFW/AbE9RBxWFmdVEEq5xQJDmLYh9g8+OKa8t6UxY+W
QaKD1IxOHIWAo1I6OIC4/ZUmNfOd0F70n5JodM8ZFhbuRrgKn0pE/H5clan1J4C566vUKZk6ZjRw
p/9U05qwgWTzdxxPys6IzWqat5PD8ZldJStJKLwRtrlk86GW1lpPEpX89nuUBtWOeiSqGKGYwD9J
Iz1+GVICIsrOBZeMIl7APBnqAtpT9Z5UTeeLJA6xOYnfXMYfZ7ldgCcrY1EQ++Ol3bh2ymolUPCu
UwjgFfKODoEVOB85sKH7pwfHE20prx3DwdHoN6aezbLe2qFSdozOmmYgQjYJ6oRHHsPUekO8ekFw
TdloGMHC7JN+UWrtObsHZE+CbBO0P+Sx79s48JRHT0AUBT4hQq78l7dVnvVvdGxAjaEGkFSDitYD
Umxup5Cbj5+ln5kjArlXSXu48pgtDp7p39t48zVWFFySYwLiBPAMpStvgCRSRUz7eqwnd7ODd3Bd
lpgESWMbtdvYzICGFIvglfYevnBXvHccXv7QetN93k9Qv8SgFs55K2y4MnxkgrW6SZKcsa//BRvP
IU78gL0pr7elYfNfZTJm8AUMBG9qkZAwCDrcnhrjlRDlbNb6hOGPrhmpaOz8vIw4e6TfEDQXWFVu
0IN7MYtR8gjtE4Tyh/sf0bIpKo+zPpaW7cQKTP6ObvRS+K45lbti30V933P81PI/cVRP/kFFG1iR
SrTZDfaH+4MTDDQCp3mZRNkbVT3kbRXKmTQ61fjJN6dOdkyy16UdzihzsLxEUJBKIgv9S3p1X50Q
jBlF4d+xOijBf6jpZQDO6NKqe7I+86WZFVQIXtEonGclDVKglqi2Aa6ZS+fOisg9rJt7/EOShaai
L3CjsvheFGurI4QTUqcceoceyhNOsayi5tisEGkxpH1TuY/snU2T2muSNoMu2ztlD4BmexfnEHGp
afjbX6db+2SMntG1hdQ5mECkEzClIMw5JiFtC90kh0+t0+oG9BsxeYr/w5sRUqsqAqqd2BFq6NAd
/NRtnAOjNs9yzT7U11UyRGYFfzprKgZ9fW+uD5KSUZKTtKvIsmfnrcPcOeION0UOlNV+I0Hnojdg
1knZRDoYn1L+EtG0GGfFNG96VPLB6si+gxGN7OSQcHArdSzgyIquwM01+8l2fAQbefyW9TD3EeLB
7LlulYvDeBrSWdiSPA6idh7pvMUSNGk8U22b4PAV1HgoDZ1w28JGOEkyNwrgo+GyfYsXXibrVYYG
laUkwC05aPJXWRUiH7yNEDnupyVursDLnljDInYxWFa67I1Aij3GVCkiETfU3e+344WsT9X1VZ+w
U6jrBauBBFvo14hPFobQR+NnzfUmWK/q+D9vWVesDg7Jqk268G9fkbUKEMtv8j/WlHdR5Fqw3bS0
Xpl+xy41z6Ukvo2nQWh4vbmVpCoD2AuGU6AD0xU0OaF+QUCikIRM9QiRdjb1YE/IowDy1nAQvO2Y
UJ51xdQ57MiBrc+0xWLvxuKoF5oD/jrIf3QffRlbRbxhUuXJPQaUNcSFbSnQdN7Lt7oT3sFj7Lt4
VrZUggzslhT9yyAYDSBsgbbFv1LJd9fXozh9n7zyXo9yEQYE/aByhpS9FRvC1YDwfkzS+RtcEF/g
SdeCSCAd44LjtdaPgVNRZLbWXHMQYZFYQWnl9Dl7XVivRJoM1UrqXVkRLY7Ps7Kb/fRsrm7aXfQ4
KbOATR6F1OCwsoc/rSxt03UXwmDQSRlDi7Wx+mboCEyzmfdAF86Wd9XyC91xDUaYYdJGXNu4Vce5
St0GeHO2MqJJohz2O52RsLVHLF+YqBZ3NI3mdj0C6SEU+ZqGCDLllKxwGELms+mQaqMRrfomx4cS
XJlSLi3BhV4saFa3azuluCzFtTNZ7MAKDrhhyfdS0PPSvDTJOqetUvVqV4/bSiCpCUi6BBtuVZ3P
oyabqEBrnUdj0qxr89dB3E0/uQeL2G95tdRtG7FngeUsUpTXM460gqjkirJDpQ8Tazmh/1G0A9zy
7GcKKJtEmXVKT6hZ6aw7ZlDIhDT9C1hIycv+1ZBOo8/wtQ2f1n0xTwjS3WfTbKRpXFbDTDdvmJsb
NRakJtfjk7zKWslJgLk7a0WwlfFQvHI4K6tY4SGgTq1XD2nC+6AN39lPhXS9M3uBieyRrh0bT3hF
MMzLuSLpnO398NyrD8nO0ncI7H/qXMZZYy5abbZtQsQ5Pn7ZQ5g5B/QgktLEFGRDAOnG/HrTh4cb
Zi85SAFlxYVLjeDhKr37Vuby9gY0ng82zte0pZUei/yRooYV7PjPEi70J2M4Ukqq2bkTitVK6SEb
lOlEONfgg11K3WAtQg9CKdYu6CqqSYgOOQxVbvreHJLH1f3xfYvrm7D1Bhjc4EZmLIQy+nUUculn
xZjOvsLhXTsN5qKR5pSNONmUOznPr6X/tYT4AOq4+uUhlYYjv25DHL5bTTkCjP2jDJWGRnZvJ0fv
lyvulGw1gQJ+c1pG+9a2Rnqf/Mprbt8+wRJoVbrQuG0a5LuiOSvpdcsCtZSaYtoC6GcpliIaK3Mg
fhWOOWZfYUv9shcxs+77xKgg8/ad+vxFno9liML0kpyWsIeIfLh3rnlcoq1vv8g/kqnt3jWZEUsa
DH6N6D4rwoT7iCsQTbjcdPF+Va9RlraTxhdRI4iSaQq0Ha5bqb3nGoi11bRkK0v11G74PEM1zmhp
/krW+edtJCH7T2XvbXxg5ZIgGH9PpRH6E0jEzFLzFu21L3gZLtV7jfuRt75MFtYeS6PysxEes1Ji
foz4kd0EZP2Hq6Fxw4FS1UB8S9O4fqa3XGdQE2PCV0nsaFw9//pqH5SSO65J4FaPfS7NBuOA6jxL
+b4XAurHPVctqiAH9YRiZXH8B2OwWpTMoOf1a3vIt5Yt1DV+Icpy+FiqHZc4Ewu6DBMIgkNoy1UJ
GA+6qGKULZBxTufKrR5JO9ZoH8Mh5l0hzW4qtaybiTu/FLkdacBbxYnn7y68rCXw3XWYIBZHa/90
YgUCbavUO809QMEsxKHLavhyXvjZ96GUP4xzY3Nto9gOUyjXd+2Ql75Pre/wzR0JAz5ivjw7WRMb
wiLszeQIpgTNrt6b0h3zQX8DaKYLubYlx5/bWXgMuaiCrP+Z9ObjB+loHTeA8jYhNu0sKyYjMIMw
gA+0VhvPmO0rvbMiXU67hfhZ+RhJrHekEvmypbDrQpzv3FvnWlLoCUtdFyMHr6LAR59fgWmxT9ZG
iNAULI5SvxJF0dETt4ojgkSY655nPfh8dsG3OtlmQci21xRh/6AhQuqqWemzf5im8XE+PtIGmlZY
BqphoirrPOfsN/5FwDDujxpgT1tKrru74huTHFZnsDlAhXZ8IfUWIY3531FRed827aXvxU2+Hdfg
4xbzwT1ej7Aq0koCmpRIVoh2G1CQkFEB0FgwdzL50sKdURRdr1/VAzjOk9Cdn6COPw2vnr9RUZUF
w8iT4j8dbl7raC7S+7mVAEP9+NynQl6bZlEPBPwmGFuH6s4pGCstAzFDUH8VqVOt36iT8ylitp2H
8lQsul8yyVU4dF4VnB2FIX0vdqmSD/d3SlLR2lzRTQklqPTF33wpMjRMepxHhjZDK5SJfTqbLyys
IjdwZvq70y8OdKgg6YsbmoPyv9+BJM0CMxlGG6P2eFBqqht0Y3iAOga/tE7LTMp40yizxuP4PwqJ
7IxZSAhVhFGQwcmiRGf8QqJrwruD81y9cemtFJ+00jinKnLvRLVsUMSfFNZKVmOtToU25MHVxdLI
NcGkpDFNiMVZAhCR//pwVQk5/fwuAu7QQwQhsYLUuSIJvurjw0w+/ciL+1mHd/D0UWgIqFSxLhXq
zja95Ott6GHjjZzEj3ZtoYb1LC+cnNQIQsuSO/f4cClxdwH1gqI+QbHP9SFMjilHzCPvAX2iHomG
nb9sQ1ZoXQ6sIznXw/jluAqALkytLhS+aOkA3kSdFYpdLS69vnGGcqj44TIidsMifOgU2f9vGNB1
bWF+9Ep+T7UD3TvCZlUKc7WZGIBKNywVaYKSEMgHx/SDYysYijGtm6+wHTUFp6Nz3BDJ28tgWw63
Gw6gpO0VpfGkDjy023FjcxdiVYueUhZ3Kcs6P5fKkkIaS2Nvziv3Y85fKiiulBxcQvJd83OyhKE1
mQXqlAuw+I2rjEayZDmc0adVCUhlTkP55Dz0QAV7Uj9NoSQVcYHtYAYlUuIzvQF0ct2uIpm5t0Md
TbrUEvBjeHFE1E9aqLK3S9DGVT53w5NK4ojfWNwbKwLJtDp1EHn6rb+cBhmBbNQFZ7aIpFOs/JY2
wdvuLn9CXeofX60h+b+eHGVYz4lxicYLPgA6Wxh+GI854une7k93UzFk/uIqWcrn1K6ehtr0Phh7
V02zZYLA7wQ8f2VM04D1VqbAhXcI8WOBTlrxNMAcjgQGGnNp48LzB8yPZBtUeLz/M6PPWOX8gBQO
N7wmrJdMRd5BgpEwwTOQhr1xuhxYnkxTsfRVX5epseQCo1nZxETVaSel2K73gao7eqMOYxlQJtfM
ffCfXvOyFjB2C9QhwO3kWIEVqHVBpSq/S6CTs9+ijMBQM7ySIVdwFfpJmGpUhmu33YOdOOBKEPe/
0zHKmALOGcIp4eDOu8Z/VyNiN7FPxf4kR8RIyESn1w2c+Xo0CZVwwW6jU1yVUi4CA6dD8+Vx8xph
3br7vfhvNA0ZNIjANYMRCCWkPR3jt9YKR5Er/OCNAkrNuoMGlPd18BToyEa0wYbUB+tdsPJ/3PDL
gc0XsO2U8WzHUOCm7+qnw2Bx1MJtQsJTZwxVe3uM2nglpfRK+04fpiioFQXSAUDyWuzTEraSjgxJ
BU5opKHuIaeAJTG/cLFvdv11rbsNulr90SJ2kjyAbX6seLMZHjguMEh9oAjad8NH5BVdlsmolrDG
DGPeRNcGu3qeSf2YcJbxLrG0nmOh7vhMlB9+nVDsQNgwPSVnLSWC9YlKm3NzV1uWdNRnhFYgzgh5
ZtvnOnHP79bAlaUcSftln345H++m/EOuxhS7dQRQ/WVNvz0CwEXPaPoQxoloRO72S0c9dv5eDQmU
/l0SROcKgqN8LPhh3LdKzQ1EZf1Olk5xmVZHLD96iOe3UEAh28fnnO0y9JTiF70yb640ProXzjUK
4mCnkPNRp0UFMnjfgwc36MN2/7BaGbnGsOluyd3R5WQ2AggvEVzgkqXeS9bo/N2guZ+BTG7jaTP0
lHQB862M6dGIYaRA9yy6bRwX1W8DKRjTpc6q/qSgqOEI4v7hxGeSZ9dPpXNeBoGYgRM/5TEG6RWM
vfz4iebYKRl9rxVgVfEXFJI7EwGcaX7xQ4bs0SmYj0cETioNr7+yttmS4p9L3HNBdyodrhVeO2Gc
WeUsIqSumAHiErJMNqdtOvtP4MWrDLs9dcLGA8d9hY8ysS9OrmrjySMSfOY/tT9be5REVUfytJva
mULr7zCroe0zEkNGCWb37I+b0agBo1Pmz7r0tZBMnIO3oelLGNdQkgQFOIhWml5vEDIUS4evaEtk
YOt4CY8OYZ7z4AHZbDqhN3XX1C4jkhGJNQNxfYr7vsXUVOi6y4uhqsWDHmt9P40BCf6W8s+iUfdL
h5PdWIBMb7atGlkbLOTWhgwuggd8gBjoprj/BO1qTvXn/5U8kzRMdyhhFqkfhc8L9uvyNXjdyvsO
nPGhNIj6aJpzffu0hxqDHhrdFd7JJizpu1QRHf2+ybMnOuENeg3NHTlCez8ZOamLk8yEycn7QAtt
VaKHQuuCPSITWm9jbn5KrX7xZzW+V5h2pmlmeRkGze7HjTUBY05k3ha/Dh2la8reru3Iy3lvni4s
CjWtbBizlO01rSL5CZc7Znw+rTnQB1Ffv2+o18u04FVVSTjUIJDJyhB7U8bvN1bhdld2UvMPWaON
KGe/7qnC1IvM143tW8xudLH69sWY+5RrZ7trQxni3EY6IKDp1Dey6ns7zdNaP27mS79qSUeRAleG
PQ0fqVGMe1G+Apn1lXOxSM5EPURpVbI+sC8xcfK3zG+ajcRYz97OiS3HtgAM9MqzXoweha7KlVTF
aoCYZmMLtUMNqvZMF4i7myhuK8P+N89kdvkhv2Ey/LbKfB/GIQKu1fbZR5u1WWWNGIR2ukjhBS5Q
hPVQ0y5SyRK3mWnFFVtscOqTAM2kHcTbtE3peIG5/MqoxJxTcbFhyBlqjFeqU56JYD/EWsPUU9Hs
br+cfghkBompJcENGhkw8sTLBOuYEZXDxnMRVHTyGY6OnJ6Suk+zG0O5UPreYUmYKn/7djHCpxE7
s3FpHP6t7vtRGVR/oriHrX//DzdbqksMs+qoYOSSm6JQrXEfDA3DU+yJaZ/GCD0eK7WnbOgCAdgm
mT92JDkav2AmJYK9ReIs3wMB0yUREt2v/EDVjtpLsTtmHJ66qIAcBvWRA4awsE6304jv+pn7wiBK
n/nsS82mZFCMz7UtBRLI3F9tOuh0eRztNIGuF8dRHYxLl/lObeWOwijrqrSTTYzUZ68FXePbapgX
2fv7pN4vDYFq/xkPo9++XawHI1YxBFHVnWYqrvWiWHev5EyNFpe1esCXYZOe2QfFXosAR3epQW+v
n6Fv7FAAKbKJKVS2DQk8m+7FpY/pdpH9e/lYqnNLhDPeMIF2Udc2jx4I3x9kbI9YEQLQ5h1IluTP
Scg3HAPmP09+sNMu13PZ/ufigVWdh6CeRFVCYi4QgsO7RjX0IFkF5/XXmOSYKbEpyZwn9DXYWx1L
Lj0Z2TWkBru3CS1nTroXGJW7QziUOfB9YBerbFG2OI7B347vZ6SxdOPW43wyCuKZObctggc0QjK6
WSQ0GlxGVaxE6Yro2GqcFD5R9lMhWOU7FXl+mtupV9CrLWfFNN92MA2+nZNNO1GQR+PELINLGIw/
OsTzXCqJY3fNYp75V3/xU/2kKnurKB1gWZDO30/cCbQnFIVrSUPOWfSNKa1Rn72dS8tWRwyVZbU3
zG2U7RIgSh8c4TZBJ4QtBuA9i7cm3lfd3SvHCfJMm1lUCwqxuDUKjvndoxK2mi1bZSzBkUag09wH
JFgSgg+y0KhvWkazcEXcIZ3GSlN/acFPOBiOv7ZScGYZhA2FvL7p4e5YmOzjeIqbt1ZiGbIGN0zH
obzK68ol9nZFcChoBvTfmS9b6KkVSoEbD7YopAThvjUZVe9BlCsrAkUpQ/iptprimch9Es+ETvF2
bfK3uawnFxU8v1e0HApy7oGi8YdoL/gbCy4hH8PGLE2hmpl1WQ6gvUFt0ybj5CBoxv0OFQNtG54a
SzWWT0rdF5IggFbbFOhxo1tWODZMkNhh9wcVeiRLaU+O48MycWHsxnRCo1IEfWTNl/pmVOHC4kkA
LqOopiNY2a9btmBA7LUoDGbFMK53bgmOfieL/fN/z6hQzvvvfHzMd6HQ/Vn8+NQZyYylxJ9Y8d6Q
wv8uEpem6POR6SVfzUUHnyfikb46zjSyZ3zBNGVvmviWy7Jtz7++SUruDjQLlsKtFRmkMg1S6LQq
D4raVr3Li0HufdIcfzNKGbM9FTVZiPKwAbjNvF7EtKjHxCN+j6a219HNDDnG9SdvqOWWX6jtVngn
RQt8R8PWyvWuG93V21kWxQ3wevfHMIpOpfOQ11aMGvcLmo/wSOz08bqqFL/obUaQdqKXFbQ0yGeq
3a3VgH7I6VNM+Q4DPM+AaJ7uLs+i0IeCycK2qvZWceXVyZgJFzwA5S6VItUxTPvRV+js6Hx9nkW9
+4I4JVJf0Tb4eUo6pAYGhS7HOV2TwSox7xYOZ5kyKd6oyA9Z0m4nM3xP20od8qjENFW//UQzVXd2
n9kx5sNw0ZJYVjP9dhEGd9Y+N9vIdA6KXryNx7ug51SwVluZX/EGKedrciH5nCVv+hiw6eR21ADJ
e7OWjOMRb36zgNNfaBJTRm5N3WmIhYepn/mmMPyT01e6OoLxsZfUcVYgySuaUJZiGxPad5PG52k1
vhoIDaSGpSS/INUzh05LXiZbT6zV44FAPJlAHqjmO9eWtQfeIGkeAHLgRJigBRhMsu7SOEBFfnuV
g0pVEuJo9GaC6xn4AdZdOXEjr6DHCgnLVKWjvrjk6Av0x2e5CvJ8z+OtCUqO/pPloh7tOxR0F+O+
o+U63LDwRSlKGoXeTMwNO+8vbeYcBK6t7PpqbiSuUoceOv+uGjw1OG+URXAfzVQEnoOOBZ7YZW81
QWWsTAsZ/baDjN2XSwp5jf/lph9pFZ1bmO25G7e+1QvB4GOtvyAuBSTkSF7CAigjNfP6qbU1tZ7Z
cQsWjh65DWGppCZgwrPb7ZD52WH++bIMcRDvNFG5S8IrEZrSkQp8vgqZeHH5PQgAxPswXj1baqHr
opOJ21nmZUOfDMUCQkpEQwRCY1u2FXhcyGuM8iiZP1CmBKhKRDPPv4X69Pf4cfui0OTTFjviDxG0
NtXTmZEtpc+uuJxTsYYEIyWVyhtpENFmJgW1k0o46oViTRNKCgE1zYXaU1BOMWkb9cuR0bIGIfLg
yeeQZcMyvcCL8yU5QsRlO/nFivxMIE+HWOxMh8dgljqY6p3gjv9jnaMBGzpe0jTc64loRDw4NrP7
IU/KybiOL6U+AVHV0gf5IhVd0dvOvGMAUsfajnyTt03VFptgrTALlCAUKLyv0X0L93tv7/fF6/P6
cRCxvY1XsZWrtxbvhOj31UK0kwO8vZv8z6Jt0gcJ6nUacV1WZhQAbnTrabuTkMWfN3yAmDk1URGn
TQmFheBMlOQOw2InUNLrhIY1Jt4VJmfFhfE14QKUqnNsOqNe0/ZumhRONo5ka1FgTEWJeNOygv5r
ZEtQfWBcs00+FbxcX6oG4LBESjEM55wbAhLEdaTFyJ9zi8CMGs4KQn6akYrDZC/A+5hdaQbgSvmC
01RIFfJlyGcr2ZoOwVpaHpBSeZMQ7T45ao8BD3MOLHlUrdimvEh1WFUQpgY/4ZJRrH193iZ7zKxx
y1xDqFM6gKni4GW0+v7kvGO2BdiCHHeW7GTzjdQVxdas8nsbGjMvQ+Zhf645pdbFZwotPqJHjmID
XBiENDlVT3Jt1RXnRiZKzOxgvBRDXnZzV7ikLWJJaN9nsHpH1cEPaRGCKlAC8FRAsXNPJvJZ+YwU
v5vxQ8XP6qH7rNO9U/OM5fWOKpiQzUjxM12edCk91aW72WOqhx+pe7/NukBY7wtMYNnLj8awK87d
xZxz50iblpFJZWkZ88lH3pT5D+xn4wzfh20tOgD5yG7rxFB5yHlmmOhyZ9QFenMQohM6OC7XRMuj
QkICUCs4+VINyc7xQ1TNtBk1y6oNpEy7LGATZ23Ab/Cn1cWNz2QmUy5QQpdZDGxxt2hyqPYfUomS
QafN/0cqWjJ8of2aFYQ881NPaO8drMHF+zH5/eBGqm7gF91RQSTB0ly7uxmcaIoIn0XUPLSszHUs
+wNc29tf/hYOUZY5wu4Vi9xZksUeLTRFLbn7EBpyxbgDiy74aSAghAZSN0SlShqclHMzb2TYnQd0
suUw44cnIZK7Jcjhy5R5cMNRFlB+dFqJrPftzk9AYmrqh3Ku3urkYYzKVhUD8bZNgwuK/kwDtL6R
yDITm9qmaahxv8vopumrcKBnyViUoIUttG36hH7nY22RLCUa7xOdxTzHROHiAqV90ogH8BJiY67f
7gsdYcs+S9f1d+riDwLdgnLv8+uJUUDNRQBqW7Q3ZpHH2yUl3aAsb956FVL4HADG/ryHkA7nWh/L
lX4KgRV9WKbcUALX3FuwnzQgixCwq1cK/l8I39IZnxQvCEYy5IMQ9qxbas3R5/2j5IGtvYj0ZGTT
+2FWKOWJ8W7yKkRgAnuEwCzU3rF/uBshuiB32Zzyq+gTRejSibik/Naj1ZIylHdCDizg2rQmZtKb
I0Ja+jBf3CGbZ2OgTolfsnYL4fHfVyRGDfwSjCj0SgaXRR5dNyd31k50AaL1FO8IzwUGx/bRn4td
/lqqID1m4r+X24GTosqmRFr9wT8pOLQ+zooPgiKc0z2ty088hzPjMfeiMbWB9C85SU/sl5AjXv04
+M4wk/KTdyf0ESVW0TYrxePXjCo27dUQLm9sYw8jejo8t6zdxbU2W/wsfd3INkxj43IizXffDqI2
vPqH80HRql6llmccyHtZnSirTi+JKgiEbKDRNzEwLKmlerYHCFMliXHoKsAcLwEp2ncpZ5tAX9TC
gnKBfzT2b/+LAhjTMUCiOHerb1JZx5gI3SmQPSbPGmtfNpRnALkRJ6BHVa5V5xM5TZSa//XCOkUe
mKUW9hiNra8rVP4o+Qn2R+JiBbWcfLW28EfGM9Y5x5PKnhs5wU51sjvdpAa2HxtT5B90433WKL4j
JIEAojBG0/fk+QoAtHy3BUhMSTsaBsk24fT64j82B7NZ5qtgyusD7GYHn6bDs8DEa2xc9H9e1I2v
OTtUtD9Bx0OymrqI/kNhQNQ3jvt0BUfj1lps3+yO0BdKr6S0yvLYlmdlfo/tK47nqwuL0IzikUh+
yfH5HjosquzAEUfx4rSHkuO9ZOyZ+vUvIGcfdCb6GplGKRQgbz7BnIwWo6C4HIYOaFpdlw/WozgB
lmS6LXCOteaKVKLPI4/A2o4axVgUu+5Z0hcMN1CQw2xlPnPMLSbV+iuqln7k4YKKVrD6Gst6zOWJ
jBXLb8iQ/dHUe1DxJC5RDfiem7gHN6xkrEzCir8sL7EGzvxbWI/C9CyfkUPIzBJO1COt6Uv2Nu/e
5xgqyNhciZhNU4RtRX5InyKeEmW9IKz14IjNwrGwSeFw0ytX4XAZ4binKIOF8+mMRWj8oJwKGwPV
FYi7Hw+xW8AlKKQJfseXTzvqHIi3t5db5waiXHjcR4JTUJYvKOk/VdKrTr6P/i+90lZ/8z5Ja6kE
DJPAvhPmwCV7D9OhG8bQverqnd0K0ltBr4iOpun+9KPOAuIV/r0FlPCAbOqhrZPQKWk3L1qwacYh
ZRdgHzNIN4i3jEaupWbZTsCe8gYnanKpHxCg4PgtsjhEJ9GU/BTkeEhcsc7cEJy2ZD1f7P+YUIIM
UMonvwjydpvr4KMPYfNVOdvYsipDm9Pv+zhQyfDCOYMST3VQIL092Bqyyb9wZlA17UQAIG6dLL+9
BCWv6zCwv47t+JCeQ5gEuz+Vv9iBC5vmaxEZsj+MeVbeMV4uYdcjPgoCNHMvZZGSYL2xOPu7frVJ
RLgQhOB2rJ7JbEzCob+cnCeJMokFKV9c+VqA5qizbH+eGARsBUK/2UYwOLxkYfBnMxNRkmdnO/jv
2aTbY0l7b4ljDhQsl4OZTLUbXYb4HRMqARZLzMGoCpxHWbylfNCjR9z4j9UeY0ZoXe9f+GPNz4Qu
DmfQ2Nsi5G+nl+rCr4XhYYe6WJFm4I4U5rLRPxpH6li1g9OOVkJeh/LZqJeL7tYv2RalYlHHtUl1
XwdPMDJTCATqYSadI8E1B8gz9kWyZasSt5JXfSEmDEKHniNMNkv+t+vZi8/1Fwqz6UNWxZLMcQ4K
qepnC34q1ToUkjgcg03N2yC7IJulWUxmcMKfrkD9vso9WuvX+ts4Fbl2NeNGSm9z8tVl/oWPcJaw
kTso2zweYrFAUOzNYI0X/P8HxCBGnuzDAaiQmmuWAhkyypWyYvixTMgSe6Yy7nNh3cuWGmjzDhQH
FuI8+GszDQh+ulPqAnc5c+RBoeW8cKggjtyy3rzb2CxrLa2qNwS3+wUx6g/JGfdlA2W4wKE11N5t
zUdvu23FpONFYdoiktRYKeYJqw8GwdOQuwRsjtsxlYE9s+CIfOltxB3XmA38HYLOuHPVbWdhi6Qx
/ldu/gw4NytO1pEaPLOKeTfAT9W0U8qTzoujUnTB9JNmtx6nK6LS4+0MyUHhXOFCO0HtM7mzob1c
gqfN7EvHHL4ap12Xp4elTkVq+vQwE9i0ZUC/DM9hQK6LUxk5daQPdhiGHrWSO0/53Y2ZW4USZmH2
YI4/ew/S/7v1C7HIX1rujWTOJqb4I9l5PimDCbxklcY+Jmw6PfUr0QvHRqT9GcchQ/OKIPOd7mtL
FbCAE73sYF6qFK6i2k0sbOpRdaIxz30AkAYkg3VqPa97LiYrLF+zUfHxh+aF1yhfa4wr9CmHBsgJ
emtC/ttzUhRxrvrN5zc0AJoWGblphEbD/aKU+awPtGBIXJ80w9uMQITvTrrTSojJOGVBkghJz1BL
5vamvQcsmeCLh3T4s6EOGMal9aAPxCaIY1Ko0/Ku9UhRtVD76a9/0CVV6sEj04fQVu28oiJO8S5r
O7XgQTz6bP8OjRtTAisX2SaMAbhT8qXTE6xZJpW4RPAXcK7Pm3JOTv+tds1UzrLzkoNJUZUyODq6
6bSU7gdsfTY6U1s3FEUqMOjGciTOSpO2rmfKEVWknGzgWaGlV9tEWeXsPh0iG/U/M9uwEyXpfQxY
keKpAcwz3swjyojXoooQCZjLuBK8pkkdUwmsjmUrFrYc5rNN7cOLxoHPxedHU44uLHINk2iF1OmS
kPFCvyAMDPBIJ6Qnb6PVGxFEekEeixzYw6IOzjCZmdIprL0nR+C4ModXks66zdY5HljL16lIvoRg
63cwqpENlzmoTDZJuUavS4jeQO9IeTTMHmAlChPIIqUHJ+MAltQL95QL4QjMYyln0Dy5hnAx9m/J
Zf2+nchosnK+zd4D2jYMFp9XEJYmwroIWAwZon+BglzQabrcOsrZFlCCAAuUwKys4xzNMjtKTnro
m7gi1OO0C5sTfh5E2yWBRKTmGIejO6ToRGPgg+3IWSjbjWgeOl3ouw/RwxPJVRdDk1aLrR7Arw14
K6R5PaI9RO8XRiwlJfdD7rYwrfw2iFdT75mRbwOqscoXW4zlxAtatEK1o4U6J+WlrsFk8NuIY/kk
tJmFuciHDS+hcb8yeSssQtqnOt18g3XwB1GP6qcwQpFKRZz/W6BlXOPylB9MjdAosBOyjqk5CNeF
fpfBfUiOk9D0xBUtSVaognOD0fnIxQAkF9J7iJAnvz3NQ51xfoTy2vjQj6mwjm6ibcx9lX4pB7bX
i+ESMQwytSYnlI+oUPB+OuCcBRjD75eYiiY6ZZkssyjVXKzTNBA0jthMDlV/sWnzYtt1aIFoN0Em
KxdXHQIJJ09dv6M4zsEHO/0JdLnhef7v6eRFylxvrKcWbuvJrW0uqOri+7v5wHdI0rTQEsJTJ7+p
nzr5hZZ6/T7arNh/6ZtKH2hFXDJjuQ39EuVOkMLEHAYpv4JpjMUJrHdE1Rj9xFT021aHsbyXut/q
gFJwl4y6L1VL1BfYXk3DKH2O8RPti/U8UsD+wAnQ5TPU3SwY2Au7azy0ompAADWwNpbCDGI7nLWZ
3WBBnjl64yXMet1r2Dkfeo57ZI98FNkFd5yV7EucaAtuOWtW2O7LU9prWdT3UvQtMzQwD7I2/aYv
Ak5s0rPtfz781TQ1ALh+Cuuzl7Fiv8hMTW9NlrksFeBlskSg328CpuS5w30JXqZIXlrhUIlpleyE
SgcEG3bRNBPlBNpyjFaWWusRRF0fGbfrlO6b5O0pg07o32pPQFcv/ci/nMIVf4eVBq8FyH86CdMC
IBRd15khwXyrxeiG0z3PO8tDTaINJHymINOp8hV9gCsWLnmYQUdakzPtghGs9OfhzPflXd5UF7eK
UrSO95mj6hVO77Ye7XJnvSTFg+kkI2SDG9Ib3F5mbKc5sgodisthjIzgUokR+kVHVo7z5fsqpIMy
xpuUN1atirUh1Lp5QroDzXh7VoAEIxcg0oZcmUP7ms5iup5VQYkp4gr/ODC3RPC4aRXtmOWD5PRX
LFe+kgCQ1JR2I4IkbkVFL9zSqZfU4+J8/xK3vruCPSaWCOoPdIcwyA9J9IPbMsDFjc9RP/aItwe0
fKf280q+0vg8gh4AqaP3+9Wv6mfET2dnBlcwntv8V4ZJpNlSIp5hRvSqfbOge9fY05iyn8gkPdrT
WfvQI+jpffkxZzMRIZ4zIQLA20i9GpUZP/gIK5MjfZxSHxuk8q/VhmVSWg1evhVRMICsrtpbOdW5
NOP5hmA2zLoiMgfrrkJl0s48zVoxrFvzK+ADYAFOx0OdpehKbb2kacJaoTdeys8csW2l1Rva8GVz
9k33v5xl9kR64Lh98erEGdKf6Fu7fs6VegH5+3ySX19mR/uY8uD9NqUF+FlaZ+7R1EEowrwtxf6v
D2S3TQ1nm3tb4BMUnMcHGr07wwqViigfeXMS3y5VwKzwSrTbDgrvOiGzUtwjTAfcR5dBhKA7s1MC
VBz/hu0Ax/nxqtzkvL2OZ77MrlUwOBaGTOACl/VlOw29iYypDgLoqIcLjA2Ch462g981/ifbdpxS
BH7dXJHRk8dqeF17sPQd2dQLc/zQRjLxTW39EFGbypY7ZegfP5dVOiMvKPZLCs1DrZwVg82EON3A
tsYrBZZpatCphaKmrEb6K42A+kzA4xoAxwn5/iZfGpFG5xOWxV6jfuvM23xF/zeXyibrU62Pb/HI
f4g6hiaVGv/qN+t0gc9mkvwkT2BtVKOs26GcYIRFuj5cKDQfe9MfFjj/thY8ACT2sJo1Pj62jwb4
qkQBSM67dZKjAChZiFQrjJaFVr7jqfNQXX+LWtW7B11hHDsRvuXixg90E6R99Y2oFdhUULFoGDPo
mqHh3q8c8fH5IIcoczZe4j7n4DUxW24Q40SGrC7wOukCwlbTv8ISEyOIXowMGI2/KYMbg2qpB4pH
cB6LwbdqEZHPk5pna6w17zUFxJo0vmDeVrJn1/ZhIiA23KBqsv69aI9mVocsBmQhavSoD2OSbg4k
dPUyRel3+3e+1AbePMiFyc+2xX78Ck3TkipZNmH7HeCTYce/CSHVJ/SaYNyDRclC6dYySgvg8VjE
R7Fw6DK2uqvIa8gmOE91tzWJ7Kzd9EY/4qmxuppn0a4sHbOkL4INkcu/LH2lh+wuhRw9kZo5Hb4q
zIqrRy+HFlYsu1qerlEShh6SIgAISFDkf67OUGZAfPeEpPEvYcxNJtmQnEtqwU6+q+WzLwKZd4rG
UhxnrTjn0NwZB/hRGsBso4PPLtSc2FAmdaWaJFCHipNE+e+PaCir58pbOYojNMSKYuNewk6YCTpP
YtLDv1yQtrsOBFOOATuJ9hhPERNkqrHYFjCKquaBHxe4CTlLnT9hgoogAaMkWq6AbYu71zH7DRay
leodRAEzG1p8P2ghd1oA8Q00CQynxDz2gUJ2VeXDE4rOGOGRUXir9ymhR7SVhE4jNRj7qQ8myix/
FvZjGTcOTVVlthE39ZAvcmk7pJynLSNFQOa++FDKnyAJGJ3lLob5d7uT6whQaywQhAlvkAFWaZo6
XS7Fxe4TT9ltArrqD07z9RKSuDsozetUPxeCw9O4FjSpw38zLko8tJrG9g0vQeyulVn7609aPRxm
QDNmDDeIdO/XTENjrWTjQucVRKAQ92C5Rk2hMuj+uVpdJ4jYdpS9VtQwOs+7WsbcjspqwjLmOTUX
DjsLI4V2Fv38UOUEhq1cSn4qrgXDee14nTI2biFeQsKIm9347S5A8IzQMx+a68yuHtmKHcVmo/30
5xKYC2mKc+/qDtFnZFTSyuascgbl6hewBBtRK8JD3tknK/lHvh0CqNR8zj7uWOJfnA689M7bibFV
3F+1a5ObRwsU0baJ7v3lRiKI5lCSnowcd7yTa/LZEKP+AQlKaw/8tSL4aZYOgQMW97KNPh/X9PR9
BmX/rIqniCF7StgpCcttO2l3rd7ZFZhEHY/pMWlE1HBq0k1jJOtEKTeR31PNZUZt1KYdCrfklnpg
UryUYkWLSZtHKVQibV7yMmSQStHRH+DL7ibsU1AwoJXUTFfJU6aHAHj5W2FQBsBU+3SXquwxD0e3
+IOBkI+f5p5S1UIUDgQoB7dm8j3cssGsunTU3rHl86tXx5a3mf39zM8aHZMOlyWIrQsEAr0CuURa
/c7hVRI3rkpf3gUeQQWoIB7zA5rnNq5HRZk4PSfotO/I0GDQEWjGYtHWgGjzdnMdnaZ4I3g+9VW9
WhWczfSrjYoxxkU9W7BNPqPD+05iQKlUf5XgeUCdZHX/I3dsNi2+S9RD4/oHH5EDyk3RtgQgJffQ
Vs9nEVTScu7j5G65cWmi6vuKwSJ6TqaFW4KlNNzqr7KnPRE/FTdb1wObhDydj/r2rD8CYq7LStzA
6fyffJwMxOGgUQPAlyb8tnt20/br7UVtovdGB/U8MSQdEwNcmFUgpN3gC49DwZEUvXDC96Ho/wo1
PpoCP1qRj79cDt5+z5CNCgeuuN+wYiahHYgUijx2HXIvZaxsgN/zxhCE3DmbddJ5PBX5Pn09w1kx
d1ZwEpCMyecaIVUPiOPkDrbgbSluU38s2/8IroxhQ2PId9zhoYn+ALKL9LTT2bQQBWzZW3J6DVhv
k8pejrxYo4Uie/wCK9f0DOewSmJb+5A9bvQ1eiLi55Q/KZ2lRX6zBKQpMOsb0IAnYgOwjI/gXr4p
FT1K/71TbMWOVrynCeqW+ATeefOcuuCRi9yz1NR4DW9DtAM+STzxfWEeQKyVIs3gCJ3Q9/uDRNXd
vK5vtQWAJoHZAwCXdG01c9/oEGBOSdC+cl2rtONtMAtaKYFpb+PkApd2dLzNmdrfkrUWBtp1uBk3
T+pgyYNPgA0cj3XHCilBKbHjfU7VU+WZnMxVmO1Z/xTUbH2xMePDEtIlZmc+K3IpzaZkrPRhqRsz
QwNsldIGEAzzoXYe4L9f9mkvv9J8H+O1wzsQzq5g9lNyG1ztWBjbxaDg5F3ZOfiEM0u89yEGFca4
Om0wuNU/k4kXTpxddYRgzCeNGb6acPRwQ17+CiWkUodS/3S2qfactSnM9N63kb2SBQ+dva5eHOsw
TjpLGmFvQ2d8Fly7zWMI07HAbaMnbDzecgH79uuPyGZVWZGfxX0Vu4FYLgqSeIml51YkOWkSiG9C
RbEeKAd9VjK6n+JAxXiBvCHkCk4hFFCJbq5hBvhx2fFlKj6I9jK1LfZjbaKa0uXvb8JEtui1GVbH
BvrJg3KHIzB2nRLJ1rW+N9Yiyjih2pbzjA94YXye/bSrBq6Mm5JTl/Puo38NDcOQEJyDOmomvuQx
T5ShqIC/rdvEsPGxnm3OMsMQF+rjwKDdc8QR3T5+AhgnrkWy1pskkFDuQYZTM1JIl1yx7IveDl4x
gOWYhLK78IuEjlXDNF8HYybTl5iEA1IHaCTBYnv4ooyzGDRJM6UNJWSpUPJkkiAaV5ILSvcWig9q
rUvp4sNVEiQLZbhWVVCeeUWZkY5Mfq1gojgXhTNZl2oQZgAtYR6IlIi1MJwUmM9DfgzemOQp1S73
isvYGUZ90p1R81vwdTS3DmiB+Um6Yrj73OqE1eYvY+d8yTSEyIq/54FsBFzasKpv/m26Q16VUp7u
Y+kf4PFIWkkmPxNkeQJg/0E7ptGQLK/aGNNI2m9NoU/xSUauMpCb3Z88fTSwhnL5Um6Qa2W3srBI
TjSl54AcByIJMEU86oJrBbFUOeWybyulDchhTudtkd/z3LzQzqKRqgRQf05JcvExMeFk8T8V201N
k6BKw75PNkbWZ3zIujUGg7QjYwTF52UdUujbN+Bg8AsmGfjeGkvo5rGxk4XRxOsYRxL80mS5C5WU
FRG6V4RYG4tp+5Y97vRBsfwXhIZK0J2HkccP8SSSNGO+ap5rVovdFXRzGw+8AM331NIK3JbJ2DQy
tIkOyhAq5shGiiW+t4FWDTpLAibA9dl3fekMt790D/iqMxJO2N3ocgS3Whp8mDJW97udzT/4dVHZ
ulxwddv+ffdQ/cO6biST2X/RPACH9DFWIDWDzvs9vI2xwsVdKp7+OCTltKZBypKwqBW7gp7MkDV8
sMhNyIudmKDV8sfxFOI3lBowdt3W676p4Bxzi4+N+CYUqrUFwiUPYX/6ZcZoxp0Q6zGBqXGEPZW+
uKWarynQ8qBRiEBlLn13mXjwkk9YyrRUKxxBH/Buujv4TF0HfLWzeIBEv8s4LInjCie7/ZWtkVHD
9BA4KX3LhxEMBI2Gz7ousnNnvc5xqoPSkbZ79MEEjNE8hRTTMDVct1BqdszL1WmgpEC6ZR6FhgnE
BFmUenuCfd8/aj7OPz8P5HK7Mn/8pWjZTdXIptZP17WaVAoVu/QVp1NpqJZvyngv1Lm0s1nycYyn
SsZu8vsEf6lIR51tDQ7E0KPkJlIgTohM/inyuJbdG1YylQnACLnAkecn/xi0ocf3INUFAZzWW/ev
46kUUFFS6/aDUk6K0+nXeHFuWHboYgP/7/7mp52zCUaAzou12ln3ez2dcrgky2Aus+aqGIeahzye
BYkxxqd4RkXZwAwshVzxx0S4Pq/SmVAh1wxIvM6Ph21V5gXUxCre60Q4BYfwAz7aWx5kirpWakxM
wR9IJpkHpg5cZz5IlIx+5byEqH7C/0IxlTI9LjtKMnJC+RpStXEjQGH5Ggien+xBRJZt2AsmDIZD
IWIVzEWAZ0wzVRgY3G8Aixr6d8YIBGkvjZ2AE4+gwf+CdKhIHlcTUc/p+5VmNb4SDjSBp335hX1r
Scx7ZXg/+nC1RTGTOSCKHdhpRFPHtOvHrlNh+1nVEbQ/HjnbyjPTNIJk1yD2EYSIAWD7ud6aACWa
dHRYxCnvP3in4kNc6PecQ94Ei1arY0kk5wUIh7f2DagvtOELczUvdgCi6y6aIF1RMTzbnW1ksBmI
h3zQekvLRsAvsKUdKFbC8Gna71G9J6Bmoc+dGvtuHvdq7pdxwo5GY3/4407rJ9F9O18IQ2VLShSY
g+3tAqcgUH9QN9s0HWOPpK7ie8VLOL9tEBoP10y0zjgoIoZYCOkBNuoVDcDI/XRGUa274JsMKKuC
T/FW3lCREvN6gvsCz3UAnLVDYRFEp8pN5eBQ+op1nkNP/995ZWEZm+VMiiu4GEumNFwoqrWUj11q
tUIa24jbTg7hhbiSL0gr7uBHn4V0/J6uA+cC0BhTgOZofxMJ1xIerlPUhhTwYw449g0fwTgDmoDW
2BhzfYujMBt7IupRhiJI3GZBOn89aBpqYXjANQLIk0CBV8h/5yeE/2JDi+Z/oKw3R8BNs+7ajFYa
A1gq2fCRWy3o2gEDyU4wKl048BaCaU9K+unVjfPqtPrRETJ4LpAXOAD//Sw7VucNr3kFeFfBGd9O
0DwmmIAD9nbsmvD80Pu1sMyhZowTxYE11zuqpHRM/HNH28hxmHpRbq/UxTiV+Gyr5zt2sQTo1Eb4
BW9TXGClvonGb+Qrohc/6L9eBc0rZOMovOPMesYxFb8QRjew0lgI2FfOIcdTy+ffqJi940TMzVM/
xeWoiwrCdx4AeFuIB9hORIyOP8oM5wAQDGWRReyChUhoOTsbmerLC7IjagVbaEdF7vXKeXihAOoD
i8sTxxF9HCVgWo47avlFlGMcq54E9lAjra1XZYCGZ9gkXUzqeerTTFBme70ImEuweDKsOzt/ObdZ
w9ZEN6pQEOGrJjHiQ8113gkNWqqw62p9/6If79Txg7IBchxKLZanxp+aWJwP6kUbmkUhKdyK7Y1P
LPEKoODvkJKq6rJjaA4O2fnB2u4ASXoC0JZjvh3nmjPzELz2BX8PDhEtt106kFy8SP2BFLplddKP
e8CeTP6ae3OeBgVhvBYMavL/4LkBnuUf2rd554mNhlBqMb30BZqyX3h128V5F5cmLoUacMD00JMi
DJ8K17lOllozQy8Yzw1nircX8gQEbssZRwYlW5qVecRwK2MU+NW9WqWyYwrUmCsZUb3DR3kR+ZGY
NHQAamvUqmEJP+tfqgrkMrzNHJjkV2mQ9IMm5BcL2w2VAYLZj5aoV3/yICzzEf9Hdbnd8BfPd58D
WG7CB92bBIQ3wbAxtAYffzjWOr4/0Kp/n/jk+YfbG97165PF3b2haT/49/5I5kdGoEMCKr5wWToq
+Xmop1Ny8+IJkB7hy1n4UIUzEJkknf96uKtuyXGDykWtgR9KSmd3ug92dXDZZQubZmrGNjHOuEBN
l0T4yHU45QvixI+hJOx8EK9YHZNJ5V3D2ze5fctpqhPZPjApUk9ls4lyo54BD8wCx+b50UtxGRqj
me6mtTv3xdpbFzKTx65hbbbNge+58C1oLh4BTyFrr9IuEKIEWCpfTxPPonSEwhfCVYa1AjQOfjPc
ZabqpP2mR6H9S1z1/3C1bpxEcsrfZLPocXhNtkxuPP2I8I1BwPdcVaHZPkNO0RE1Axxqd4gEgqlG
ZI8I97BbARG2/g7aTvDH4If5abB6+EwquT0NPPOgwTC2h0BR2ncc2jFctXbEFpX0El7ic3NxR6qu
6vSo5NzEU+Y4P9Xs9Cz08YiMTm26Ft+UBr/9FcbXL7d2IqP9E615t3cEvua0CQx2oVhK3gR7mAwF
Nwn/XM6PYO30x5MEt0U5brTQkTJAnTe47X84iyxNj2ZzWM1BtR15fqlg3rX6uGoN4t72Gxpxq9v7
LAnhUsSmjw+qvigTe76pp6iYRpBKakkBwSGDwj6IOnXgICRDmKI8wQcuyZ/h0Py+sVeTD8pi2phj
cGl14F/RMEh8lWC4Co/dqY9XZNJTHYucbjD2flguA/l5413hg8NHp8QEhxMe+3BG8MxJUl7qz8AH
hNQZ3wmsBZPUsxBPFJeY4tGoOCB6e/eR6b3i/WWuWLZeW9aKJX4ek3Vf0Vanx/VOgfDU0unYclmu
Ql9OjKCRsCTZIX9FxcBzUN7wACdlzn7+dNx4hK/KSSiTIhZLjGPY/pKklkq6TMRF76H48h8fn56s
867djjNeP6CVH2GohDKzONmNWCOn4t3DA4jPFR+4sdYvujpTOP42N/U5pmzoOxD7vCZwiA7SfIcw
nEVLrXGSm9fISV/7qgyFPx9LIIZOe9W001xldoCcvRiut77p5mqTiBqHvgGx/2oNdvTMVbJWBwFH
gdi40NlkEJaJp8EZRbCqHFOtNqCJ6wXwPHXw3CSZgcFvG4+P2G+k4OTcTJGAHGaARejWSw7vbHmH
AVSvg3UnYQs4PUDZ2mfZENlyqyRko9JSvVuuCs9NALZfMQ6NEiJPq1AA+cbcA9eKI8BwZ/9vRFZL
BMZvl7q44K9IPa0l0rX4RfdPldQCZQuomb/NddReGWGQVMw1VY1UPE0FOwo0eym/7XQrACOtqlJm
7Yb9xqqPimM0GMMceTl1PPqgt0IJWYJEz5Ekcd5eeCZ/+C4M4yJdyE73CvO/BIN6UNvXR5H2wmkI
aH69DbJo6kBVKYfjNZC7e/IE4rVuO8hWU+fUblbSkghiImLThEuFi+CfBRAM/CDuyawB1iOoFf04
ZhOf6bq0rGxazFFE8RoQtRBFoLty25SjeR5I19YBD4B0aYN21P4Pt3r+zWvjZBkYtkByDtaPtvkR
pdAnOr8sure+omLJcg4Nqq6vg/+xwQF7YAfo4Ulz/Db7eKGPPPQMnLDDSa3bSPWNp/sfK4tiOhtU
sKPzAvhf16RhbBxoN/RwgKRK+/V143UkQnAHNDyYGDw6VxCJi11Q2NJvcgQ1AJvMXBxGnT1qkiI2
5Mcz5WAtjE9vTvCNDa1/kre7kRaJcnX3SSzWsyE+Ji7VYOJOWojgpaNzoXJxwMTeBYvAoK+eJTf5
qvUSX1mgpLhOmmwD4WZlOCYL+RsM/KBrBSxT1ioPEvhxbbszd7VhaXE1HSP8xE0Lksrh70JKtOSn
OSoVrE5wnT42mmCWmuDbD9ltcmlcV97Vf+bjw2xxrfWdgin85bTQhvSMeroYuinAZ1tyrN/hqPQv
GSUmveGYmp3YcnwDu7RE/cGBTBE329GBVDQfX97OSSS7w2dJ0cnlx+d51sKrj6UveIpV0eGLaPkj
62F6SrZll0y1xGeF8ljIsRZzbIlQxqbxF2hemu7rO/RWwVwxntjIt+kOkPx5RQQfdjQU12oq6GOr
NWgXq1/6QFloRJ0P7Uxy7yWEZvYcdmRmlJSwGttt6NcUy/GzbJQUjQCkCGzkQ4ld+lSXPfDh7Enn
BQ7dwJ45AVAuOU0y9qMjDWjqyE65W3+FLIGqNP44v69WzN8ImqicJgpyH3vFAOA/VjNJnZZ32jqp
dmLB9ioSJFCc+bnQVphXfyZLM+Am0nOxgSY9eNQiR2BjNn825BVYScDKpNRN8UX3pJD3LwYik53K
sinEU2TOqdUtF0rtzAgV0dj3TF2IgRuZCyWGFUSCMyujG+sHDtqbNfhk++o8y3N6+zbfxXs14Rof
Fbwb188egWxtE8ZTWMejs5k/DyLLH/QSnTzRGBpMA0E4dsRBu/ACs7+nWEhAQoPDJyv9XBKRTFx+
Bqxn6wn0u5IVR6U1hvUT3GIfQ4cn4zWw1cz8G+SLzfEB5mnUZiNz+EdVu0WRIUOWO8o4irPBIoKL
spbgR7rDlFoXfYEFlMSCV9HRwpvC9uob6EOieY6EpQWpegeJvqEP81Mp3XuoQuhh2l04i8Q839QX
MiIUDY5NAwoRqQowlVe9Q4SaebU7Ce0UZgYFZ/qO68XipjoMQt8voetnNiUoApN+lW5uPhQQEXXM
LjpgrnOi2POmZRmnbYk2EtzOsl+OAiNWGtGHZ/3fJKjNKSn31PLkpx8NMoNbV14aoeraGQEgq7gT
TrF8i2MJNr7uoQGatP5bHqMoXs9IJdEZFcDr0fOlR5iLmDmWkpw+n/Xv8UhWPyrECQ5AGTXNXMx6
Uw9oH47BwPsc4CyXXtPgvbN81P1bLexZYVWUH/H78xbrotUhoqeBcHlz0jwSfDdlvoa+mZAy6CNg
kVLLwqWzA5c/n4/4N1DIuhpSblNwH0ixFa6gpllUCEpKI6qWUNrWVhIyhl5dD6nz643OdyOZS5aT
HHcq27IhvU8Dlpfx75ZfzYHjVkmXx+IxbKoC7Es2H3LHF4DRnea6wuoou15MhL85fgvQ5vXz+0hH
iXPAmeYB0+twmfrmTCqIRXyb8dHebKgxVytJrszmx8narCJXxda2gJsV+z8weaTfXNnJ2Fvbf7t9
+RnsMQfNUDq7JKi5Yu8cxjtAhiBrwn3Lfk8x2v3ESYoPWSvyM2t97RZs0IwZuy7VqeKrbFp3iMXz
WdCRnGbzRfdVAuUzrusF7p0FDfWeiUNe6BGe85yYp//M2vAhWbHi78iVO0YMWJvb9pOWMgqVBsL/
liS3abGE+HEMApVk+JTtPDfTLG/o3l0CwEZgzBpdN+d2nTDm0g4dDPFjVX9eBqSOzKA21v7EyEwZ
oBmTFbI5Wr/iCSh5gEPx3IJvL2N5yJB0DWNHviFtxuSabOelztOKrYmMgETQne6deTqEBPzfBUuA
66sO2QhaAEHOVBipatsmgGfle9mZE+3bONJmJnVIOvl5uG0tabEsF9ilala5F2nW/Xz6sXinA/pn
gDtiEHcP/GYmBPSwcWmXc+NpKSKAPrhNQ41tdcBAayojEZVuR2GMaP3FB8RvT9GU+aYsH6EvF+eO
cOXRtL6f7HaErFRFO3excp2ArHFb+K6JiIYF1zJa7dYIoN5CKoFw90etPzVKJhU6ls20VNYupDdQ
SgWDjI29LjIIrxMHx0E1RtGx11EpHcbc4mC8WNs6mnAFFo5xcRTPnT2IjhtP/+3P7ZsfXxlAOAH6
ZNl6qcLEGGl6NWj38YCggjCMN9+gwHTiTpz3WZBY+vpEgikXICZkUhQepL/Wgg2soLUBCArbfYf3
WyOTmNi0kYK5sPFsFtPbbQcpvAcKjnpG8ZnlbGnyaV3skRPRRahh+H5ZF3ceRUF7X58UMUUJ7a6n
mxwY98kGFp/bygxVG5fgXp61Icr+JQiD5wH6xW3b0EXtRwqUlLXfgOaz4czSRlulP98tHe1sMAVE
x/4jzHYBSiKD3l4+1ki6gWbz+lbmTLKheXgsnyqwcacb1A/91cMtOTkzjQ162FYcg/yjr3uusvXW
NzEh1UgEGq43b8mpKBxWQxMYghqGtc0InPZBZ+UEfY0dXTQwSZe27ZHB5Fg59JY4oI2TtuPfRIdC
ZrYTAN2umJZd+C7ANTM9yraejjXo3YBS5dxpcg9WhTwkQDGRCE2CH793Z9XQ8mSpg/3avvgpxCKR
ywyqMKGjKXpWTaHAC4VW9SKLo/lbTB5iNu9jgkELK5z9Wcpy5llOWBN73hrmgWXwWEODB/4bir/f
FSDSQWPyG+m43K17g/mLD5iavO8rz4ybb60QLj84aBLywbDHokUcRe16Li8efp2aDoGoEMqgm5WB
tloFahXhLIAIePEWdbTRtUpZBqDKX/iAvuHST7bolHG5C8iEfhf284596zRnDesTICDNbuMz/ZO+
pTFPMfEGZ6A4afcACC6WMaoR8H23KIRQhCeHJ4pvwTyUP42o1ZFEI51PSDhVehFxs2LNhL1QZh3A
J+srBmfFsnwljmqsui+5EUB4seOkBWyFzgImBbK5++8/lXOUxuzW+wuticJsv/0FwfbUHFU0R9WN
gUabUnY0ZMAYM9Y254GM7xuaKQ7y4wESYOaL6Sf8NOwc5zcv3iXllca2mLyc9Zes3cRbvYgrOU5O
c1xU2BbN91FaAZMlnRlhLrA73TLc9eRD5sH/Qlz7+uAYUk8GR6Dej4JSmqI6I50EbG2ZHwpsTiMD
4xUqlc1T/4hbOH2l4KeAgBpjG/QtoLDChJxIEQAywhXDLTflF9p12E9Vbfr8Ir85tGnHRROhEZ7J
670hP8D5XQHbumBDwhcXjtkQ4rRzfKKIYWC88hoyEi/laZeoVWf1dVyOiHuZePiGwne6583oPILY
/3E1wYvJejYbNtf9h/JEKw0FhYZGhEciFvOF6wki9v+s8c0BbvLmOFI0ezKvgyVBY6laVXBVUSaW
GFZc5Jqkwpr67ITfVu4aNG2EuLqRKOpKkLyYm+/0kN+MGbIfSGfk6GAPwR2p3MjJ965KzNR7RXzK
gbH7sRLfD00unFoIcbxLsOWHrUitPaPsfVRCYvupIUdoTT03m79B0wIlKj8xM0btFAqfZOmlT6kN
rrq9oXTGLN34u10CLbBGy+Hopnz36zdyCRUpWHAUFxmCrXYKRDkDssbfqp5XcWtBLyRh4AXgyL9W
65bIA2NsZiP3Mw88m5Pfzo80WTch/nEskM3egOPdI9FBu8Uiqm2tBd72snca4Ntos5wRlQml8XeR
M9bvdhb7bt3Rc+/4WBX6KWu1fxa+374H7G/27yhNlurw8BciP+NP9+0YLKf2POMZq0OkW7YwglWf
Mh3x2K5u+FKUZwUGRJLQ0nGmrwcDSuS501fMr46PhKu/Y3zUSGzVmy5Yi5WxvfOnLZp0fMzT+7j6
4Fw4yDLI2iKFPCkBPCSgQVE5i826qoH3TzRnj0uMZ1eND9RNv8cQMtq42wucDeK6f1cgj8Jelseh
TM0GNXJEn3tdKV2xElABpGiJisrOpBCj5LrsypZliGR1FIvRxxTZ6Hr0JYYP1ezj7LN5Cpc63EIZ
GYRcsuVYwjiKrc2IpEgyH/BPhedrF1oMldURyMnBq+7UQ973ogBpGHPlZsr9R2ocRQecrCTkYEO0
mcnWnviS/d/XFZXGEe9CAEZ9R5Iz6ZT947/z9JBa/KFWFPrLnUqMeDMZYq6TkcsxNcBLUdwEP9RA
IXNHV4cJCdeHC1LeAdo8T4a54L+S3R3npMpTEk1ZmBG+N8LWl63MLiBLZ7lS52LYAj2KAgQcykVg
abPgiHSlzdnDTpQdh/Qax+EvGvt7b74wkkOQUF00eaa7buYmj1B2DB3d3nyE7GvM49wTNU9Pdczt
hIrguyWRo5eme2pLxDmf9B/mjuUyo3tNvTuwAlZmwcFco8AcMlYTjtNTAIhbUJQwDWZfsQcbEki0
+F7nS9No7qZlByIoJArA9BQrO91MwKjeXReJj6uI0m24TxwKk+hry4x9JJoUBXUewxsFq8UlymaE
NSVo8jlPXLJHw55LM8e8XSrjoGCmSYGilndM8zRwDD6cAqx5ScKlwTijPdqW4PCnYguK+UpAOOww
DNn7TocRLy/Kx3V6BbfgI1HVAFozG4Kpk9yAMEPKHGvFbZ1pLMhLRgyHLz6KQ8OLM3ZwEK6jW/f1
vSHdY6cNY1615SlIrdZXiA5o1pQt4npaW6WKn+DEqHI3GKqbRdvcP0pSMrnSCNW9FXh0lcd8+JKe
6yR0XjOeoDjkUtBHPGtxRsM9ks9B94/b/KT8qAg9MIe7EPvtOW18l7B1gHv+5pI+iX0UbaHLzPYW
lZhl89e+Q0SPCtV/yMS3QODbe3bR0KfxC6D4U6oKKPJDN/pp7J4/5xbDOKUppwYPXE7+gZ10Hqgy
2hTOFVkIpCulHdpwXtNXuHFcXfBw+e+XlFdhcVwTvncW2p1qqu07kA1dSt6OpqM2Um085D+1oxH+
EBfPXxp4hPfiPIAMZ2vNZX0IAD099xOjtYaFJFYjqv335CuZRLUmPq4sh5FBkyLYn2Sr5qaOBy+j
1hFxwvw1OSdW+9i/UEY38kTqukj3xxK8VEPWSvQKK6+NaNQSXhQ0tTmjz2ysOZThlNEFjv5XwiTh
ubrNJE3h/cvJSfrrRyjKoZxnr6dFC/oemcdLSbkOJYc8oMYFV+fLXcHXBaodyHlvcvxr5K14Yopy
aVu/Ljvi4G1Ap5Slh4TqqpDd9j4IUgyoKZh2+JHdH+NNH60hf6mPh5TjdtMoUdPuL7g8x1rFJ4Pd
QEwbpamgRUfsYJ0SpYmuUFRF0Xt/OQwtkXDaPvSuVCe2Ht0b+Y04LoVI6uopnehOr8w3Sr2axTZV
4iUDfxqx+GgCSauajtzymkPuwyRy8B2WWdu7EQ/2OtEj9RdnZNWwwZnjU+PtTeFh2r919zSdHYx5
nBnVtSopsjA6ZoDhIHZUzKd6ezw8uwqtx2s+6xwAqgUnpiqVDl1Pppb9UmiMMHxwPxSfUeUt0SmQ
NiTdLNmkmOq9n//rx4SxX6BVzqnCNNVTXVDXfNm7lEBm2y7AbgCGYoWDKyPx+WhTed/eTlbUWqT2
kN/YPgIpSU6IpT0EHfXLry8RsR8PiO0H6SdtYW+eoFFc1V7kuuiYqWwIDkn8DnU1FFnjP3uC/QLS
OGeilUop8O/sS9GpjlyKSbG4ceSUiKA1Hh7bEFUlZzheBrwa/az4uQ6CYDu1cpVgyva40K+9n7cN
JJcmFGRaCvWpVOF+sw0QYDU2YhI8jzwL+d8jq7dTE3g2lt/OmL13+WpvakaSq1sPHRDJNr/sLrVM
cSwRyoGCize3x+zvD2aD/Usq0fNCUAQfzVUexYHyWy3dzn7GoDsUqk8+iyu6jf9AJULWrM8/Hkp0
VdbXk5bMP2udhv+Oixt3fJ6Z/nvMM3LsIwnIPn1enO6AkW8USQuyyHgkaBSn5ANMVvXlUPkwRNbO
mPXgkCfXmity089L2erTApQQ1QeEOc9V9bZPXsR4pRolkAcoitS58Dv30PHJ/YIhy3Ef76Ou1WQx
mGhkFsUdtwXPPE9eQ/Rsv+eFtYqrnHgpa6Qy5aF/82+qi5tfnZqtTXn8pPJraDngGkxdSOWDzZpV
5Io82wNM12lOUg7sdbeImY0AaRF7iQGXMQsLtbD7zZDoXuiZ/yK6GZCJDVd7MQtjfF6qNcAIdJeM
707KxoJBx2uLujcfZLp9jwV0T/MJMXBQzkK2EZFn1S3ts41itBA03RuvkVPuAkLuHdCPOzw/WaFa
VkqLyL6Jn15Dnw6Tge8Z9K+Ku5g3NY7/1U8ovnmiv8/YVvTaJgza6LCfLeNwMwrNc0aKpXL0uH7c
jUC1JFOFYfzLlUkJyXwBTWaE7Es+OBt8P+QHuNKzxKzkB3BnfvpAdRObHhhoA+I6dhNyM45Z98De
m/PWoYsNYA2cI7t4ejll9lGENxqO3WiRojyAKFI0Z3gqQg3rWkph8tcOHduf0Qoj9Gze9LsRb8V/
b8D6ahqW6EOk6AWzhIDNFklILpSr3Vmjs2w1QZUtRRpW4ipuMpT1cfdZ/CHPaGDll5Gz4i1Zdw+8
pb4URX/f7gbnCNh5g/1bGgWUjHAen4ksprh+iUsS2CZPuR1mJV2M70liRdM2MovBaRljS+2+YG5C
35OCKI3Z6zRy8WB55VKSUgiwq+E4nrRR9HxLjpMskzBMc35cj49oYtdUL8rxH5YpSw7SbpkmUFIq
pOOkGKmkHh8b4xDBEX0VrYe5z4LJ2ZY1QSlBAxEHdrFF4ekfYPKQcs5dJiL2l0uUG08ZXGCnBk/9
52hhsKnjVUBI9ALkvYESwuk5DNxy0k4pp2btQ8AEzu6AV4XGoc7UVuWRwdDEckPi5TJNx68wqmkY
VaeK3ijDimLLMg1eicw4FXcIWdA32aHmRAs6bXfeKFm/cUrPWnO037qvXgHy/i0P7gThPFl/VJFg
cvU6oEZ1tWyPZKZYv8wvYoOffxrKUWzsOxqLkV3jkIMq69Ei2ZjNvtmwO5aJ01vlVWOt27wHU4JW
QiS1/PcVLQLsmwL+PU46naEz5Xj6l2abBgZatE+Pb6KE0YwKQ02pC68sf2gFD4BC6kawbuacURxr
34fFl7b29uKAPxZEvXSAsxJdeoJ3OJYgXgsv23/UuTrB9NaTxaRrsdb67eSd48dgt6UXLb65Dgbj
UfEYdI5YNvL2yIp7CJfYTA3CFg3gupleKsKrmrtheb+PnGHCR44dx5V5SH0SJ8mZoRtop6K6b9zd
3F//gIjHjcWfv9ExlQa+L/BZwLMYwejId9wxBKEg49WbrJ5e2sHUNzMe1TRL7FBFgVqiHGP3+49T
LvoNxJHBUuthg/UARIfPICGRQZsEwiSdpLUMAusY6ORxE0X1tzrFsekfN22anLf7zPLuHeb50vu2
9mSy3fBSL8vG1h5Cdc0pPvEqJMDCZH8TjwMCx/NocUsBCRvzr/4NtycflWLnAitVNzkZinrD+bBM
nMphdyWbtkvHfK1TfX+X3alufEOTgRNNPJIHoY8CE7bE8wBBSSxy3q4S81NdYhTQJTenhho9ncEM
eP7wL6bsDtQszwMF2kha6RLOTC9igf/Vz35sdFtYNpOXVBIzQ7mJgQPTQ78pGL+5kSm4XftMiltm
/SyYMKXFUQfwyJ/1qA0aSnOJfGeQ/xKAUvyl+pXSQIS5cPO3SHBPh6SEg4jQ6edX5nI2tjAbLx75
4qtigfBaooWY0waauxghDM5gajt/vA3VPg9/FhsUHE3FbswvAhkV5XFSfvDJY7IUwEKWESSvPaNd
O6j9BoRMJvR4QRLa0+bhZQFbTdwNATRh/jVwYU6rJuxtkGkjcHB770DPtEISQo+UzVmG+xoRs6Mh
3lZcig/hJ0EcXacoh8aAKLCxjE4rZnHIKLpGCa0aMDg3XTGDtKwmQd3JoYLvyJ+q8NcaMOsHwLAt
76V2WtIwwwkY/AL/v2UPr7dx6H9iJy9t7AONcWFVqyMwtPgTND13HCW2XwqnvJwJDJngcIMkjNVz
pxJACJ7o4uZe8fR5dGZ3Qn1VPuUCb5rzZ2jfh5glZumvxt++wwlux9Jhs0Zb3PhNI/ZGo2tPeYKE
iMF2tsjN7Xi5HxchfgFOweCIHUNJc7QAVKsjhKyrac+1sr93Y76r6zSH6ecvxsim71Su9L2XS6C6
4KnGq7hGoNVnOsnhn3PrVtyTMMPEWenq+sE1sCk8KgXJfLZ/7LhJBJDpNeo8pJmgY3NJbo248sqR
VhUyM/FU3wDAAJlxkeapq/vr3IdAyhaOyowYGk/VDIAU0hxa+35zsZGku9WiutyuxTRgURQcIzU9
AL+eJM/30W1e4ER/8olQvwOmWnftc+C4bM3S2MCytMKolgbyAHAoM8eojOn4Z3MBksSLnfbLP71/
PCRxfWNJ+/bo7nxlP8wIIKJ6w6CpCC38MiD7e8EFWhsZU2pHgmeN6qi61XTOX/Dbj76wnJTyodKB
4XgYUdVWU88OpRQxVQDXVe+vtZ+c3q9M6sU4uyNf7Xky2nZBF0cDMwxVCwhVwD6yfggYgDLVaoCt
56TN0dyi0ZGyA0r/TqVqoCIPqE1npesnQ/PinyOG6JDGvdpyPw8xPyFXZbZuPRkRPb8HxXrMUQRV
aTuw50oQx995PS9Xn820lnf3EV/CsNDoTqQRLYr5KRtrmOCapQWAtgfB3vhLuaGG2Swf5EbAuunl
59AnV0J007miymG/DqkurNV/y+X+hElssOGd+q+Q2pJEjzv6ujLnnqnxe7Y51GK9lnnkzxswQpBi
qlEwuA5f91J9rAQDscFkr+I+t5oCMmxiqtTT9xJUeQ1ARW5/vpsdtgC/NHDGEmp7w9CQWUwfgQ4n
KMyHt3mdyUm0UQGDy/9Uujb9rZEcOxrHZffRH6KZdf4mBSfj/Z0EHw4hhmJJjFWZp8xhSSgLAdTc
Ktm1maNEFBwj9V3GEtkE5qkvH17sOZc/ri1UQmvuU5Iroqwq39gIjE3RcCRvR/rhxRx88R/lrP6U
0UEGPk67/l+2QamveJkrt0s5mo9YqHwUJRGtsaHre5CQVLsc4gf8j6gPuZr8nkMGtxINHnSMFiaF
Eyho+OT4nAJ5Xh84M4DprTk42xYJuqA6vXf/agO8TtgpLoWZqJ2NkQoiBufT18sc25p7NNP9YEA5
X4a5giu8CxwdXhyOpqvqwRm9EHYNRaB9R1g1JfZb615bV07WQAvBLWoUnJeJVmzE4OWT02KGY1rd
l7EKFjL8YzWK67Nn34uZUl1uZkOz1yeCC6mPIg6LhDVNVe4PZMmCyA2djBUlH4EvU9Q+ryi72JDN
SCeiSEklMv0d4z5ENe8IR/mBMkES8qx8o6xllBNMUN+WvKrWaJ1Ox1Pf15yN1X+g7WSsVGkeeRPW
/33UPt/Vvyqzn7XBkM2f89Z0d4ylpN+V/qG8baaYOy4gGueCY7SPSjZJ4IqdeTL0aoDsWb1nU4/N
tP5PEBXm44xZgwLHxtdvPn9Om0VWFcdFNjLXukLnozKRK13Gl9qmu1xAJ9yf+pbXCvRtyceQcI5T
DsYfYHy+rxIfGB6Gx0FoualpJ6yTBs2l/7ateNTxT2SR60lm7Ou6QVvN/mdw/K2fXec/V92ygpdJ
irPTDuQ6hmRrrfeMRNJP5pDh7eoUERNU2LoOWPw8BeeDDK0zeJ9NWO/7kzNJLU9B/s9kFUzPhTqL
dnotVvVO8eQoATKb14WgZ9O6mRqsgobFEhyT2EXowh5buN0O1848K5xSMqFB22Xlot/lKA72SMco
fhO/OkiJegPVqqIk1bXfA2tVYS2jl4JAireNs8hHCEvktJOiwuS08EjMM7Ev05N5KX1djyistz3D
8XTGDYN6+Yz8MiZhhNZYszOyOSrG+2O7fzGoVKRz4wqvTRT0y7Tk6ybup62KnPpPijnwPmS9b5lb
q57+8TAOA5eHLGWhc0S68UM0Zi/HjOnyr4GRB/8XVWjT+NIvFRK+pAS+PMZ20mEEZRq4+gHcLRx1
JsIwQL21xstksfoM2UfghNHglP+vxe7KSj4DJE2Q0Knio8hxUUjjg0I7dVDEmPsfFwPRGThSGu7g
pi6XTyGBNqg6GakXSjG4pKHg0MEGPmXeKvI1ZvUsIOyJgmM+BpIhFKJyOJ1OkFx8R/qsMoEpGDn8
Z8QSNnpNvq03d7JbBnqn9sb9CbtisLIWJNN8BS2Mgtb0ALNOBhgHudMVzQ7s+MViboJuukVuNFeb
D4M0h09jRMjc9ukT1XNVLDaR1NX6ac7ej/tKa6bUZ6nBOFZFcsH7MQYnHzh1jsM5BZiHI3A02/pr
rrsrxax7Pcsz43NxmABhiYyGJQ5LIwxNEL++zNCLAKiHD8tHLjxlzEf/vt4JGMRHZDi7tnyt4CNI
ZDNdViauFz5KEQVIsCq3DX45jYl72UlH7s9OCZU6kAaK66B0YZI7W/RlpNOxHrBYH40fWD7dT6Xy
SMrZXeJNkiCL4AzoE2MYiKIGmmGvW+Bivun4uTBFRGKHt8fZuUAmptS+CZfEkl9gEf4mxGDTEYf2
S7GGG14FbRwu4de9yUmOkBgXK46VH2U1CtBR5/V2cVfpaL3Qoe+rwPwmTgqZA4wMJe3l8JoyFDIb
RnWyB3Z5jspFif6w8120aee3Tp17oUk1eAsoMWVslrus58q88ucAgI2CIhwj9LoMuqC4WQ0xjTRN
JbRl+4LCvHJgujCJoHS6ASfC/Nj+eppgfRoK2BJxzA4ewqEErMoH/AbTzR1maJM3JSyEc24z4f7f
DuTmNS9qZZ0mvINI/Pg6THsKxOE2KmIKwDLtlCJzKDLM0SIrYL0FoUOb96FqJius/W9EKgoGfq7o
o/RxcKhaIjnF96Fs5ILocVhlTzXSILudTVLYLX/YJf239OjpSOXJVKHyuEY6KWsAc/JvQh1MiEiU
8z5boHGxZ/Nh33Nty7juFSRPNQfpY9tU777kivBqlVQ6+rXzH0bkihN6lYCiFv7Cj7eSVeqK0Yhr
xmbX9vypXrRLYLHPf3ONeGGNuUYuBfp5eFkcb/gTXcaWqFkAWtNcqi+nEKd74KuOomTI6b81Mvcq
k7j2q+X3tMjaObfi3eLCvjIWRgUk2eehYxJsuaFQCnpBaSQMb1M+cxBMfCHei+Hv6NDie4CRyjzn
5bssvdyraX5T6lw8nXM5Dc7DsHFE3RdVhYG/iKc87UmJpQhJG/sywt5coJAp+GY7KP63X6J2jIMF
5xbkw8BPrwkXMPGDQ5hJIKzp5wfm6tPOA2xZ4XvLnk00DEuuhj18ysXLsEdIk93li7sSSR5RJXdz
imXZmUu0BdpYkVTSG5khpUbCKMUdxnZ0JR+fzj0rw3pZ8njidIukZbeEaX893bLE6nszreUhDk4Y
SobAdHCaZ04Zb3OKX0BV6JQNw6ecHVgWppCXAOd50eRpUdGd877ewTyVzGM/xbX2nZlcoXKjwvx9
PnMUi/lMDSlOXWZPPQLr29TeawV3Fe9CcuaqHZLgSFJiU9LZOE2PJjNvO7maPrUsCG70krzeC0W2
kaurQzz6hARo/qre5cLWqhMPpMqknqGpmZBgu+dYrf9pBLRMWgoopaCPGe0LJCDG1Gj0xVsHeLpd
dyVkk+9PTVHktDNdAF4dbihNPxeEnZM4IrMCCM9hjw3kEVqeqhNyta2BWSrLMaRqltmeEI2NGcfl
NCJ6B4WoxPDunnkMIN1hIwHEuMY9o3M7GCDhC/ijYWHs5ZIpf6W8U9p7dIkGQ5ycBnY/WbqY7IWc
j2dEGfodlfIZRN6B8vlWHNSFC29mGVuROLYaivbDXWyCVPiuNN3LdwWfjmIzaTD6708c5pXSsW02
2UnQjRgrpMl0bi3JkoA7d79ZPI9ttVQc19NSoHumxy+D+yK1VJidoW04+haUD8whObBD2vkBz4Pn
r0MP8+GBVQ0gqHRHoga8WMv8uSa4Ejxd/ySktS5ziWG1QkH4YvddnVLurxlsxy7mDapeoYfNOI+I
RkSrQKaEQDg02zVYfBcFWO4QTmUCamlb0lsuex9wQid4Lq5t3SqSjOsudKkpXIZUKfHDIOQ8bov2
PdRMBvlN+0SstcwGlyd9LtngGjIxLNxbHMYIjrM+12iep8dES47MImQ8ODfB63v++p4jtW1jjkg8
Yzae+CfrpEgSz9DqeSbindIT7WUt3A3n0AP3uWPYpmi0Dq0n/nXuhrjiHlbF7B1ruisuXkmhH80O
e6r+LWHId5Sim/UR10+U/FPke0RxxUbDGf5k07hEKpDC4WXBEUj5gD87MRUO3rR1uYipA8UdymSI
pG9vpRaF51GYg8K5N5k4KKbJk6WcN3t6aer7N6vt1svCMTx9lavSNiyzAJnXMyrKiEAsZd8ZOrYH
dUS7uZ58IVyxUNc8abAFM4/V0e5C4QqEurwmdiFj5iNeqh48cjov90IbM+bB8gqlFOI3zssxNtx3
wH3AXR6bsVFjReBy0hFwcIdKtDHWhl8dL908AbYqaNy4rwB8lQDAgRwUlcPXLDP0HgpgXaALowVS
zhAhpcoCgt+k8nQLfP9sC76MXefRVR6SzJzd3a8hilU6IlXAsZ+S389ulbT8CiRJ0tm9qEHC+LRT
OhWQ49IIKHDo54QlA8IWaxRpgh9WAqAD150BRWlhU0eh+X1wu2jjebE4oU/tbhdLAsDM+LlG7qNB
vpOvzsXvfOPNSubzm2WU1xiZqOjpZDQw9oFXh+VGe281wfkJ5Q3PPzpxgyZofRR5z6Qkb9QV/7Wy
wesXBqhoGWgtq8yN1emB6YfGao2nIacxXyJ3ok7U70dcVorbXQIgGW3rv70CBakhoFU6JwWQudww
7a6MtNx87Qm0WhrkBNQbYE4PTlY1hxg74lNU1iDq2TJdxZy3mv1jryyw15lliEQMXEZTT8PyPiC2
HAgBi6/pz4LeKv+tf6x9tfJMswYvBdkVdxYNaiAYwiTJPOCA7K8ksLWJ8QOyhtbQehCz2gclX0Jz
LBK1UmldWT1qtspFiF7eMsmVOBmYcfEfN+CoPm2DJWlO+jOaCXFTYxFFAKyAO5kCEry11m3+3+T3
oLkDMVk0meGjnVeL+3kGrIJflqHBOsvE6SmQGTDdOVwVekCQohVFbUpeUvNu6xZlPUZvR2u+lvzc
bFm5zRGSyIE2aAo4dIGW6jm50koma0wTuG8fPTuq1EOVEUvVa7dcc40ml9PE7DTlUSI7NKcGGnQo
XtT6rM1vYpwVJw2Glof4187NoE6NJoYQtmv203JsOtG1zODvFn8EMltkNDpizzbeYDyFoK50jFzR
aiceVlEwGdFpxtjGbK90BO0H4apF3Fc3B9eiLJtn5QxncOzhKDUpZvfMJKWIWGvuiZvcIfq+kpSG
zHKDDi5q5u7AtBxoLkUOJ+ekQhmlIdvynsSebbOxGvXagLaMQw47IJYB5HRqUFdzg0CX+ssSmUNX
kKgvZ4LmQ15O4Z1pBDq/GpFG296TqEWOtXQPkcZvLMB31XuLdQi8S6JvbPWCxzPTsqwmKz2q1jnj
yD9uJDFK7V7K2yLNt7JD9SKG673sPAGhfpahUc9RywDWdH4MITwi+y1NoHamIl8UCQfum0YiQ2c8
G3D+rxrhVtBqdS38AGa1XQ5qF/KNSJquiqHJ7fBDAhkIareZ4u3IRdshFImzuFfCzFc5qzL7JB+M
/iXaHyv37e3dPcQx4XiZt3eFi3YvTV5R3evTK4vRhlhZ2n6BthibMWoLYsGdSuMWyC57V0vZ6iSc
uFNKa+evzHeon1AumHes+xnA/lIPVR0oqQlWvGV7SuVT5Fo3W8U6Z8oUTOVpKfkcN13T9ONAPxhi
MEZigsm9PFy/vx1cyRjkducU5clQMV4CO4E/tz8QEOmBqutZ3efvb2fXa5NfQSZcrEsPErUEB8ik
zzLam+HaxAkYKHeYNsmR5TGnSuW/z5aqj9NoGd0y26oIxpgVOvmMnggFLC8YImEh7dnMSyU4Qh1y
gfKQFaBS+dQ8qfqtaIbk6nfcTiTug8tBAqu2APMz+SEmo9+op4RefjCvWLBGlLYDo+8kiPd+39YM
J0Enhv/GQ5qKwEjf3nn77meFEh0kXmiibTqFvk/o2k372ny1bXuqhUfZczJlRfA3niRF1qWkfv2P
RmykOs12Rfy8sCcZz4heTnE4oyBxKmM9E05nj8D5ktOQQLwoPfnGyj1aDBB2FpO+Z3pXDgvR8k9t
vHu4VGb9oLS7q8BanyZgknF+nzGMu6hraP6OS/RIo1cgJ4UMOnHlm/nfQ3AeftF77jiCzKkvrEIH
UYJqM0dBg8uBbNmE2pOrSDWYAJtc7gtVqOIk7R31e13ADRQKEYBiCCuN2xfFv/HOVKW5MG/JBfrn
Bf6cInXHGyVOCVSXGUOwCFlt8f9yqq25xFSm5CIE+GZEbfnQc9oVA+cv6C+M7Fa+Hx5bxagTtsMi
Q96PYv3KvPmjewv4m7VLiuUly6PtlzUcjEpAG+LuQ49HLmy3yeY9m7P94QNc8sTY3rK0ftGKi/IY
6tNLMATXtSf3gcz+E0lsW3UMtwYP71ywZq06ei+II0Yo53TvcMtPYbvrE1C9whJmBJPIFUiO9RQo
MuwzKxtqgplKplhETMNGUBFezwC4rebNc4seaY+rgY0wq7ZI3OpDRh8oSMq60q9bqj3owrpdsMnE
F3kii1KZfGlWtXu/r/bTRkiS8pZFP8LJ0/sT4xjG2Brnn7WdNK03I0cD5rxsJdFvBVxyBsNSlHYR
0mP3QMcwhXB/21pOaFld3DMi9XXzqgJ/W/GDb18DMaBaQ6XJHafU5D5TdkIwFDh2qPBymmecX6pF
/+NdI1Ch7u96kfmBZfyOo4GqMgoZcxMGQbewk25yl4eYxBnpWTeT+72+q+fvzxBffJ5i0xe2LNKo
RKUW3gYEtI4IBEcLs8/P3KbGPL6WfcnByXnypM9GSOVh20hy5a9t5EctwTW4+9nU1dyrrV9HvOHW
lHW9eIHvOKkOyf/YTQCMDkYvWGl77rJ9OriJ381gWg6AYVssjd2WFapWTvHDOeesi264E+p6NqKv
vZY0PFJSt9OAKs2g/8nMl68rnpT4jFbffzzEpGxZfb2ENQ+tHuuOnNxBOxRh/rP4W1OWTUJdVUFo
NCcgzFjPbja2uLhXt6Oi60j8Pk2l3V3GUxepJShc5qNDcBTCXZWnMXGPlECpZGK94YDgnBhqxPPz
bYXhYcsqxdlnKB3UO3xgYSw+43AQ5LcJuyt17YpWvrbQ2rSsFg3YAIz/TiLZB/P0PW1WZsJNdORJ
iV9jdSv32OUm6ucvKhXND81b/M1gozSXG+xKB2ffWAkktsFRp/MhElFF6HRyQpJ0QV20SjvxgL2N
IEvu/WyD292PuDFVv2S2USS9gsnLM13g/++3kUPmLwEIg+CY84rJLmx94J3bUgULd5/TeaspmN9j
HChPwhQLBcNZih9XbzrAD/iFZT6/Z78sU9EbvUPyTNezhJxwfBbHoO5llGym5Gr5zSI5HREPjLTu
ee5O0yz8Snl+hhX5ZzssOhDr+iHHl+Lpjrk8BM+c8MC7MJdkbWXT1U1GPuvAvzaVBj/PM/sD1A6Z
fSqwjluDMGpHDIBc164ekylpBZW2/xgJtbp+JsvllKlbGRFrZ9X41ieCsRK2EMfj/+O8UOX0hSUI
NZPY0qBO2T0DpCl+09QnKeOzr/wQyKhxic+N6pqL1l8GW6d8TvpjboRzeNZpwc8J8nVR9EhhhGux
gmDRNFIRQt6FjWdwJyM8R0XDKoQhCMQ9qgW7i06vOvfTuc9gtRkxxigqlA6i3WlwB8uSi4FX9+w7
sZ/HWb3y28PFBqdcTR/FdolagtqCYZLjcmc152z3efllGST1BnQnzAfvXLACgD7n+CNNZBrQSLJJ
WUAJHAs1gDGWlc6biqM4vQqiPeHcHSoy6TyURdlYyCMMRgSmozXCIzqFLlRsTii4u/2gbkpjXLCe
NY4WwHzujTOuLRYcYyiDhYbNLmx2KPAZPExHQPBIGNOYgV2/s+7Ur4XmOyQnEbIoTMefcPN+3ikQ
LCfp11z5F6torvXc92I6ov8BE5JiJdQqHA2oGfLAY7gaUc9zSfKyGBT8aRrJ2LZBLppjZtxliPNu
9Q5nTMtG41qv2xxWdsRhKZ8lsYaBc1kwRf4WA5s0Ej0AJ0UYQGY2cZuWh4t6vVtZo4DZRMqVf5Y7
eauagNeBTuTea6wHPOV0zJGmToatUDsozFKbs0sdJEpR63rixH1S38nuepfO3Ba2jx3Qo+MfJYft
ODWqFJufR++iUNnbLiwZJZIqWJ9VhPdk1yQlbiV2pHjy8+GYPQ12VPpNHumj2MdbpUK8PCMaGsil
lWCDKB8eZFhA9h1h6w/jBNnHSIt7lQuCIUysa+VgwmUPCqnax6rZe3ccizWoR2akkgRoJez//lch
AT2meg1/0agbE7mctR2tAEC6AiFLgX9OpjifGV2GxWCxI8yUd0OlwweGe3fRUEmjkJKzPPI/A4yi
XRiYhaEriHQin+D1N1/FYE53WrtM+jy3MM2FgaNGtrshHRrEQqDozkzAEd88YvcfcJyHDqPHoNpe
CG7hRDNYnz/45mFz5S0cUCcaC8THTg4c/dJzOABin0/LAWcktCZSSJJ1boPO6ToL25+F7gSdlICR
CmJvrj2XO8vDwT/I9Zr1ih0z5zyhP0g/433M+IbwdQNQWrTvN8tnNUPjnLhp/5GbY/wikfkxTq4M
nM6771bToCIUMaEM8M5YToVjv0sS3f84guZw0al4yyLCjBoOBkuan4omsVsdxhaFYO0F24v/+mOa
TKL31sKwSyDn9AF1sI3OdYgLBSsx830QXrXOdzHNhJpPAASRvRUSvGq+rn+Hcx2Ltl6ZJAVjj9Gn
T4Ei0VL4AFK02izR4AapO6mv7Jj2uc/4C0gMH9suzGEDvyBPmxWGtRGROyhJSUO0lqveRwgfcBAF
53KHfboTA+J2oYSg+aoAAu1NnYRPAldW4hOrxYclZidyVqUWnxL9bUVS79nPfz+CA0powYTuHt8I
AGBd+VaXrgxB1fOCCcERmcbztUlKyw0WOw76iZyc3Bfr2wn5GY/5mNchzm3Y2cWiQ6JyDYG2cq08
/gE/TOb3KYoHoIrXuaTOOoa52+Lk/ENdRlp1sU8enZ7otyLXK30cv/B9SY7TcCO3woNe6cNVe/vT
uqXqo6hbIILN1AzuBdNznqoi3Y9P35vW65o81d0EKsE18lUN51xH/h2PXDjTh9g1IakiA0Zy+tsP
mAdsxp9W6K98uBR68jP20UvgrlcMJaI2Ye9r+SO07wVj4ggr5pPdKQIZpKqSy5ae5L1AdyuOcy0N
ANWsyUgsyTsJ8Ld6onpwH3LXj+pgYGSX3VP6CjUtq0lCycIjblupZS2xckFj2bgVy2tcH+kz2qLP
zKC2ROkag0NefpH8vpUKyIlODy8AuJI3ccabuS/GzwAwpXcN4BQ5rP3Hw4QCV1BqSulKNgPY0FTE
QM+AlHppnkrlYi/ml+DNeSzu7SWD8hwlyS4++79sqC6EmQqODUUuXFxVNt8sD6FIPLBak2XCp+xq
FtInJOnz8uTZHxKCNngPUcphYfOmS2QG8Yp+mIjawo/TTb7B0Z+gQv779vR2/aeJ7Is9Fwep2+ET
/x7PKeOOM/JFngng/kqXSa/Whziqd04vBXM7HZLUB7BW6KoZMwZLKjrlHJQo1lqeO2Bb4yPP3hH6
rf9fz9/fvrYWs3mRIjjoovX6GJF3UB/VGqdi+p8OfNdOam0JmZLiPvcDfM3x4dVVIl14aGiASpO5
MoT8NBxsstUW1XyjLszyn1ijKGU7Ys8aGyRD8QCsP+Zo/lI9YhNAMV4Zv8KK/cw9N9b68/B9hBlG
ZCaNPWJyCPeWTX3ZcbTJD1HhSleq2yLuBEiWg0qAWIOf9DUjVfmLNK69Pg6ZxglahO06XIehhKwQ
QL3s3ZCuFJpFmDyZ7mxk1M2MgEGcMrITl5f2HZYyHv26i14lEZd9Pb4zOSCcOausp+kQbxOduUm5
wqku4QdnVd1J0tpMkIaoL/R1J1jYeS7F8O7LePsF7ATVZIKH/i8Q9cQNfcdBlRRj9uQRDO1A51RZ
KxyoPIUd4lolavl01CRwlLoVSWNO0+rEMfX18xLHiIdnT4Yola7ZnQc8SOUOxAPxj0wPOTR/t8B7
KD5FxOd062tOQCD4EE5CiFy9vrVblP93o7zlTBbG365RKVvnKVaUJ7/XO6t64CNgVZ23EtHrxHKg
aqWM7J2jZTM67TcD4cRTN+Mn/jiKgsej0o+G8p4KkEhr6kQo0RHPmqy9zXZs8O1OWOmfByBKllXX
73MZys+4RkbeLessuOpu6EcDUpfEQ+AWXRcqEVBm3DewhNc9YvnPGwHAo2tfZw03pGJPj9mgSgsD
GQarMjquzo4n1GCeM02uOk+bGPJdAk29vALITgZr0a2nLuld/V9e1R9eULenUcxnyqwDR0hOu0z2
Pfon0yaE8k5YFh5SANr3Km7x3w2CbQ1cfp/Fig1+NyUI9+Wf8gro6LlzHnpne0SrXNWvjHAIKsfp
6qqIGr9am1Fc2PkdvBz0Xx9qNUL8ANWQPXOHJvMTzrWMkeQ91WfQVyE8f/oxHILRz4NkFzQO+wRK
JjejELuNjtpqorFdhMFWQ2LkEVRZDkQhDszng0KG4jL+jMgsBphVyAx2c390yrBj/ec20UhdmSvV
7q7nfAaDiXtWOWzIbTPT7BihZLo/AzPFrMgYZ/0hnPQDuU+w4aiSinmSj1RrR0SUm5V22iwgrQ0c
tMYxQT2rhhGvfbL1RVKExsUyWUcoJ7qO6x4P+AmNteEasGxSrPphw/9U+dSBa5qe2ydB08+UMqrp
VvKpixKO3n1NAngiNsOYKVckYCesOozplcpcMXIyYw2GYbt7YndoJFjBCaG4B0kq0LBFxUebiCrd
o9ie58DULvLLgDhCRUMDfUgI6RJf0Ux3eJRHszo8hvIAAROy80TVGfR2lR7dlbdK7Gz0kKh5QlQq
DlHQfo+XB2nnLZMTBuOGVaC9IjXXTHpZZDuaiRG59Hptf9HP7ME6DcLVV4h3sba4eEgjuzVU9pj5
X7osNKrYpiTDnkM8ikm8DjTDUE70oCCa23STE9iQWQngbT/rmtaHCPxAoPqZanvRpIcAhXfm5kMX
SRCuGdH5TC3wmw3pKQNYL8AHfZI3/zGa8X/39+iDxhd3Lm0x0O/lsN/EW4Yxo4KNbIOPsJZiFGT1
gKrg0sji0WgoHXHl4EbFRmkbLFfd6nOoYG8WeKlHKaq1lsKuIj44uHdLynODCABecmJVuu3gPrDY
86mubqorv0mSpy1n8s8+T6HC91UqFcd9t0Dk6LKEVcWMyx66Gdz3o7vtVw+Wz3l2tnfVqIM0pJwA
AJbz/YlfitIdtEE1JXSIVYeXNPaifE98kq5XoH+UuRBe5ZOoB0DFypXLrB5wkUMlrOre2LH+s34R
GBNjk0M5ZE3Azucae811/joRB2LQWhP8ByJUb98UwaRJA+9v3fZoyT87BQc8yylKyQH84SybR2Fv
HkI+aHf6wZOswADgAGb2pJX7u3WzdYFQQvNh2lPhXss5JTUTg+mDaHY/xMuR9hlU9TmGTkb1pwkE
B4t4HZN8iW5wGvQ/N1Dbebe4CLLm2vxjC/DBrzFO5cDjTuyWApav/oItdUc4BXRuSMBsS2ZARE9r
Vto8yHkS1PIESm9Dcaw09q7ro6Dvx2Bu28Hx6k/+fH9ifuQzrtvS+3ss2zUjG6Q5aLjKLfPByC5H
ZOCggBt4cWOwWF/SDef3/MXavGBRmjT6vVMkcsWr6ykieHcx8TDNBOw4JawRFFGFRvJeqgjFey9m
kieYWwCHH792YgGjioC9F6OZp5Uj0ILr/abwgD2A94H0+XZsIiroNTFLIngQF7OKSQq3Up6/KW7k
rYj76NFHeM10GTH6cDyWOUXKSUynOxFW3oV2i+rx76Pv/HfDUcF3OSVpoyF5WduAeKuHZZ5jWEeH
ekXm7T30XuHgMctaaqlk5ezPfsTqCuTu/qwYLxFefhNxHHrcMK8vrRKW5eRpkPip49OVvE9X9H+p
lYwg+QlzYqZWMhRyfZz6bkYIIHCvni+R5Rhj8jvgXf+v9obr4dWZSTFVb0YE368hbzKhdQCvvToq
VlIe5UpTh+YYfViAWDx2pnChvWLM/+cJdH+qKRDzXFYhEWN7qErg/kHkuKRc5uYeotNaPE5S/Cce
GVKaIZ97rP+f5Veizc1khacGUUcbj3TVCBxmfrDfUudxbZSJcyXFsfMoCGYTOWRjZbMErrlUQVNM
HwwDzje77l8ygTzEi+emd/vYYKx8eFIcbwmeu4sVoWqRr/4xJRQohIRXDZ3c+ZxE2c2Nhz+zoA8E
hyl6aaMJtTiVRIA4R+QI4Ndf6P6bJ8/xvR5VJTYYYhrznfWp24Cz/rCvCIYOB37LNlz8Z9DbfyvM
+fTu2b+2KfieZwqMnrYpWn2+D3Wf/23rE9LArSb3SDQnWJ2zI5rDCGB0vkPu1HcVTF6LyKbky0rs
oprc2Es4tmxpe3ogoiD9wSwV10yJmR8M0nC0f1Y7ATvYOK0w2je6X5/KjakW42CmLOt80zleUylR
BrJvc3dXPLyfh7E+s+PsmmYt4gxllnckv4eo6Na7AlRf11kva4z3Opp5SWypEFthELb0C57rzcQE
hDiT7vgyBS1JYJqWn0FPAZeWKrcgLKxPN64dwtyHNuh/tf65c4zrGvE7O/weMdJTnNuugCKbYJzp
7hWyhoYrbb7kcn1lFtWN/I7DEKIUrL3b+gn25hu1udCO4PDxUAT7ReEoqvgxX1NiNB5laHUOA0U3
eip6QwIN0l66i7Ls5rvAKhyZq/wpxQMa4YKFmR8O/emVFSFsFjhxGc+yLjKAlXYCA2rSDtLoIEcp
uDg5HHMsztIPXPvVXAWeyiosSfdBvmeFFQCOw7WYXDUGPid+HrP2Lc2AdW28VpYQjSCsSSIfBren
dx8B6TS/7EiYoHTUdTjQm3lq+1fNW2ksmvpKunHaPnyhTZcvr9qsC+/xgH7ednAsIAEQxrF4F/f8
idPki2tTCOOzLhOC49KxSqrutuGevdB0gQ2p8x0beeOlTntEncCmv+lwmxn3l2+tJNwhYjohop/y
GbCN+2ouLAw2FjOwEMMGudQqS2NXDsOsvwrVHWUTCjjtc4Dq3b66bOvB+40wsS2D/eZjwKs69QCr
zCacu/eRsiaMc6gj0dflLiEcI13+uvMMxF5ES69SwbIgOjOmPCxpkjAYnFG8rYSEWu77ejigg5Gr
A1KPv59jFKgUofG7Hw/Rvouuu2DgZBQbZbp1dZheLkD9DFyuWROKyK7y5Af63BDqfThsshW9agfN
OSwfjJ6Mry9l+dTMTBSBi40bGNLx52a7dL6BkzB/kq/PGHL/+fMqshKsCJE2LfvuIDzZ+X5hVwMj
67A6idSciDKGM3kEO6HqpxNV3+0gZwb4dEXBj5eQUMFD38PkUq9f1/Vu4dSukA7zsKkmmJ5T4b/J
btPCgIqgHWMKKesLrTk8itVRDpAywTqKMq/GDBL0esS77cRT+laAgqrzkwCghDACjLQTz5rCJKpD
WVCp0kXyuMfNVMcKv4ToDWL6soP5f22JLWaW4v3JB3ZPQwQf/iydpo8W88e62iZCfT4+1BSDZIN5
Q4KuasIElDD5wDYbd3js2ld7JlwGwgoACKYQm0StX85gA3Ux7loQt1PlHo02bnJ3gkIDhi7p1vtS
fD0JBbBZ5+VfTd6IiIisKI32uhHnF9vbhDazA4gDScnBb7ebhpIBgvA+iLogcHPCCOf8wfdp4tAZ
UZ13H11Pvd1hu4BtFmPqLS8Gaep13FQg/eO6bJsU5EUDb3GhWNKO6U6+fX8S2aG1lkB5GmmbR6l/
rBgFNmRJHU0E3dNA/APVMs8u/m6/74CfBmWSxtMFbpDBGhHOHsQWTBjVyx439K2GN9b5ENOZtKPA
MGddHlFeNwQll/3o1t2jTIqootma/hlmN9oEjVCIq27Datn0oHxITM95DkRsqSK9cfYyK90BfEuS
X0DV0byi7rva9WM7KjCNzSfc6skXUrUixmIkAu9PNSXoWFwbZrob3Ztoikis3cp0wm99CFqQpoBB
apNNF978Dh+CUXuhjsaMOCOJPoAeWNXJoccxeYQOq49Z8IYbJlj1vBz0ryLWiLbdajig05q7LZ2o
12kXCJPj9xxuwK8mRXf61NdVlDpBAcIFZC5NQxFRANFzF07BXCF+9ev17rPeFNmu36bkopQCIE/s
LhkbPE5vXrXp5liUvO5F0tO+fa2iBBYKQipoABAHEL63FOTWJXQBTbIpB5+H71YtZp14pgBSVdXm
tjLDQIhY2c/Z/eJ9k8j+gx4Br70jP0UlBA1++P2uLw6PRtilJFdh7DT7F4p5f2pRKcl8PDoLzsrk
yo8soyXOszjAu4HGL/8XmrXmrXSf0txjcOtSoZWgSCyPUpGURDjr34d8/2mTCbVVrskh121xjVyi
HuVr3gIEt7EBJgnTYe+oqgFOMjiD47zzWuL7tR7g0miUKOw1JUYc1pvEr0jptUdddwJAtOdpEM5Y
MIaU4eJoteqVr7M5paeLABQ2D3nlomYFFHuH+Q3ER4RLo8m/Mp40+EO2yj7N7E4m7SvVbU4PwY5q
8iB13KLUsA0clyCbT7L8zjhjlwUktuP6plQKAvPjcOh9itO4u7dm6GW+yUMiJ+WyKs4C8t9Luml2
28IMwW96u2ksHDldWVjBg8+UXHU5p0icB/jpFIAulhe5LUjd6aBPAjN7pWkYbuMlN5Ixfeo3kKiW
jlwsTRFx/9iOWfZLYRNxdmM/XKwttZZ2nVC+Xu46wMNkns0x9M2Q/dy9YI9iBRAT0d+zfXKuKNT1
uGnREfhHRpzgn90Y8M/OAaLpR2NhXQZkFoP/Dm9ixjJaiYGDon75zaElC/6+fWyf/18LzmmYctWq
n4ybR+ti28OUXhB2f+vBZ7VuQ1a533+qOxSrWdxmSvzPvxuznJojaIr7iGBMlDQXhxKaJMU08A3r
WhFujog7J+9qgRjUQeDJYZC/WQxJaSLwXEPldkBDm6jt+EeW344d6KbeZVrcZtY56sVcFQpA3TgZ
J4+a0LKLkmak58tfQ4BOlPlqPU4cG6jHudxCrW1UPnNPb13+OKBzaMayRpbHS7A23YaZLsEWGHKF
sdq4OLKIXJ9lsvnZs1JMG8Wsq6MPfklhh9CupgZ8rD7ZvAfFp2KOU8eV+xJ2ymcxRCPceTwoa2so
RDf/2rAq3Prdc3RVHrY9oBDyUqANLXG2ilLXSaTy0fx0FJluf5vDEKaPaLXFsfUaWimiHRngns5g
M/XkSsex+22OFP+ykDaiAcW0F+DyrOFEcLlyCD18mTsnMakzokAjLy8OB4tj8fIuXD9EHJhUtu26
fb/FIkowhMfb+tkzau8GtkCVH5gS7zbR9PLyVoadbkhj1zroRkWD8TnxKjXXc0STUEAnxlKxmZdj
88hADeOQrExFM3FSJCNHe2OxfPJWcUyGoga+b8JtU7G+MPAivRMc7wEKVDycuvr1fM60IsMNF2Pw
HzunOOfMDd5w17hDNZDThbM+UdoM8eQXFKdN8n/URhh38Nj+gYvAvf+dr1M/rG01MZGtW8SWk8Nf
algHYf8daFVqWwRWz5gAwkPk5vfM3SofqQs4u6HTKt1sHcMO7A+3cTFiVIaOvIB/dJ65iDq3eokW
G4KVb1p/R5abzX5m0KLwNpy+basG4OMjGPw3U8K1JKsXYty+De9+Bm1x9VDohckusLvN1NsiGwva
9OebT04fbMPKb2cw218WL6qzxEhSJxjg8PuBmwo6QYGWEXL6mYoCDH4ovWzWesDzS2/IXNYM3ifl
d//oseE9JqK682nVPc6tdcatL38+52oT0vkiUhe4em5vmp1ch3YlLNDRvl6eFjOL6MB3eGuexjOg
JDC75eXX4DArd3znm+BLlAQ4aHK+LROutIdR/mGAKuEw2RjTSUOoHddoa9HS2eHHC6mILpFWFkEi
uVp2SYPeGzl5BZ+6MnAWsOg6vx1Ox3yZGWECpWsXSvMljZZyWwL7wA4biwPCTvi0Uaq7ZYfn7fNo
W9Fdr5HznizhEdQ4a+cQ/YI0wre4WMGiqI0f3vYvKaXM2nCyrS4hrM0knAVB9NbeTtIKgHkJxoWo
++cAFWfRjLlFiG3/j6o8r6UZ1+MZq0rKMFEqBhOSusCqgmyilDM93z5+a1jQNWtj3pF736bbXX4A
QnyLox63XktKbb3qmb0+a328nUy8hzsC5hl3jp0C4WYFAWpazkGKP2cjpGwQ7sANoIFmIvW9qx6a
vECalU/d80khiYRZtKAFOL+aqEDiuhdegc5I4vX7q2t4uurG0Wfywg+YCQYlJB0gY7iKMrvZv2vm
bVZbzgz51V7Jw32ZnXcknZ5csiI6nzFm0DwQHXbORllk8r/1a5sN0op0dgQuRsuxTdhSUT+bb5jA
BlNtXoQuhonf33nClPQ/17lavNzZNrn4ieQGU7GyZbp5WEACSy4/W571TO9PWdy3QdId1RjBUco8
qCuleDBfyJB7rgFHHvR9ReR5fq87u03HzSwXqmdfxcE/JJQXsRwXxeKjikF8bI2pW8Eg+eB/ESwU
lvWpravCjH/rkjpuHZNh7e7pLbvskn1oX0mRW3go0xtAhIgKhix7NgvQJehqhxkUw+ujfxtiE3CT
f6hJWU/uadUIkT2FsElpINsTW1xVoVv4XqD2WVigzPMugFAESDS5LGumQlqkwJNAUPNyWZU5LOI/
9waVaGj3Ye6StQZ5YERzE/hYSNR19/yGEgYIW+adB5NUfLKZM6gqQfb21ORbfBPIVZEkqyYv5Emz
E1qMu2d9sPa1rHwQIRHfqXL6Pu0PtD3hdE/6yIYdCSWoF48EMTZ666dlzIuOs1O7EEdivzO9vF6R
/lLCpiyApZ6K/YyD9m9oLL7uf6vymZ+KUAjp6FoFnV5bvSIrlShcXwetBJWtVpHM4nOoeKEv780J
5PbruLtjW1itrXW/TVzcpHUSFKCXRn1YVIyEkmgEsfkRuC/Sn3EdSGzdQ4MnojSg9io/4hmZCMdE
4mLipZL/8OnqNiJPPga2SJ1KfkE8Hng+8IEo8btchjnj4dMOaSSFkv0wcC4fvh+fPxElFNRUD5Fx
3oWIGsuELUd3xqHYZdXPIRq6w5EumpHgdkd+l7gtzacxZQV9zJ5ghilhnYy5cwFtsyulCjTzV2g2
nKinptEfiA89+whL0LeyqLxZEhv7LAZe+8rhqh5UIG+QR1XRpkbE2dVBTKVRni5j5e6irNM8TJH3
ibovC6NI9DFlUjOXaYG5Ju1h45Bt5dHHF5sVJ0KZClEbCH1DEZybh8nB9Gqfo1bQMuGDfYvEDTxj
6BDVco3zTStRygaTiGhDwyBL1HCLV6ZvaTrRvkp1KpqmZuqb5k9Ly+yQ00qGBypwiVMBsfCfteWI
WpKvLtOjccGz6vgg+AY7P57ogGmN/xfY4pye1IZ7dA40YrMlbI33lllbKD+WJ66IPqkjsn6c3f4t
X4T5hODnOfHRoWrEEeavow7epaf+e0gzY3PL/rUJxDbIPW/oSbTeXbirk39VvwB1OEHlS8HXTYZy
sUQFX5XX3ItRDTbhKez2AEUeCQ7WnPJ2SpOBY6drGdbi97g369u5qa+ACv2EQOSF7v6wu1IW8LSE
2/Y7N/0cbtTmU4HCYUGV1PTtuKMvTyH9whVxYLyvKiEY1q/19PAeRYlUG9dhEK2D3RP6eI+egMcc
kRx3feOWA407la+4vvW4OE06Kr7Y5ZIgQOcc8heRnhVzrbup+DwfT/6cRWUHsz4n2Q1iwKPtYt5W
eqFYWRPlx8oG/7Jszyn8mrcuglPqgfof2kuNUIc/MFa3tqMu8dKHki3Up7az4E3EHzkPn2qT3uXV
28ycIhZjkwMtqKF9PGS6d3L09+R3gi4VPNx4jOJScMksT/kLs7djDXHabiKoUzGIxQOq1q5zoarl
64+z61ySvS8ITPVMBuL9FiQz0DtxG3H9mJc1gZtwFc4wQA7kiufZNrTmNNh9H+grU4e7UmngsnK6
prPYBsXtyBGiNMRqMPDy1krcx4wbNdqEfbWwI93n4pIEyFHaE84QC9vp4U8U3tW08Lzg0Wxh5LxY
ffUmLoWBeSAL+TXHaFMQDs1urxxnxxp/981mKN1fUDh5bKyaPZy5SmKu0XHh1Yihjwqms1mni5Nv
aDJzz3NZwb4AyZ8wPaPNxdOpaAHSWctxoiEmzaQJnF9IUS82QesK9I/g4Af4ggxzeiGmg9SYuYwT
Fr3R2KUjQzPn1CUZ/9HjMU83j8VZYnQtw1MNte+0XdZtpnaY4UOpZnCjSL4tnVp7mRe2Km8owztX
JDiDziZb6xv6BzoR+zRlAcEOQu6/ysENWxV/R8iadlDXyIU3WM/C2GNDSrNVOAiFKCUS+nJW6wTc
ZHbOUo1PxYH1kpFeQvjRlOX9WXcABQmywgM8QCnAFauHAcZgrrfNmyEuxno9gG6OA7tghIYAvkWT
aHYBM0ON9vLtTAPD52j4N77Wjz6tcQxHsMvF5YqEIMDzK1PwuCXnRxbyFsJiBpnvNjbV7HPK0hjV
kyKa3Cvy7+el6HR4eJE7NPgaNkQab1eMxi3IdZIeg7RvlSNv0xaSRtbnzB6IcBa+6UKZm9NY+cGO
xno8ZKv4ePItitfKUmUQw8oqD/AnfxqGPAuqkke6oRhfb52eQaacDialeSYWv5/n0XogNMrXk6JV
Z8C3YQsOXe4yrWrGxrnPKLW1wJO3WOLrEctxZ7ZRdh8LADDhtbadSdFwCnaMGDwP+a1Z5SbG6348
RiMh5vfTCgvI6vF49Oq96dqKTwqV1RSaCmDIr9RiA/9r6FxLcXZOzmeBcHnpSRb7rDWNXtXfVILZ
SN7wruz0weP/P7t82qqEhNgJMGfL09pwDthxIeTjpo2+Z061X3jDmyTCCg7L9l6fj2Cg4nemWGWb
HrftnOiGyJz6CLDC6ND5R7nq/KzK318OzUgbKWV+qjQS+Y9m5VvBeNhUGMloSMWMajxhzNNUEi8R
13XhOMhyBOIZTLrx0jxfWLI1RINVbfNEM3QxbsJlLY3cGPGNUngQMStJsBmHky+uTdN3pdN0p3AJ
yS6zn9FB3a1WcIDB9j+ET1ByaaOTFVUaJ6GwKQt9OLVcrVsG2aaZyumdrBSg3Seq5LgDUfOGp4oW
lLzVNVk/Kqxw3DSNpUtd+/W+q8JOB/hYVj7KPl3xWcj4v26A10XTGDbtFFv/PqmAt3mPNzGXzH5E
v7t/5JHdG6f2ohS+7RkjJPGTO6Wsg+JfSKK1RI6gassyCUfjv6gGHd5RFL568HWEaGzIcYPo+b58
A9PyTBcpy7hYSOch7BKCpoamhejLxfLT2M4jx+A3hhPEqpa+67SdMaLt3w5WGaVIjaM/2eOsSYpe
aMcF8OLFbjZWmu1r9iUhBK1uihfX00jNMXACeIInFe2gAHZfr6ZoUb4asS2UJWq5D0oGRfWXDS/2
EIOD0jkaO3560/MHzO+0M9e7sxlgNmrfTM1rTK/E3v7+bS3o/DtQcMzQy7sfelHkylRjzmmMbm1x
8ecl5D+wa1NHHrgs2YoPOZ0s25LBLYPYKT+40U5UXJsE2i4u3zBUwEPzUOQ8oSy5V54OteU0aOnM
iiRfD7HW5dPHNXdPuVxATQ4X2++8PsLh9fhWc/D6QhQ5DWijwpsp6VfOSjlT3CElQar/AzaAk0p7
dLqFD92pDhaZQBe6GfCCauRFdF398DGWAgjN7mEgscun3BxxxjUsY+5HXRtGPerRJPBaHI52Xwi9
B8DIl3+tdmSDmQmPFookF+ppJRuBRzJ65iiNYh4QqVV38KIGtxaIcemRU/jyhAV0uWmgopKDgx3t
Vmkvbzjwk6DTjMUqBhk0XpvCFuJwftwq94JTz/Lj8z33vx/WlLkSFrdFfd7TFgmbeLPC7MJTsZIx
e9V4VXBmwxJW7GrxHzkv3KNx3LX7NVVeGdEwlVK5ZyycvRzP/av4wp7Vpkm7ZOf0f6zJLU5vvCVa
2GSOEWnKAgjm+3JZI1bGdPSoec5Kv3BL8C8UoY83fLnzqz4DIKn24qmQo/ic0rql03CeYD5MiZEj
OGQJRLRGHzv/xgPNB6ovMOP0XB5eRIxrBd4zQuvYDu0ObcWJ3WsPai2dPliJ1jS7DGFsZlsGJnCW
s+qXwduJvYxoRSjUBcZZ7813XLBeFkTchj+BVoNgKLr/mgc4Fg37u2D/IPvwQ2nQeL2eZsHFiYht
uGLtCHrmkTgKphHs4PzxWU0EsVy6eBBN3tssN8TK9VXrQatY3474R2F8U4aB6F43k77ZLRdaxwXz
bzn4i5XH4ngK5+7exLLTI0jBrD6oMWiFCXJGUg5UoGCm4tC41eLLrK8ja0QjdHqH0KQettkEedPK
vgFpunSEk10JpWGKbtuzSWfhQYSpRUHZODwiZcyVTEkTvfKUoiLUY6m1LNmSKk0wfxMmUCbzYXGG
Nnbryh5Q94O1dLS9Dm3pA94CfPEGmVyzLecafIq7fHutGyrIn+AuNoP2MMUThX7xubdIAGG8E1wJ
81BH2+ah3AV6AfDms7w0YG9TNCMuF3ko/S0WtqSmLOOSKc4QqJWJLS4Kh44z9EPiMEuXbTID2+SN
CKT+q/s5RIC4A/4AQxROP5JTIHfTgWQpYK5CwGUX2CYl7dIsV6Hn4caXqgj0oXH+1x7dwwhJtdLN
iFzudlur1wpTm0Q/H4Y6bssP9wXGFqSzHOku6EpQ1J2rDXxDF+oKWhvXSgayiFj8rK3Eokw2KZed
xRV6vW3eau0fLq9cfqfQj9uRKb8EVXzBS3EOgVvDCxJ4LFhzK35fUFFwix2NxWWT29sjVa6ieWxV
AQPGbaPOlvXyKqwQcpiXc0LJnTE48PlcOB2Bs89pY0YFBHZYEeJIS5fQifrIDzEo5mgO3m+0A+3B
4p2mCCMhopbj0MOClD6xeAyjsYCoWUCz8B4Fvg6GxKJHKeqF9ua3Ac9WQlCgbkizswGQAUgsZUco
Tj09wb+EmrgOnG9biyYxE207TnLjElZ3qZfF6mOhj6bPsy9tgQ00/5psVNi3lqYb36embvHCezFO
QnNn59ablgsdjNN8L5V8oAY2m7RV2Pu1Tw6vMfuHQbQz8G5msxw6BzbDeOaKVq8ktO9byO9bp+o+
kkiApwhsqLD9AgUCp4vV/ZnvDjdQnGcSNMRzOs0RZT2jvAJB42+pJ9q7xy1KbS0BJAnt+HUFXCZb
yQWCgkxsCCnRAlkBd01hMu/VGXBpGW498ZzVcCOpcBbZlYKEWL8d3VCWniWT7BZ4NDsQ7shkenvX
i+2VymM8yZXtXwFTwWvCP+e/HL9Zg3TB+DtawqNxhgqKuD78LmxkoI6AMfmSFER+h2EEFAcvBXAo
Myzvy6WNbUaZpgPfJ9V5LCRiZYm7JAukVOoRoFsp3lzhupcruIGSAJ0Y1PT6przNrsyi1cOaLXHC
liMDrXrM9pvlWtbCD67Qaoq0YbWBovCdXG1Y6FYrqeneHhksFTIVkrQIo6pwpqebABGW58MdI0fJ
R4b1v63dPAZPqMGM0VG6TbKQuiRaxQFP3Iy6vrOwhFhgtnkqyDAg/T3Hw2RMi0qoTyWxWv8lv0MA
K+9dyAtdDrRkRWVgRvKrA3UoLfyplIGvK43NM6WXlC0/fBH0l0FANNxO0k4PpbkbRQ0pOFu+KZxn
EUrTeiGk+T561OqCj0GGMBJJKZGq+j5b3d5PYrQoHGjDXR/rd2pNGZtTzUAB4uDNicO9fXI8SjxU
8HpoSfxEBLjC2cmUYScoBczX4GvA1vF6yehUi1D0920sEj64Nff8sWwoJAJE29z3OtbNc8iZGJpv
75CUMA76zx5y0KT1gjmAkPWq0/XQfpAnXuaFAlaMkPwJQS+pLxmLiRZiEKcu1dMtSnSar6GwvFn1
sSnWOROmJuNdptHpZe5Q0EoBLySV0L9jgKUofXw/qwA/A/o89/NeLOc2VhqU3aq0ScvpU3oFYHOY
nbioLNuddyNiVSh26xvGUz0CaB5Rlau8uF9DC1qUPQzy6XB3qXrGgafLh01R0MhLMv13l/H0rzVO
iX0C54pDBl3cxtU8ssy9qKHwziS6VFWmQJdEja+Bts68MsvqaSu/FB8NMQ69agV0gdT49Q2nuvnR
/wtk6a9aFendUTITKlWMZTR+qnSTEOHhTzME8A/JnGAjPWAx3yFO1y/uoE4D6dSQOYM0MNJ5CWFz
JgpUVERSGVv839wVkPzONIufh++RFuUOu7b8lSKD1HLn5TR4w/zI/G9q6FsqTSBdeo3gHNhGhSFV
sahnK2aSB7m7VPETXz+fI1FQ9u24xffbzlMI7Sj9B6s+0Qd7WneZpXkHm7W2J0fd/jvTNCEsosJN
wi1nBEzmmashqRc6+AU6gXCHPQO4t+kxG8kkFdprb8xls04A/UURCtfuJFGTDDL3ORJ5fk4vncm/
+y+PgJsu9ZB/BNidguUIV/UbZN4oma6mpc8iOL1w6gkX3RHsm38p7VOQngPt9puJ9TMNBdVoFSRv
GlZvNItIZfKF0JAwADCkWF31Co3vf60I2UN1WVbf7IYzl8Ib4Bh2vjkeX9ieSyqZVPaBHXQeLoTq
DaCcpIrUwwUYJFaRG+wIeibsyix/hKTTmVCMpN3xyylI2o08Fovc3gNRLQPzHJfVSmPLjgu64FXZ
S2vGrwvovjKWBNwTfU81VpgsQ6h1veWJKXCx22GW1pzjiGDPsln9zc4T1A7PI9FmBRmq+9DQTkAA
UDCMMs3MZHGJd7EL0RnJV7l1b/TmI0YxDlFsfnWvr5T0hjipVsJe/hdVqC1SRliYc0YCuwOm6IHj
FnymPK9n28MhmAe4VOccYbCA5LuUuBQybbc2MCRiccjuN1nBqucW87ClxQTSpXfP3vNTJU4cEsXr
71Lbkh3woxrB46SO4vLOc2Z50BZvQ0HJsCrSEEtreAlatdJF/D18wGlHE8IggrPxIfWC1LjEJKi/
JvyZVEXdr47m/CQuxydy5Q1AdxJgKnm+Y13G4099Y462W4++G7pjsMDaDW7Vnhbp6v7NgLCr0V85
IPNHf7EaW88ulX2wxQtruLKkQ7HusMDq3uBNnLiycdHBA1jtcui5m0PUL9ZkDrm4MnordQO4YQTI
jXHNE+vVIWFo3XQ24jmgbOoeqlBa7/1kIguIRp9MYeLRrFJBt2Trguy0kTEa2p2z7LpO0bXbtUug
RAxsb0f2eNrbJ1g4ZEb+D6JKeaelz88lIrU8yuZuFxF9+wwKmmugTqBb71kyQdaCR9qoJXfogsY6
ME9JKGqSkpA9LyzIxCHdnfp55+ZRFnJZZcvorDO7a8mFDvqEgtuKV+ywKHjDnZ7guOILOCf42e7I
rqmr0eWaSYvsC8BmaKaSoCF0hdJZ0PaG2ZEJODjcbff7cJLx7Fvt4ycF2yHDMkxOEfSMUst/ghSP
UVBNeFXbLnAsE6eiKqgyOO4uxMv389WYLK7eZ23wWS1wz4HdV2wIga0laYgPtyPKbwYdwzbB25np
w7+eMLK7yiqJRGl0cyk3fXjSRigXWFQ8cY74+v5aYMWpvdT+HzIeRsS1VnLM1NPIqzaiCGMyCeCs
vrLiWcdiiD55jbDms11EFqjhh53CP5/cfKZpngKYLyengz6SpfBESeQRCrneHum9q9LcLFr/qMV7
EpHTPF2J/dGEoG5UXNSqmIy+kH2B4t9kjhbFnueGapVURMyoao5sOHxg7dQ3WLvHx7IOmXLMXLUm
ovomPduh2A5GzobL+OJpKRVXPSrBN/DoPyj/fVDHAQuPGFWBdKfY5cbQK2sRFTT2eT2EtefOGHvf
bZuyMjCQgOjH7VOEidEgoEXjRb07s4ei2izI45LdG4T0m3B4HcOKIwirg7yMd+wV57bDf8ggflj3
St3gOfrzJgxns1wUKGXvEs9NOIjah2/ITf5RCPMBYibESj39pSzMMUWGNJTq7ZSZ4GWfhVQfAU/o
toHmf/zbfhUZPO3tfAj7866IHgccyKWLWJhXf0Cpbn+E6G5al3HIXXgH/uEOVhaIq6gIj122xeoV
w5PB+8OCWY4QVX2BnE8qiL+jTDpJNTqViNqzCyEemLAyc5I0J7rqWHPHjDV7T8WSc9UPZuM6zrV0
bxSH4662QJeVbSAMp2SK4BAaHIktGjEeY/sNlO3ej/+TEJUq6wrsRcZ52Q1D2CVUM4lAgxmBNBxA
A36QPjD+kzpf3sMbgNIpnlqMIckVnVwS39DWK7Hi+ok7cqb7oluQ7Vt3nczm7DYh9KdNCfezH5Ge
4vaeGgtFZJPBBdZyITRKoV60bj4PbsgNpcjUdslwHCNF3m8JviWVmOsDgi89bLxQiG0qKtiFnZnz
3WhvhMUlHbZQJ6mT/8xrfbmeBO64Xkeqk+Wd32PbFP6v7W03ej6XDQam+4H7VCuV+QHsjiAbh55G
sAujuSq6/TvxDjVluEPUXgZGG8OhASWCYIWkReYA3HO7kwYCAHv8dC6Izr2IfjSZ0VWpbh1nV5Sb
S0PC+L6NQKb+LVcUlROyf3vRBefJX5n9zDviksTMK020G12V1jdixymPkd8aZgAAsIdE7NdEWUN5
OYbRAu+5idj/L7J7xnvekQ+cTUvBW4zTTaezgLQhULqSr6GcrqjZhoCIpIyRKQ7CMmqajlodBceT
uXqMKJsH50Dc89iKTZAGjEc0brZPcBA0gk94s8JmnWWZT18WYA1SRwFGNBvo/heKWFSKIIkbGa0E
SWt3s+9WD0bCF3r1qv7MUWY+mEuMW8moy8xg5dyJSfkKYUmZfTKYPBUyJtI0rZ1MNY1qjQik8qzi
x4g4i2UYi5TCCnoZYj3bwi2RB1nypEpE6ta7lKLi0hZKZASRoMpCyNd5MBIBFHHumBMRHpEFb16B
4V1T58l0PHVjoutM/HqM3vL6t8v8GwBNEQBiQTnNcDGvzrc8AvVyfqOaSdKAAJ4eD3Zo4+lcWcWM
2Al5/I9L7QaX0Z+luL1VSPxzfXNYnt7GzeUKL8hviCDb9PBT71pqpNJ1Mfh8ApwFK/97mYk29JF2
WiNkf1FKl/4UCT5dWlcyPz6Shaim+i6MOTGpsmhG55laIvN2WxNNNa51Zdq+NOz9ya5VqMAvuYvF
Hu2FwMkkg95UdBgM+g2o1eG71t72NKWaYdcMg9oW1zGpeQSbvgv2GAW/yI2sZFe3WCxsue8XnAjG
metxH+GY3Z/rfs+tE8vjidL2EF9RNmFYWRH0Lc24eaF1stMZvl1S9dOm07theeW3W+ZAFmD699v0
crEVpboLPe3xkEcOBxJiij6/LgFYxFjUs4BYqlS3bKTAkUDQLov9pfZywzn2kdCbi2l9PR92Td16
zP4D0dpS0KWT20rwrcEvYrIPjJGDYmgta8rbMLfD5NvvqCl80dbM5guDt3WnTxMDXBRruqKzw31+
De6yUdtHLqXzfR2YTE4YOcjBPgpoyxZdUInr4kVGpOvNHLECYsD+Lfj9+Gptf8QRweBFPFdkXjtV
IB+gCzuh3TlHRUow943X1pyhGmjobhzoHdmPPqOLEjMqnqhhOThGBaBNcgNAYDuGWnwT7RNL87pz
rscqXl2cgv/wfWSjBYijhRrxGsSOPT9x9kXyLtIgowii5QaTcqqRcN1W4RSnBrHOO9h6A+fsWGPm
GZ8ZtouYegpRIz3lpt3LGX6QdfOZ564TspO7y9eKWc8PtScMmloZRMZ/Q4drtVm4dHv35wkcP/I+
H3yePOH6T4PPcdi/s4fjCMOi/rHOVhykUW46PQSSW9Uf21tEpQP8YQGttDp+OXXpqRqnFU97ecJx
kpwl5LmbdU8zy7gJKdqvY/eVcmSIHFIzZ/S/WfQ2DZn5aujpFHa6gNfMWJLOau3RT34z4j9eVVVY
4znibjOFEL7Nq+yRynxHnuM08uSMJEbD/p2NQQsE/joO2hnUKhTp3gBBMl71o2DKQyXuLmJQ59DY
AY250mX++4jhXDcskG6Crmf9zE7NXZH3ahHWN1KXxsCK8uw9fTqjojbLTknwBWSQCDSQkbswgCtm
qX41LB0LXf6a8gQUSBh0+c28Ev9rhklGtFqN9ieH0DVGPS65E897WvxxYOSt30X2l0LAUGwgN9++
97mztN+qj8l3vs1MojwpaOae0OGfOjdvqix3u9GietIPLZv1RNB3PUKcpN4PGxl2yv9to3Gj5PJn
q0bfSNBWot664GOKXu6HydwXWwdiT9oLjPsr/TlDxfryhzQYQaIiyMCjJx7+iHAjGTRoNrb3Rfrt
TqqrgroZkP6BH5IEAQbo5FBh6PnFhEnDsrFSsKD9S6RiKqZtQVy0cVkIPy72L1OmgYQa7Yoihxv3
Jfu96AiL9NldUtUR4C9KseMq3egl13Ih+d27jfZ14LvrRBb7cThqbi60TUBlU3gVfLmpMN0MC9lw
hM3Dht3ekO/KAa1K6piqSFQpNM38OH8O95yP16htAUPVchIdTJOFgc0quMcYVfvR0WfQ7Oibv6dt
QDzi/yFlItspFVqs+oOx3XSnIyBtNVzDizKtSlZjwWUAc66vvrmpVexLYL/Htb+PjY8ij3RtiHnx
/zSR/KoOzCA0cZfzUayVMEr77ywISXj3PDlb2IPrsp4yomH3OIy9HhUQNnZfuHAp73Ghr8J+pm6f
Vi2L64qzWRqiiYQqgXfFz5flKPa6WoWuww3XJMYzyWYTex/YIr95t0DI83RHINiP2ZKsZdpAPNzN
vr2cMyQJ0RiTrGFjboIPLK1OR4O1iV3Sk3t8JMYgoT4tB+ImRZklJ9BX9wYh+29pirkSV5W7jpix
HADQ6rUrLLolL+9San4+iAIKs5ocGV03/gxvLQ0Q+vqUFMn1D/IDGSC6j/wLkhdWeaF78uouBCWP
wJSQLWuhjrD8ZGzIfKNp7hxIT+CeV1JwzoY1PhTy/bNDFwl3r2hQ+BktcSYCnOjsOgNXIpSZ+d2c
hsEa2hAbpCjAF8fjWRyyK4lLg36d5OCVBQOs9m2fhs8UylItcdRrj8icwOHgDt8Lx8/H//ZnBLza
GtySWRSp+jH+5D5rCYdEzwtN7dsrbFYHhXJ+YWXE/zX0z1m8qKc1UEJLtVDTzE4i0BisCsuLW7jl
6TVrXDEdzIHWEBVwUPHQXPsuPjhfLcK3NVHXLDQ2zeQ8uk5uJsSuFHhNujRwIb9ITTJFw3n6taV4
yXd4YUchPH+IcnvqVliCFMyPsVSejsyJRsF7A2kvHTmDjjtbbQXJvlTdTFTYwXBUm2y9tRh4IW21
BP3SKtRa8/VRGX1Z/bLFD1krmzZOqz4IhuIv08CpazidgMP38L4vgaXH9Oo/+V2kdqRu4SE8C/FF
TXdofLqgIX1JNyGsjHKcd5GawTi8WZLVRqISxnIA6IrabqaSYQV3xL+XHtaD1eQNQHmP0DQ5MU2U
ZK8w7jriJhMrYyqlM5VaPS9geUWiAa0Xeu1uxpF6iYLRConB5mYYEuF28JWP83HWW6GkcXSD8IY8
JzYvYq/p6BbGGjJG3LdyOwX4vP8/IPjv4Ajr7xHfdiUTIjeqVFotwW0rpDnj/UMpULi21HZMpgcf
IuzXG/Qxg5IHslIIrrurmNFUvbkojMvSwB/rg7m5fXGbfcEAWcYsBu4m1i5uKeV86+cHbo5Z9+HI
K+c+4Qban3fYVhPOiYdukOAc69OFM4Rgp7IQsU0ROod/h0UO9xKdREzXprlMumieoLmJR374QU4Y
XsYcYH4iSXxJsbbctOou8sKIY6O1HivKYP/vYTAMGQ8FjrdsCpe0O8KGOXbLyzRd5Zv61+U3DBnX
UCiLyUO18sXSjJo3yCpD27kjRMl41kApjLX9UZQdoZoKPr+VwBfVXhfbTYQKeNfCJiEA05x+j/2K
uQ9tDqwMr6uh8dVEXFmxMnG0cYfHdi7hdfeehScky+JyoZh17pdaEwTZdhV+8p0LclKPeMQ6tRA3
uIaVcWa1Qg4rqgSBsgWskh+es2fAQOx6cI7fw7nHj3ZcQTFP4pIkWxvKWA9FgfY9IMyKPO1Zn9gy
8YK90UM4WFXAZVMxQ65FsjqGRQormyAE+N6itfiGGfOsnXoRyxHO3s4q3k7TKmWIEIsCCZ98KBnX
R4uUtgKJLHvFramBBTyUBVnZtwntczkNGoyu1PCzZwpNf6qwVQqX0iB4nfFL12l+HDC0lVnCgHa4
dP1fEhtRIzI+pd3Qg1OiZlds4sA8z3Lt71blfFdWgfb1tqWBHSuTPZOFl8fqmR5/vr1XUt7q3o76
Ro6NL0E7NH2J2OSc/qzOvi1YRHUUeoRNdbC9HOrl+DbWLBfQdvO1DaCIEZtNvpoNUmSE06yXjutO
ziel0nGT8OVuoALgQ+m0BbFj6xOXqd4RReDdZgJKTu/h3e+cp8zlXzJIOinQMdDy4EEWWqEgYz4F
oLhH3hdEL/LpcL8QfKyP/umoJ+s+vOw3Sx9JQDPPnulNbx5t3q5DGWhh3XuF9YHg7r+haut6IPLM
gPSEoL0Ob1GyPSR5SUaxuisl7mUY1VYH6Ge87S1y7pj1nm5wTlLiIGbhhFhuu2qOFWiUG8Q9wAEq
FfSZ7oWKgKlrUHGguWlQ4afIYdP47jwA5m8ZFYGB5Mui+fE8Ztd4awhoErcIPHA9Ikx9c9RenfdS
vewQeanxc8Bw13546pZah2s+7T3NhwBfOTqqqmx7YsAev2yWEkR1vbjFzFdTOKjJzxlSWwH3pKKb
I7gX/R8qVRVax9GgTnbyHb7225IFKCBS0IEkEkjg7sxRNW4s1Qo054fLB0CK1c3maKyYXvvgr37E
ucPpLEL/hqtVo70ZxPaZkbG3/vgajXWHUydfntcdKHkDa/nRh4x2VbbgW/noq52MdkGu+7UHdfPS
WT4RWcaLdtr06HKYX1CFU3X63HAdLmH+LEf2DQHXEMWwvFDM4qq2ZemRKuPA/odtWjg6qE2UoY8r
ra7Z204GywT7cTJG3U0EJy70udRm3Zs37PUT3dIKnLuK2Ebq/AtyjkPpnRht9DZZdDBcUjzJBaKd
9l2oyRycfrJJDVuTZeQ8pdmQxOzN9Kx6+UtD/2/QLQV1LdCWvJ34o/8RJlraPUC4553Gg+E6i3jr
sgZ2f492LQ3F6no6yZD+NMkjNk2oepR9dXzIpyYQs6J2Z9wIjuMe/pcTeOM1Wk0JyJNvnA+rXhU3
njczHkCdv5VR+e4R9fqOmerjvaPN8dabOgGU45SHnOP/Fac0yVFJiHotwQG9Zd3rQoXVqSq9opQR
stpTyTT+pYUl3uxxdlkEstggUyKdYNUp5W2zYFGOIdsBUfTJiA8nyWp1UK+7TCjMjKr734fcyfZt
zXBDTLo+FX4xIMmzVhQicPlJ3kl9Tv6KS3/jpx+2xM95R6izC7oqlGS34F6DkR7AoXUMF+O/WucU
VCuKAozAWm7LDZ4Ar0tmNMKF0wHyeljr1kNsgK79P8WIXRNcV/JWpvKRAk+l871/W91RBRUv5F56
oHCduAgOW3O09BytXZ84iEnfVW/Ew8SIdExHpikQuwwTNKs6LzSmXByZN2P7bxqA/ClAZ+Pu//f/
t4a65efbkZIujL+nuCWqJxacv2QiOQshbP9nJBOigdyGYf/CoovTqGNLlVwWBZoXbfdkBzvaDlYm
iV4juaK4z1yflPCmk6CoReL7HRtlYbsWPURiM4DbKSLHd6M/RGIzD/2sAUBU7wZ3L1wZmRGplHv7
zMsbBuUHuGFfg3YMP8moCJbi8QgYphDaBMsY3n1YL9iey2Hb2GBoxnfWJrRpkaFegObjj6TRtsbp
2pHofpA5iE8SZiM3ECD8piTUtXI9ABRQl7sP0whHvpmfEaN0KUt//PNwHrGC0eNpcdd4DZ7lKqiS
vTKK+C2XZ5cW58dc1tZn6QtPfVDzvQm8rOkTB9g43zpcuLa2kUu4npi/cyApst7GoQmICqRBeUZH
Dxe/2VKE0QLBCZfytgynGkr1iQD1JLa7mi5varMw9D6sa65ON9qGmmDo77zNLv57wmSuFi5z6HPA
VNAE92hWBXQMBOMCL81z4PZLTtmePvbfs6EkCjkcSnCPBXEQglItTkqyy4RvRkeomAW1xzwadveX
Csrb3xEHyM4xduGc/AVpD2gA3l0H9dNeCIjcxE8PNw+HG1Qxl9Wr2rSmjwvj1O2mz6F8xPYp/ykc
N8N/jLpQmjKxvg2qIuWqo0Bn5t+6FERBs6hkrLK+vSicjrTAqj27h6VFpSSILq1yEy27oNrmu9NI
2tGCr8mfSaKtyrnhNuUhpCE7InMkE49p/YMIFCGIgxrnKXZ80u0DZieCeRn9S1INkjdMSnIAKgQ2
SOBtuIgnpqlaLs0gaqEWb7zfhzNulOe6coqYZ5j2a6Gl9aGMU1T1EdjTu9PFvPdRaXPFn4kcTNKj
Lr4VrWHUQIBQtpox8ww58Z1HU0bGShzeLuw8B5z9ycrkgPULL0YYoqliInBKsMXY7+bHDMoCSkzN
dYTgyREad978+LFqq4wBx2CAo2cLY6kD8YBe0xVW7P89sJH8LDPy9rMGDn4EYUvPwv5vYmD3scwm
ePUjOfM60JFy13p690Ap4aDfGjfkGpcpbs7q4e76Eiqt5j9Ese7DR1niQsnQn+wR74GXy4LyjJsE
XLqQ7tGYtbh6Y1IJ5hDOdlsDOMv+Z+HI6iT4ZtQQxZiUF0Sdo+Ia4NDsSwKNps1s2VoAN8XKYwcf
Pw0ujWqZ62dQkwfM9timZAGFi9bSb/0VIYuoz2nKRuzPZcwmAdpK4E+obyFqUT9lu3TWNpOImaLa
h6CyJqHmUtQ7TB76bNgTgApokKUuD43jYQofvT01SpXyxgyzb3Tv+xBn0OaOckHJ0UAJzmxcJdkT
dJh7iEr6RlRTCR3CqGwD2BxTnsyDHGLOUmfrsyBw9JHi2CDK0gzLZD/Ud1MXZDIW0HAKHabJpnm7
kvdp16iS5JhFU1v/4xLcE3BAZarF0ur7i1LxOdeqySsMaIl+U5I77WvAfD2kDEbbQy/ms9cb8bkr
zsZSwourqFRdHl+sMeYIy2owRo8IPFum2Tf7DJrWImKc3bmZM0hwtjoZs/VsCeXbjYzOSBukOlqd
vzVrp0Ilth5dx/zFwkDJoDC76R1IWZ80eLHkYGYiO3xzNsqMI9oX+2FEbPd1MyKar5DqOQ1RxGaZ
NMefoBy2aFu+xehjdkmLBzsNTzTPOmMD9qA6IEtz1Gs++yVegjbVXo9vW56vjwUWly3UP7cD+bBU
y6sD8roseW95+FnfZKROBlSiEZ0oaDkg86M1YR5RJFwY7GT29GGdLZiMDjtirdFHgfQB3Rg0842Q
mkJ0Wza+Nll/7ZeKNwQz74ZvJl7QNq0e8XLDZHiJJgUNWu33tXcYlAwJrHy8pPQf9Y4rSRZxMOn/
S9lOZT4yejQozMa9Qf4iPnbFFLoUMXDGQzN7VFMyveo/qtHZIH68ScG1AaXzLskELJDV6kJZV7vZ
9DV/zO1Akqyz18BFJUapdKcDpflWL0nVGaxWHSlq4cNvI13knxj1Xgim+8YISkNyiiZ8rn1ujXKX
Sqdsdc3DeihwVoKVEUEFkp1lB73ySQr3IVcBOPIsCTYIdfQdudHzKZhEG9VM2mh2AFrXHSbAJoi8
daa1YsVmP6msd7/drzcAUieezuFKP/7iFEytm0XfN6o0S3Yvyr7qTcNasCInnkYXxIXcGL7H8s+i
BoXVSyyfugXgQ1bv8M3PvJxakmHxqW2e6UZeZxPgxdycmWLUZ3nmhO65CkAc8JGUf6KH3yPClf8R
GpmknjCFr9a1Wggg9ZlDyatowawbKo8Jxj/zxnK7GSIYP8WJ+KjSzTsURakMbTLCqqOsznWgLYhJ
dbmeHE2WwUI9shaBJTQ0cNx4qQbiHt/7xhKJ8gMOgb9Ib5YP/JnqpGTyMHgJsH6Q9V94fyKtGzEc
igkSimsryf8tyNGvaoDhIeyeSEOrcNrglz7vGt+hOGW6BHVGVdpcSroq7hXaPhI15KaQqhVCwGrO
7G/0k4bVmNYCHD6YLuh83b9LzksmlziXEAqdnvA6Iw/6Gvh03PjHlVdeRqCW2vVhIQl9b48bg21O
RrAIGi6wizLa8dCretis9kogftltfaQjNnwxCuCOcxwI18Lq32/JK5XN0vfvscpWZioSkCcTa60p
PhSQ2koYs4qZI7AKqqdz29y1cmqHzjELPjdI9MjfVOFNsX4eni4x6W0r9WLnvxVOYbSveBZeTgIZ
XPpWgqdcHTOxBH7BCd5/9mROnXXtTt6xjJmydS/lhR2UDb4vbjdm6M2KgjK0vt2gqbV/tO/s5o/d
zoVRBHUIc++qZKNfWcg9KCxrrMyuPAfGLLYXEAZWd+FfKPJErFUfKAv5u35mWPLmL/v7wdfnYS1x
cjuDA3moBamfg/bXj9d+8zhsB0IowMJ4aqCK9m+/fzpLZz7zUioQkuebfNLlrAqVk0gZyZiJhTH3
SrL1DfLAvrLFXvxIQZAGse/GB1vVI1iEIXUy1uaZn8hdwsdrzfKIxf+dvZmLMaMZfnHo7Sx6bfXY
JJil3Y/ta+Yk+W7sJ/CIgJPv5/Ho8pzCUujfctndP6Hwapz4qJv1/D2+C2vAVoLCL4gnDmtcotaH
W1IYyvBu+6+Nc5EVCYuAY2ANqH4tNDpCzV4lQMhcNauI3TmtWz3fKKkJgJ30uLj+plyZkCtPF3f9
YEujb4TBBldv8EVVHmTF+iEtQH8crOub46cwpOmWIj9sYWbduYg3ErUCsF0Cfointv9X8AeTBCN0
nok0vY0I4kPKTXuxHt8FQyfXcrbY64quy3cpJgs7WGb3qKL1ZZ8CKajogRzrpXHN8EytpZpEVJAF
Niia04nKkfXE/xt0DRGgvZeG0nCxz0kgCA88O0ajeq6DtaVKDv8oleKapVqu2RU/zs1/9UUgWE7L
oB45mnE24doChR9KTWjMd2ZbzxTsg3BfdM5LDXvSYTXCIkjw8lhfFJXnXuDrOAfzvYnevetHL84D
Fai/+xcD+Jqhvie9XTPbHCeLHzyNOKJ1kbj2X3HSuLMgX/9jLkf1BfTLSzRyYoboVR8S8+ysGBA8
fWcIyb7H3UotG160M6aXx8r7iKoYdOV1ZAACT9EIo3A9FTGqS1vbFMIeBbAOTn53qnmxw/ljHgPe
wCqxbvt0bXegORjnHFb0K7J74+zgJA73ZOYTswnc6E0p1CU9YHTs6vWCojOBVcSlkEhPyQ52bZNA
IrBlYcQ4h3UJcXOmy7WEKeZmfMjaAmmwcg5hBbnw7KXDR2d3S1SUPdXJmj5qWd8RPFO+lcmbj73M
sDcny0ZXelOlPOq9Q3TNhntUj+NlPBigEuFCDr8tdmTYywRfohL/1bdoUHXY+5LptLZB9dEfYHUL
R5BKFxAdYuwG6H5y995TbMdVPe2j7LaIGuWhbEWnRLjA+qxYLav7GnTh8i0QO8Ofc3nAVx/rjtiF
JctVTzAO0gAvVZnoqJLAumhXmLT/PiyV50lXSCPq7fzzLSRX2v9QcSTNX6Kt525t72WTBR2JEy+c
SeDoCnjuov3IF8ka5XFs2SlfbqYsefYy+YOXLyskcwxH59qxcOK07GEMcOwDcBP2GmlQEyK/qx6h
lnrJZSeUOr7YYLGuwvtQq9L2ciKaGvYrQ0blmmfnNtaCWpTt0VclnFd7ntdQHqOXXUkje5ESotSO
X3N4mYe8keOsYsGmo5wianKLh3y8BuP5kFHUnMMUkjkxHGA0XTyCcKq/RpYYTMGovjeDfEwOHBgy
PpIMXHkRt6BJsYSQxszcbq+LoHP2IJ+rb1cUptB6q5UChd+uYeSEfHs3s+52ecjSJzwp1k46jDoo
jQxOLFL8fmktXZ94RM3rWJJJdAA2Q959X3TKNt9j8gLmaTdF2gkKWhowqiSHnOMhosytQu401wqn
IYI/OkImqPh7PKvXP0tcuWUCoOducqUeTbP5ayStXg2y5Q8oyAkvCNYK/bvAn3EHYVyA6kJCb9wO
pdd2EVGM9SbjTGKzT95u8DWmCe2z7Gm1QJm5cWVR/d3xHlDhkGzdzmPGKChfesBBYugnAbwMUzoz
BJlRvanhR2ubRJ2sFHugKyqxVNpJ1vq8usOvuukfQBtbWWd34J9JNhb7SEaWg3DQQfjDIM0EN4Ff
nf/aUrOn9bQaI6fPdy0mqdBn8+zTqv1rboQ2ryIGItm447wUZJshrxoHybSmKdP8L6YuRYLRpaBw
JJRb4SzwZ53sl1N++x3zXO8tORXIgWYf9Cvd852cJQNiTL4scNy7gqmIu3iMwcUI81Wyy+28IuEK
0u1E8SU8VZHa/aKfaw6lCKpJydsmF/BKf6W7DbU26ZofDseRtVpt39Efgnm6aW6pkhp6KVfnMVMs
xyVgqQFkPX4ul17vL0yKgn9wB2F8/O34/RViZDQklhyvp7xxzkHR1EalCNdHbjAZtcG74EYtNQzy
kEqCVqa4Sewn0ckoWQH84mTzHaDaeo9Izn1M97bl6WmHgXN2gG2C10jv6UztX2z1YKodY+dAiTvv
illnUto4AkoHeqpk+8ClEa8RnrY+FykHDn5cEXf0phnJfSuynhM88kfj4ZAhmvB9n5ePUVydNpkm
L0jujibs7ujOMFHuKvx5x9nf4iqHW7RUb0EcwzeRxnV390JAP+nvsJQjHIIw2DI/YUyYkF1ztwFC
s1htOlxXWZrTdtFu9liKnJokQPziqbaJvBsEItB0kfoUZQiSKEm5tAdi4yP36cFplzCgZgnUo+TJ
UDsqBrAKTOX+oJbCbg0TgCCrZJU550cp55Dt7R50PYEgHixz4gzwYXO31P1OaStQfaaTvTnai6yd
X9ChoDWkiv8KYfwohvRtmoVwrJ5ItlA6dowq1qIWXJMT4LFQ7+yF0R+OHP6U4pzdy2XXYne1hiIG
PavHVqYYBfmZxPmfybWnX5HHmrp5w/KDDKP8WP5p3TXfgr313yxswEP3haUm4knOzC1N3w30y1gY
sj4xXvLNfUVXn6P6rAb3BuYKJaNUxLu6chcsXez2L1BuGL4FHgsAKhpqHDfvFeubzAfqswBRmz9a
TEY3zktrTb2QSKu6hpH2GBcbtytV6qXJ4dNKCSIZiQpccbd3qusrBAx0vLe7/4LZvzbG43Y0TkFT
xZJE+r7cJrxgHGjEk6fLQ/grsGAWKzSYK8fiLFsIxzPbL5ABscqVjvo4sP2MoAkm+W2GmQKCDRpP
YhsB+cJjz0Mh+nZtahNUj4yGseEB6etva6btIHJuXyiQWtGUTeen7/CkFYGh5TUIthJuPV/jCYpY
wo5Mxq8mY1MdGJo+F3JuUAQEPUZaYX7Ku/n9ZgN4y/OhYO7vvgQquWRIoweYp+lngLKCet9rAXfp
PmX0pK851owIhPh6dUUmHcO/I95VYN1oGwSIy+pAslx9xtb4PK5gJPUJRo42cXciO/mlgOYqLI/q
PZO3pHyIp1A1U5tc+xnICn8NsNzKLb9tGm9QFJ6hBFkDoc2I3hNs6iJ7kab1O/Ywcp9SbAEGmKwk
QJhE/ViUohz17m+Z9KmBDnreSKD1scoh3274yL1O2W88WJZ1eJVamAyQbeymODqVw+08FMaMWh9/
0eu21A5r+jDe1ENrHaouQ7kslRDUjNlPPWyfPzUNT5eFaVsVMlxQRTeBrxQ18/DC1SdjfPSq1lur
xBg6jk1ZlQHlAnmysdMLQutl3I2q3XUACOYY2D1KPzEHfK4Jpwj0W67G2tc01CaFmrSqSDhh9jqQ
99JrW2ynVDwj3qj0jNKBuYUVusawad6Ub0W+fRDROP9pwGJtpX8KkE0RAWpupyKbdzvS9w/7jTp4
A2lu7Q7z7sVkRiTkaKN4tgerJ09P4OojqqWlr5SSNLW1R61VbLtuGZ88p2pk9UDLuRCiMCPvE8f8
nDh5SZJ8Dc27fmHUfiZckW4ma0hgekGNcZ/ukZFOT6J2v8yESdswNVkxotHMj5zWgm6ubIPzjst3
g5QwH7pp1omtHWdlCHaQNoKfxfDQBZTkQ5Ht2yLAYoYD2AY1ClK9/EO0OalrG1PkQu5mMoFfUjNF
x1IzLrQMWRJf05us+iUNOggWEkJP8rSFwI2dfBU62RjgW4TQSWbP7JgTafCgksLezk5Nv6VbC9U9
GGFO7pkcqyewyRX6vyvjHBjkxt/FDKQr+noK9n5Ri5qA1vQIQOtgF+ONb1cFTgowM2Wm6aHjsce0
oYr4hachVwdbxr3GgPeNIKUZSAFfpmi1EW8PSUdvEQKuc10EDBlgkNg5i5Ofq21xqY4tIwnVQXNZ
z5AswzTRhLBQzS2mhUlkRYcUNcWufJvNmAjjLiBaYMDNUoRrcqt9RfnI/B5dbhJOxrTuqs6lhwfS
VMfnQ8I+0j9mk92To5THTLkccG9YWmK1rG6nlHJwVMzZ+Bh7I3A1QoS8B7xERlwG0jUPSgkuxvRj
qtDMbLFvP3Y65SYrIjaIFVYFfPdbJVDx4Zm2CFqpCtc/Wdpc8ijOlJ4QTyfS8d9dpPpB1gFtSiX8
gLRLA9Eqi3H+MVqV4DPD4GVvGKAOxC/itNbpFHYcWT/u7/ZN9JBxEiQxOmn7V5qSj4kI1ADje83T
sgJ5o3lSLilbkhGT848zqW1NC5N5IM1Ifsm+WDK7r5MIuPzvn3++6j1vbmvy0DM3/SRWkApJlB8f
FIRdzn614cQ91bLvZuZ2k6tdj5GRu6ShX4MnG9xvMt1X4WjmApfveVHJeNxUSrgpkEqy8rc+YAql
vcsTolbq5JnJFUUdt1sQgKL4wGe83oqtsnJ2xEjkKH6XtuK6GTqHrfxLr/MR3FXXPV8XEO6Ya1Ry
RDQI5oYyaUApTiwP70GhvZrbWP67W7Xs3DvQsm0/m/YkQW9yygl5VujWCiwjCzH74UCd49OPCXbm
WqB8aGMT5jgchYAeWQUWAGSC6djoncDAbSAeBSS/VDEh900jrDuq4ltrEIcMH4hl9MPBPmZuFoKB
Skps0zoJLGMvQegf6F2pIz5/Q4A5qvXbKlamC6em9sTw/BYpi2e/x931TtIHomAxdaV8/jZXDB1+
kPsW06r1v/D3tkJdQ8Ul3HIpE+R7k5cRWDnJjo/37REEvjyVkPcP0FCm10hwX21SH2F69Z3F1Yfs
WUhQ5850ZMN3rntJxatmENKLOI6CyfPSmYpj+ftjbGh6k6+crzIyrflAz9RthUWv0bOV9od5Z7P/
EtANakwYEwEfLvBSDdI3xZwqien+QxKiv0Azwdbvmg1LibWdn//ZxY0O/EmpnUzzClHivewIAr54
XnoJyp/ByUgmVeH5ODLPHtG44fVOF2AZ0P7/1piAPx2WuP6mz0IeyoJRXFjRi/Hfwj89x4deaxUT
8xJRaDYHIITosU3cjEZKrWuKn+pYU/QpQGPyPKRZwrH3dowRR0HsFDsvukHnDjzZLQftYXiq8oG/
y4ts0mrHHbaGHR/Bt+RaeRxjLiBuUlIKXs8KG+QGW1/TtyS8EuaewkRlSnl4aLxzWPf2jA+eKqLw
3oMiG/oi82ycfl6HgmF2oWrhn/9dOQ0wQFckV8G1TOwczGrf6m7NnxTrLDefs23UkA2ItKnlETDP
Y3Y9PKWgfmAVLsO/2s0yPPd4EfghaYhbnlUsbZTdisp0rg/MLeD9qVGvmvwqadE2A9uJU0+u1qOM
AibPmGmnWkFRsuXGKXQCbPaDpN0DgD/dqQVHRrl12R9Ldmd1TEWGjF5QBQTrXuXDlHQ7ixVaNuji
lGd8LWiH5iYr4RJegSTQyjLhrMMbebvIuUE/jWsQisG5sSOsvHpyynM8RN4TleUxWJRw/5ilPckT
AQiO2/cof/vu0ayCVjeivrz62TA3gfCmw6hiQ2jhCLJu7Odiby2L13j861CIVBYm2eRS7MenIHaA
ld7tZNNiG9fpdKysHuIKSm13WDK51vA0sH33yYJ1NWYR8xGLnHVAKiX1WQH02EucXGTi/RSBfFC1
sLuFCrK5MfE+BkHi7uYhVEVqIIlPuzsucmw5XS/PBlg5cu5iIRlUhMTm1GnoqLSdHqYKKDUe4h5k
auvGYiBM1lKWGHFYNArEBHFtVVlmIjO0HRxbNpQL0LS1LL2ldOqsdql8vTwTMMeDhyn/+YNrv/Sl
LNhZa6gaMa+7y4DNjUPjrSHokn3vcz7rahgkeH97FFylJ3rR5KouI/FYevFGdqsSxaYLOOnJaNFb
7xeYK+Si5Ug9hpVVrqwW8G3rjAWlFdSMOJ+aHzNvK/q5nUXbGLcOTPKSbiQYUk6zbgojCpXuBQCj
/9WHAzRSlnx7svgi4SNAll91GGlNJ6vOhNq8ejDJL5vUmFqcezVOlZEYk895or8nZSK5n9A3h7PJ
sg89b0ayrPKu4vbhPkou035f97QofEkTZ5LctGec1kpakxlAVBJuVtmkljm7e/p8Z94GUMPzRqom
2Qq6ffutscWYdzMX1uqtgLDHOReST7An+ZD/fC9an7fjiXLzkqiLT8FacWGQ7j1pFosjbH56JLLU
A68YrZQxGG8PcJoihTnlpCu6wnbcA6qGt200Cif9LI3SKQIuL5EHHOYqHGv+aZEBYQNlGpBXqPSq
K6Yoc1xHmsskOaeQdZjNFmdq+zRJu52WoYwSEfYSST/06nexoZ1N2JBaUxdIPl+KcjizA64KeKjF
/BuBIz9FPRRxatYChGswCTEmFqj8FoKDMI1MT3PNEws8YiA6RkRFbsOmSd2RzSZaCXoPdkdABDV0
NXxZYXVWuKTzwaerzeuB5vl9bYYNg2ltTNkiAP8357o2X7wUu29Q2tjlIGy62rOfEqEnyQj79ouC
2gw5olCetFaKb8tQM9yeC1606C3lkqBP5aBRpAaX0NPwQXNvn910yuZ1H/Z3Qo0PZIOb6dHxHhrw
6jeADOqlktWTdvy/cJ7TE5GRJpD9lraB9WqgrqBajCOpRrW68MyFd5oIePAdiqE2U8MuEbW2UY7H
m+hqhhXnYHrjp3JamwUsWeTs6cjY5sWLbTBo6cF+exs1UcZHJrtfES9K0qpFgfJCjR29v8ut1rcd
D49Q6O2uUq0NEXqPVGpfo220KtCt7cCd95Ghllz8/LRnlvWjKwyxiTQ/brb8g4BU+GmHcysz9Ley
dMaP3ckACtQKYicbMljaHDJgcXjjWWwzQCQR14FqYbtX4NwVmQ31DCHitCXkYP1w4YmCQJ/zuilm
5LDWgHkiDFahsDD1j8ndFuVLtoXLOHoymFQT39vtb2G8RBu4Mo4sdwIc/GB8WkUECqPAB+s0Gxz9
tJcqyw1oIZ/STgTqGyGEpIdcCZQqP0z5v5NteAp4SX+COtcs3h9e6cScxXkgXs+64mZxeEIpC1fY
YsX3EMjN5GpDWUHLErGPETivXMA/q3oarNzJvyW7GVtttJCfHOdr4T8hUCPuc+yEX6VsDbUXIdPt
6vcb+tJZ+M2VYduVX/5NIsj4mllVnRk1M2XuumkuIyzMLK6yDM4//H/Izvvu+QipYkH0OqpMpNwq
jVLkalGzFP8htCNdN/Ns2UL/7HlovRVsMw/0DPRFRseaTOqlywPP3tPjZgXVQlWeI4iXjLerC60T
0HdivV9o+MsQUUWfCU9io5QMEjXsSURH7NG79KHsxL1BczjjSwvmaxLRciaHBEMsIYqoFqVrmVph
fsrBYh9pPmBuGNj8TKmiF5A/WwiO/wzeV8Y8+q68a2w4l+2Z72KTgFqRPjmmnEDXNmO2JqV0omek
CyD+xRqoaeo1BFth8awOq1LVr8mrVlT45OjiqlMRxH1cGX4xTLnOqhW2nBliMRW3ZFdIEv2bF02C
Xa2GKW3BG2Cld52tnRbcV0LYTSBlCY9Z7ibwZVlTj5TBNJILsrazOVpwflSBjxQLSa5Epj5Pok9K
7iadOAURfIU+OE5y+aaJcrXice/ulGPs7mZg2zUCntz8edUjtlXkskTpF2Mtam1zr1DL7hLrVFop
TM3LLyZYUThMxs1xC0CuJIW1NrDnSS9XE/EJKqEpzxOJ4rrnnjTv3cClVJdBs7Q3497HEzF25WoL
EV/mD2tNgloKvxm7DlgA8FGDS7iHeNfyUOjvScVF7vNhviGhYI+K64Uh0IfzZoasqb316t9ged07
LflPlPfUWcdlYQ7a3WZjb5avD9tR4Z/FX/V3P5BN5a1CrlmX5byE4cd/RKlXf1WZ4sGJYqvrEb+Q
4LYeFBUm6jOTGPcBmEg6BF2YMQEjvIZ7SVd1f9ncyYluy8A+ZxQCkpZIFjE+MzCXUQWUH1XSUFxI
CflJhYGVDbkbrmPZqcHOHhcBqA+5YV3mjmcON+rTdXCDtKcADVhZxDMxMbSRX3TA7nloUsqOFLsj
v0oH2+bCeYIZpC9ee4PXPkKSO8jaxrEJI5QP25ZoBhKLCWkuS/5ev3hT7Zbe2ULH1285+4LtQEiE
mdIIT8cmhgt11BBL6rV9O4liFgURWMB0GpPtyXnruJPZnSEr7n3UE5WPVMTjAOlhHn8q4D8HWjff
7kMXenvJ4/TEVkAXmDJj/pUue+71fZ7+G1ElUz6GDdz07HPldt8m7d4aDLxIHWG6VkwRYW0NdDj4
UF04OoWWkIRDEQfQCcnidU5XPf9x7sPMgIZFraQsg9hb4zymEW7l0tvc7Rn4ac+2OpNdAb1FT5HI
LnwPJnY1z1WZRP1q6ZZCPWrDRVDc2yTbYRwFWZqWkU4vB5adaf8GyBAzrnwx1QMIaFQDveOrZcj6
dQQ0vENV2wdevSX3xD8vnS8UpP6YvxiMvE+3OVyGPWoFQMVCKi89ZGNHCh3s19eYZYgN7LUmPs+C
NP5MX0IhE2QBUI6kDkga5xR5QTB/DX5JKOLufBa9VEXlL4gZmtgabpluX3zyiIzXYUFAzEqDk+q0
Zitne3Y5p21nVEqTFWkmpGhqMdnl2EMeo2m7pLblLVU8l+ivOnqBVsCvBcFtXBf6JVYPH+YfPgP3
rZ5jCjc/6IJIxBolb7XwWfP3DViA7AwQbrV1P5l3n2KQ5DhBqgVu/JZXwmefnQktzDeQNsaI7jVb
zOYkezizvOFa89J6rNUmeeADg7uZCruk+BsfyJWKfc8Eb/ifFVpLIbAAvctedgsDY3Hxg4Iul3Mm
P83Xk+ERdmr+GAAXwVVvjsCFfZMpHuR3CaFZI15i+ZzsF3wgamV59Mylxa5lyf65vnhkLE+Ol1E5
ixKajBbCYvgbhskCegHDD9GmUx/61lFiBprAuMasDgcgJyicfOFIun+8xWMQklKhiXCcnVc/ilTM
5xfM/kVbxbjAucx7YmVTagiC4Czg0AH7C8pn1tin6pE5F14XS84hc5qoPaX4+ZuwrqdLVk5H9/Sx
9QgqLknlYWtjxl8KuIz28nIX6iIyore6s79rAxQ5mDJlHlZ81zfylVhDhjJcCgG0YFqR9supCnsZ
Thcri7qHYEXqRcXpwZWHLfykfhEKus9jrTKIrtTlugvglzzoiLRV2fEsS37qkL8vuBkFjhijoBT8
iyRUqqMUDnttADuYH1/mW/mfaDKqoJmxJyLM0pguusJOyOcNf9rcYjsc6aHmBUZ8NWDbLddtlS9P
qQa0vOwDqlSnrYO2APq/+GG49GpwPHN+BNiGFYNOeC+8OmAu0O44PX4RoZqUU5rCZiXaHhmZWX0W
cv46prRJF3+majHdON1oxb5fVD9Bpg3CBvUrodugTJkb9ZEV9B+JzVgbQjUhsC6YPJaR5/cRgOz0
jrEZ9eP5rKrkgCXas8zXnLPLLhSE5jKnRWmKT5cMtQswBjbCed0Wtn6wXMXrOKQ4jXaLbIGuKCRe
7m/Ku/J1b8PQNW5ehwaP2LfxijvDrBWrxuuVKiqMLP07m77x6YDS3UrIGnRsqC8BChhVo2Sp5QMi
g1tAS0+Dw3K0T6Y7Gd4FOVTS8P2yRLIwFVuo7ovN7fL8VAYNbOPRi2Yq2tFDeB33T3Go1WowwrO4
5vpcijD3E9tuD+Hvl6RC8ovRAyhW3lnOhr9boW2/7iKy9i7TU3YWTO6bDIpqCiGWu9y0KYNRJSla
0+SaKQwmqaMHVjIUrXOTYDoLKtF8D1wEvcS+WZvAkpJ10YUDd7Wu3FdVQ1CfGgKOL6w2raywdQX+
zTptRQmPASdDw+F9T+13m2EPPVPFWGrbMrHat88vvym/W1qdj/z5Pyjf9JM7WqRuj5GaT5rm/Jq4
UW3OoqDUz9FmhwfUuCjyDiISeWi1TiK28XYOy9fdsqCyUT9SncnFUH6gPnHI5L/gziTYjqlFdo0x
Uqu5XKefCvncvOIIROz23QxLYplTqIXrEDCGpy73Ij1VTLOu8MbrP2jylq8LOswGhHtX4dzvwww6
TMaOujzIalXXxq8aRzUJXNvMhTp2qsRwXmg9kMarVLvOoDXEiZfxx+R0OOhANSPI2ODtjuD2N/Oe
fZoIaHwj4YyZBq1WfJ/seb4u+yzI9IPfjmcTRZE5PeIarLU8gsp3Pap/EghiswuOc8Dw94Wfx1d4
RkIbxGilrE7E0DbgEoFb9AFA5bB+I+6M6E+IW9s3xoezPUfIAMJZ4ZfMpHjFE3mA4vV3elxiqJSs
4jTlWkQwgvZAu/TG6xRNsdwkTRMZ7VP1mpgBaYUt+fSGsQIpUSZ8LY0AW53vguuHbbksampz57kv
m+mg1m1blqZ6EZIgyBpd43/NSmMYUmbMcvIi43jzBZy+KjCPdQPtmsREUP/Olqbd90UlRtGzYbmk
gXkfUQ/d+649AvnmT/lVoQ4sVRoAuCmjuWn3RWfsdcThW/kwRXNrH+RBPp9fPQA/gJAcuZrj0Vkf
bs1s1HK+BUXC/Qo8mm5JvJ6ZoSrdibdCrAqrVCctFO0ZwI3X3Rs5WuRH2A6CS090iDE29Cs4nbDX
/i1EW8yP29z5vmm622Uixrg4KjYth7jHtO2vy4iO56mljo4yhvPtnXtqA2Mx+E+r55iI5mcc+wS5
3UvCyGOzuHPY7MT5SwQkkUO+DjzzWzAOM38f0jmpnzf+GHWqLkgv/r1k/WrU07D2VONks4hgNSwy
g+H4IkpwkBtd2yCEXlKXgNyqFJyb0EI0Z8+gmgcIOQSn1ByH7YfmQcHs3TqJdd4hNG/tftMEkapi
zcIf6mdscLRb3pLeq6lkjmogg50OkHpF/MY7Sns2wHIFSykEnlGL9POPkt7ah0BFHXGS24U0ZEYM
x9JO9VhY82LJzEKMUbXYQVQnEj20NEG8qHZ4HhLjzxs69YlS4prLUJV0F62sWqgqaYqwLl9Fswl7
jbtIACAa2VCW7ZchjFT4nf0H3vjtsTl30aodxDf/uDOSCaacK3Lc9uTNS3p8TZ9JhBzl/eynXgMe
TkSoOqfb8MT2RGO7DXJltxkPbXq3us2p8AXbw5aAvx2HJS4cxJyMipYnwSeGtf3nG7r+WXPH2VAm
8eDl3fBd/gKEVd4800FgYgZy9JZ8KhsYhc/FjOcG7zzYUrPFSwGC8v4LuzagEJgA0fDSzBs9DKEa
et9v0dmswTgQajCoIa25LoTqAPY+q+V4qoCIR0jhEeTz+5koURM+vJcAmlh8Mk4mKjg62sRgjwW/
2C7Av3L/RZpB0h5f4HUr05YGs52emt5MUmMJgdg1On9if54HhNGN0f8LaUezygbzrsUUg7gxD01V
TUAfrM/OmOyEhTaDDHJ5HaJSuYObhpwHRc4g4dcX+FMoFf5NixosM2Rl1PS+B2kit8nIqEDydPFe
G1I3bg2Lf4R/Po6tn9tDSsLRvVaXf+JxnMhDOaw9IENNTLOTWXWh8VD+BYgim65UoH6ril9u5Rb4
xlOVnhhqXV1YXSdRRX5WqJK+NhoR8ppbc2ewtRpwihOQA0fDGh/8BKQJo9FpjEppuSZQdNzsbI+T
+Tpibeq8eKmkV8DBThGzzgf0DqvGE1bzOadtIxbUz7DhYJnw5i4wzYLivu8WFijpmKY0t1YZh4oG
UHUEqrpA9dhHEx9QHLwSYiLSSScmI0ewtxhze0Il5ISMaVzbk3i1cDVo6vQvqMGgJ96p5xG96dH3
4+GuDn9Ke3ePNAxdhptIpbStM/W5OOaagUM0Ro9a8O3LKMhJTcbu6nmh62PJwfPTSJBG3lpGv2dk
Qo5aE5Jqnt3dx5gJUPMsEM31Xfj4sT4H53xRjuW7PILyZVmulIgQgHevw9oksqwSvv4gY/J4rq4s
33iHaoHsgWvf8IoIu5wRn7qjtxWiYrdIZp7YCjps+0UuAc7w2dSqyski51uqnlhr/DGihFfa5NGX
LXv66yc2Dsuax+L5gMaNc4t5iYhs68Y0pS/w9S0duie8dcvH7nBDbfanZueJqraXOmK7usRB5bA1
r53crwymWr/Bz40cNvDwmH5MyRXTlsgJfGSrRWzJHT1T4JQ7juxzpSCJiZehPMJgfs76h6Ls0SCp
gtbEJCwh+zcy9J09xSKAFaYxcBoHdzoVh38umnoG5PT2ODBc+0Is4UeGZPuX5ah89WTeP/h2Utbl
ELobYHRQ4PHPVNKOtcdN2fDVjOMTMoEYZe21YxYZWhfMjtsiytX/Lhiibiw7Hqu34GImsFJAsspG
JcX9Z5uELg9iNhp3uBJe8TuIRlsjYrOGG60ZaA2uUjCvYwaoCj9gKyWYzgyg++i46jw4ZRUw9CO9
Cu88AyMfzo5qWv7+eOtJqrdDP6ehHn4+v+y99tWkCTTN3PbtKgpR+8m0hA96WU3Ugm9Fwtw4iXyg
v6XJ2K81u81ptSJRXpCi/KFt0CwO0yCltA1SE9APpnZIJ0TOQYBOZB22SaMrWCRO6R+jL37ptvou
a1l9wihVf3f8vFH5uKtA17hmuFLyDr+S/WM1uzairLCeHK282V9U9WAfb78l9ViwiEm++lNaRwLr
l03coGUkceoQmpxBw9NbmJlzHUodc5qTKQq8tJsXlFePD9V6ZQZY1qtaBDjp6Fw6pFpOolTQvOMQ
gwGYC+Gjrud2y1TBQTZGpGfdj9Yq2l1gE/VZ/a7a1TmxxDPgdUfPEcskqzbcwpAba4FwWcuBeVdr
MrGP1e2EcRO/seZ/WwJ9HmCXNRwBKr8+zvZoCmfUWPLGOQA/9f/2+8dCA7ie1GH8guHVe2zotCko
7M9/Wl0Ph56UDzlxvXR4EgUdXeZm1PSwH09gfvMVl2PE18KEmxKrEWoK/C5BHLDUwdU1W5ja8yna
A93H82OHNZpOG3WEiVrOPeILjr2sc52n3GOdZy46SWShPz19kZiait0rOe7EzIlWkDlf1Cdwevib
Q3hylSV63Npvx9A6ZhEGtKBxeFX5HTSdbyPml3acsOTT2b2JfmQfvvi+GzIxtYWAOI0VWml0nljK
KXzJdAKZGr8sB6V7HZ4j28R0O5acIPY9BMd/0bJymN+jWwlqGXUbwstXWC+jJmp/U48ZeqSJWTFg
yR1C99qXd7QRtSP2YMFssLX+8aQaD9i4eXCywCXleAy7gDHC6WOGuLlwSuvQ0hQK/4v5UoF1diND
0dpE/iOW7LYjLmkhsvGq/Pybs5tteQla+ziiVGLCU8iRd9WFJ0wUdKylVbjOx6zsQFLy3Om+kW56
pKvyGcQaHN11vBL+FwHAur8HZtYdTdp6BnXZ1lv17EhZCzmo6HKiGWSJwhiCpoPTsM64gdM8GmiF
QMMXUNffe5+si8AR3RvSDqN3udDAyz9P6TAjGDqfGrpJK75nUFBTfRYLR3cGTqfx7ud9Kf6s8GnU
tWGddpsAlDQEysAiFpk3s/Gcl27aHOsjnfxGjhDLjBZahJLv22Js6YDP3/nAvoE1U3Yo/PMiW1Wx
JlFuBGttLItrzY5aR/tcZ6O7zpgGds+gw61eu7O81A1XPanzF6JrEExbz28VkW9bBSvr/WyNHh89
5Bm0+E7E9xoklLGt2h/b1qDJ6vtubWAqh5taBXm8OJUKqwb0NGW96CgF9OvBn/e0LelMZaRbJf0c
uMHYlZUx9Dw35sqgr6b1keADhjNya2fVMJ/XnWpkrceFpDm9OtYwicMnSbC2k017yRi0G2QXHiC4
ccbprevQbqPKH9+NgFZLPl64ZWZteBoiucqwX2OzfkKdIipMbVplOCId6V+2MpeVhevjjR/U96Bm
9j1NRlob3+MlPOHFx4RohhGtVPXzxI1CYFmK/ZN8/MQ8lcyTmE5zm9Lr0l7GwNsNM0blB2ZfGMlm
PE010Q+y6fIxg6JFXQG1wT6JCt76AWOVFFDasqYcM7iAddp4Iz5CLUtoM4mmyDGNHjOLWMkWIQmy
jT5Cqhvhy3Xcpa0cSAQNc04ZlC7SeD50Hgdzbuux02EB393xHW7PBa7CBd6d2d+uYMcsqGayOXjv
sbvKKh1Q2adllNj9hqKUldzQ6X1z1IoLdSdsvx0EawZmPkJQGYAprWZxtMqNmoOkkbUATHE+uPpz
TmVpqqqSlrsyyoiCOBZ3/qyZ38b5d/j+U2IaUrOWRWxwd6XCtCsXNwryNcV8cKr9z4xEofAdJta9
Q1KRfTFDa1qvMI1q0cS0rlW0gPALTCj2ui3NwqYuY+SoinBtzjQObtSqqSwoitNaf1BXEAfoIinp
Fk2YdlK5R6fczZlU9/4ZNFdJboLe15KrNRMIGv8Ar9ek0UpGjd33rHrGbRLy9ctiX99lfGpDUWP7
g6EbvceUapTJZ9LCQ2oh/Yv0Wb2zg3BwehXzqj9OYqxRTZ/bYWByTleD9n+6gtcFDpmtcc3iPzvi
gwhBUghlt/KAU2BJJCHK+ijUXxlCP6fHPb/t19T6K2s0PLc5lDqqUZtH234IaAolsClAC7RxJMwC
lVO5cZ0W6Q6gePom4SE5H57ORx5iZ1BMfCNpXFJAIoBNwsd93VXw4QUfCuGnEd85SJxUV91Evz50
Yyc9AxJAbiE3NjKf08eRnbfOSZmMtNyjz87OFtb8XBYhFbkGyx+hEvmP2zN3EraDM+vtypC67Dng
/l6r/0CV/1OOfUn61h63bjwNUZHzK4OiEsqGNrJpbRi4I088VS4o/ADtowXSm9iV1DRCDNoc0yT1
MMsF850nBHjN5x0v4R4KQIaWLAt9KTBXedwhpiwQwh5nfA1xJg9tyZSiTXr+RR1s29ancTfaY84O
9hlc/ZqePTQNtsLFKO0F8dyYTPZkpbM5T3L4tvvyWU70wzHWx+l75IkpD+Bl6hWwhE7q5iuG6d1L
lFolylqfMioQmoYuE3nb2ActOqOLQVFMJbaCg5z7b5CcYq01W4s//GJnsvM4FLyX62gmSji+nfEt
CzIyMEuLjuF4+Fc/HVABH0XQglqkH/IttVuuPryFHaJTpgdPPX3jtPruRi2gIBIG2IwN7zBo4q2I
yTB4a49LFqCmZDfw9nelG8AebsnH2obVPIWv5eB4/jDE60+Z6whbS0nUGHKKVGyCouKAu0Vkcg9i
FuzadXKG4Ja92dl3kCk8cyeukMKKiIze+z3theMdKi6aPsi01WPRMDCRJBKrb8MmLJpopT86PuvD
gSfOLmokixLna8+tP5JVjWmpiVBAAzioLbGsPRIL5wrvEhAk4kWdgXEMdbIMJc+iifkg7oCqJBPV
7JdazZrsPlK9Y5IfYYmSkDXZcfXH4Kc3KHdz+erc5K3NYg72ju9RLoWQDUtsd/9hACoMWlF8BYPb
rJQB4QwUSHXSj4fMDESYB0tczvti/DMKzO61bZUtRUAc23bcerdrMFhNyELLj+gbF8PjUs73k4pY
7+g/e8Z4kMW+02Uma9OtTpUnm3eC8EIuYsbcjnFCgdW/kSc3ZBvMZe9Cr8UBBA55BMxW/Mn0zEQP
XDtD5ysQKtKxfQpd6JuSVMQKzxV1B9P/0wj5k/amh29JSu3oXPxcFrMLfgLxAg9SMc9kS+sRfke2
0Bd5hvBKlI7KC+MXXeU/FRNhqMw6PZjzLBpo34foERoqFTNXrDoW9j6vvceFF44GAjO4wl1JqcKs
D84H4ivBRGeZuDzpcMMyPWHnqYYIpFDmXIfpsqebJj8eksuihyAFMAWqcY8Y3f3H/vbJ2wBSNDFx
k+IAMNHch0pS10VjrdtsQDNJ1sjRK6yqGjhkdTBG4cZqtfRnLLzxGSZG4s7qTFCFSDpYtrV9uOs8
nKrnLK/W3SW3gsR66YxeIqOnsnyc3KQRFmASs8Qtw7o7mpL2yijlYpVaxN3mB2o25Y+Dv065HhHH
ccP74K+bslmeUktfW7/g62p2Qoh8sqkgdz8sUUhT1S4kGsVnwKvFttBcOPodz1qvsaa0LFPzuTN4
TNSc/YPdEvdi3zV7BfZofytWv4piho8VcZimFJ8kHT+9X/Cu27P8y+Ei+ji2Odfa6lTuVWPNeQ+N
U+SBv5rvz9CrNriXXYHXzhHOl0k7LKPH6oSBaqkErqUdG4xfRohUtxPhWLNvR0QI2tRQMGqsGQOI
f9ioRUjnUiwc2WeLqYNXWHK4qFNHODWlENUrw7yvdThedJi2+AjXXVHlANcWCPoO6htzwHcly7RH
GLVhsok/i9k+yFI0ejo8seVd5jk5jnPF7w0UsT8SE7oBmBS9tvPn6aSvMOuDXGx9JJJ/yK+Ute7X
x0YRUjbGrrjWlpZum4pn4AC7opRQ8TqzFLNPZ10w44g93YqN5VkAKUr6rrja3FFa3T6pECTizkV/
hI8J98CXwLkwDOUSojWj0CRvdcSpmCAv+R+cox2Qnc7mzSMdZOExif9f86IoqXoNF4lI0H3Eofas
KHD8mplvurIPomKNJN/M7TftxMT+aEVLAEj0B91TtQ/Bqf/Rp09I08bNEv5pXovpSQ2DkY8EEyU9
9W99Ps+D7CtjNu7Ko2dWftoIZ9Jf8+ZitBNvVY3WUseBEVwF/cAasgJj6xXObocC8pJldnmWS11Y
SwlKhtHX0jdJ1eHbv409fq+q7S6BZJ81NbGq3/1aKRyWa5504B7x9QMWlmZMYrOSxDBnj3+aGP4o
a4AEY5eSVSqFCBfdyIIl6Fp4z6R+4X+OEoqcCUeL3vhIYcjVcZAHv+9q5382wb88d6khKzIIbrEN
o6xjVSuhLZRrJHWkBPf/p6kBozGj6asibXdBE7xVsnKmpwmgE3JVTNyXhQDceRsFOjpa06dh/Uem
8UFz5bhirWh5MWhCE5bHPhllD/wd7oLKOl+Y1hxEDNz7Ks58rNA8xyGqoZLhdVMJpkv6li2fuo+S
pO5AdmC3IzIyRgYuGXvYGe4pDTCYdSrW9YWlDJH+JQ0Lp3AeraUESnpkQak1BwxU7reJ5xicd1Ll
RnhpvOEe6xOnXMJo4YqfXH/di7yKk4kOfK3X1U0SwF5B9DyE1YvzK24Ve0Z7DumH0/mXazptn6wp
jgR/KCHEOaOyGMGOE8sNOAwFt3vdaTE0j5mui/S03dMR19XF7mbFa0cpxRfid210GRIXbCHPJsyv
MHuZPdvPIvurZ9grDE6Ui4QIWOwYm5rYoYQBanTo6EnfZ18NWFxx7CKgXgqMY/cuvOPNBfses02u
pWan7z/4uIK6azrtYkFa2xCGnANwaO4eMUmvVpGa7hLvq/Nuq+DBkgzKyy2bYYkiuChC0rOBIcxQ
jk454Au57lZVr8Bvfr6yW8yODt4XRp8THHQ8fwWBY0W9MbVEfltvoKVyrnXSl4Ixw/KRu+kkPj33
F5oDr1cWMr4ueF27GImFD5No4habbsscG0Wl9CHsr9aaog8Dt1rhB0TJ0MoA/JmFC1gWklPRcJ5e
IrdEqOkpLZ/njhhx
`protect end_protected
