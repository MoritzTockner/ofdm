-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yH7W5gMet7fcnuJ7WhO7Vmpw+kJ3hrT30mVMRZR2atZfWR8Gc0rvz/aK5x/9neHu0N/HyQK/aQj1
PMQDWU8PEhH6NTgwtaIZajJVovsE0rlaa5/ZiIzRSku+LOV/IIkZZWDiXh0Pd73ntoAmDNtU+xm3
YTeM5XDJB+wsjQWTiw45SGkr51D7+0kqvj8hPscuuAxatdi1XslzpFflyVrdy47oRlxl3MXHZz2F
Eb7bu62KLoRPzDq/gH3SetWmPzy9WoSbfXkAMortFcK78hPCzhpJSiQ/cU5TXaTdh/3Yr48qEOwI
GLawZWA9WV5pLezebyxc29D8OHHfpAyw+dXsfQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114272)
`protect data_block
x/+aRNtI2ZRUXUdj98bmqPOn6SglWLB2MNThen4HvpoFTqQApiuiMUe8OaZGBlQUwP0ybVTAHzOU
cK1vq5ETIj35g1XG8MistLCJn/Np0J9tdWa6rYbn2PXkaMH44Ba9/djvTYPwktRfSgY4PaP235Pj
aXFwSTSY24oTGu0+nJsZ5+24ZHVmghH1Filr39Qgio4JHSV8tG9ka9ytEV5lBccCZv66T0u+I8Mf
tA4iFygKhbpk0w3ky3t0TOeS7FpappMnab7goWslQusVPc0z2I/oH67hULXHE5HMAKr3FUSs7y5t
r2hBVcR0BDrJAFtpxSqVZZE5oLYonAgySJEBge5KmMyakyL7rlTvBjKuwj2RqWrpQfZ7mM6ZdWSK
nbB6W2R535feyTXY/omyH0NcTRxs+GD6iPCyf3X7B33KyUlqm4MKEoxl3PLDnbmKUYkvM5Gn6td7
JhEgP81z4k0xYL8S4j7dPxuKERmJrLYAK5zUz2OTqYYfeQI3Tzpy6EM+i69hoHsZwiESgE0HPTMI
8YjrMXi+a+GTuIg6hik1XBYOmRYqFcdBr4OJlmn70TChsqgDXhpEF3G/LaeKTf3orveYA4QxHBRu
aa2AUy/lcRZaXvC3nMVIE6ZsXTAXCERpdu5KW0u2U6Nmdo6pnmrbUUqcP44xkU9onqozwMPlo496
4QYHOB/dKKyYDrSRkhZoZguXybEtahJB06QkZNe44AGCrU2seILbYil2hUQLJawU0Q0emVmE4w7B
xx1NKkeK+FUNV8oPxtNuZRM7skYtvnHS7BBmDz6ojOGO3Ai23/GSeeQzOCqIblyTBs3tB4lPkjiY
GG3Ou+ygYuKcDQU7CAimXHDcOW2z4c5czZWsBq86Qh+x5UAtweWgFhE4YL5fxbFS/pE0KXyo0Pqw
5V5BNicArBKUNW6Jwt9AfVjawXgDvgom0xgxV54ZIkz6FoxaAxRFH6+tV7KCx8LZK5QnS3fkDsrm
1Y6mmnZucmKFNnJS2c1CWgbOz4MKfFrt36t0QcV5U9ImhpH2ZWnHBXKHQNfJos4/grP09a8nZ3HZ
lmU0FM3/8X5S37EO9yn5j5sMir7OZVIjdtojADJUQ32V6W5krw+qdMOHcQr8CtIKM/Qccros2+07
ZC1fP4k27N7ZttsXesxShwzCRsoW6dBpfM+lZ5t48D17uIiO0TGvxLAPzL2trZodL9xbi7xx/W9o
9oYLbnNfIcVvGO3HE4GX3HM4pqTHiCP0NmKem+JGNf0qCy7O6ros/pRF7Kisx7iP5ke/WmKBdLOd
ID+QBql6X113F6sUECog9n9Az44iSIGbzUylMfe3LpfbTzFXQwXA2fZtgu9Aq+V2rfhWev00kHgX
h3k72M3+3/B4TD/CgKOXc/0reySJ+obuBndG6Yxf4jo5ooxZ6pFM4yMAj3KMWeeGMgpmldOsh7iW
Dn6wDRae6e5bDbOIhL4lVMohxR8sdbR8ZyUFhsk+bpuWQZiPVivR+T9QhJfnldVI+ozxaMf7g+eH
fzoZhFlqNHgUpZqX2Ml/6/iWFdV/+kgapwFsbqYx7O8mAy8nSePByPVHEOHfS/nalMXug+qMObBq
2dbKisQeCWGx1rij+Di6psKBFLW5HHBdZaKUbCtERJUVKz5QcB0jvWgQC0ZjG0YV+vlnmC40V5U9
AFYVRlQK7nbZPONOofoZK+vdK+cvGvvjQG7L7kmbC5EGjSZg31pOGQA5CoGzyifeWOFHtlXyVMWk
UVzsN40YMFAlTKMux37000A/oY6HIZArjX7ZV6kP0E54KU3bX+Kp0obTJFzwzqUAC70IuygirG+i
5A4d0qw+t27S5A43uiEbcdT8tXWiPpAEVwV7DutVX8C+bZX7YzrpSSyGvXaW6n2roh+0py7NCbjS
W4mPlva5Q/xML7tKnMOwhadMA2jhpgd7EjLj9oior54BvcmEZthSv1x34U0bPV0GWTrXwi4Sp1sW
l/nEftfTgnSd4aVz27Tgl5iIVkHHs7kRAcnZ9A75ixW30Gl9urlnZg+O8auDmIm+mdcxgCmfmGR7
7TmFQ628SXvNnkq+JBJ2OGw3goUwOA/gF8bna0d0RIFN0Qv/gCEkUgd4P35QAuqWTKYpsnmW9c4j
ngPr+pACQAMuV6ZzhxvaHjUhU9q4cYhZn7ceocOumEjugDNNHpwTX2QJlWCZrSaBV2G8UD+HuFrn
bdZ1naD5kF4e71q4gbETc2ngKO6L7bQx8Skdqz6DADPs1NChFXvgg4IVy76bSZ7r++KXEP6Lsp2Q
mxYl48ppj7VXmuVQSItxA8SkskXD2f1EcJWkpLPwYvwj7+HOXKnr38XiNsY45vPPJN8rD1lj3uCg
Cbe25BMb/lfeYpZKQLMZ9B0oQFEsfTCFTgznA7csw2aoha5168cKo9eM3FW6MFEAlRRsMONtVouy
o4pN6HBFFbPR0UJgkgP7qRr+uKU/2iel9eOlu/Gswu7BElWnI2vjOchNpWo3soBfTNUMlGgfpuny
Um7DaApRRo1jcati2sJN8sq6nP/O5rtjjKhJaXFQGbnS8XD1Jm2qp4n+Idxre8oviLeId5sv+nCS
2oZ0cLngXkCYK8c4a8l3Egd8E8zi5wRYvaGFCex6Co1Z3rwO4FxmSrJXLRVn0uD/dKYIMTa21b7b
JjPgVnqi6nyeBob62Bfk1qSPFeLZOGD44XL2LdFbl5/4lQLu7X2VtRsomCeYYBJzZTzOB/oZFmQH
XUemQlss1ZYfKXWgA7ClEviXChIvUA5isyr7TsQB3d98Y7A3RN0EE6SXx+V891RU0xfF4shC2XCE
2h2+se7Fl2gyIw0suklS94d7rtDrTNWiLtRCHmlcZYLeuYnVXUulR5HxLpLD6Ixh8BIHnxB5Dltr
FdsuX0l4Cy3kW8SEbn0xnW0uctf9z76qKwpDdTAaBTOT5v+a5K0pDf+c3Cbd7IMK6t7yig4bLsun
h666IoSwqHRnd+CjalikQDHRGtiq25u5mbzJp0hvrzmXv5VLeNJDUrdIhUR2J7Pn/NGgDru4zRJ7
6SkzfTLeIbgNy98oe2Vk2s3QWhVpSIvFt4AZVUrsd66Faz+uVZXiIzWb8afZq55J7v7Yqva47bLv
niHHJE89hVUhhm1QUhfQPhNUE/usHed2IjcEtX7FQ1R6LE1CMzdvjEZe/ceFLaPlwEhYkDEDBlME
7UfZQzn3SzZooMhK+D5iufTR59otN+wI0Ss9xy4qtkMg20aMnKWW9cSM50M2Srbgk9nZgIgwKQjM
YaaFyLS/LQVerw5Poa/irvBHOtEQ0SWfwlEBPyO6K+DSTaBl6ft+Fr51sc5R0/9g9xm+WgdVDpm1
WqEFJJmpXIP2lx15Rfx6xfI1bUdj+PbgMuc6CD/iSZ4CZSvMPq9/GrM82O4qgBBBkua4ieGz8eX/
cwM6Sbga5nbsW/gtU8ItM9mB0F+R696Rq3BBVbjJK7j5ZAgVw4T+G26z9ymMZc2ehwXawrAJU2Gm
WaFZkirab5xnP0JInDUYFitOZZBJKisGpmu3qqthztlT/LTcy5nsNXEeTefjaKA4khxVVvJykjoA
+JfrtilbMc0C32WFXYHQy3d+SxRBmKETOdddAydvpdo/Gxb4MWG9z47oRKWPnbfcud/5aLnHkE0A
ljuH0fhClVO0pO3FyKL8sX3ijKpH/kyNCnQY2G2MUe2kPawmSjyrBQ9AmOtfCZT8aLFHhba9aRag
KPr/SjDdhcT+LH83uyA8cS+jHRV5JXcpYVac99Kbitp9PGFL4gT1SBn8AQyHhHTjacMR1XIufMrm
2lGvFiBNzwgmdOrobkCcjMOwz+xIksE1AhzENdrSi7OP0oyqPfOvlqm+zpUGZ2H/Ah4MyHsdNGD3
upK6qYrdp2bo8YGEixwWpjCFJ/p5LY6Kx1DBu2hqEidgN6x8kYoicJZyNjajKG8b01E6xLV2+HkN
R1oJBhZKZIBV+DNeLth4zviN0qsYtIdPbbUa/BdSj2YLXWpUmRCaYxHAMNvIu4tbckL3YDuCXju4
eabID0epSmEs8e7RDckP6QYzVbjcNhIVkRN4k9bFK7jWUyMiuZDiLaTYOockIOPoIckJg1FCUHZy
6eu1RmyUXcB/KN+IqDGKfI0Tq8a84P4YPO68FjBpW3yWB3jHb41fm+fuG6grbzOCmmQqCSbI+2eB
k/pu34g8jtfDBOchX+CBtp/VeUiYVwq755rQ//ylOnxSXHJPqh06Dk6BQmHLCdFSLFWqPCzhwqx4
GAaBe1i0JW1tgc0bqp/7pDHMnnVhKcPsy8Ag2lTA8dgaIMAp0efSkzeNOVnuoETm1pv53Ri48IuD
4i39vC5ROY2ny8scIZ8gSotwAVEvV4XrM1RIQlRI6eiabSE5ht2Krq8wLSJKbR5eSH09nACSNHR9
gfuByRFQC7f2GuyrXY4G/I+dUw5ryDLxv6UEj5rNc+Otk7FpgQkZgROVon31mjqwKCtrLmSm1M8p
l/6PD53FIZqePawQPIphSbodD6dvf3TRTsAPiqwkU5ObXb3YXlm46Z1GAP8VbRPLnYWbg2FpsvmE
ngOiB2R5vXYomt+KgjHeKUG0MPc7LDwBgtHv6JD2iFir1J3SVsSNyuqP8EvZ+yNuybFSvb9TaRQn
qvPBXjPtX4qzgPC3u9z8gL9q/EnTNe5U80MXE4ZDXdV3b6MYWRGV0dSg0mpBGEl5YwXvA6tWd/wZ
v+VMtkr9eLZW4NCb0GYqud1ZbP5SwXz1zgzKHMLx5bIO8pkM2qSoQYsCnK6OlUlKzUtFppxsEO4d
eHx1sqOScmAKA/7ao1En2OFXY7gVEOGUWYAoFJ/lEi/TlUAukgm/LTXEvhe8rJDCrCC8RRiSqrVd
CHwFgEtpvnyI6AscxDx8OtbiNBpBMsFHnoasFZDyHW3uj22OEZmfhRy33xWPtPF+sCay8MI086iT
pWlmke+tiAsdVEah+rAtXqYGo0H/p7wU4AOgjnqnEm93IJY5JudMu//c1FPevQewhSsTHQUMw2DY
ORRdJGd2nfpVxALB5Q3GPvT/4x6ZgXdrY/AptMr7CUzb1nX45cYVQqBIvRGz7rpMJKQSb0vQxcp5
sTm5RTc40s8tI3p6H/wShzc1dNloWjfq6yi69vXN6YFY9l2nQ9CihMo/0D05y+N7TVUwlrBFk0Lc
xbFzw1ihAQw2hCwbJbHX36TrIYggwnkuuEfYWiLcnNCwMeTLYga9Pw8d38BqOr1O8SP4bKLV5LAD
lqHp1FSH4XGIkL0SRdPPtHbyFO6BMKWR9f8tiFKgnyMtxaAVNhIDpJ4lrcZT/7MYhCwWmlqSH/tI
E3EdAd2XYJtHIhSoV1MyBuB0lPXLzHpa/73zbQaxeMzkhNYj25TKWGFpWRi0E7XMNcAoKNtxYJQi
1doC66BvPZN/obekX0dFJnFkX6QBKeq/B8TxntCQe2nzHKo8q1PdDzePAjxZdPtA4r8srJYHMzzZ
gIKuS62dzsDJU3BgjAElxy/E2vz2zAEERCF0/UunBh2L82NFu26lZDq43g+kmVhiNw059c+SdjOK
s6MG4/wO2N2YuINkEMkho4KDOnd/pYnzr/eAhNeL9r/DiQv+ug4XPU5I2+VbzdS8mUP4mLinwNWn
Hb4uD+H1HSzrpfWO9vFcLG0sWe8fYRrx82YNGccOx3UDxTjycxW1/n/uRezDVyg44fXHYRg0Tu9+
Rm3hAoKYyLA8nW5spsci6hds9r54z1D+X2jP2k6ML+w1DuOGiwWOWeF1gU1SSQwKWhJGV2upep+r
Op5GvWR54F5y5D3D7DESnAjc/CUsnyQmYb4B+sNrix8MRzI5oSb8A8qokaks4SAX/xiYe+bezb15
wMmzpx9WnOr8567JL8TmHDOmvpiH8CPUVZuehTVYkaQuR8H3Lt5i3sGe4gDGtjh/JNIrOy8s3lOg
HNnMiBlBycilekl1X+boR0qc4UHl+8DZLdrIE5kpnqCZkf3neHRu6Y1hthU9R7Lsr8gVhJnkfp1a
Pz42Z2TS5Y976tKiCfEjXnjvZtAvJFBZsEgoCfxqHyoPLyz5wx+qUgC9muTT0MYSZPEKn7sBltGU
qWEblCkbccuMIbT23e8oOhqDhaxf7VIVfmiQ/LEOGlIhjjXC357j30EczY35WsG5nitVKnls54U6
rpLsfOk4vxcSoOkx1i7BemAYyEi8mXvKontrpWYSWWrpg+afDEDywpo7nZDlbA5yWGj3ENeCp/mO
a2cXmO5JcU+TLAyAzHNiiM4IanfMtgd4Z2VR0Gvqd3T77WGvcfk+/GR0shuSyTeKHNM6X+DcnFgv
J1c+jTFGM404rv6xdUCCPnoSIZQb1bXzdzhAgm3mSjrNz0MXUFkrJcwu27XIdJGw0syO6xelT3Yc
pZP45K3Gnf9balUti012Dsv1wbD8VGVWrCmsWWLGU6R+SFf8VQYjYlBs5u+nElP23BhTz9/w/lcc
camp+IfRT9A0SJlgiFmuU5jKon8scu8YWFq6K/ZF7UnolSkHDI3ukdYzScxtrKs9IoTq+9aswhQF
I23gQ0018+Kr/GtH3jJQeOa9zJl0KlRXLDGOLVeiUJOvbF4bZedZcqJpun3Dqi4TwnHEFDMejzBg
okBy5p82d6iUW+ptE7qTpJ+NOPDL1d2+7Lgj6yWcKUL2b+ay+PFH1qq2Y3Rrm5WtMIMk4WuUYs7o
F3l1ted0jt7UYWTdk7YyjesU5yNQtM7CuWM45iKbi9l+F4t5VYMwCs7K6ZojMU9LP0oJAKYMDFA4
0GIhXbN0KPlPmOl+cGRvHjrk7HyHhwV8QQag735gqlZQoZ0uYo9pIx1RHDq7KDH/G1El4TcrA9PW
rgcEQOSKbxaeps0bI2Nh8dHsZ+CaAl0cB/yh595cSP47xgHsiHSFVBmAtdR2rr33Yf3Af1cNJqVH
UHdURwvydlgDxwWUeFHi6mq1nDTOkIKunYeOtiR3BWNvNDbhLkPqDV3mmdQZ2dOqEpMSoRGh4K4Y
Xz3j5KtwOYeF4vu1JN0j3W0P81PWVQtRG7EHugpD9WF0HyyJbmji4fQq3/YrtPWVn42WqwHwhcaq
Wb3TweXUuB+SNQ+3SdnOe0ubPMoKEaw5J/DB4wyg56tKj+mWHyr9KT0WJm9e6GK4CnXLZm99Nnu8
MSq7G56mzikitsmwBejAsgMZSGB5mzg6eQDr9gzqCqdv8DmVAUAteO6NIOOGqLioD4hiWMK9EoYW
F82Xj2K2svo+fObDSEnxHppg5noTFo2S2MssG01Crh5z0g4+7vigATShO0YAmLR7YPq0qSXgli5N
HtHZtD/g+fFB4VBe3a2DRAcPLKfVpnAgLhPQPBYiZr7x1+X5gK+xFWuzsiCtoPp6ecfpxo6Qoh4b
mZLAN4SnC2gsAFoKQF/0hktw2qLX77OztBZwekggdgKJxPugngw+WlMAH8PVrOt+lIoCxof+j4Mm
QDkt5eQZue5e/Jk+qOJO46PBRIVFcPLgvI90DKcxsjOPOErP3Ln1KrmOpfHseLXaq62BfEEcTJdu
uxzna5AcrUi9LlWGXhLcm6VRtuXiUNkDxLC94DoaBFVo/9KGxlJ+qMn22VpQscqPEyyWnsTpCIb0
aGP6W+fAd58yIym8SydU1y+CTfSXe/15mRPEHzRdLjEfTABqqjqEUJl2FTxg8DKnar58jGsnn29t
q5hKcdbcLVffZ9Vg9Q6QFnS5SluDU5U+dupXYj4/TtvZhIfWeVvTj8Q0kCZzyhWIl4es7CpBx2Da
3aJEeYcLKwhhGNFSuGlBu9/Zd9sJup/toEMlT05MhZ/1Egey2gNjjW++383h4SPdvVheigq+cw2h
Do9buA09hPKEf4bNFk3LNsOvutIDt0/33i/wI3KAehw2NefZTiKY3PMZNMzqWlUWKPsmdxqotTRl
mKFMogJWuZRvtYu23B3Fg+jQ8X1hdK+Mk6wJKLXI8Nqw/DzehR/0cBrYLsdCpQUBcrikRgCWyhK7
y0h8o1nKW8YarL1cUaXfvR1C/09Y9s0R3NYUb7aPA9M4TNI1Y3JajQZYOUu+9QhSOKGSHtuBDA3F
HJAx1EUIzaqEFC6AGCk08PiYaLRMSc3UnmbnieovlAKdilYTXckYS/3W9ncAPsd16FzlbOzEghf1
djCIl3DMNQbNzc3TqQDtdZ3NiFZHN61CR7KF2SEcJ1cG9/u/rp4dfdSkUX3U/0Y66Lbs/M8YodXu
JumXffLsXm2QSyfThMAxj9/iF1Z6/s8tXVa8ZfWOm00hBYGELZqjflonLBBgI1R5xJIPEiZEHmGw
e/wkYA7IoUWMiDd7bWDQllXcSc7ihxkvsR2wMwbzlljyOftq140vx7l9SludjRM5Z7zv4AHPh6pL
hEqvmsSyrRSv4MqkjQ/K40n7gyts37KZTMNPxGH1BkeTlJM4IjlOU6GaLTfDkihcwq/S1VgtH0ad
gfbgN/p0Ygo/y5IUF4R1rsabPXiQXzUMynR+tAYo1MPd8cZXHQG7IVa8DYDrxbC+kQM3oko+pR3c
dhL8vkuup+V5BSc2wQ5Z80O6KBd2S23hcG542lgaTh4dUTmoxgNGb8uxQn0k2VFsfl9/rwA9Kfva
8R9BUkYIx3DDyZmJDOC9sVDieYCVNOFv1GuaDcFSmA/lYrqqfDXZSO0J/azuRvvqRAV8ml23nvTq
tn1bVJG1EMjef9BvoMJvsGxuU4ag7vOSf2LRy8XbGCYwc/M3gQsowX8CTKcx7qM9sEeglHpzZHpm
dEmmYRkZ8dCTps7t8qVankLb/+p7ShL/WqjFOIntJEXsQZ7xcVHRA7geI5d4VyQNUIuNIi4jv5Q+
HRlD5hmaaE+G7pEaKV9GrqeXOagnvEdMkZcPczvNCh/fHLvvIoOIOwCv67vHnRSlVEffZtjk4LQ+
fv0ebawzJOWEAAiv0L8aCg6epWV+gyIItZNzvN0fNFx2s4jojJd0T4g8ZO4d79bSXtnwbjPmr3kI
vp/6i5ZBY4YUrWLNtugKEdl8AQ9LIoRJz/PP4IwZEC2D+yfCXyAa/pPsuqFAL/XcoRcRw5QToX9L
EoOTxiU7KEQ5wWPVDQB5kMth5wdJh2knJWZK9F57gEc0GNftPuD2nhajlsnY3Z4ZgxFGRWROm2pF
eRjdREowpMeTudHCeB5t1/9pPF+LIGcrQLGm2+NHFO0bqXCmZVYVO826SQEJBzpvG4gK9hbaAC6g
y/m1k6z/33Ivl2We3BL43aiTOhMm1cGKuejteEZClUGx/W8LuNrHOJZVdY8wLLuxzJV1gPe/SuDK
X+sfNJLeLdmD+x8JUuDbZzWG/ujz0FoJafFy8t13us6SYAgzHxXtoP9lLryuHGCrqmMwELO0JTWt
cpJpjAygOt2HstuGE6L6wkCQw3U3k2AkFKIiVxhPGPA8MBq/Ff0xWRvXhUWIoYeR/uA28iBA5xYx
aziXkZTEuNLyGuMGCNWz75os6DVlf7zclneWATUcA+iisQWiuZuEVQ7gMzY0yqu7AEcIvBB2UL8x
WHeYOPlGN6A/pfQF0bALt6CQsu4Fdux41RsTznGTOeZseVtD6aCOGHajYXcd9QZKIgmZ7QfxXwGo
Cc/pBQsVumTtC2scemUkul1NMfmSXQRJzHndMUlkukFHE/NqTbqWKKILIcHy4T6LA4jY0sWlojjn
WNmEyJggDT3hVjiouJeJB1aH+MpRWCcy/WIrWf9k0tdX7Dm4oiPluEYDB5hsDWR7OKSAh45Ij0U2
mX5gZu6CCfEawX+25DMfdvlFPYJ7ZTlwwhJ8jMLQTPoGIUgPugEB3rEBVEVSZmcl+0K6rqbuI9Af
MVUZJeAO41obYgQHeXyLRATwSZEAtteiBU+lpW2BGwmXMtigpXX3/rISB5BGoRV+/hB+IROG+XUZ
nSebYL3kSHz4w99v9jRfGyxXjoRIFu0qaWOj8wdD+WBz/u2Ve2cWIZfIY/Fen3Wa+fXKykX8wDJo
+WIHVQzyNBF0+khWJMcCH2LNmyyCY1V/ULwIssJAwbD3JHFWAPc29+CjoKakuPmb0TSevwjPQ/R9
kfN33AWkFogga60DOopG1YOG5t2R2DfyGDfA++lHTEdQK3sR0GiZq9SAzdxc6aYhDTPXUk0u03OT
NlnZ4EK2IUq/dLnirhhw1o/0i4wvVmyc8ZL0IlUifOUhp8wNq+bBoftkvRsnvyUh4LHf1Mi5MQEz
NDa+Y1VmHC/7YHpS9jEr4j3YtWyBN0Lb+sSPeAIG29gLvCNe3Ij9vFe6okBkWhsDy9hSD72Hu5s5
Cu8wl4AScmZfAPkLlr7kRzKyCfBLSXswmKXbrLiEaCU5hReWjWSBe+/LB7cjloaOYrjXxQ0fD6Jw
fhbk0GeRi0jVtl91TGnsiejkD9Srn3W3f3qnTCePxST2+gmTmzbfq1nQoVqEwCjzVcEuCH7huIfb
+ovav1Yo277KM05QKZXCrUeTRB0jEaf+091TqjHAW8fBl1LCfaW1+FOG7gPDxD8g1n5c/2B+5Ld9
ZNUSG8t0V4Gy14aEB4GKwCFkkQFMn1pvNUPtbclxU1Ha4rz4MGrgqBVaiXPCfSQ7PjkWueDGyhDj
Bbt1LDdzLlne3KJtw+aKmikChINac/sOVQ1Cq8aaHSB4VCxhYabhV4uEpHfM/C1jhwclBcxj6rKI
09HJTv+KBuhBAtLm2c2jOxHu3za9q/JlnQ8OxSAaBLoFKbGDTCSBgjUTCQTF3RkXT2MwtilhA/jb
HOsaDljvceG94JSG7s9Wjffg9jW1Hh6FSRGg045954bKYvP6+0V6DXo6HuYbAnNEeuywwJgKVTNq
pkJrQIigCaQhh/C7olcKxbOcTAma7RqY0meTM9XcWXpRG+6NMa9gVdQW8gs9HKs+RWe/BMILQgjx
BwZ4oEM58Fo7vaVR43t/3R9HF5oBXWDfZx/nyyPfdwhzlj2k4Tc3XHTAGQh6qzu1mMXeLrGOF1Dz
3c6TPZImkhjoy/xhbrmIabSRKzVQ7WrXMkRrhAtMn4FxSNTVD/Oac6qHLzSetJ1ziwyHAaaI9BHQ
703E3rY+hMXPKdwTrdpPPDc9r+YDPG/tb5FCAYWpgJEba6D+1uHjRkSkmzrQI31TLKNi1DGX/XOm
6cHH/B7jw334k8HP/azAdAEJmpWbgnkYskF7TTpw9YrCTJqvaqVq01A4xejxpSkeutBYXhcjBx8z
3BsYeHlpxpKLViIn8hwMtwt1c+yS4pCv5T/Bc10iMET0OHOkSNneUXhKt1FsDjdaYDHL5rzPOVNc
gnlYukJq5hSpd3UCdo9hJMzHPcak3Dnskt1y+bbngdeBFyjyaCGw8NN+RvY/sJBW4SeiIGS/Ddzh
fxzoGRz33luBFdOAnhs4fZrd7ZobHCevK4U1F8M7zTCaW9GweYTC3gStI4V20GNlub7Er+Or7gMw
VTR3NAB8kN+wtUrVLoay2xYGlTd+3yz5gWOioi/GE2jFG1/bsiP3SFfPmsIZkBirCbzDpNKf0WH5
iq5A5kZ9lwz8Roa+vGeMxaeO6l+n5xdvxhF8lZnJFGpjwI39qatQx5wGd6HMHzhMiHPuvuV3EEZr
KWM5JdIAEXjdM6ze7Sv0Yq2MGbivwi7636ZzEfCZdCAvTR5MPc0gFfBsCaJbcNA2yg0rH85tkyT4
sWN0jDHQ07jQVLpIvkjaIf4kJvP0eHBzKdUaMxov6pVYoLZfAI7Xv4OAE4XacT5Y/mOWC0yKS/AU
d1JcPDZJQZpGwngEeUcp2lD0MoLcss/l3HCZuDbZcitWu1L30BRPO3k6c0J8pam7KiGzaQYPkvfN
sbzkQ8UEVtEM/pBiU3dFTkAhpSZu3u+iKK4ISuUJTZIKMt4rZ27EEOm9TBu2AkOjUozhJFnQLWf5
Hff3vLsZH+skGyOPCjKkLMek09z4OJRurDsHe8oiqt08eLG1H2H3YBmFvbDTyM0LVEhxovk1Tof+
+uweS1GqJk+6MbcNpwr1gX5k9ZSaAqZCQ5tp9YN07fxfapvJzVwx4HRd7vAn0RtuY5KyD7C7Tt4f
N7awDNW/Xpm2T4s5ajZ6UdgZxx5Yy11H1EAgb1OXgYiwmyxzwLxp5/hHOrO/y9pBgN/e7x29ACqu
hH/9f5ZUVw9mBerC/c6pQ5oYfDWKFo8LrDDiVD/f8ohYh2A6xnCgNvzAOyRihoxI3mQKRDZkpp3z
kI3CG38iOeOZKGM3iVltBVXsx8vp2cAWT0BibbgybCXcE9ZL20ibrzjBeVfsRA9g4FRL5NairXQr
qoKn1rCq3D6IIogdmpJUUdvdKLrrig+rScP086llWBAwQti90Y1DK8OWGVYpaxsisNs7ZxOnjqTv
q5H1vIWcIOTkvieTetXjw0+1114rcQf+//J0PjR/lJ9tvZdoDsSz/yvQjW+iIRBQB+UiNjZMnL1e
DI2fDZoqoDuu0XY/1yDLgOX/chF5j6s9aoVgON/IamGVXQ2XbNuvK4cBBmUh9FsSl6YqkRDOMSfY
ESVOoF1tjGDTiW0+HYyagNjBcmoBd6LDXERW7MCVLTD2zpOnlFiZ1pYNL1olH5edSizGs901ZVLf
aHbupIIG2+g9JcZ1/uNZFD7/7IqUDCo/PeQX+qNIw/rJvs0N6LKIf6o+x5RwSSe8sSFQ3j5JOmoL
PxE50TiDgPGO52joWpkw1OqKgV/VYSy8srUz7Usjo0ma+kgpEU8SNr2ESb1Pspbbsug39MVgTPSe
WZXeoT/7kv3msXktqcswaNvV8ctpiregqMN9cubQh1D/6PI/B4Wf2eqRoX2HmBTWOCWV2RdANByl
Gtago5fX+XjeTFleE0OMD7rNOZziWbBPLRy4oa0QNIJTA2m5bsg6nSKjd8nw0WUsDh4NACImY27W
bbuP1ADyZM3xsN2V+8tAA/CHRMOvlebmgfPJR6CORr4mQbnH4zU977ajXL1AnklycK4seZWUVjqN
rw6BEwPooDl+zYjFkki84JlL7/XcbvjawOx22zm96RedNnteJkeNXGWxnzBOK/rnbTwMwr9Zxsne
GPNi8I3xf+Wb2DOdmoMhykdTysTFy72Hdxx/wb1kfBwtxbc3YHyOSwJRVmltb4aC0im52OUtb8/r
FUVIBqEfetJJvRJXW/WX5cTlabmCJ9b+9N32S/LizvR5vsrbgGiovcByfySF1tqVeVPKfoBRA838
ZoC6B9GzwH/A5b0bb744kcYu90bKeBpii7ifso8xEEFlxqI4bFiqD1jyZMxdhDGaMR/vXzMdMD1M
MTZ/LY+S/UaHkx/UoncQJnN+oAbJrm7hoNgRRg+4VUSu3Rq7Uqr/OgwRXRlLX80iU1p9c9Iz2cCv
7PwsrOFLUnYTjrNxeHhUdXXLJ6RaNGxXwD8kl8GIytk7GoHyUi+vMrzj7fi7jSoDf0DSAL+lsivs
WbamlP5UACddCXLruW4hAXXm5eVFilKrsGNXmg5NgQWt4NhRwBOvUhlc6z1Xrs3Z6P2Te0wDTrzy
YVzTbt7/KuknXvgPMC6teuu32Xmk2t61K6uEm8+Aw2q64FYU3sEfOYFJWkBL7jbkDuljquvrqG/D
v9pCNGAqTwsoK3pdl3q8PV7FKmCysvo1udcQCqy5mL2ROy3gcuCaqThEQ4QaGfWZ/MVmBr+Za5uU
uf715kwQzU77GOkZ6hTpI1j9zcUz4oQ8PLk0cC4RC6uDmmFLhc649K5hTxo8DSFOAJcvqCh96Ef5
GG/YGRC+sb6P21Tj91Vmt/7xLQDK6tdwKc6SH7k94gDZ0o2nHEqCEqausnG/G8DGz6U6ynJmw6zX
VbKH7xD7Tf6iQ3qsLEnhIyv+pnqEpnoSUfsNyrc8nDioMkod2wV7pS8OEA/I/hF3OOYSdOr7/REl
jK6Nca3/vqEScwwmwbemJmPqCrQSPAuEGdd4fJC4B0c18MwgY4QPMmZD7Q6iT8JwcxStCjW1lsI2
TaRjbM91wGW1J08vO66wukcGdbpBi7fHgrX+dgTIYi6e0oTqwR75Kd4kwDo/4Cab/2zxU94r+e48
v0vezlilwFym2AUCIzSu+MVN5vxxVThKOrGFnkrenAXfKfj5YniZNKwqhGokh45YiWeODry+cHG2
CikR7A/PLGLudAbcrOEzW/xWBztKJjKCryyuI/NDHKNRfiSQOovYUaFuEWuHhYsKXZbdDJnM5CYJ
PElYwrJH7icoWzzlec/UoqGGuZZoc0Y9H5xlBAIdY6RfvjtpY23INaAHb7DKRI7tWJ7ijcg7lnWc
fIT+kHSsV/q2MNc46Q75E6X9hCTaBrybPuRw8tR/w9aNFlUS2n5dwbCT9rTZrnWgBqUep3p+MiER
+EfOWJBJ4W7jycV5GNUjw2Qx/jLjN5V1wnvYvzxDFi8U0qPv/siiRp5Vy7KFnaFtGKlL4uTW+6k6
+EacOH5kx4OI3xvtGPOhGYiKjSY8ronNWcFBRUuOjZ5s92tE+whka2YYfmd5+IYMycFmkjA/RnaJ
X1m7Zx8fajt/1ly+7pxqEgEUFIvi1HJgYvUWrerHBYndlSXhR+WxkRp+jor9IBcxnEsJc7jBW20P
Pz0Is+7cFZK8EcTt4a4c8I/VolT8i67mAaqWvZcTk2Yi/r6MYTVcsWSGbfcCMKBWeLXKyFbtsRsb
0rzNjILzklXZJdqYtZ2Z86tEK1CRJZhrQYrUUfrLykzPqFK/wBUJtNK+7b55Gs75izkS7DhsHrTp
hLzh2tdiLCwDUdYaXdHy7HFMUL/qA9sd7woPLbyFkQH8QQApzbLCEUg2ADQM8tNZKQqi8bYFIDbT
hVLOJ7niNbqVoB7+dTUzNbrEkt5veK6vtCdVY2K50G4RfpinUXpGs+ec3ICzzsUweMJaV2OmGcTb
gONuyp+foALCgjAmBZFXGOorM64ELEbHymQIDB0JlSfk+v4q6jtx0VMlAQypqncHNUGJFYb3cgBO
RjZINyO0OEy1IjI3klAFUkpeuU6RPErxFhiOpEXUq7TDwLsQQMTa6jBUT154qrHUJD2PQqwdvpbF
hbMZUyhS5ce+fcozhhmFe6XBUvvw94beVb031yhRRoFtGZesrZsZBjMEp5A7yj32VVlhve0r4FZL
qLlerWQjtUabFGdFXvJ2S2xp4Hj0WvHkqIeWOwlmqOaSuul87Kty3gwSQYr1gvB6UWWf7MyvnkpN
NJvHdIgS+yx/OHNs88f5+rZhD4UWSxpqUGfzAj6Q+DyAZ33D0psr2eO6eno2mgFOe7WZEKrzREzV
7B0XqFTzZlupw0wZwwa8QTuzQ1fXSQSTzBDxuO0GAH9T87k4KV6uk2r7bocLrHcocg+tX/4ycv7Q
w+Sk2xc/i6TFJka7vcxHTYpf0V0dRcoqHrjAI0qxC0u8RHEwZ5gaha+PRh1PKxK+ZWaXwtw0PVVT
JwgreuNVywbOVLp/CKs5mlTTk0DX7A8auYyUnTPR8kjoZuFiIegA4x2JESPb/z+EAmoykRKduNDK
h2+WCdnj22v4a3fkAAAT6NBNeXR3xV0sR/uojorIOyPNV0Kw5Q/05T0R5GFW2R3ZgVR8cqQqGq8r
62BOE9NbNZD54YQHoOrNl36AJxQSBVKXgSvc1fk71ZcO0Q/o4LScpnWfhlmX975pVO+grNS/e2k2
3bWSwPebPyshvz4CVbXlbwn6C8PQYPTifm+mr8qvqMuJ5Sk1Kp+u1egomM3knQ+KsMimM1TWDuTC
RlLs308Sm/xZwhLlh0AjBhYPEwQW8HCvgC7hLcZJP76ZSR+srIelGe6/FIS/Ih99TU2GiLm8iQvv
aMeHnHWrbJmULNSwErRoOIr5ah/pHj5cyzTu4pjoxJ13366oIiU72NU9+CgyEGNdpUOzKI2h4qJ4
kA5iML/mvTThWtebdaHcU6O/wImlH2/KrR/TWr1VhwdxN5WWBhTDFd8svtOXTgLon4aYptYkM0pS
Thg8POoULNnGxN+xoBNS6yGesCiO80ctxwcSnsr/duQAijODZHl8JjtCU4KO6YaQJwOt5zw7mY7R
se7dGKVhue4fxEu8tmYpB+RGo7bAOnDHGFDCepUCpPTdgVZ4gENMCd0P7wUjPcd2ySyMQMeLtsQ+
ulELc5h3WHhisjHzrmUZgLqAlTwhEwj+qx6pJRvqNsZv5d0x/EhQvMCyi0cYKC6X3Rvv0ybk91jH
s47WidOwNq17E4lftiSpOsnzRLtT8ApThbSJhuWcJwoYBjv1QL9XM2EktBdUTYm8LmCL4FL3m6LZ
w6zR9SRZn2fr6ibsz/Dgx4urIsaMRKyh2zJrT+Mipuklim0W4Rq1h/mfCoI5S9emAHewIrZxMFdl
dqCg2VnQ5l8pqzhh2ypQLBg5zts0ySvsSzlFHj8oAm6OLbt3JlMQ+AesZj80nFk8uT+6re5yBFt4
Gz6lCnILzwdzIfEwlzv8rxe2w209ZV1WZQ71cVcZzWU7Y4TnSSLKIGIlrQ7EJNb83jv0+IPSlxOA
N8xq9Z0gBW60o4RyYe1yXPtiQsCZUQ0lYHIwBKuAqL222pBrakE+gvXlY0qGuN+MPYtMZ3mxjBcJ
EBTyhauojUHZyrufKcMYeR3vtm7DO69VkgffjtoW5awcqIx629Y8lBI4oy2HQ8CqKw1fW1P66uMW
OTNV+BnoplYgM9eaxrA1tPcI0w3QTX38mOL+XK8+NvlncRGiz2i02uVh7Q5O7IyCrxLjNo5JvauY
ic1zoS9/+vg7vlTDXq7xIPP2zvO++sr+FNaFO9lACpODjOaWHk+rlSlT3Nq6KorNlWiSCTZcWNfH
986YwcpoG4RXf1gcf3ALFeskIdR6R4WGDLEta9/+ccBnRt7Cz7i/TP7RylBIxamYSydcPpmDiCwm
ejd9mgVQJ7NKw3YGX2MrT4tB9yC1N5LRy9kxYw3zZqOj/uTtgq7zzmvHLE+0RNb1EdQxcdv4g5BU
se2bKHQqdF7h65FitcLQ+I53y58vAusXKTjsVGhRpax9EdD3KWW5TfUZWfwSAVThiNFmYpmEEJHS
zdwF9VO4On6dk2TjnMjs6uuv/uyIFuHXDsSM+CR+9gnH08sWKfzxDIOJ9QkFEOvNC1T/XlViOqVV
QAbUPR4xy7aMPoXKMDpfzOVVxF0Wa0XbFT7rDTqMxtP92BR284iMCxFi72jfidqvgWMKDxC7GiFA
7UVjmxJe35CgQx8mT41RTcxOOmgpueqi/GjWL6kDGlCkcoKoU0aemDoe5RPB9aI97htdc5Bm8bwe
1UmWS49+n8P4pcTEejDWZdcSHAOB9O+6T2gDYOAJDAARrbQ9dlDqAOALbnAz3z6TCnxbY3zQd7VX
tJdoF0IwLz8hpILjD1VP3u9J8V8+QUFSu81w0Y2JEBfM6TE9L88E+NxOsyr3d4nByf7Ol7gE+Yxv
HG2C8ZWY/g9gOC3hyNroWa8lMq4FPlXrrcXW3Gef4gwuhtZGZQvtNAW6LoO9l3O6NDDre1Z5u/Bg
71FPaL+bYyie/P6olhYncLjifNxiOzPhIGOfB6e+n6J/q/1aN+vnJNa0kkJtl2Igp5t1LeV2d+8n
cX3feQtx5Qs/7bLvKKFy2LN0Fzx8Jyk82KKu6eBKuvgcDX9kI+Iqq9iJ33kWpJI+J/dwVCMpWnX5
AdYyum88s27nmKSMH+t8yc1kYah37Z6t3Ek1cvxt5csDLESzyv+nRYzrmo2I/1MP9dMtAtrfunBv
ePKR3x9AcIG7ys4QWCOeGnvpzq5EH6OUPusBm8jxQbQ6aRZfngd5+8hGUkkZx4qwMcQZY4K/nHmv
aTu2BHT8uyRybwLb22JcCbofiEYWJrWMtdC5KTAO2vH7yikazw1ecVvTFnUdqe9lZq90m2CIYHWv
Bdw0M9zVuOC6BbsNH+OMP2HX8ItEkC5eWNRrGgEYttuM1aKkGX5dEsssvsFpIES4G1LBE5Ow4wZL
Bi1rypFRJ3BC6BTrzIdW7ZTg0PhT7xH0on7GD3/FVuuisfwp3AxT+rfww6t+O/FxyOc1aBL7+bL/
/M4lrZguQhPZpnyWaySQJ+LiJlk5nW9OBsZ7lGdv5POoXNpaLN/CFots2lhrd/BnIbirifo4UNZX
HH1u5hQq6ZirAJVAaJGEQZ0aFeuQqELby6lLoIOcF40dAG/W+JylAK7AN8YTpw6yjUtJCe0r7fgQ
3zSFbmbHmHqChIh2iEwGQmJAYkOhI1QiRnQXLMI12gxSW1tPQtI0N/Upm1qVziLpkuLlQzGqJc7p
02iRoCIbjWK+Wah1MzSW5iKCyr6SE9zH3RKLuQ/9nnUsccqXXVoUHqe6kWzrCsOKa1Ak3Tb/+E0+
xDtQ67jznFpIgoSXRT+Wqw4R6O+OO/ibWwlj9zOgY/3mK4CV19q/KZZdDh9HjpdNMrBARm8f+okL
JEPbF44f+ZiI9hizoXx+3AE26/REunvw8g58YSP6zVZ5wzw2sHpOnreicVr1pq88t0gcVqf/pdNW
YIzvcDz6EeihHZ2ZYXF9dQ9Pz2NPeiPXqm/lvEE+ah8x7/ZkxYyyovDlGn8d3uptqLA8/k4PhP6w
0hLuoFGb52KTKmHiUvpobWp5GZLEebcXEt2qgHyqwQ094LosIRMjx8jkLGz8jm1koRqdJxZLOYIZ
FQEhMZSUXoHv8iW8Pay3DmXEv1LbnsCfjjSenwe409oDIIkKWG0bbVqOO4S+1rP4+BSLHusdlv1I
gJjG3tRAPQHYmQYuF8meRt7cZwsrV1rxdlQr6SVOEgZssYjjiJkalMfeOEfMsjwHH6qjd4v19rI3
t0rrY+4t6dCINgG6p5Zbghs4UpVmFCCPoqdF04kSwBliINmVaAKzpZOXOCH8woX1gE+12lnWVbli
WEUTh5pPdjs3iT0KXRwnjbraUxlvtsR2t9oKTVIMtAsVfv/el6QqXQHKeQhQzyllUXB4pYA40GJi
Jz69kUiTtvuVP+gpxnEy28beWfTWwbVRQi2z7Txz0kwyOVzYggvTK6ZDsQybyZpzlFiR/t+wbX6L
5QfLgHpODEmJfoZcwPd+Rn0fEO2A1Ys6GQ32LSaWqk8nAkIem0LVjqGpHzFcaImr4GkdmY1wiL9Q
FBa2bP6Mn+J0LZIRac7T91p/Sw4qIQjGmFM21nL82tkwK6GewBlr6RQjLqlvi6uPqZZNKtdQqrxe
Ozj2I54dlVUTr7cJWq5XczkVfb9GWET+fi30EAmxb4450qMWBBExjcZQWKLilCDbUmyz9m7uoAZi
hxhEmb51vJGc3RLH7L3BEufufoooE7mif71ILQ+me7Us10bEOCpR1cglRgxsYppmRB8Lj83TIEYb
qBMY3vp+CH0l2d1jgsJ4E8lRo9bhFvZUGn1bMCxlFt0RbgWQ2JAjL4OFwn8Rb2bzR9xP2zzmxB+U
KrZCI5CqpAAprpmocQiTN8G72ky4svYecprNW63gPf0XZfrh53+HJYnuJ/tYXo4sU23OEHpwvHfn
NcT+XmId2uqVQY78AwfF0ES/sWfuZBUPPe5JO0Ln6EdE+5g8s258nmduC6RcQVN9CMg4LQwJnlxG
Fx2+53//zG2KctNsBlnLIH3Ff6Bf2gcZffhKuu2esUBX7MLTyXcOSrgYJiDl+vloAuRjCygmOAjL
EqvAu9M/v86LvP4C9YP0ZYsreM2Q+RdzRm9EEju9Bqb8P8rvaSypNdNaGcqZscXbgjYD07ofmhqt
D4xPYugHGBokUz5vADfHezIL2kR7q6MVe6mrup7VHSgtHDiTqlK+WahJo1FVEfiOpmOJVdRLaHL/
Av4qnhMHEOoIbKh5zVeGmSlGRDMGJqnxAa9rswEkC1jr3CqZLPieos7gesEiRWm/NWaanZHJ4xRf
CUdrcS5I0sjSTYi1ycvfbZi3PjfEsQpuTpFqeNx2DiZnD4wpTLN/KabWUKL+3v2bo6iya5li4fWP
k6Ga1mYfxNIEZvyIQGPXPRM//GOa7bquwDlaLBpdImvrZVkUwzWuAIp73dolHGKCyYspk/lLyo4Z
zuN2umO1GzvkytFCr7NywD3zmfF5jh6MAPA7v2atJvliH7Mfa1Lp0YvMUjTCf0naKNp4x2TlwGL2
6zikaMQNYfjD0h+eLQkGfxxT+DRvxdgNWHgtWMSbRBAfg2PWmc1P8mxjtG4D/gaIl9xqZIJf6vge
BQgm/XOeaCDTxVJONsoxwkxkNpBiSSdSqhhyPj4zOY2gK5gRheCjw3IXenphl1soz0Vt6Y/gLexB
S0UgmqQNFZILeyNn3vQMEYlYdkSRlS/7wpqcbYuPF/Z5lcNkXrB0XlWebq34TUjB02RNehPG9EXL
b3I2yIFs20KL0d0R+z1EbpsNITmHVWHey9A9c+Y8Ez+XtbaZN8VmZoVC44laFVseqnoEWo3ahMCc
vnXWhEpRNTj+G2rPxO1w0i8GQFZExTuNfD6hmeqJgJ+EVLCCqSki4QPItIcit6vSSbu09v0HW31N
HlTeI1JukuN8CBE8fmjm5ghNVf+saqdbgDEIApcQAfpE1fieNCEY8wXGmtZaoEw6Cwj4CnQOlZr2
rgtF3cYDVUrZaaazippNoE1lhsL/InsrEWYrpxWOSKkbpqUNA4llLGmQM1az72+jFynNuzTZo753
glScCKnN3JeOUK3zvf24NSaKSNFPVSi9DPiJitI09OT25jaaT/GS9TFRfhtLbdozI5uWHJoOo52/
ELTM8YWQfH8dmXyIsXCZ58wjF6iQRKLm4KWkv88Ap92+5jmDF4NmslfO2SzTZXqvkER1tQbVmqsE
B9eNUSrjD7soNFIdGV5hFTEPE0KdfdwEgDRLymlgCsEL9v+GoUfx5amX3fWfrYMQ7yujtW5HSuer
7dAONZYNO7sDJsqfSkq1BJsNu19iAxa1HqHlH+Mo0rO5beV7g9Xd+fY4/Te+2KoJ4QEsOUmtzk3N
t7zgkdXZ3IVeaiKG4bxRoOzbOS0D35SkIojYjgh4qw4sEyYs4GmOx2eswdz+PRXsl3Jd+drddQQg
TYOx9plWu7iilIg7WmkQgcis6oXBMSEMc+2h3XYIxTc7mNXDQkGAGvSRdoj9xcrZ8DVG4J+ikPcm
gy28/QQJyaAcujajZGIbaQEy9FddOFDXU0zw1qo8PXyT8kbolKqD2FnLKd+r4reaJmK3E2kH0r0b
qk9LiDM96iQlLZwzj+hKD8wDaAQykp6CMSL+/zNo0jGOJKim2GP5ToFUbibicOATbdaH2kF/7TSr
ci8wRLnp6nbU0tAoGPJSUELuVYKaXETB+E8xHI5cJ6r+HbdTyOXwEoqNtz1OTBlRu4upcK9b7fe1
8KB81t46BFRf6IlE9WZklAhyWLG1KNds9uUvLpbJSFyLntwiuxzqmgNhoBv7xBrrFt/hHOwTbPNl
eaFY3M/2At/LQQnaqb4nfg601moLDOYIeYmb23wq1I9EHMBC+GFmvMv8CZTX3Ffpak+N9CHBdXJv
4jP/HGtWF83UOPMvHB2vCtFArCSU4/r2x37fMfuVR+q7oTckakZJe2J5oeOF+P9YAaSxaqqZLhTV
edCkgPJIQq8r9NCjkEmbVwmOLxgVwSoEO3VRGOh5CdHEAoIK8MB6FdL5GB2wKzcuhRBdBXOTpodM
VxuZ5Zi57NyI+tGJrL4FL62SP2ddJNE91QUwj+m2h0Em+Zzx8Blslj19YQZxDAFUfwZVRi6HdWvK
lsBSU1aehCptS8tVk0+2Zqi9DPN3Kd64I1z9UIXwOIipWPZIFrVWemI5aVU8l/9VRCcweYJaqHoo
8HSqyyCOW0fE2Sh/ffI+5ZpSFef3DMiCaHHc06YozMnDbNxNrWvEipcy6jNK2W+gj77dIjzQcp7Y
LPu72QqAQP4EA6ESWmqhhe2+PK0VLv6kEoN0gdP2gXuJwYVSubesBSj80xq6B1f9d+ob/j9FWnzw
qoD89f5lUk5qV54s8kiGH8QfKigwqMUo4yOQZuEZqGINOnV2u9qETBaHdiRNTe93CP8idSERXh7p
kPvEug0cBy1XAJRsfn1yFcW06Fv59QBrBqJ+qRMTvIb2u41OV0aK+Bi35b09jflxZueujOyrEmq8
0VlMl3f5jiQV9Xl6anxxbTDlFJ4NiGn/pKTvDQSwp0PpAjCAjAIyJzC/HqBTEGtxGbMV+rjT4QU9
pikdaC5A1nP96GWQBs0JuHp3AcGWrksKimQgDKZIWOSKxccNHl5s7JASUsRfzEdxvQffDzK+zrJ1
raaNbBeMM6Z9pUKe7jLd4C2CuVIv2rvsfGTn5K8M5rc1rnyQW0EhI5tSNIIvZOyXg4E0nlv6nkYi
wfYQ77LOLLqIy84O+qXpX/iogZgbABvRVZvNdkoElQ/fhxUGOO4uxQ4Iv35B+LFnq31IW2TohB4+
A5hJabav2AYkzI8+Yfz+ljCbK3BBHi5KbRwWCikwy/SXwL0jX5ugYaPLXs1hB5JRFDMrIi5FSnn1
ZOcbo1ZY5zCRA5gy1rV61TrbFjSP+MeQOVzhYhwmAmd2nTqVlHrAvXsDn0QhNcFhtyk/MbNQ8/Y2
MW6AIblW4NrZtCIeSpOeojhty5yUnT+V9kYHGpqAIGFzaUTEGaTYpfg5WpC+mApVqGkO3k8VRCos
bC1wsggW86iOA1Jpvy7EHbyW1vruXD5HJDaJu2fSI3x/xK5hX0NnIIAFzVMsnx9TO2R62Zd7oKwx
XPbv8Gulkz8Jjlqsed0iNcZl9RWG900c8AqDgbg6efqwkh6GBrSnuvyhCmLf+3++vWgCdQ1t8Mrd
X/fh5fCHXGnUywMj68gbuB4IJVXDm4HaBOIKf+7iRELOAFrb/5CCDtYqPAA5sEZ82RtZQXBYQ6GG
qj81lHAhLCIPPOzZShZPuG1avU/Q9M/7PQpS2AReEuBY2jj2pM/OkZWjPg6KQGxP+BgWF/za+lML
q/yxyqHyNieyw6SGpvyCtfy9kqXI6qIu2JEUGTBHMv0zPSgsbxyldcvLzUw4hHWbxjOIrqpnQSzI
mt3MwGTaKSI/2uQgJ/806hfrf+x+qWBLMeGTtKQD+zdWy7yoVAP8VHoatsvxBiAUpbm1Gihp/W5B
E059ZaPuEZojhCMJoY4rTBQQcF0rQB8qNHfZtnND4slc1mMWtMAUJlN/hXo0oa8DvMEazfsgkU1I
cxZZYv7gDRb43EVMsy9x1tbYC27AHadRDd0bqMqAWhCGQqIY+LrsVpd/AUxm6iWyIxvk+HirJ/IB
fsAzRlG9ZWSLpaLF0ZumU8LmzEYX3Ra22QXrcwIl1vxJsUlb+W4hC0TnWfrUYu8XScrLvik/lHjl
Et19GrSoK3hcaobYu6c3RHyDOEOE+qFICK32jfN/LEeyQqKwCVvgi8D0bTkGeogoeGEZoGk9bgSj
9UIs6b9akPUZoGoyVsl5OrYN/OzKPddyAcby+hJDDZISk6rW3gUEIaWRIgUC1vo1mgMjGogHHWJd
A9ftnAQfym8vBTPpbhd74e9OT5MH8dQjA5VmZBfF14LYZ0xlthCF18PjBlGlRMIG41xnTsaeSoZ5
PUS4IBCMKOujPGUN8rfKxIZY7a+K6DUes3p6v8LtlbsxoZde3l/d4cbuucG6Rye3V2b9ANJTuZ4j
bFI/Siz+cKLyiJ3ZMrKKhgvbBI1rQMtmTKp+ksosGZHWRpYTn7w6CdUxvoBuWtC53banzEhZ71uz
jJ0cNnwpStna1htlsNJwrDwIyXGwAoogAdBswcgC5xeDDWtESPYbaym3tpnSk64CQr1eOCKna6f+
JwpeUe1Q+xkc/BUsoWzucEoywiria00XPGcLa9FCJsAD5YOTcBDsfityFuBL74q4cNI4Q4w3PVtU
SPtV892srcrUSiIwqtelHT6mpm2bV0MGfhRYcdWh+rJbG3PbO4jfPIPMOqJC3YqcTwtIzvjFul7b
egoY1y+zCf8/Hud89pMOKIhnoID2ACp+UitjJ6cUrpjNumtjmGPAQKFlYmhbG05l29QjYx24aE0U
WsRm4wZ/oEjEFYuRfN5v4ERdgqKh903MLQ/KVZ+HDxOM2g8zyY174/P5huIUYqXKvf5RqIeqgml2
JaUdFa0k2tIe9GFIZh4F21qIqmeWKVDciwNqUnPIWrkXwMqKQhfVjnxlfeoIhvQv3AchWlBGwtLf
wjqD0/cWp/bCd60qxtwmgc/Red66h9M9M2DaVq7sXl7W8TYdtwMTVAR5mQUbvjSQ3CGMbH1iA7iJ
/Sc+fcv0PKE5udGlQ6ncXMT4L9tbvsRocm3/Thp/mWt/CR7SemJe+ucQua8iWLyL/jfGZ1SDxi30
6xX2fjlVmSNof55OWq+k1olr6Tqo41U7QF/kl+t/CpI4WckjjjIbQ6qQvU1HrgV7iSKN9vojw4kO
PJcCh1LhaeVoiPWCnlB2YRlTA/xMSyr1J/1sbu/7e5xl2KQOAtAKZp33C6SXL1iNGQNc+Kj3xYc9
izqu0wJNHsAb8RM2qVcQ/2Fvzp05Y4R2DL1+hlwcLHiwG10cU328BSoE1IaJYzD6tbd1tjYx3VYo
SCPTqfUHICWIRZZIxs9I2jxWNdmRAIFwHp3OOm5WqPNXPadtK13KscmChmB9xBdngd1l6eh/cJe0
HLdNAjgfa/Wu/KeqBCY+Gw/0EZ0VwKV3Y8MqvE54KqbNB0KlTRuh1VIybk/hQZfCiviiqE15Tw6M
Of8Tk87ZPhn/4JaCRmYoL8WTSiXrMi7nWvQ2pFPhK+f45/RE23UAFVlhLqTBy+yLqc/xErjMTHEk
VPsFjn9m/b0tuhZpNTWteQq+FNscnflqMKIok7eESY+oLTSLGs5AwHee+AUlV+aoD7TgtfxVCM2N
yfA/q8qvwzfjFtTV9GyExMJe/Mm2HvfhGUTZoFshyhjGuqsW6Kwe0BI1gI1uWb1ch6I6nxNUEiBQ
wXcPg/XQbsL8BwFU5/omG39KMCgj3a6S84LsKfgSI+PlyZdcsTeJQ2xQDWqhxNm1p4tF9i4AtCKU
mUVdnZCMYHOW6Qn0woVspUKAJ8G63LXTcZRSzq8H4CkU22+uS0j4IqsihuLlIjo7X5iDMPbUvUW+
bpLZVMdatuI9thGbQVKxh5cKs2ucAY4DhS2l56Cnfej5e8ho0A7JyxBQzu00CyMj41SB6DLas79n
TSgMDoGb8R5tlNoHwcsH9aGTX0LZzV57siqxOG8FVdPd3gTHhydCC9PoGrVOkGTunX0Yuzy6rhwU
kTtOAk1cyYYCP89A1T/7lbi66DMpPtLy79AXSg1FCEK+uhYJyu6UdrYJ9f3QmjLgebyrZ7iZrVGS
m4hlOc0RCo3apbFGrndeMR1ZEJKz4DGNX7Tj8e1OiGtnTKIIHgJRGjcgoykEcFdv1qH2p32IOgtt
IJCf1uBZH7b9gELQCdROyiRPHtdh3qjzW1Rayz38lJ29OXgQloWFGmkwM+MVpyuTnTeHfbvcwBUE
zpc+Rhpx+9Cz8Tvpt9XYerZGfSLHoup3mOhbIXMBFil8HHROapiNigq7ChvdD8yNIEOVu7AuoQnp
vywdbnF0YCBkXa8CE6y4CWgTIbQUaCAvVaA8f6VBcmY7f/r7NwEfA+lzXygLSbWw2MDcuVVvHgus
2+vffADBaYpMf22J5MD+EKbIOsr+GRoZg2suIC+gUhVaD6SSAn5/POld83+Q3LsHMMn8ylwSOlP/
PYgx8N5bWPrBRk4aWUf/0ER02niiuKedUqwrdvSQPplDTtcYmrIsp+KbaX08VUPrX+FQ8+3g/xYl
NvATxddxR+HemzqqA9Dh/y7SBkEkYzKxFfW9TXqx5o1BfvEdDKUFc8ic1C+Vwr6vKUNa3YVi5ZGl
wEZ4sxsluSL/kFoBEdNje+LCb6cKAPPCID1M0A5my3c0COAPAUu3KN9kWihezf05cYIjEQUQoTJH
InhB/r81Ine7Z1pq95oSc4IqDdLXNC2XoBnuElpZM9CoBaCsAXLo3Y+owIA7PcTzguN3zfDHAcma
8K4j3e/3P36OJKqVKDd/H1gpDNgU+aIkSYlOmyqf3LQqc/xvfJf8Stiijf8qCYvWfnCg1BC72Kn9
LB4+H4/7YW7iWEyO+9QMPwFOwvFbc2HvcL6lQmNKLSG+0LyecI5yRE6Hg9TbMlzCM2/3RkQrPQ4a
aDvaYtlfwEZ7RXF/MxaHnda7sCZ3I/dx1kX/CcPmwCxoEsW+yBvRQUlDAmVl4tLENp8IpJZxkVP7
E0xocx/uteP6PAJtuXUOy764ZqeH0KSnTJUT4F6b6qSxxvcjfMt2StuvV9EdzJACCbRXZI8bjK9g
RcLP496Q+mXWcCNwF5sCaXwanUr2phWqr8QLOK2mKAZKLLet/v3e5LqfAcFiZ6sbcdbGUsJl3SkF
pm4lR+Aq+LVmgSI2YNqU9a1l+RS99Tx3JtBO6v6+lPkxfRA0OtPBfwpDmrG6b/IWft3IKGFREdGu
4nGWZNOF8OngK7XjBkL2HjzMegyG408YqT50jkU2Jg1/IYks8tDz9B+FE7mNAdmf+UUCC1Tt9EcA
uoUV01e029t1u7Gt85qRwiRgsMO5ocMqcjWE9Q+DSGzmqDGvAO5eqrtYW5tEFE9F/UCqteyxxhj3
GAzLCCngQu4yAbfevhxN97+yOjcO9qiXXwEjnnRItge7r+ktkp/gWPngKxQUJ2mAD2KQOAwb172R
7GJhK+7xfuyClgRCncYPMZ6BFAYG/tFOD251pll/p5mnDDYyamNBj8JD/LlI8OmYKQNKQxNov6pG
MIi4Z2n/CqYa5jt8+1bt9H48FOu2qoA6WezUQVuHZbLbjAQ7Y/kt+Bz5BUr1Jt/7w+eOU26VPDK3
5Zt64u5zoUoPPxMX4SYkI+nGdUoYNN0oA8TKXBckI+kr6M7jwrqaj+GKHBPW6U5kmvmxLPFCf3gm
LjS+DXlHPb24R3HfOhBuSdeLx6jzZ1R5l25j/cE7jD4+Ol/gnHflGtYhgT57InFUPhqwFw5F2MVR
7FZNJ0p39dgX9Q4BGW1y11MVvgeB8+BVhHyRPyc6CAYyf4GbjVkS7y0AeETtG0DFF0qGEn7JXYj7
tt4kaoEV6Idb7mwro3bbuHIRjICboi1Llb3ninv2UJKz/eOpampYF5FtCXUVDc63ClYd47/rl26s
qRPUrAsHnvoCiwl2G3MPR86A6ZMDiNLh6FNi1g5rKnZqUTYj8xzlRdnNFak4mVTK63x4mdEFHSGr
x2/kQixTcOy1/bCC6QEsf/Pp0ZM76CzfhdtmseOj/x2HDqPUN22Lua+yseoTsOpF5SziEvJKJo1f
QRAqvSynZOHdj4aa8KcCISeNHEe6rjZ+fgqi20PRpAF8yqYFzPa9Dj+yZ8m6lmfltHArTJhhsN1q
FYieQ/gTjTBTmvjc5LgExxRmDUdfe/fKtX7Rc7H+Itc4Mc50dbxLEKCEBnpwC6Pt7aBjxxKyawvT
WtrffmDrOuQXTyOSkdtja5nAStdQCbxy5W5abqvUD1SN67MpogMycUMEYWj9G0xQLI6TzBLjHmhn
OH5XqfQQgSacYEh+64w/4CCF6uMTS52BmKuDcI+g77mq8MGznx2OFesBvdiC3FXnW18OOMZ+DOv4
v3qoGMbrOCSsBjMlGLVkdE5Ahh1+E971a4BJpjFjxFTm82owMdNR0IPrPXc+tzolfIzc/CXp22Pf
XDy7t+0gT/gBDpMkN7+9wBKqQzKi3wAgUfE1rJCQNQkZ3sG4HZD1BPr+nSDHN670tbVycROSfpBm
22nOe+E+NvvQUFv88eFdodrpGUgVa+BJBDtXHjcOA5aqcNGehqT0h38QeT8FidmwD4oYvJjZ5mX4
RFHxVTEkZKpDv2MTmEdeqGMvnb2OWMjwppj33baL0potGFoGqCVQBJSVN93qHp5bfM0+f98UWv9w
jaST/GtxzT3vUxHbXoLvSsBGE3XFDqqh8ryQQnFNI8p5h2LU4jLYp9X7BtbrSLMe2X9sR9UStI9d
/f6u8AcBXjkqsskjRA4h+faDWpuUNYE86E0ZbZWiZ9jUVYFcCb8R1clrLI9ESKcE4UmAYnPZKqA3
2sFV05DDPBnKfS/XJLV6LkDtMu/gXYkoHD5aFBaIOCWrCISmjf7YbpspmQy/Eq93xy3y9IwSmMkC
GhlYRF+2EMuGshr+hM7LHeziDWUMTafyq3BwA2EbgQe18ceMfrMOTnPfqvnZeE0ajchgK4YZ7k5W
A9NbhqOw+0SDlv2CIwO/pe+FsalwcwgtO6zcG7caHj5spBtz8Fvk+15L+R5vinjTgtmO4hkpQG9v
QjF5MWgMmo/k864yyFXRy/0GhRO/VhCzWJsTgdDt7iuury/TLBn7H+ibtdomaJbJQZAMMZlpqA/V
hDIpMbezf736edGHlcX6yDkwCAhaJUWNtHKiD9ZWJCPtQTMTUXCzvrvWulaLVmQPJ5PqmHtqrUJ9
pOJQQDRaQBonsLN3jcsjBcZm0leRfDhnGsWu0AW5E7Noa2crSN6750JxwJZ9AcGH2rSA613mRGBx
1MkmAxiSA9NuRQFsx92o9YrIQ3iQ4cEPAMNUask3qp9WwBs+K4xYLpTN8b+2g97FXEdgRUsmISie
lzGGe7HfqxBLxUODBGBZXEebaSne6HjoEPCFa6jhzS8+2qhxrDnh78uOB7UwJvLIQEPzwkVJtYpt
JaV/gjPBRtQJFYR/dJmbq4pDaK0jBLoI4hUIm2pYjnay3y1txzc38forZuIJzw5w/4gj3XDgJE9S
fCduH07ApYaflwdhwmi4GLLRooJ6NkQvLOLbiYn7W8abwYyMx511OkfCnCBGXYiCxSZk1Grzio9x
Jp0r4NKmhrTnzN20Re3jcjAZ/v3j+9Bagt9KhZMiDuTJ1rPhK79z9kZ2o8B9IsBG7sZhuJhnQfj6
pKClk4bcb53WcKedcTb/hhCx4PpOhFr+d3u/z/hzBAHfUXWMN9B5xKixe1HqRHTbTsMZe0LjN2hH
rYsf8wWviKkXTG/K7XyHOUBlfjujjYZRY47pXGmjWkaHYqDOJokuaMxX1YBo1mFrew7IuzitXoxb
pq//P798fzYi93EERLVvNXkJq86ovfcvpakWmerTEOAZLqV1P7gP/fC11xKgHn1Uk/SpAOyXk5sr
sj0kpjgkrsOe1BcGbdsQM01hL+tjDOkn4Ud/EUNaJq09ImJBWEYe3FygRq9eVURS3FnBY0J/46+K
FRGPLFZJSFCCLH5QvGMh7ruiAexnmipscBb1OtyStOmDwdYVdLBF+5ElSZUcgOtW9RPaYdKKKhkJ
KfPMgrK68nmI79NLWOFR0JDWbYLLbx7n1vvfcgathHouuXk1pOsm5j7GuAYUw1Zjxo2aSAgoxAlP
UIH/EFTK6Nr3RTGHLV14e9D/75lkqDQZOxEZsKLgslcpBI2qo4SiWU8LRfWlbxPJzYB6Esq9hrSx
TT9q/IX4nuZv3awdof7O4BZgbjTJitoGJjAuc9CxypM+EtLVJl/LC+G9fodH5zJ2j4BxDiiS4GEo
Eoe5N0q6bMuFUvnLmBarGDZbH9crSXsvDHmRlWYIlc7P0HkfmHSOwDoV7EUFbuxkFdZPS5+/42FZ
rCeohVk9zQ4tES9DPknb/8r93pS39q4kOAo/2+tM1GoN2suZPa9IVD/xcggM0yTyTIcGy+QZiZvx
yz6zHzzdCA6FqQ9BQHuNiDKLvweRcVZXm8TuZ8aqbh78FYsuYBk5Z7NHQFViFlQVG1Ocqmk2fcAb
TfZY1xSUAV5mqPLYzoLIbJjpgkQ4Ccsh/tP2CKqOGC9bbBgmtxRegbrpnwhfoFWD2hA0/Um3IW1j
K28D5GksOiiREZCXeFTlSrqvyjfx8tKBQ2xxQJrGe4exHHyUw4dUdMavifUy1gcagKnnQHiHMDhH
fUzT/tF5BkKd/dP6Dla8tSkya7erSimG3sFEnq6luLiHFj8HHbeklIZs5mjs1eMws5OxkkeZtBBd
Ryu0i2f8FPgyom+K5zWhtnfybvf49VQAljnOEMKO9f7C9abBS/0rwIDs1T9d+0kK8I45kMFzj+UQ
VQVUjGH2JJ1zoYyonueVDNPUEbHLS6EHvRoxHOtJvpsU4X2UZMTSbG7iFywd07XqJ8vFkU6e1ESS
g6nrYNSFYHUCEAZW96R5AwT3sRd/MbRFOhQ5ePyaR+jn+V5VxU4U4hMqpJBe41Oq3UvYtnU5Xqp2
fkf+SKdTDduw8lcUIyDW3UVSFZk5E9EHAqtwp8d6QoFosaTI/ess251jLdiAiASCqpkg7xtc9i7n
P3ubuFXSBHls3hJmxFTDI4flmYTZtagLaLqyrELS/LoxmUyIAHOxk+bXcgXPglmo1wbr4jmAmoCT
5redSiYlY24OsLv5Jf6b1fWFTc6oO/5S5BtH023Gq/EdWlHdxlJxPOydcNzewuDVfg2YyJhdCsbV
RUT9JBIYeFetHiTv9OyzRD8OBuxQ/PngSUu1Pf7XXGR4wgvLuKoje0LyFvDN1ErtTVmQad1r4aea
5QJHlHjnGGiv+Z8vSqCiXwRiHaCaVyIy0+RCO5l/tn4yhuPOzui2n9t6OACC5VczE186Gn25TtV7
cuTZ9KK/j7zjXMLJKdv/OrSMIvsdPmh/yNouytC7OFW+fk0raOl73XkkVOzdkxc5pehw5iSz0XV1
2f2BnsW73EikNurj274SZq9azzAkn0O+HJHByPKOAUxDKAypheg5St3HvKYqwR7jzWLQkkeUXQ+g
ozVEJN4s2mTPSj91Q7WT9XLY53o2wNTpy5s1cR0HQmFVSwRYoGvTFwsPBdH6FH5X+i1Jpy3TaaUH
5Z795kC/pia/Ym/zH1j/tPBD36pBjn5RFE4cf1r/eTr0N0gEHrWoPvDBzKJZrMUqmpMhi4jPcVF4
Y3ub7MREgTIVwaY1BjKoFKQVI+F7yymEdVjj3jUk256o5rC11fx5W8pLhui/mO/kA0XwJD7my0K7
S4BAuchVB3NHzF7ejUovpkx/5glLAhSGxUx9W7VdlHzbCl8cyrhIs/+DIH5N/n0gCu+ZMOjD7/fv
CViqJbhIuP4HPeHTd6uZo7La8ebwBiQ+9v36yMJMWsQmSkr8boQNS0QjMs8QeinlhWlBuzWNO6HP
6gE4jIS68/+7+cac565PKIjiGILy8CfDt7kR4N0A39qh9vbNK8nSDgPT4eCsr+PQmHTYUzmQ8lZC
u7EgY2Mxxzb7gpdWbOc7u2bmW/KdaSHxp1tAQRLecsn2WBT/sEts5uXnh3yddQ/fe9LSrOyD2M53
dr8avwDAtc7gJyGRbMrwnrXa9v+ixHyZkRZiNCKpdCP81q2WqRDCuB78I74USoirzJVCXFlA92cA
k+0gtmwH+kwG+IJ4fgnz0wajuDuqhUGJXTYNCVzPfcIKgfBLv88Tr9WxGnU0Zgrm88yiJwEnfkr1
k09/dhIBo9cY76rfZakAxb1zg8ROw8WgOUn0bZ2nzbGtFoQrYqCJqXnrUp9HPAoOdDqTrFXjNAUN
D6V5OEN/QbLsblj4BDQXpf7bxZb4u7+5D+fSrmKRnDdQ6GN9FcbY/AjLjUHmb3V8nCe5dO/6E2Dx
IAjrW11toFXp3/l4TALKgSOHltXZG5WE35+8mccBj6BhF7qFTXWBmpLRT6B2xKhYAfgrDRw9uERu
TASnoeg/Nfxpsx4MyW8yFds2oQpFEZo9dZBmszmzY53rGNn4goc0u8czhZayhF41cxWmnR7EWSQf
Oq4jbYk7ywOFYJ2wQ8gyKA+EWQX3iwn0Fu+87yRJPas2v8BneByYTkz4KFzn/59A0+Mxva24ntEh
Vcx+Vs5zgqZkUpOouBkIf9XhYV3iP8rKfuF3VtfyAIsA9gWALyyWnPFaRDXFhLY1anWPu82Nuq4d
ShVzUwz+4qfa7Cvb3/upsnS3PkfjTK5lkhBa9wtgrOWteFiweHAlcVIHHPc8HCow7OsRTUbHRDcd
Kt9An9h596bCcXj8qvWXGHwa6t/P9D7rT283FdjPwwR3VvBE5u6TfFAytF1QlE/5B1UAVQ+FFQIG
rC5PrJaGvgK5TXJelMA0w5u9p0qQer8gb9wyrm5Q20zLGp7jNq76IqHdaPO5rwpVnKBQSmPHIAZ9
6I3Y7LGIgAzU5SMpKCHcAMncTwiAux2NGWUXtgK6d7/jDQeGY9439cA6i07b0FbzLS/MLLSZUA+J
5Yjqsh21t92Qxda+if3FGa3Xd7dts4WOgogGOlWxlpgYCJXNFbxNT4vrS689R1cMfjXxcJ52MGRK
wgBugy4F/xYSf/iLzEzJtypPgCkKtvEJxzYaPmYjlbNyrTiN3RscJljqsmWgDDK0T7OAoDrSsg0t
ZKlM3xBco+WUJMuNFAWvDUr1Lm/WDLQlxJZaFUXTyjeJt5SncBdn+//Snj36aLef807sVfAX/pP0
8+gFg0qMSVF+GvRErV702j7ul83IRKzbWyTf3DQA0+YvYq88eRL5eS0h57Fnddx+1RqI0jgjKwxW
rw4JiXGpVTZrl+zEK4kAx07UsIvxnUb8dGBEI1knKeSOqlR9OIh476WG2KENYK6MrrPk9qCz1k8p
CQtNtjA0mcGgh9Hwn0E1N5JXE1c/XY12yzJpaGbjZnKUnwYmEgAWjFwGFMi8UYpNYCutrouQ2sve
Ts2BvhiDQ/CB44JZxzkWLWgiJCkDWclY7ZG9f3RiLV4L2jTb2zpXRGfohFLl3kmfVTK2jlZ3e3QC
8hqg6bXf4bL5lrKSLXrdKLXIpyOULPUQ493M1Es37ZV2xFvpoOz5ONAyOcpesnxod83GeaMEsMK+
6TCNuE14Jd3r7a3qFfPEaJmqVmgm/2/AUKRWvdjsC3Gz7OhD/2qLiXNmtN/Rql4itDNLbeu5P41T
wrqMpKAkiwIPaTCUS48iFaiO3YvgUpNFW7ZeXRrQzXfMXAs6hKImyPgSYr3ww4TvUgvzzUnuWGFI
2GEoJWUtP6nK3hwHFQN8Kl+fWLdJYuHonvZJHnlMklD3zCytAt3tTnlY8L1bRlInsqnN0UpnQNot
0fOPNfn/rCPuF4WsGF7Rvt/IRGR1oHXpxj4ecqKQ8KV25se1UipaKikEikE0AYcPg/h1CTpU+zMC
PZJHX5C3ZrgAS8zp1kbONl0RlZqN8yzS4MZWSb0xQMZVaAXTdU2MS2vgv5fxfz5xO55vkW9xxCwk
ii9SY8Ryio7CxjooxOe++7nRUUupL44oq61mL9YSqLrN08Wk/iM5Tw4uqzuUvAp9DLPl8W+PraSA
Oy8a3BsV812nqgXzPDfi7t+CmnzcWG2AdbSPleWYtjGn3XnHGn+skNR7Bh/zqjCWF3A9vXJttlbQ
8/TYhVqv4PApC+YMvmgwLwZVc615ulXaOx1Ln2ZpLv9Ln+ZKlKRn61/E/hZ45V0448Htwv7PXbHP
Tmkbf7vJ74tZKC1sUmaA0LQXPkijvTVCMl/4beUNzsYzIWU7PgymMmCA3t4QMTkjHPCHVi3jkM7s
ggDfEiWEsDRbLIB2Icm5EWiREhkmkXGfsX0ZLxOl9fVYMDP/67YX2cVyy7xVuj4OFMbyeUdPrd14
FUF8Hx05aSdQXVqj04ZJHWaWC3mXTTSSBnDPP+HIaYk4A7poYV2moSuJhKXFhKLfchuenegvN7jA
3zOfX11fudENK7H7mtV9GeuokcV//uVgaCTUamJhSXjXs4GgwKPSbcjyzrCUzpi9+3/g61s3Qoxb
sMONio6MltH2L1cBzk7UQhIQLF0DlsNzcMf0iQNZKWvznMLop0/bWmgTi4uqBnAvHjKvnxSHuxvx
YLEV71eBBfXad69riGxXVM888bT4zz88lCin/H5xVFxPvAZRJQNpOALt0514/endgHRxBafyhjLx
6agEUDzWbdVoy62pk/Oalm2CcFtK974pCg5JJ1kTpBAY6R53ttwskRF8mb6F+KyTESmuLx8yxncA
oWcKUccFuvyUwMJybrYBnlNJedfcYP1+i4iDvuBcGVm1D4qLSvFXOwVgnPu9UcPOhFhEqn7aeMsf
+eT5hpb7dDnwp/Elp4w/rWLD1D6eSHfY3IGG3Os3MMnCg8ah0gwqeIKOcdEQd1zJx7CzwHyZiPNT
0XltrOPN+63izRuHrUdPcr58oKXw6lcPtH8unA8eyqwT4VKdjPqNx89aZIGZ1QceHJesBh5ILuoR
+wmNbKOIkObzkq09QYUnhbDKnpRJZiKX8Vg1En/h2skvdmbzLUJai7Eck2x+9ecbCYAXdWKDSp8F
nb8FOAcwaR7xh3J4x/wVxPoYmHHxFDnUSjrAR6+e1CVrXiR+n7DjERwrka02NVeE9WTMmX9i/cPt
bGE/8TcvIPsiN/hxGtWJvcgfRJre0D3U4iY5fYX1xOBxCm1naoIviqPVhSZpbTjosw8LrVv/xcuq
n8Aa38JKESLi6lIdFQHvN8h2hPMcB9GGjHWgZ+6barGBBrm/lSz3DpRbpJheAozrJKD2WTDPOLro
rwh5txAjZP9ZOM2LrC/72fqavyQDVc/+XHnJM0vfe/tYTTyyctWnCmkvZhVlsNO0S4ixEI1oZvTh
8LOhqmxqu23shf/SAnPes/iX9J1VN4HwPDs/zO+lVJjfg0L1k9qTZy4XVg5GgOVek7O2ubvJB5rX
U6MuU9iT7lY44uceDAEAlK32qNZ5YsBXKyWYnoTYgYvs2D0Q5SLTIQ+kxWZogPR5W7LhdT7vPgun
im8Rqlhxh1waBt59j2pCEFx2+VYPBRt/Vn193KH3XzgPndQEl5onxwfSM5CzOIUxuBP+89XFFrwm
/eWmM58a9O5/15p/U3SFKEkjJ8sft9N6jXityI1ICa9gr6SpS99xHTyF1IAuf0nhkll39K1FfcR1
TXPeI8rA6HXPKZbLdquyRFcoEAmCbAyJLRBpPrASS2EBcxm36kc4GpKpVmm9NnKcjgem/LcT67lA
uFCgmBW30izgpqDfMXgLVoRNFapXiXlK6vJn+L16uYOeIz39n26+eC1lqCDA3yVtVw4u+eDM9Xy2
K99Zf/W+fPtZX/0BCG9g7X98f57LLkO2q8fUZWwF8uArDeaVtnKM66/q99T7mo/XDdjqeOsiVnA9
y7YWMoqJkfgvCr4iSA6/TsyI1o+MKdwApLCSxLa18O4tYMW9/8v4pRakhp2UMDLkynxZxK7D0GJm
0TUoGveb3sZNyyQmEz92MTcdEUma1y6ZHCsHTmZrm8LEa4gLhEOZXram1T+Hi01qALohIBCgDEg6
sk0LTAcp1VMESKu7yBKzLm7dbTeWqjWw3uB2bVTGRk8jIl2IPridaPnv6GYIcr4mkhqSl3cCHPL1
XSX3Z4FngclDrrZ2HGlcmvNjlg+tk9muAYPJv74WO5PMgy174zksR6K/kKOC+xeDKNedYrxGMfCM
CAtjSmpkwNEkxlWFSmYeXPaWJfuy/qixOsosFA+e66LlnmdQ5IJsFx4T5oQDyRY6lTHZm6xJq7LE
GFFMfOOyq8yZLKWIB1vZHmijgGrRN0ovneNeEFJBddOw8P0sdV2YyusjhhmEq8lnNeaJ74YClArr
qViC+d/O/xzZ/sqSFWgin3XCHSGR9RDEId7vNR/UfKwIhzBmX0HHA+vHxXqovRisIsHKNt1V7uHy
W6S0KcLZjSK4Tk32qMwr9kG3OlSIR/1Wr5LDaWAwD6O5i4YxmIO9YoukbPn/ThmK2m1CHDMV0Aa9
T9GWBy+rbmix+QY5WiGl0VKI/KFKhzIIs7x5SHk1HL/Lq4wj0li9BEZ3bXeTbrhyaunF1GL9ZHF+
eKCr3Dni0k9gDmgRf4EUyqF2omL+E4Z5nW/TWi4RMMKI48DEuigQBsJVQrO4g8zeJPMhGB7oK2he
w0Z7Auq+BVz6Anwmfk2HQ6Q+3/3VOkqYdAjid8hCWNhNjQFq1hajQHAyuhR/XQRZGJViGkokhfHq
/KHlmfQjq86WbecfFjpUlsSjTBXchy0PC9qoHy1DS6zqjmIQG6fiU0jP2bt1uTh/WNLAlz3saKUD
xhtbD+q7a9VElFVUo6sYlT5AzK8T0OkjEldUytGBJdFKY9upGLDyoXwB0jrmjOQs6+tZ+GlL6nsH
kDDNXpp3XYoHzkRvQ4PAOcoAJ+Tx5O+Ga0VB3Qi9QykP5Jwvsxs3AOsEZvBplD74Illjnzi9I9wh
NkNtQna8Zgj3aISphCgUnWPvRGd3v1DbUke0+pCKOcgbra22pn4T7ybAHK19oPFfA081fB6M7Xr2
Xmbh8tMDfpg5CTSlMPtwR+FEq3qJeZ2UT1UOTRrnGyONzSC3eGrixKwOLwkgOnkwSkITLzxEzSy2
OrMPPn/GaGYtNRwLWp5e2n/FOI+2yfcIJTPfNKgH/uoGYedEp/T9zCRdO9gGiLIEcn/rpxUjI9Tw
UgW7+vWlqed8r3UlczL5tBYnQ8wQcZse85vtElI/OVN2stWlS3HRc2JxbJvfutV/2jjfksAOs3QM
ODs2MkrD4XCfajXD7N1lPJ4ifB5iK4+C97dN9wQefacDUNDHMG+fR/6TvEfZ7wZ2v/fUSnxKVH0W
+x8V7pycsSebiwxpxy08ESoOBdh6OWhCh1XfK6KMDcicBbbSC+A46KrStK8VU+EJj92K3LYzetEO
SMbM+9IiNnVTkRXuN8irdZfiNE6btKtVmORf+0TU6LeF44hN3Lcz9fA1VjYX4QRZcxpONmaZzxG7
V8YmY/WvN1nj/356e+DvUwPNdKmQYTYb3X2gjVSZQN166rt0HSBmWuFJ2i64+jHxbE+EEKQlFFBY
Qcgxgakk06AkC3ki1opcVmcTE3QSY8H34nRJd86sTDnPRFGvrF8chIWCHJIWEVt/aEWMc+5erxHK
zHKCmYyiC+xLaiXH5i52O4kPC7t1JscsK7IpOztw2WzuvhKBXNxEqfN0TjMvZ1IXQvohBZALDzcd
XgPvbWUUKNngx2pmR+8Jegfenp7RRjiZZZBUcA2Hxt8p8GQ5RCGQ/TC0XrZyRVscAqaXQ6gqTpet
XxLEeUjVZfFNbnoX9Moy0TqbsIBRLuJLZPEEfouZlqM3dM1Ay4VyHiFDXLT/5N4Jg44I3A248CXd
7qI9e6m33McBmykVLqaC/hdTRRZ+c3LZixhiXt8Pw5r2FRAkvJ+y6JvpoHnFYC6wkCVAHkWkraiq
UVMXAOXk9xmQk0iCzelFAwy0sOrH56jRPZ8OVkqLR283HR3C0KFihQhi2hNXPijAxw+zUffn01x1
iu/qIPh15xzUXWGm6jjERjYgRdsdjaxx/TzlARyA+GmQ23Fl31V15lJEwHUMHbWPWc9gkml8JpaH
5btCeTaLN/9b3pNFLP0upulT/Mn4e0GLXEfMb9HOLPhPYJ6f4Q+aKheoZjk3zM3KS/INm+FjyZL9
ZO6NzlPL/y8j9DovI1SLQ/P/nPV1lUrJamec58pvMB9N78WCYeQ5pND80xZ/PhaxjiffB4Qf36J9
uaEvI1MR0bXLKM2oGvaac/DUIZHaFgnQFEOy0GWnPDu4GKbhElKUnNkm33YF1yIyjGlKbCjurAJT
x4Va3sjC2Sp1OmJ2ZzOe4p4bYTuCmgQxR+qPU2az8aXgu3eiPEOToo+IlVDnDf+XzCNyzMWkC/Ej
gHRK3+rlxuliz40orKP0oIHuO5mj0ezzEljoSEaRoVOc5az3Op2j7s/rv2ladw/iwqCenE5FqhZH
uyhqMMS/f6j3yddFsz93OfLw4kPbg3V32+vGJ8gCwoMyoqL8xUlmv3XduiKuLdmqmmiQbhJZ6x0O
x1OxnFCByuhwPnPGkniAatECQhTachJ3QHJiCr3zmcCgMjx8y40YcM2JkOdjaAYMrQ8QymeCfvap
RMtVV3IuhJ4OS+1MsxStTByr9BpZu3Q9mf9cXKbyJo+B8UAy2OnnQj18QpO6IphB1d6pyf687Hvc
gaG0/O74oMnvKDiC6zb97VMUia0MYF+XZZ5i0ukGOJTMPCjcRugi1UvgLd78GaTGlq3bpw4oc3S1
4FmtLkkXDhosRMfe4/XONuoEmC+2dd7g/OCxZlyXkoC0gxFz08UmSDG2xNJONp3ZJEHHy6C6iOHf
pdQIAKDolwiDsqQZCa29LFJ6zHI5I1m49n9Gr3O5wRtLrBi+vsbnUMDZcl3HSFN9JHSghzAryfF2
Nq0fej/sXHFp+GK3xLkc6PRZ0Te9tfUVjK/2cujhbJTtLiuZpSTJcAwRS5OM5E1gHyTY/zt5Dd2g
NJe8ayvELRBI3YUvasTzPeccJHFKGrEQimBV8XDc49gxbjs+DsZjmM/opL3o9L+PFvAhcH5aATMi
E7Dkt+2B5ztwF0h98HUqWfXEHYlTz3Ijj7l2P+x0GziVJSHiaf1GMfcdAgGm1ahGJwOQ7S32qjKQ
Ln7SgGUfkPj2Jizw/eXcaAuER5SX1J/itIawaxLM0aDtctpRZy4dxnW3nqc+twlL3+HSlBwWpvGW
NYNgmVMZXnbCPv3BgOdax6+yD0dHyJUViFzognvIUJ1dm6rVywc0ex/eUHuGw1Vp+CBxAezxzFeZ
W8oznk26y1h4GMUF3riLNVYd0lkKSjux2Zm823qCesWF1FSPeMixQLBu3tsSX8FPjpVA9u9+BfXG
fPykKnI9SfPQjjVUY6TrEnwVBmtbJRwQjzJtTEI2IWGz/6utRCMDc/1xwBBM3etyTQjmPoUoGmC3
HSUS5U94AxiYrOkwix1SXuxVeXXAmoWO6izh0pKMj51EMxFGDL06b3HUiiEYhKvERD+Gg7L4yj5h
t1kv/J4nYf+jMzIq4mA1u5XGMOnF8KpbqheNX3ZDNnz//nrrndeeclSW3sosjUq5dUDxw/NJcKeS
c4gkFnsFEjg82EUf/jwAD/sXZf4pl43xyk8MHuOOHVIUGC5+kcW1j4a0bAPKhESreL1Yq2tEK4uo
VN/Il495jk2oxgrrY2OWc2zt5V6CB8DZlG+kkLrcXHYJ2VIxew0/TNgEYaQHrv/4OWSR25k5QTL2
kaib6lrqgDKez8y1EVPqY306gAtBS14IJ8ciuWOFtX9RGa0Cjr9Izax2HQPWLuW+CnT35n5jyEha
D65qtEH/KRABCcyhWGQMILljxzZTeb0yF+Udn7ncVS9Vwwom4FQtIaQ2nTybZYzbZBwzWexj2qTP
X7NGHHFZWZQYwDTYKryw8lG2IZNIVgRF2Xa0/quGYlEgoSdfBvFRu1ZFHjmnnCpxEa0zRTjvGRg9
J416+d7RwQIqMS4XLRXSQPAuKKT//cLFCVCdK/hhT4bhgeZ2WUzPvQIc+7doFQKhohQQZrtXKd5u
6ouzR745pIL4xPqp9YtZjV78X94VEsuwbGICcoOkQrCbQ/d+1BEC7VJ5SJ8M44y+vNO/Xgd5pXdh
yHQYdf+P5ZEKIB9vNzDUM/dQOPf/FOLhZkQR0y7NTCng4T9M4K80A2+jpM7S7NGLYYMpuXrm8PnY
lqWhweymP+TOo0Gr2lZV6TwQD4KG3ftZouSIWVkzEKs/SYUwX1p1xfzqwqYshPaV6lxh9VeFHD7l
odY1QhyaSQjqyrl+fzXp3/SuOI4VdO8Sfxfj/rJGm8vZPkVmUlKOieCa7josniK32vpZ5jQJseqI
Q774UQ8cb0HrLV1cSY546g/+y/JXubF8bokUMG4R3ORTjd1qpBgcfnr0cgf9eViKlA7r3PSYp2hd
HMyjTdrJRmysAqBJ6IkVmC2zOtcyoKn7+PNX8MlIfzwaFp0DcUDiq8MfKoJxoDEgl1Dw4ZyLokdF
uWjsg/KXhl/6BRRd9pcas+yC446MhsCWdfX28UYOpv5yEsZE/0xZtaqodW0VQrfXJkU28A/rE/pU
qWM9E28TWt/g5pw+Ju/S6/N1zBWpaeVZEZVqAv5RQ0In4/8w66Lc8LJ1F6Ri/r/+uIJrmMZTE56S
creWqCM0aU7EutlAA7MFKvkKFHhWGuupJgBnYWq/ABcBihbF3SzcDn6W3vvJneDo3Zte6sypColk
cWj0qwgORjukVN6tAMtlKVWd0p/hKPG8sd9DnjRX6bzuu++O1aOVdQWVAX0Vjt+2WwUggtgKkC8+
axc2KOm5Pitm3rff0RtgCHo8tn/ZhJfCc3wdc5gyAd78KX51whGkOH6C5J9oLBdluHyeVFpA5Te+
KM7zuEFcV3OhEJSSoVZOSHj0kXtSqofxJWITK1JtO02ru9DdjHP5+M1/+s36W52+wPd9GRNVA4bg
/svdNQLYwsgBXFDuVUY6gPFHvunGPByiqd+UPwxJd6wHiygSichA+QA8WQ435rBRMO6/S2rCuYmc
oieQPN2lQwfztBC/EvQ/IWGrGydXxOr6U3Vl7i3b6SSqQYHrWUqS26n+kxwT3CM6ds+1LjB1YyDW
i9mb7fWQC2WvI0s7+2hzZRrr11YarM2B4RjG5dBYDKzYR3AQhHei6pH2E7u1qfUiLSqfqtufYVoB
83ZqzhF6DMDJxOdyYPuhz6WYOkoQg1kdcOVmbtcGbbPHzRRseg8rTszkodHY+6ixE1SCkXrtaWVr
MnYFwilh0POU9XBBmdpTsAa9FpphLhef5GNUGPZAOWE1NQzePJ2HGo+dotZwl/EIVPWd4fRD0VqP
4kEks3I1oeI+iiAsuzKnG4F8/5fvV/ri0J7I5RsBvDM5fEKqUDrbMjBKXNcIQgPVOBIKmPGgQaf+
wF1f3nMal6Wd3yHdmQ78KBNXB4N0/JZJKvLdLCPoKGdqdWNRZmKiCNA9p//iwuXlRwytm3BvEE0Z
OryWb0iPtjETURcAPB6jbOIYM67fyO1/FOct6rhoEzNxpHk/GQc7vuVMciou3PvMWm848Ice+zP3
S4WfC8w8vtw4X4pspUuLnJhVP515GuIAZCU+j0OgR25F8fMDmjN1REgC81sDpewm0H46UB8I7VY1
kfhO5LhzO2X5sIpfPL0y5WCOSeh8qbieoAzVaay/bebKeZrQUE8Xet5f8KHBJlVnD4tH9+MrB8oK
XuYZFVfIlKmINYSV8MX2auvRyKwEitMfVxVMlda1fxJasgppwHiQztT8TTEN4xc8CpYqoKsit/1L
Rif6PgedVzvj3HjKB5W4z51dJs/osdrEuk0eulcn7SuiGnCDUyvWZx71nNEli4sSgE+3+Cn1QmNA
3eTdAQrjbOdbXlWxnk+RAwJEY5dM8dylRgwBtnN7Vxvfd7DjoEfPUZIMOzFFxeqlxnB2nW3MgYkZ
wkdXS59R/wTACeR9fLmtslmZp4wy+aWpiSZ1gvnBu2SByAcC6BjqMmuji73MStHoMFI67ZMDp7oG
ycf7NNZASRpsZuOjpBxTejw6gH9R5oTjSJO7vgcnXevy7K9CXUaynKdCNyhS+z4hzXGIxbLTUbnQ
I/IyEbsTI/bjbGGrMP9+2NDzGZJ5FImhYVmcbrSrCuk9XTDi4tAZq3+gzkGuZOdQtIg7Xd8QwWHQ
NClLrEi9usnV2CeXSuQf3qk48C+cdpyNFYqTgR00xOujrdyRTLQV1tc5LnqTM3qZVlnM6CPTPxY+
/rvpfHxMEO3qJUodDa+TvYG0EcviZEW9XIe20irHXyD5QzTeAMYeygrycu2ZsTira4YEv09LnAv6
eJolLIqRTKihvLcXd+PT+NZ2v3gsN0GDPk6AAoCxVJYTn9NwYUr1PKt8vSEDfwB4wKnQVGLOqvEZ
lK9Y/wyTPPBJ0yAfOILOHYE/+LokRc/N1DUgSqrtQwd4b//Bxz36/Q1ZxRF/6XkpceqvaWLHmJBk
QEXto9xiSIL9yfKLIjA3O1sXYAsgawWZnFD5Zn5NNUay61mvQkbZQy05aZ1uOOlLXHON0wdWPdDj
SCPBqp5KS8VCsGwmy1+YhyD9BBGDnBSeSYTjFUAh8Lr3ilSOLuiHB6Q1j9g4cUICppLv8FnYEVC8
FUTXuFFdRbOCU0TRm7Pkj4OnKeKDxcHwG/FswZFVJa5rtxDUvpztK0h1bAuQ87kzupA+dDuEBscR
nXE7gJmxqVnLXUCnXRy7uq64OZf+Js0gV2CwvvimtsUnkLIJ2j0UTGrgMAqfh+PHBC6aH9PKvFmJ
oKf0KJ8/SSp4WrKoTWLUY6mGGjz9AxLaHOD/03EkelO6OklK1F8sI/QxQZv3ewGUlAlg7vSBB6O1
+VtdnNW7r/BMGaw8OdbmvYncePx2sRLVdZw+RPLZELpfN4rGQPujiuIamBWWkINpTmjTDYBbzC5L
wm2YE2mXwI+affetk3nHeCbhABnDW2F5ozfW994mW1KmGLD6oMmQ5rGNiewN3gHqO6O1KLAPjBbB
HiHZ+tqctNVLxz5RNdgWl5UgQ9lHRUryh8YJrQq3hX3knQwtFW8MjWQzYPWsY+qcJ2K97F9xqlwH
27FIFj9BKaUAoiuJFezi3Mo76saBal63O4qO/uIErUzKNfzZzif+7jQ3tCPekrlTTyeABXCCotVD
UCknZQeu7Pov2wMoCPV+HDmGwLWwinteWNxS6d1kj2M9k24OeHCLq+K7quZFuN6qRitNX26wyOF+
Vhq7heTuYjbPL4HVJn6gpwHFoyvOBcG85UBcLpmzK+gG35yhrWyHe5jZwPKd4ysAPpbxBV4+gEV3
Pt9TrsBo/f1MoktsI5rlWpQ5qsZ5wzBRSJbawYFN/NlYPfVrzlznOqY9DH2XxqKJlbPC8y8kZYOd
oAxibDheLAHNF/ctcBvLoco82P6FnHuhgOxuUH7cNrX3Kis8507oDlElauuiS7pZhy0shl67s1uJ
tSvIzoaeTP0jswIrQFSqDzZGAvI4X+jtOAP4SJ8cpeNJI8+6JenZYLuIJZ1YysUuI9pEhOX7k7WS
wUG7CbPkPxl+klEVxy+F+O792ONHnLsDngnMn+sBL8aOERKSNalVDpdhS6Y8BSK7BBAsA6YAwOoT
lh6Oj0Uc155G5YxbVBwtdubaESH01Z5o8BWVERx6D4PDWFwgxsjox8MJbD0ggTit0918xtdcBkYP
dzQANv/qla2L5oy4ZqffCRyV+a/bsrZyXYMXkbQKAa5gScKTIuqZpMwhSIpEXin1lU0bt84o/dMH
YAWamR39TzSdNvb0pk/BP2H0hrpOasSBYId4q1iTUe9W0kwE56WN553UtP+rUSVRcBX7eQcOVY9M
Vt1lTd8Lx1yiy0My++1+63mU4bKlN5TsSSEngz4KbPnmUuZoyAIQObMTvUnSnOZm++r3imGpyfei
HRPZZKw4p2MUNJrGrSBuUA1n7F72l9hjeAri7aPkKv8aVzwJ24NuCw4+vkcxgF5RAO/DMysQLA8C
c88JQdiw02/bhHExiAShkDrsF/i0nQNPMWP+P8Zr+YAbv5HgGxWX9wbVk5cCEbaqjpExQtI6+FQ7
dhYJhahypTPU2Ynn1KlPOVJjc/XRe9uZ7ElE82SS1SQAa1EmC6Ocqv1kH3mulF3y5kBkWYdNsrgu
d4KZYrJhWopqonBBOCtUWxYllmTpVNuHuBhYuUm4k3YK5eN+Cx9nxOyYH3OdSwyvrmWz9oTmWjVT
pl5q0t8ALfc96k+LfSLcv7YR4zwKPxIeThNrQ9MBWtil57GXis/knIrTBGXawZkxpwQ8Aywnrac2
l3RgM2WLSLF2Od7PVhhOOOgo8iGe404uc6Ig/ENIpEgh5y6kYVknMrf/2875Z1s6zjr5YbfyLLp4
4CvYnE1OGAjuzIixokevFtsNrJC+YQCkPMFoie5Vy60YzyBloxlhyebEceyNmZ8aAJLmewEX8Vd9
wQiSfdLj8ON+XUIdL9uqCbTZUUwZ1hwL2HH1FVGlajxf2Y21arqj8vEYDmKrVq1guxrag6m5hxNt
0jFLErXBX/6dcAxQYnVC/DgqDUYaeaa5XACwTmumRVCpUK5vc5+DmRXUHIMnAF97PcR4DDB279j9
hij4mA18Fzi/KmLYzzOMDBc5c72Iikmb7Fmm4ifBUjl0YmoGgevrXjNLTZ085qrhxCoPkUqBcMGS
yTdJaN5IPZX9UkAdzjkL3f5/hnOfgFDsAP3r6GKCAmZhfMthG++JGun25ItpR2lXVKsTVtW5XaBf
NwRUVbaNUlJCbwifkMsIm1b3th6kzSA6GKpL1zRjRgk2YsuTLOoMbnbeHmba/4BEzeTClmraAF4U
gQqjv8EDu5JRzWUfrt/5p3AVqjJrPFZMwLLf5dwWId/qAlhIYW84/56Yo7oI+ZbdXUzJbxs5zdrD
Z/mR9vddbbinjd3zn8zgNelQb+Nb9XAHffrLoXOn8ROd6cibXTI5k3wxZ7AgavEf10OGoTP9Qcu2
ynOANaqEmZ0UpBaNL6NgU1IiJNU61jBh1u+zeqLVoC0RU5brEi0WLrup5RKUOll4g7Y4ZXgiITXu
OKCDO+ui31DdHc9iuM5SUpTPMz2FzpD/Lk8c41MHXxXveaq2LBClmi1nmoqQ4e2MSyZg3P3h+l+c
2fR7jwEkxDiZhRO+lsb9hFf19FYsICmTesUpBxIEd3ZxkrCsAKSQgfHBts8kG0ts4wR0z5fVDVAM
mFGMkjka2jFGjdmtwKGYT1ItO6K9NlZoCWr6/mnsYk1fkS5J7WFntEMMBZVqeHXnRvlus6Sa35fp
11+ZcHGJvEoRaXg+DHNAA8KEjz9kyZSql3tWcfxE0igIor/mHq86OsQQnWQTPbw+OohCQbr+aOiB
I5+BMLVCSoIAZ3BdbOcFb1PjneDMRSYO2wYg/z/vP6Zy25xGWZHUM0YBEwApYtrcx28SS+VZ7/mw
iGb9Em7cU4ZhJocNhWwF9lJX32k0HOj24KCpKlRggZMbekMACSoiKi+RUqMxyIJsxyRdVWuZDQ1V
fXjzv8idQQYjHLZCoMpjrBSzfLR4cQmbgRnqWvrNw729uK78vIK2FycIYse6j7nU0Gt/Om5ee7GU
77b8ftb1hQltqLB4A9HexZQjy+50Olx1O66qlpHEq+HQzNNaoThemZOuIrMf+23Q4mUzH2mZa9XE
nN2++4kf3hK6hQDhMPwoax0ZuWnWNdVA8sfzl/AZGZ/eKmC2irvoYN6EXXKa/V+xB1lp7ZFT+DLG
qzIicz5O7AtPz9GDCqbi+utH3IXlcivU4cmKW/eyl3cITpkT8MMxcuP+LqPiv5Vlio9wYyY97QnW
scVbIb3BMo+ymK5U8i8B6zALxI2MWjzEK9BkfpEoIuGiupnUUwC1xZ7UPZFDhIhna7PpVOvm2Jpj
xEbJZMwZ+hMCgEr6SoIlH1pIcyw2zJKwi/yEPiWud+Qn6ez0FqQKWO80ClZVMGKIh7lLUVZm8Uak
HMhzkVoo8auPtmImnwNazXOelyhYPKh/nb9DjG0v6NptEX3ER0L6IHeg9e7hMsiY3poH/F/wp5T8
B5WWaT6Zb2Q/uEfpznCjR1DT2wW7IYQ0NR1TkouGpGtfwxc2KC5zvXO8oQ9iVXRFeMyl+RkAb5hc
ZMbxh9xzcuHnEZNWdqVQoETpQVJUczc8jiZTWoqhotxg93KZJ3wYglzNQhTKx8uDJmQbIYnAWJsl
NB/VwSb5XkSmPTGzdOUf2KMNito4i7oNsfhX8svwK7duAiUcLT5FZM0sJ3poBWM21+x3Dr5g9Ffh
kWpxQ/p/qG97EZ89TOBCzDekuTVVUm91dCaOtPoSxjsSD16fDNww+6oZZJNoL0T1VzfFxhP6Cqdu
if9PQJwKTbR66jomYOIL88ZdirPmRs8e4Trt53ceiBXea5Eb0Z5hlYARqOstmOFpH5Z6dg8TVFaX
Qo74LY3wv0iDANX5BCVl/bH9Tj6AyyB3l7cZWWPTwvy4X3szz3GO5MgFVvj0a6+75W/00UCiqo5Z
gECkDX032mCWOdw4mZvTwT+ohz0b3E1A5J5+xMskcM3C6NvG8iEIBQ6DKu3dHNPZbLvHMz3FGJ8o
kbX8OOzGjsHn2iNyqixNNEq5opLeDDPVb4tPjREvMJupmK/Nstjrbt78X2ePcTytBBJUBPSmhmX7
3Xi6FKCoUaAhgJyVStGJwT9QV/yTpQUkZ7H5oj544XwmWVbCSY8++5QKIzhamzRIHDOTIZ0Zsrvj
L+xbdSFbeC8N6a7oCZxdMouezVf3pgR8KbsRyidBePh4A07j5f0prEoUPaTcW59TbxVbTpTl8IoS
RygVG8VUi4H9tGY4MJ9mU46g2uaVV/c6WEYEHDdKSCfUvowl+Ai4yDATRa995J3vA2mqmjD9Vr7Z
rCySFujxNe2x3Y9msFqGOeMHcxOR5JGxvV60wxDJZyUJUpy68ldH2idFDrQBEkODp17uc44uMQJo
r37ifPpNQyM4xWY0CFnt2HoLsrRbjaHGKAl5x0Q2vQ2kSR73e8UAdk/uyNQeJ9IHfp/McI4+XuON
BqvqIcbZewZ60o13u5msCQJ73BaeHmN4U2/2AqnbLFfsCCsHo5vjwNGmcb/D/5uKeVfC9dyVzcq0
Sqr5QhpTJ5WcuBy/cfOgcAt3SipnC5Aje8WaXwdl4swO5cuXZ2amIVqRjUvm7cjupHYpdSRiFvP8
rp+R0S+cOvlBV6HUyb+UYw5K/t042MTtgp5aKuvdaHqIOO9R+UKKV6eYFIinWAU8vhgf4G+uoCtz
0XyGxbk5wfXROwpiew/G38dmtLUejqs2EVazOhvxquAvgunOqYgltAX4viDjWotc7UDD9Xc5RHdh
YQqRQuPf5KgfkZxI8TDMdhIEk2D/0jPq0pXkUbFxCh1988d3+4m7D5Gsc0BcPVHX9R7iNLxvbNll
dWqSRQ0Tublz7lCgdITXBQ3yTD/efJcPtKr77z4k5B+6JzCqn9TiTLg38qdWVSGuHuig5Sj7XNxm
7m2WCAEE8IquPAnFAVToB+KcGjNi0BS7M67YrfLQaIdmHhzo8hbOhw1OdBH7842HHudD8JNI/wmj
UapJ6cKheYV0ILjCS5C6qGgKm9CZ12maenikR2KK/dseri9cwu57DuQcRnQ2n8ckg7NVemwh1zuu
ceJe/H541cxyVXL9XRNDSMqRyJmgt/OBri/K1AQIVVUNl2qlZHBYwB8Y1EB3qdFRCtvwh1Mu39iD
NIfypD0cLzMhEkwK/0cyniUmlInhLwZMOtfVaZgkmbpXp5Vaxtkk+c3JlfnDfz5quZ98ppscghaX
td4ZZWwXXsytFyBqql+ZFu3j1060o5UNNX11zm7WVhL3Fyq1tBY3JZv6s7sGFPItjOblaUeTbjej
lCs1IxuNcm+GspSmMSRnuQww/MIcSM3WjrlcQJZP0JoRMzR9IZ4BAG7RjbAf7lINrTMFVe+soASs
jnbErzadOMzjzZgaqn0v6hMgE98dXr7+pPXdPQ8mLCpkrOF/PjUXr46yLYLXxSs3tlnNYUH9J9bc
h3PurSdXEI5rRPhNxLDrz4ouO7I+ugo3mxrR2RJw1lPqMjbbwm1K3qp3OGhAdZ0k2yEbmcbLknJj
y03qo31Tvz4+UOex8gAxNn7TrUm1co1mxEjz/16BRHPHIu9PRCdmCg68H0V/a+84FFWnox8GJxr8
LKw1NKKdwFhqffh87QEuJn3t6iufMzxBn9J0+idJgaI0TJii1jOBhyv3lH8U/yYyYFzsvDclDIo/
kCUErZDl+g5Fl0/9RO72RW2yxW1MhTm5hysTDvwfeDmRllOktaDKFcJyGasTyd5kj96FrvCWNsw2
nyM4429j3C2oj1q3BpxSXW7GySkvU6NZ5bZhSHpgGyVSH3+K3TDLc7Fosf0srb/s8+r3NAX+Fktn
POXbR+ncsFRsxqHVico3WwtfCACnxnGWKZILGMr6kHBP8wkMyPatOsq2MvdyE8AtNKgOBNOjnox/
C6pjr3IL3EVCVQHDCex7Hwm0H4o7b3oz2SB7nz3KN+HlHOQxOSmj6cbTaDH/jytjA0jj+yXBARpn
Ezj0z190o4A05Mp66KjEKGP88AY1KRw4tka/5KbCfTbR1KoTICyBWx68Jlto/QJz4veUJx6qmJ0r
XMZwRqgRdgnmIU0aT4XbSfuXBHk3qAh6BKBg42tl4iicZX9jWQPUzJnBqmwS7nKeOOLt+VSensf/
VCw9epWvUyPOx3ajv9wDTIS9QHG+em9yg3xyY2FM6GIPyOfFY8rgUBPL5EDxwrZ1ef7atvajmL5L
gxuWfoAwmWojk7139s9VjmEkyqbTB7Tz+ICBg32ETDKA4qXk4xpDQETSNrEdT1z6EHhTJUOQ6+jm
fUE0irO/5RMPPlEQVzGxChULjwtY0ZS5W7yZ71UHirRfjY84mCgDPP7R+52HtVknt5RKP/wYGpRB
mCDEpts5qb1152c/5ruvsmTb0jB9yHEvepM/3LRVEvqldQv+Z8fToy83bYp46jyECT3KKczztrWR
NOwPWUNptJ3X2rtLS1oTRwr+83sHkPec75/r0sBBkDDuvThfePRQoiypNpjjAoA2jgfjR3OBKaPo
tzLaMOkrAAPx4Bd3SXOs5wuyvItZJr8j8fQdfRDtUvDZ83QBdpcyAUAvR2Zx99dcvGH+kJ1/PA0R
eO+rAQb+FcR4gXm76uYSB3nJOzMcG4fZjNRnZomNO/V5QC8NuHUNwuJ4rhf3uC3WPmesuexlUmJm
yr5W3soq6oo1rLACAfYnz8C+qh+S1fdApO1KD6mEIc/yannIGsKDW3b9wVCICzlT8pAGL1gFNBR7
ci/6Tmc3UdtVy3r/te0rC/6Z2ITyPRPTn7lQHO2CWtavywAK6heF1f0laWV5D/hlw2cZAlgABFHn
V88hL3Jkvp04EGaw4IdkkRxQakinaKjcXmbvquVYhqVRtefc/WNz5k8otK5/hcYfwIfEbwPid/6+
5dVzYZ0U9z4M3SujWOPm8cCMIB1eda8RH58JzgZRavqZh96wD6tpQ67gGk9hy4EdEKXNNDGIOyFw
7yFnytzPVlbfTbGoqxdiEArRQy6xViSVh/Vmzf81IFfjETMW7TiMGNaVLmCJLWmmZleYyt+g8JCQ
/MsaODuQ9/+U+xO0KDmG1prq9jtNbmcwfIhOlGXtqSim3zaeF378EXrXmCX2EFN398RhhpVapAR4
weEazuQGA+gdtEbcMK/0NbRsDwMFrxyZDhHqwwV986gvnJ6pl9PjtcEmVt/AFOf5eiDqLkZh66gu
AiMRrl0A8y6yHbDT6Ju5SeLU/d6Lpd4YnOtoKy8m0f4b79T6tTjvhFsI7CJUIkjGG7V5HYQioP0Z
nYTWQvtG8Bm3V7aQRNocnQeA7WIVt0MnNIJHbS8WIiB9M9lZoqyEw6t6fNuQxq0vM3IxrlCfphGK
Bokaehk+xQNsw5jC7H5O1iQLS5KusmIupEumFDhTlAVDUkBZh2smblQC6I3kQPXXDYNYGixBkw2g
ipT/QpTRNSy1jp3udTeJFBVsMOWdBFOaGbA826zw1iw2zB8h4B8Cg3M06N2uLOR8/JnQUM1LQOBc
l59ISJN9Q11b2GgDX8E4+ParNpkJybcwp7H9J3A3JYWm5Q49tbouwlN1inEgGkedB4pwZ3AKoHXp
CFggrJiJ9qyY03Wj/y0/wgGWVmv9jgkAUjbd7IuojKWFSmSvkWI7AtJQm1TJD6ZzWnA+kwEV+2Lb
SFW/McCHrrKcAARqsu7kdq1qC2MKqXy6iyIj9bmZgrRG9K8A0Cb6ZpecOxL/K2bafykqCQYk9X9y
Sa5TBP00rLPYSRHyqoJT58MC3MLfjSjbkfLQVsWlMu96rvOr/027PuIxTtQ+1mWy359U34oBJMQB
x6exZDEJICRsVJzS8WYUcSEQrVNb3JFJ/Ju9edCbi6cqRO+7G0nsWM887QQ+HHNh2CvVXvzVe6B9
kUqvffGur9D1ImeYH/0fP6i/am5lf46qC/IikRnhYmxumdctMgtDTm5DLAEv5y9xXSMiTG0f9WRG
oZZfo4zPh6hjZbEnCzSLNwUjwiqT8TLNusWAaz7Gb4JPHqA8yuBV5fteGzD7NAAZpRht1frYlJMU
pdR12vvokMztX9u3gVDibBDQtACuU+OjfftwlsGPoAHWT6PYRaIMz6or34A4jnWASNNdnAe8Zjbm
28glIhX/Da1wyhBl1+t39wMGsR7K0INm8YI7din4UnFp3rnZef9ks3+2wHIpPM+o1OwOrQvGbvgk
cEJd77in8poNyPdNEgX0nnz76hYkqBBKVLy/J8jlquPGXVVKcnpxvkjzoJFWClaDfVKk9eJrZMSf
ZAPM7GloL7qDAyFgCJgIezIppTi0PTb0xGCcCzP3PIWo5Ko4ifgLaBxg/9qXP18Q0K9wMAWNQC5e
mAUnIzV6QcDTWt9LFBtqKZlkcVXioAiu/RB/E8kTfqcG1CNSKnjgiByyWa+QSRdMBKrU6TgmpkjK
c/kxChs5PTZxtaxdrG1WfI0H2S966blUYADsZHKGk4nksfv+pd6hT2yFox0d/xse3og1PnGm2kdP
kTswgACTyg/F+CHW2e0dgbye2V8fxVBkjHWFQH8TAfn4JorkLsabuUx6zOy0WyIY8aoBE6Q/esz6
wkK8GjRMxGr6uxNaZwT+TXe9rM7hgUmAWH0sG1obYRbwu+P16c4hNpECODoQV1WlkA53CW0VUMPs
9lNBmIe5fA0CsXv8RUFCLVZZeNhgRuCeSdnHRkc43aK83i0YriADbGMapq+m2a8yHATAFxo2so+w
7eLfwFC0wxd/02jvl5KUikVv3bz+ncRQy0IZZYp+kvoCui3P0xg0yJaYizAxPqTQDuxDLmuvWSLv
Lafp6jiep2UZf+2ecM/Hz9fZJX3d24A2VzVnN36gcOEOPhXQw3fNzC8JReVYHejoyX6Q3TKWh31H
k9fwyXgX2Ekuobnay2y6pcb+2oTvqmSFXk7y3vkNVt5wS+qRG/u7Sr5scHPTwp+4M3g4IXi+Rf1b
VQOWL8oH7zSLcmjkT6FRlA1XC8pgv2VI+vjlaQcUlITE5u81aVNeaaToQTDiRzY2MGAW/VbxBDNM
a+xlfvOP7l3FDEJzv93svOTnD78SZgOr8eo57vZo1ETVd5Pojr958ew8Fvq3q2IDhgG1/0/JV8jI
pSznJ/YmvSuhy2EtAMq7ffnbAnW2GrwgUOPGCCV3ZyFYO+3YA6Ca8tV7A3fB++t4R/5HioRY8/PK
dOwKuqQ78rSxU/PDjFMV6hQ+6P/n+KX0f/DVBd0zEBzDYmSEf/x+tv1iHVWLV0ywAZBr9C5M24kk
w0MU9lEgbLEUEgLNzO7xfL/iNCAYthgn0fjx7mHjD8LruD6sggxUqIhv84s8tq0SwdWjwf8fyaNG
YJwRO/DX5UCLjqsJt7G7853PgfgMJkXnJWXCZAWrcK7R1nPiUjwPFotiB7jjR3e6mIT8p7IGWEUa
QIWz4kLHfD10QVhfM9Zk9r+FycZJgR/Miposel3tfEHXtETzaq9nJtHjL3HpkarJCIKer7p9Ki7v
KgDKlP48+2LgtlluoX+doreEV3XPxdrp+lSgWRDFvbgk1LbNoyMHNRvrM8aicHoW84HkSQD48NYz
U53Nm6fauR1b1h9kZVdCt9pFKV3bwRC7+x1mQoaZJ87iv6DrHopu+S6LCOZN8HbrgNKjsAbPsEvV
rp5cZ8liI4fkR5xoQ04mOCEOLLNBh/WIOfMogvPIyB301uNEknfgWu8CjgjyQddi77wxsymV5/U6
8zo553nbd4kl+Ow78DEQdhrIBmnwUuFvei+eftitC0WP0Z2OlPA4/5rBiBQ+4NpRD0H3FCcz0xd/
CQamFZ7xuIr8TuokB3cKVLzGy1gYuMuy7h8S45fF4ahr6xTkITxA8ahzDn4D9uW5d208ubHUu9Fe
PgF7J3/HxRlonuQn8Gaz6PAHIUub4BSt0nLbIivNZxz9mYN6zj+SSSWjlyuDNWWCoFXPnzVW+nS2
LVPbXyarEzq/ObN5Y6Fkv902BFvcMz3VECmytsWdUhYPP8LYv0P9+Htk74sb7H/CyEQGVVObxe01
UWWaqzus5HAvYfskIAUO/j+l2e+dpg0VyApeb+sifv35QtW7Qx8aCtP/qgDUh00cE+CoKg8oxz74
im93aYQtYnwykfH942/UNYC89xuS6WEPD5/R5bnv7iGrKjg8V38WewWJO12kvgAA/eHtcCstZpm+
cRgxtuLioAkZBSofN+mTb488Qzx/aY+iK6BAybMI6p4W9Q5h1NFc6t1YDWV/7yNVXZ2P7oN8Xxa8
0ubRW+Y9iwQd2mDqVHSju7HByIE1JfgcW3IPKNRyKngCTl2vv1paPzf4IA5URQEQqLYFxkai0AOO
A6xns5Gj1PTfa0m7u9WGhGHKbXBFBxoli/qbtgh2fdND3GZF87Ijyh620DWX/QZsVrqpYwNC1WRN
Sx5G7vsJ93RHNDSxaE0KeKOlt190H7Z0hOS37p1g1veSeng5SshKHL5bRDZwnf/teBJFL93bgvjU
a1B0+vdskJX7pAD+CCD4BNJkAJNhd0/MK+DQbcwH6nrpQUAQDGjkdHjxNXjrtzgcYampIbRAYCCV
7t3cV/Rwmdfnj529SE6aRJ2s4HlihZ7HWRpWUM2mFl293ed52ugqLU0eJA2VdLSSvnrbcd3P9i9n
70/s7jRYcC61Mn5RqLD6hpmjjIQzuCu+wML1eHO+v9FgaCLsPubpldeccizLANjdvdb7KAfpmaC5
Tmcj3zXqJtOXZMxgbK7MwekZvvvxhzdZBR1PM5WYVlGPrh0+hv5/zB62SsTGj759uNdnxhVf7Vmo
QwNqsEc+Sl5eCUi7ENoQGZnLBoSeY4ugz3eOrtIM52aCAHI7VfC/og7AoaZy7w9fllPYngBwSVqN
VZnKkek8zJWM0OyioGwGkEVhdU4DWOqkyom5+cMzQ9rpMYMxTmNgfuKU0S0+9pZWA4bsOEMCA9uQ
EaivYv/4gQjMFyRHbEbO3ubBdD50PGaetKEDY4FOXL+NDJAlRvfEN8p3Jwu51KDZ3QniFgPGm8W5
zhsisSJTESXwM2XamfVhNXOar2NMHu3O43niMoiLDXf72Oh+Lp9EBEgfO1oGBUXdElCNPXmt79fb
0aA/ChhnrIFFP03FgAADddZ89TpG/wVnUON/0LCIC6wz6ilk17/2gKiSEDmj5MjwPEyRn/aWYhgz
J6r9NwWsuki34efXmIRpQMg2mlg4Br9Jh3Vl/if261Kv0H6CcgLasyM/TapwrlNABQUlgWYc8E8p
SZQKft9CdfwtzTqt39Yxgt2/6+fWLAgN2HgvIsRxxhignsvvIjTZd3QUd9m7Oi02McGtwECDJ1Yg
626KbmH3naHFNcqEOp6l2Dg6aoK5aMlT2Ofm/GDNDMPieb+JKFMcsgalCv6OGJKRPMmUjxB6TdR4
x+mWVS/650ja3vL9eBWBhaef4xIC/prXc9i/WpTP2EeIBhULp1TAeI8DxKbDL8CbMClckOsUL8ss
5pNO6S4Z7Q9EWyVmkvzWcC1iJs3DAS37QtptIezzAe/moNrqDA4jVYSilvTajTQ26xdKIq+0Q9+1
eMI35AGqknFFVkS2KxQA1AWaOstAEcL8LHDwfF0gPvEdLaqVcnw5RGJ601n69wynbbj/4A+q/MOp
kD3QAI2kEu7vC5upcbPSov3+ex7d9f1GDuKPXp1nv9cy61YTfEo/UGeC1yAEDa0Gs499uRoJxA6k
/zJJVeWig+IKU4tTQAFtM5y/WTnMyAMXjakaazrOHRPX1YVQUIOFXtMmMi+GgLFoPgcfICRDJqLN
QytOxCaqLWPm0pWuxLq1y45loiqGE0TymfYLTLOBUkj+GFsy7Bg2KNMG+c7RDVk+ch4hq77Cx4CF
FZULPorwRUOr4hof+rxiekFwCr68aifXtF5qlez8PqMbr9I9qyUH6XsQQjNocE7Eds/CDwLItxzj
0LFu8wAUzS+ZCVAHBaw1Y9PLYMgWZMAj6UUD+HuH42tADV7TBUqX0EcxJd0Ld1AEhLclBs27R9zL
ECBLzzXkwSihA4endumFoNiW3tlB9btdnWZAsXM8BKXnZTacnlPFR0q9/5dXbkwemHjI9o4SXD26
YBKf6X5mfSNEoTWf+w9J0dVTvL4eCQKhN4/INNA4dVhys9hpqabYmuF7itIEDCOmOq97O5byaP6K
yFqFOqqryF2b//EW4syD4Ha5bxmDWUrblk1I9dXCAZDDETzjonJbMG5lAbhfi2v57o2wseq2xIDD
agiZEGXnoimsvuev+nGnu0O14C9dOAY3azJ33/X3ruMbfdPuD4v1/VwtYCUW00wTbD6XW7glu/om
X0RHCTT1UPlIE/O866jaMz5S+i+8qgNtMi5GqOMnEf/+DyAVvq413MkSxdhGEH5NyR8Mxomx7qyM
l5yE1N6cgGUPCoDrhd9xvBk6BpvuagiJSZXedwHGPzgk11weZPmJMgAM41/xwLIrAoq8+JIojIF8
cX/F0uAGHjQMQafxZMxqovq2FRRQwS2zdtuPw8/CP+DNoWHp5ItqIL88JlY6CrpKSt1bAJhDA0Z+
5IChE2e4shrigkRCZKMQUMYHf0dznGzMbqMmP1QmaVqw54imlkfQ7anX0PagrEPjO2j9camKCwVS
EsrbWhWdeeyEKEOqLmLDvlGLdfEcrFRhTFcqJAyDnTutc/NPs3XZgepPrJLYf5TlzUexYBwgLnJ1
vJA4Rg3rjlBeJ/9HKUQarFsz767c68xBICd85LCLhgLzxZXZYLr4dt5G3TieN0rLhuL4gn8/KpSX
0L/if2not8UAdfvHvB4Z4kYzpse0/0RtfsR5HBzj/zxxIDfPoxHPWk9Qc5dDgRlsFp0O3vN9XQqA
Z8VbRFCNj9HDLV254C288PTYzaWBldDx8YH0SZ2ROAeXGZtep+y7vA6USuULBo7Tf247yn4Mx5l9
L2+HOfwpWmkdjzhRvbUc3izOPCLknxVYAxTbbYt7//jpU7C8X0N3YsnB2D2lbeWMXdjYP8yaDDAH
zInGGG0ARDu+Fpi1kVAugxSr3KtIAmP0hLIGJnGWvcPNOELzHXN2s0VvEB7/VlqenGAyDsRnAt8H
15PhTk+T0jgavsSL3TnbdQoUBvjMYKa3fnbmxEADFfoTTYbijMWE+YGtPyHf9nzc0InfwShwGkjS
TppKtr8hPTcPNcpAwvruE7uYrpoisH46x80ARLWThQzTGjXEVAm76V6YVtf19XNX0iM76ZzMYTQZ
VutvLPXbBDfqwvNcj+hPvrBsCJbFcPw0EKjkvXDIpw/cemtDocmvkdT+d8eUW6NUmCsDlw7313hA
B9Cqt4P6qDB5nBzunVSMMZKSKbHcthB8UNzJro1VeRbY5ZjH7dzBlzvsvv6KrhkJS7DwbfTTsKGS
Bpp+80az9Xn9cAOh+BL3exkc4SmKITqiYAW3og+XboMxbVi5VKpvu6nN0jQXTwP1djxwTp+krc1E
rDZBLQp6RuFiR7Dj2qsN9VTTI+aur5DQwMkPrYb7Jd6b6KECPJ3rdTWPndR/AajeviISQD4SMMhn
FIdywG0RpliidpQAHtRExr1DcC0ghbGwWDfU3rNeFEdyCs6+koMHlEZvQ9kstej8fVQWaRx1fdLg
9GuY0ROhLtGQsqFllc1VChPNTff7+DASoTFH6Fdzo/cR3Mu9xI6V2txgMEsccCCmyW9IUps4v7v+
cIkx14zrVwVKqAF4JfFJ3/Es+tieVM8/vNHaGrTPAiuo+ACijVHU52aX0Yu6kUOmV4ByOCzyHnJq
D7nDNSz3Jp1vlGGHE4aEpr6DdcnAyRQ41gqAxrH55IdS0NqonBaZc4RslR/9e8Q98risKEW3SjQ3
c2CXk0iVDPYfURQYH3rb1MO2r0FC1mQ5QiWpbw4TMvbLWXwNBQisWhkCexA9LbCmjemqemYJqqbP
lUnHFaBJe8wIkuMw6OhX0nx+fdjrLlrjs1L5teOyAjRjgpGZZbvFHpDzBGiru2R5/m0ekwvXmMvD
Ecru+QV1hIPbSZe6YTpTJmz0ll7qLtz0iQZhep3Pq4tplfrqTLaY7JHfHwBLtVdLLM3kZ3NW78mi
itNiJcXKQhe9LJMa8smjjRJkrVU6QvC/iddnq9l/A5rJNSfjp8pYa0UpXak6ahN07v1pPZeCPiEm
faw7d+eBj5d3VgbqTk/Nx2ghiv0hXhhtwaS+uksCXByAuX34CCSBcHefv/B/gkQPkeoS2rlzf2Tg
gbkyAE2rEjQ2LJ71lWrtwr3WO8B5x5CEfWo7NQpo7obBtL6D/A2SZuILHBQU9lGAKCSTT7VcYuq/
EtyDFLBSgOKFNA8oBDkmI600qNqQKktrvjCyJcnrQaDjXyh1Js3cvXWTGYV5Bd21WCpvv5/ggg44
tlZk5wdobyAqlRjM14gydIT/tMLQzr4cOmLoeYQ2M1PdORZnwm2xFJU+Rxs2jTd7YvGdbL28zlhK
IFoMuB8kYGMBCBJ1vXjWGI+3NusiHXC38LxVYV3W5Zs8OZrwKVlP+JmwV9QkQXNu+lHq5I2JQgGN
3HSP203O8UM5tviQQxijz21sfev2eAZua+mW1BEu7CDIBfXyZbZBUdRBAacUVCI36VzhpwH1Ecfy
mqAHfRsSEV6oSofilV345AF5neXXS/jupM/Z2jcnpLU1nce2W3Ge06Zyq8YV7D46FHPUnZhtsyP9
UBcZRS1v4+m9o8Ft3UILMhkt5jY+fmYo8lSDXjNAIus0dE7ybFQACrRy5h6dzy5+LAMcI+KYKUcD
ddI2/WswPOBR+S0uBN0MCRE5NDA80H6kW5PfooE9b3+8AZ5lsXnzCLw4dPDOGiIIj3tXIaVt/8/L
G6ZfToh1fUAPvMkLsVlFA0vFAO+c2IP1CFlUb4w+IxYvHRETE8zjEOPADQadUPNMhlYFSTSiV2IO
cjprZ4+O+ToNs5WuDu/23szZ/ali2eEwAxvKSF+DwBytco/vjNxcFkiMCW03Rh46AGNfw4mV8Gk4
LxI2agGPaDOWvRpw7m8lXSAeLAtsX54ciSkp/popTNO+5Hh6Ia+/yZBwiXcTbPdAoo/0uUPRDO3C
JwVzKt4UHFlFiRuAQ9pZ4IiOYYYSPNmcRNPpUVoLXxGx7OrUM4BLJ31sYtEB6Ha5W6Gcxrcmxx5J
r709i8j1ifedRqE2HDKbZ0G0sfxy7+7fMXuEtZOYU97SMaCvuLznY5yDq7TGNUXIvvcJZk4D+trF
nMGE4N/qnOg258mVlzy24u7MoW0AHWAanDWzQ3EJYjcf/AbjuVt5K/vHKyZeoPtlI78v/inwxicq
IaJvSltW/Mu4BKq5wH+9bGCLIizrHAxd1BKUeupB4mDNEmj0TZAUPro7T70j0jp1HBFZVn++we3b
X8myGJKTMnMpAjBJTTO8hRTiealOFLewNOMLk40OIBlx3J/4ElMyOTLWnGDixz8xGzxH/ENrATJ4
UScM13yX04PciloTffAzH45AGtVzSb1uV4Q8w64H3maQBBpTY7V0sgzRJZfGHQtR1CewXnbZGNyM
thtF8/EPcot2jqJq4KuCrJh2XNX4ybfoKHqcC5U/0WG4zBll6OQ1eENQvDrOVZoeZvs9at/j5xP+
VpMinzp83ECji96QA8UbloSnlxh872TEFm8xQWVeaKFThOIAXD/lDsjbNJo+OGuZH+UIQ8XKw456
mhriE0tQ4ZuTwh0kdAZ85UZ2mgrrtLL+1ZzUajxVgRGjW0IbZoHy1tSHg9cytooLFeLc+Hb6Z9fc
1RZy5hiLnsxikfwBYRzGi1c3WdaX4/fSxvYdurP9WzcQtbawwUBM/NM/sFRmhDkvae107TbGWhFB
vtHbCzJv89T2CE4maII4ravR1QqBtkLiEum0NlaPhH4wz0XN++5dANtcmBDeAoiRRqz4yqKbxvtW
/5hT7Yo5NrgAZgBEd+rTmvxhkqDlW8shGaW2sHffcX5l/UdBZ4TrsrRlFUG1+BX3+bOWR2gtUAiP
B8bWPcjJZb/zkQvoKgH2AHdvyj5brEAsmLb/IHoNtozuFpUG2msIToXNCcQn9NJW3X2XqWXon3pg
Yca20v2oNgSZKjeoQzb0CtJt8DpSPptYxL16AF67mQ/tWYcuy3brFWh6VaXowoJN3XsTbVQxITi0
J1c+P6RWnrNLtfUEvaVh6qWZvA5Dbj+szZajBHMatXRkfKAM9vN8mYb8SR9pkqUuDDRVohuSpOlB
d3Up7pYsSV8W1Z0nL5vpfyOWAnUM9cjvtODAoT0ZRW+AHJyC9xQWOK3v3onLju6qWR7wAI1xEOe3
l+SO78w24uX0tw/xvYI2Go95JroLjpeSoVRgYzKbAdyiToRkoKyeqibf3FAQSRu+QSPu92rmLDLl
7guTi6oCfvma5XWa0H7Nh7g39/OzjkQrwNjgmrVZh5lmh6AXtZR0fsfTJtnOIgBg8aPW1cijMIGn
9jOOE5GJr174DRXHUwxKB3oXjf5iFrrQBhyyTTinaRWZqoF48QRUc23mz16sMusyudQQmbQOGl1Z
SsrNXFhxnmbHLu6JPIl23vJkpvNtcu1isJpsxhr8wDxVBN4SvnKjS1KOtOc1cGOxHRLLio3pKFEh
XSOCjwfRgYb9TP5YwL1jGAZCLY5D/XFtk/CeYm32oZaYxn+SyDxumBJaVvwKljsGmJE3eVCaY0VD
Cuky8yknnC16d2X5ncZzgY9GCOdOLZOx1gnuXCDONRUE8FGKBdfbY2J4n/BIavcwUsV1RqoSmCMs
M6nQi8SMyMKwCB8EWjnEPNavBoo0+OrXShVFBxOz0Zk+se9DKIN78zHLVsJg/HX8QWGlZRzzNGm+
0gKJNGotM9fuzWdu2XyB/PpWLWKtHn1IbJcM6l0Xk5nTnl1s74Qcy67Ufz0n1BZN17fcDeZIZjP+
QTQA1T1Vb7ko9g+EofmQeUMl4RNWdJQ71mzKRyUF9taDtoFhfrqe/1O02U1J1JdcQWlMcHO6TyX3
1F/Cc/9ChO+E9CyKMxR14jAslclgT6xzMSkj4qNfiW1Y1+vlY8VJnvAZVZPGvmcEmQS9pspQxQMu
0t373GLHKlEilurm4Sr+4/F+lGHZQtFBW/DIMXGvmk6uNcdQwf21DldO/3pqVr6/wF8H1le73Vp1
384ZV/P4R5c7j8c+wS/Ll52zgwwk1m75oJsYTf0btpO8VQw4x1D3X+qlOPQCyvV8uTSyxOxbLwut
7WxiPojmFeOYikHXk7x8LNKUgXWmRfDllUNIX1hMynxCEMEpnkiyYP8ZWjqzhm1RuN4+fkHCxtlw
PwSyymqT9pfGiLOGW3m3kf6Eto7eCDgFYP/l4kUHxQFp1XSFh55ikd3pCZ9vndtmLq6+SSvNvKpu
UgTDm8JHGTRZhVv2c9cG9lcDC1Au9k0EkU49Jwr2xooQY6I/K8USQxZ2eFXFho09SDan3zidzKVs
tXkhJ3rfZ0UvdHuPCwaL7ahiejH+wWEnFUXsMLYjmNs0V6J6G0Mp/0xcSpTOSH+ZZuHFPxG8/xcC
Hu9xP86iLcCtfNe8wNcBTHmuqp1UP1P7rgphfKLr04tiv85Mz7oEXbGGUYh6TGdVNXlOaKFuQpW5
bZZYP9mPu5MBJDAAaED0hl2ckHRE3e/WSN/QEHb6z/ENhTwpItgrOVmrJ3gJBdQpr2arzYhtI4YA
qKqgdypaBNunEIDkaTmYSB5XugDAUvrtMMBTF4OXTiQsPwjpf0FgGGqCmgYE8lRYUAW1JhsnCvH0
LOUwQlDYy2BZKjXco3ci2BO7G9ezODlCvgmpnJAqhWAK89QlV3xfwHXRPc8FJrWzA2atMHTrP3nY
YMVdFifLKGrBVCdW1x0fZxl0kb62+pW0o1XmQsXNashQZ23kbSzaZ0HQ+MEsyAXVAe9KqqD94Mot
2jnFNeuY+ccp62vk09gtE00wF7tsUp+4HO+3il78eIS4Ah5rLqf4tU+l5sa1u4zG+3VUSrjH9jYF
DzftPcaKZatjBZ8CzQQ0lxBH/zbfMn3NctOOLbd/aPeRQFlx/cn73xPdh6ELv67L/kTojuDXo496
vf3ZFsEBR+Ku99PObBbgsIJa7fS/fqx31IjnnolY72RGMK46u3sSH4oeMvwKQtoiZWdzBQ81f5iC
J2a8pRt5kJ/9wgKibPzLh+QsdOp7MIsAGIp++vsWFb5dHAHPnPAKJvmwmWyrIs97PGmL+vRqwPtX
oHPuL0Q3tMeO+hVqRo+IZ+/JpHz1r05kHekSY8cpq3fgD2WiHa1ceK7sNjaYtq95U6D9F/F1CQxV
Ka+QiRXNcxHcTrkqx9LlsH+pUNKGSHO/DxvboKtySBdrNYJDY0kpvf9JSNQ+wDB4ik91EGhTQoeR
wPzziOEzCrSWQknTLM7uFJqNw6bpvA64eHDHLU4G8JvT7OhQwNDrMuNJnBunO15Hptn4ED5mHtZ/
fGDQws3mUteCMDczSCqA1ovDI+IfIkOwsT6ATDf+gMSb7Wn6rn8172A99oU/+X51s7I2c2d7DczN
XKWLiL1wldryIxRAvlwLeI/FS7EgaYXu3s95FvSF2vRkaawax1oxdglLoHkU7ODDbvW3Tn2FVAXW
pAHzHly2jJe9xErgrmI5Wrkj5QV1CGhOe5wmB5IsRF5f+zeBW05MoujmT9p3HXhqsrKE+oV1cXwj
gE5fgQmy7WUtyggsx/Qjj3eoGs5pgz8GwW6g80PSGeiHWj8JPgNlUk+9tcwki98S00c/cARgzzjY
yKv0vkMCtpVFNaHcnJ/LuA6DNo4zqMk78nRwHd2D74A4ZUynS8mltkW2ij0fYVHdBHbfRZVD05+2
f8Y48XgivDxgU2bSmwNuLQsHBOcN/6MS+KORw/9vT0bDztgtmMEmbTrp1LHTJgT3LVSJ6docg0Uu
R420BARD5+SeG1QNSKz4WpAZ5+l7ZkfQXWrnhkF7VKnE7VfYy5PFmwvMc4F6k3wj0Q055KFOOlpI
v0AhvArCQaE+N8jeg69hHsI1MRpcYpsl8G7cQaqOPHw+yGU/eDQrf/RAURYZbcDVWUw55DtbUhnk
pbxelunXvxPF1FViagF2rRl3X1OX29xVvSxmNIWjHGWSyihU+DNCTnObG1ji8s0PDwhmRFd1ty6t
hADITVDLRJv7vfVKsazU95a9bP/Qt6B+BjBl18wjoAsfU6O2PIyfjHS6XMxEJIZLU7NzBv44MulK
ydzPTEYWcwFDjKuI/55OHpAsXqaUgE/h13LFphdDa7fld11eqN42ffCy8dc45UAGIs7kOAdyLfGm
iKfj8R06eo6MpRb0UNkM7AwCu7+SnKwvSaK8lih44SL08DhHzozA520XzHbJKuvx85WxInUFOfew
DoEgb/3Dak8i8DgtiKUuF44DVGUFeJHuqL8FZx5fD5Hhaa0Xju9z01qcAVxUfm6LcWPkutJ+xNGv
JCbyOeC53c3nmEAuG71o4QItltf3WPMnmvAeVtr8EgTrHZB7xfyW/WG998txfsDh8luB4FapGCWo
U2KcM4kSJda0VuktG9rO9Cv2H6idBHtgojxLNjJ38Gi3ptDl20aeyAIG+XJJ01+GM0VPvG0sdwoY
oK37/fXr82pQerhm9NlxXkpXlAg4BmJOleq8a4EsGjll6UvBFB/MXTwiI5mBbf5jhhG/wCbLHUrL
LGjnPkJHUI2PreCgSUl9/U1M7cYyZSbssQhNCSzlqL+6lFsezKTcrmXcHJCvk9p2ESt/OJhmqNGF
eB1y1JJOwMhWy2lzWbnNVhBj04ChrbKtE5j5rl1SPYX5kuIUHM4AN8hKCwkn/nvwyrKSMT4i8ZkK
g4gF5OfhWnTUN+QvS1BqXYaKpHVGrhi5V1vpUxhONFihFJPw0M0gsy4UD80bZjJAdGrMhoN786Aq
+idJ/s6zLrervivE/MmO+66c5TOINKRi7IapwGfOuQd2du+NiL4iEv4TnOYtpfAc4J+wsvUlDc22
i/7DANfJpj5p9pvPj2mYiia9gOaqvVjbfIg9/r5u9aksPCgEP6HM0Er/1AD0G1YQ462tGMOlYCh9
fIJZ1ZFRaeGWBS9eDc8YOZ00zsm2OTezPbSrwkMDIGUJ0woKxMYGR9pK77MsIwkmCgZSPC6KVt2S
1qt/qZsrup3b0jRsOkNuzbH6JLdbL9gaQ+BL3LKv6Jkivrpf0j5c7D1V5/YH1WZrisTJccs85w6N
D1DChIY17H5sRqV3CLervswo2U9WLFcMIcbgBKiVCsMY+LmHHYXaMZ7xjJPGVKTY5fbWkpBUyVVl
GX4xB4SK8KKcC2mK1idB4xDV2XFRukZ1QVpGI3JQKDhjCvoQZwPuMGQ2IuVbWBoBp677HPRAwWaU
124MwOLm7zXzt9MhIyx1q6vbyVy1CreQkfvuHCHXzNP+Jp7obPDaH8GWeqiSaDvuP9j45Uh0yczh
ceN23u4/5wxlpHC5AhUcAEwshlspfofJ4MTEEdEqxrab8iJTLip06k9uL2qoXwia0KyZM10T2KIY
TNXwETXSxU6xa17z7cU1FCzx1VvX21+SLk4YBFpMjfrGMIYSx1Y6sESt54ikf/wAv4v/l/hK3i9i
h3EwhI2WLFdJxeZ1FSr9EzR8eT9QMC5E63JWPPhpAo6JAJc7xgFhYRR3jmiB03dWJ1FQlwMHeKxD
7ie4mF8S0NGPSbltYKmwPnJORxGPAH45sE31s8LrFM3jAKOfFL2PyTPZO0txr2iB0/WdqWhkeQsz
3vtm7E9I6ADq7oerey/8ibQCLB7lHqQrXRk0hbzf+cl+whXoO53wOlGIuZ54H751UeuIldntfS7Q
pOW+ili7UnImvOvaIUxgB4GCIVhG2qPLSCRhkAERjUvmVZOA0QCc67XMqQuzfxkViytf5AGRUf37
I/bngIx29QptiouRQxogNMIEAFmboXf7RE6XVXuNZUjdt/rZFmu9pkCLr+hiDJoaN2EM/bPVvzUF
F9s2UTLUa2uXo1F3ehkbe6vUFx5HauIrAE48mfAQ8Q/amtN1k9j/6ql8hiBMRobPr8DHU9pMjr2q
LaPGV4OY9Ylh+ICE2SyWvsvqCqdRYEciBHCzm6/4Ye3qQ8LSR6bTC6tdge7sjX4u+bdZBiROk1NG
/NLOw3zqFn1xUiRTDwzc1EJg6loupMcGhHdZ3UhsBm/DFkPuazgGuPoX5i1uHytl8TdNh18A7JTr
WxT/a93lAGMD2rLY1VBSqWUpDeCiwtw9QELb7kLXws/yjydF8H3WVK8P4gfsiVpKJkovG1Tc0eDa
K2dkza4CYyX84ow0iAYHZ5ZwoImV//ohnlF89WuZRSY9wP0YRDK058YjQMY8nzCnyVDSsuzzXlHF
ZhugPAHMRVznJCz6YBs5bHOZeyMj+SlYI+5Z/Orj8V6vzQAp6+E+AovCVbp6bbT8o+cw0rKKBJcG
pug1BVIhQsHm+tJyGH0/Z9PYH+VH8c40M8sCibs7TGU/9ApykfFn4wbxGv+ks8hZjpo5w4Tj+1sA
MBG904inh9+f8rme8U17P+4ess/YxBZH/VZmeY8wxJ2nJ92To9gtTp4fOaZ6gtdl/J7UhqBhbSi7
uLCXT0Rk+n/Gw82sxC5FX99U/1WoMGn5nSEI7o/kxpTWs2LL8OBpvesmQKdWDtfAqJUPzX0MR8fP
lFxmlLNX5vxmI4ZQS1Jx5k+2GWsgIqGC5PtWp1w9mImQi2nruutatDPkBbXnmoeK5OT9Ikv1aWl1
K2g1V4PM1TOyf1O7VKybFaFCiva/ZPi4FewILnKBu3S8/YiaBYHFYR6MOlttb6aLq79SmNmfAuay
YiieXsI/sctAn9Fc44Xs51WDfKElWfVmq4AJk5KvlLAm9TR4hFNRt84E+VPEZtQppQE4PjeCVn50
Proferpg8Fe9Tu/+eTjeASix2q7sav9L4uafBKs889H5lMGbVI0JKFAD1c7v5v6jKOiQSkun6GCM
5OwUtblzsJJODcBZa28BhECnnjWb+N2OA5mqCOfXLLbcR0RwnvjuHhJAiTqV1Q5Il36brkW4KDm5
GBdX0JVdCKBqfc6txAa29w3eqFuQr+xnOg5Bvoz8imY+aXAFEq3/5niqq/GURXJ1jTjVskD/OaqG
/8/IpNBiFryycA8tIF2D0EwUSSjBz4V7uZxmlI0RNsTm5jU6LO+9XYdQDjblphZTM+OLcfjEI5Hx
87cxXN6OgvQhCXuxk+vxkf6KFKHs/U3aU/1GIbY5qtr5tMQGiTL9qcu0PmJKGKuFHgo8xehouvZQ
4Gwn5iFRZMFgmoLVxKfvwGDkL3ODGnvfl1ofhqqZezOB1RcLgw1pSe03QhXvEJnFzuNjzvXUZ5mk
tK5p+4eeAN5sAIB2pyN4l7RCX1o8k3+mOnvpsF9Q24Hnc6h5NfJJPTDEZ4A72aQWFudnbNhONIj0
HzjaHwdktirYZHAjniVjbmyjpZ8XiqTciOwhZt25l7XKeA0fXGc6P20zC1XiduD3kPofmRo8z4TQ
WBQFOxfTv69Z1L72jXPL0R125m2LG4lBhGjLq0946FfUg7JJKsMxADAuTtIRobyB24177+fhAq6R
1Ge2gzTSWIKwu2bPl4MXlvVHtT/1lQ3C9HywPaUwearpTfcrxwxzPShrFiY1ugzu9e9PA43o+0Tg
RTICRSszPStm7sAb0ojEFxp/krbndbAJRDn/r3gMHr7hSkxxLpjx2yXj3Ng2VMDYUEJRBwyUEHYM
lPAMIzLwT1f1kbFIJcImUDhO3oo0O0HoqyyMFvNk4MpBjHOdFoHTdh2TYljELlj24XTHeAHyyORx
6djAt/rHxhx7exo/MZ4TeBpZIh4o55vgnGcPmfzh7we6EmmZWuaLSbVP39T3NQZd/4u7yYwL52/H
WDl/qur3Wmcbj7q9dOwU/qxp3rjGxY6wywGc4nypYEIK9lLr3QMwfz/gXIgyTHnXZbpQsidYaM/M
dP2AMZ95Oh/saDsbVeFxQO8Pd/kb9oUwyUKAg1AqjiJAtiOLSuwblDSSA7Hs2Cm7eemsiy3v9MdH
16oEfQuAOFil9B0Whmh24EX5qiwWrqrL/+e6vOAeNb3HNFgLU27TZV+HUl0RncBNxfGKGp2k0EC2
BCu3R5si4aiKuO/R2JLEdVMrs9jud+JAiG7tgfGpuYUKTTOF9rwhmwMk4jDOYqFhOF90hiQvOStL
NptQvkItQFdcZaYamOUyAaE7ZrARcaW2eOOhOiMdSRcR6LGdkmX8F0IVMekpWySwt9CwYc6zAWgx
lT7sR9+gQCMEd2FPVJMrXHA6d+mo62OmEIP5d6Ic4yqg6iL3Ba64B8bXau1K/G0sxCD7+DaHpS27
ZKMm2roG5AlDF7QhK7kS1uP0p/onRg5EkRVa2iPJnE2qOU6+lYkDio1xPfl0m3qwXA4zewiqujDm
u2P3inu67SkV8h5VPJ7fneg28vvRwLx0iRlWuPYT2ADl8E86BXIPuIvWkvCQHPOu4di1txAsXB+f
U1l9aWd0HPPndkrwT4OdfFNzEj4SwEtV4qZo/oLmI0qqexlcUWBmXy0fH3LikTjzour9PntyAy2J
GZPoc6IlqXXn6723aqUx+hu085phiqwVCWgn1bgTWvdMRbNTRf8/VP1YpO+366vxzl/hYLqnwz37
k4fulmSvP4/8TULtZH1eHO6Owpot2CDjBsnc/7RXVz26wFckk78oEntD5zP9NZQu6j49+AhMvwqe
Adj38sCdjcrUZvzuQzhZrDXbIMdz9i44TehFsPsZIbZZaDRb3jARQdQ4iVfESpgWezPJR0IWh75f
sOs2+mRIST3dww9Liap+vNG/4moAXwjf5+VSM3ebzsV+8W5KIpkIH8fRoYG7Fh3Al2jRQyVhqLzC
rPKxR8qHevDOP6ccYOaXCT4ZlYBDd8N7fcpjzewj6+uhopsK1R/BFkiEpWLYK9kIC2+Xhzv2RsGg
Y6pwXb3u3vYU5oXGfnMmunfBt0Sw8U4eUySEetdAHIxBFT/B6TfdvKTHHW89wKALXfXz72h2GQyp
/MWk6QWLtbQ7rmq8kYIS3DWGIYJQEvi1E+bu31OdM6f58lSlaccCq0yOeA8+BhEABz8kyYtiLf1a
hRxuBP00rM9CryyWR0FVXYxpPK8qiEOjwcTppZrr8ct2qCSdazqVeUs8qRT+tCww5tn+k+5/vy3d
G1Lc0lxKw84X/OPMLyFMuoSDg5KHt30Grjjj6l7HWZtvrkLq/pURj+UkCXx2qpC2uxARxsZ7/35y
lXRoRT0J8ETH+yZUStw3f/VrM/8bfSWw6Ky9HYeLfAOa7mzjjS303JRFzqrzq0QcsmGZV+AmtgZB
29jDnfRx9zqXQHntNmve/f31foGA0JW54qqrzInUWWYZ9/TyENR/vwlMOyCXpQBhjPTqhXJBnGqa
LK8Hd/yrq9PxsQml9CszVnBY9yAYIfTBYZs63h02OuEskKCaawhWLcfOC5kk4Ki4uMW9fNIfvS3e
SPA6GhWAX4n9b1GCk3z+bQNx0a9XiwOOGvEAFPjEcxQSgwwVAgDt4E5rvKQZeFnUbmpYi/ri8OZz
2VKrAX8anFqQa3DNnMqwdAFjKf5CQXmgEslA5O6RvA4ZQdorINcqT2MQzpbV+EDarLlic21jv2LT
UJaQMEk8OQPhTODTbDPKOxPdTX1uXJLM7aeXxGQSTAz4i0KONyLquwwZeWPRNfApGGr4yfQA3pKE
nWd4Jc0/yxgwUZKPNO3hEc3V+9kgaRI5B17H7791NXStb3XAdIkMsxO81V2H77tXTojPQIcgvTRN
PDuMZS2UCE/ROQ5mKmgBFI8wKc76QUYNQo0nBlHSc3GDqiUAPxTBXlC2Lb381KSrOP30JDs7q0iL
ImigrV8eiEc/1FpQWr801nCj2YUCYcOGtswAnQwZO1QdSuNv3FDXzzW1ZNe6EUvOxraqPnh5t8kE
UboE75sxnMYRSvC99JC3cOJploVSMR4ezlyxjn6q8TBY0oJEuXKEXNbo9vsldNGKrP6gm3I71XkG
gseazSypGN/gGnzBJ0YrsUDgfXT9wiEOvIu2uFbG47SDUMIjTRIbHBe5OgMkEDINnKg/MEOiGwmF
tsgoLN76wzQOflxF0v4Nz/r6KGDoAOOU5Td+peHgqiBxHZH6Pxv+Fbis04BMOH5XxC7yoxDb5osc
X1E+as20V3TEPvhRYgXxruQ15g9o/wTg2U3LKoGs4/4ACzbzpREuWmlqH7KXvEuqakVz31lu90+0
Eko+gI25qHbXWoo7Em+GwGLZNktdB477KuwSxkBZBZmgWhlufrLJitXQVRdKHUmkWzioFi7FCzy5
wbqH0fmw14LBbeyWVVm+f9A4bj96Mii+vyJ1dENGgyKQFSMNP9h3DQdS029x+omt6+ueB/kzLsZp
FzKDdxlq9rfSQ5bEuoJ05xhG0G9GMBkt14/7fAxM8oHo2e9F/0qg4FIpeYMtSLw0z1GEbkHZu98B
qtIywWkUQA5Ap/Ua404Rwq6T+ndSo2+385Fzid/1KJsZTw1oVpY81gmdiAhYUv6/QCALCPUawNL9
xoAUWD7xqq5Zc0SZyExJy2z2C4eanhO/VnXBKq1BzknNCfH7LVOUIoVHAqDyQOAgzTtzkFs78URm
bR1LdeDf3O+zpVklcEPw4tOJ2Lmhs/bxXiKTSBZRFwBGBK59b612Ze9EdHzTSl1uPwUTNlKvIX6m
GpWKOeS7l81vgTdoys4FI8MmetXwb0RXbvH7XZl7V51kLZt1QQzieBqM6oXosNfuuoEG0n1tPwpd
1zjtVK4tnZD5XrLmed6wXGxTCStYKho/lznde29X1sCFpyXCSMiQgw9mHMaZ5y2lsUW0h5JgfXYQ
CvWa4dbJi/QwLUBJ5nP77dIlBJHUDUEEypgAFGSpkRShEyyLHMzja5d//BenCs3mtp7Rnm270VQ7
RHKi9fdHVfNNbqg17sSBNkGHiJo+7b5B/Q7aZ5TFYpaYuIbrYkzprO9R8Biq8GwisKredP/2c1E0
VW08yMHX60xc5gmvoJJmEEQ8LpvXXJFh5AuK5qSM4XWUbl3/GMcZV3O5yJu8pr7cECITCBIu2sIH
HCDueFwZFZaxJUJ39RIRDFkASIHpCfhtfooYomgxUPZgzqnvsLJhVN2i9W5mtd6cPGcIWCQ8owX5
ATpHmBwBcGyCJ2hACjNDvvlifFuzCk3VSByhlAIJB1O56U18D8kpLxFMbmdAocosj1Sy1PLsCP3X
J73kUoDqHokT4a8y5v2kHczFLTyobeMtJ1eJvVteRcMRjWot2OlKmJa9qvrOlMEMJWBdDLRnimrn
BUbNItUmuy6rBuTq2Weus95e6cg7w3adAbtKKeX0iFW9Do+L0x+Un0wwb2HKdg8qDteM7v60NekR
h9u7dbi8G6UzP8y2sXalmw2e/Utd4wl5l7jURyMi8XQxUmheTWKLmhGNKjMD/1tJyur1MqPYBTdB
Axt7my6W3vkTtMonMukILlCzrVwLwGAnUqHllxgQRKhdPOfnWAnM5lNfVFByBm03C9ZEcI1qI8Je
Q5dSBW/3aAFGo20rbxudh+HNH7l+FXad6z9c25+SfF9U6/haLDqpuzHnXgFz8GHS2xsMrrwjVs+l
64R2eBf9Lcpj2yq7HQflxn7YHk+sHI7JLNlx7Ho9aigGQ2yE5rOrhyWqQ+bD1qSivoBa1k/+krSu
UXc9XttCJd+xGvUD8Ywovm2R5ERrKKXoEuab+fahwL8AtGTBYRCFkL50pPkxUl496nuaL6lKNnlz
YrCCfhxDKejMtigYxoBALYnG2C6hRQVmXN60c6bahU03nyl3E6ZGICoRb/7oOOpqSPldumBeRdbj
+PUhtH6DAF8OPxEN0v6CwFERJBvXzzm11bu89vyuw5GfIKh1HNNvknI+ixmG8RvbZqv2wxU6lZTp
OAGMIWYC5klNYVQSk3iz0dTLAfLxQyFp/pJHTTWiXzjO+7LOVL0+KPEDpUvn3IL78R617+31EPU5
yMRv7mPVhj9i8iQF5TdPJFasmgogqsr239g+sKelvbr5NOurIPxwEc2zgeqqmu5b4SCX0W1QbAyi
9aXdmXxrZ6aj8ENB8Br7g7hEQhUKkx0/Zej+5J3DK/Y+ibMno6yOHgHVNCdAIfOnKD67kgp58vZL
rvP7IILUwy3Y/0v5E9PAscP2WqC8sOgYOD40xa3LgLdGemPIGsCwn9zMfmuy8nBjW4inGpkKVkCj
7u0PtncfvRf43QEXisRmP/+cRElK+RVTasDTyRqH/qMgpz9qAjY+dyVlC9m47GnHz0wrwFAvj1pZ
5ANyLIeSzHMwgNXNQlHUjQraiX09PTbpMD1CfHV5RDtPrvoDe+Zrp77l6PrmYSNdoz6vM69LOH8X
rQo5/caRVyUqPwjA8D6WRHDGpwZ9rY4jDB8WHpOkQ9/e0k7aK8KSW6JqhTP2f1nEWjhJYojJyFyD
F3cqFp6ptlv3PcM9zkMATHvD5ocEZWT1If+Yet03QLEZ81AYzowFd2k90bbAMEh+jjSG0D6UFH49
cpYMpfZWJuMDxLJ0SNWzP+BgJfMYdEWG1zR/Qrgqg98D1pNpo/fBZfiHIuNOMYSbq/VJEF3c7d4g
PaiAJzlijfxTfW9Lg8PP8ODNKwtP8+cAVC9FZrDnsMOlJVRXZoFpIM3AjleaN43SLiyvL9mIZzm3
8cZKH5Pg6oCks+2qBbNANPlu9RxIyVaSBrhPNv2shuNpugeMUFuroKIejTVq/uFQ0TgQap4kLZPO
bTJry4/bCxEkEoNmyK2W1UQ0cMARaI6z+KasQ/dDgTcIfbi8s+f3T/m+d2+GRsnQKt1/Fs7PAIdC
fkoNxcDxOapwEMNVUny44UkdMAP+hzix8wts5ERypSlL0NkKZ2ql/KsfeRgH5hvjphl4PuPHf/2F
d8/QN3p51EBu4a1YEgVX8dskaAzhJrK9fWaSP8nmECvKRM5NvfqXH300HoZuZCgKR3Zy8gyzU6TO
C8zwozkrjIHLl64wh2bQ9Ac8RdGeQYXlCgnbuIoHw+g4vG9Q4t0l7u9aUHKoL5WeZlCJewjFuhnz
vn0G8avEIocY0grozM/bAQ0uzT3h7+KK6baKmtGy59mgZoEr1IUq4wBjiswJbH7hPBAUpcJ2fLz+
DXSqDO4rdAsqazIuoXp7IU+i1gVVHDma/qq6DhljDI1nDnTmRuo+y4r/fqlhMenwpsMHlJg0lZkz
ks3C6kNp+Dvg/UDfz196r4gqd2+bQ5ejjOSuFR/j0sAdNNOKYxR53m7buYjooF94wircv0pAP1O6
meGNaK1ay4kfIUai4l4G1hfHkKv4NzUto1ae90otsmYHX67qvvO6CYBf8rhVOA/iSym2op9dd20z
pOCFCqHuuUPq6cK8ouMlsg7UAu8ffofeHc6ddWWzN9fpBY66fvvlUbD71hUwWHTMFhboZOEqR2kB
0wpYBPIVCO2hTv/0ZK6pIu5Oh+UV6RhexH2K/0AJESm3FTVV65ULp7ou5zBOYPQvi6PruTyu5rYA
a5p/TsFevn6rz+B/HN/ctm8rvjBP8i1Y5HBBt5qJ+rXLua5E5byoQlLG1urgIQI4XmtfS1E/yw7l
0J9T8kC6AOfzwKCgyVjJ3gcUHBLEgjY7Xl66UhfWIdBLvo4IVvuoO2tPGCm/jxTFAKp/Vm3bcYzx
LMdejo80wcAQiaIJocJGDkR64d5Yndz1NvjyP2VJFafr3CxKaXOW5bTh7dbAxtO+4J48qI5u4kcS
OZIdhIy2LkeGBb5BXlLUnKwunYKoeNWsc3aGPorfOocnrOIcc2Uoe0HnlJT1MX0zeI4Kp7PF8Et7
VI/ghVNEzK6zSD3lxZ80I+FHpgSkFLaSxSwBU674wWLBuUB8JeEnxxEKFGqvA0E35U9WOpknQ3JO
TIMHQU62mXwpYwj+KSHUig4zjHul0Eh+xrMZWLvwuPHjgI+tAuIactA4EfHVHV+qC4W9+HdypulA
IpFkahRxVlIONDuiZoc6daz8UZbAaarFFvfE79ajAXwM3wmco47QxUQi38Azf8EPpopjzoJZOixK
dnTfUhYLxw4w4vTAZIk6dPRum9BOfuzOgtNufkzsglM+mwuBfZdO+J63XWc7kBRPKsvlzNzUPp/W
TJOdK1pyL3bWK08RlcV7cp3XPoN4o0dkiBo4tfxkp9zdeaQphZOd5ZSerjii9LFeJsqD7zm5qhJ5
vYc/TlqAjLWKupS0SvItgmZnsebGIRz6gpmd+RlGjW73/5WlllPb3KxEoD6rc7mJDnMAoFjt49FW
7dJNNLLFF4Ixpp4AVqn7wZQoMouuYMLx4KQt5AqpEomQfhlFXG6tzHfqYBfct9/yG6I513U/Kt32
+mo0W3NlDBercjjJJeV8L0jPs0y4YWrBJtcG3BZLQhFRhp1aJ3Iz9b5tALO9UWeX2IDKTMeNsrTY
sA9ApLUpDJsLKr57h+MzTRuJ6JFRYWFIDDx4rU/TC3h5zCzW+OrBFK3HmjADsUg9SQZYZ378eI7t
zGQy2GXrtcYpAPh/GQ/UH/MJsHAoqslBYiroBnRIfvOADj0xF60VYqCrL8wAjsw/q7yP1cVgwJQH
n8fXMdthhO7Gk16unuv0xGPeBwncNxsVJT+SyZRES2M3v7bUBmCj/wEBCVfhoWZw8Eyy1InG6CpD
5Xw8OIoYgVfnfQ+oiU/JoPJunidZTErpY2H1Pf8nQ9OdooqOLD8dYqvcth5ZbrgWOSmLcL9nsZoz
fQyJ1UeI36fn9j2/5y4mWq8l66Rsb4/5zYSDlCyH1mGfJ5jUg6k/YrBVG61hVSjZtIgiaqeL/7DO
WLmy9+psYjGogm/5rzAUqxnn1wg9R1CD9U8+ncz9JQVDCGI7nF1FNLu21q6SHfbOT73pmHT2gJTI
l6xvJSkLrykix7oa/xIHW0zsjVvf0mqQhET67Z5RdBjf4NU9A79AhtIfQBQPBkClciBAq2Htqx/Z
igkl19WklkawRaDiPCt0VhPiJegSifi7yRIJR1xa4VEf5Pe9KdGwiW8Ej8DBxhdrKCY92U7IQz+1
fX6z6W8Jp/hkc32BALuNWnnvKkiuiD6FawW4NJg3lKiwpaguxdzO/v4aO4HKlwYtq5pVgfGfA8uU
LU+dKJxnCimVDnoFKknuLPDhWMDW+N9L+GnX6TKXzd21qhe32EYWJmsrAlOwNnzCVBkK/w/dG+e7
lyEpNgrJA1yl8K2tqN+fLV6NTTYx9Q2sKZQZYe4f0ssqNk8/8Rnl8CjZqPF3D0IN9uez//wMsCYl
HfZzXNw9R046ulbJqiyoHGG5qpQKcbQas1psqt+Sj6vWMM8dV5tajsaXO+nYMcvI3apgAcSeQhzg
J8+TMkqfnMzuDpELnB63Nfc5rpQHmMimVJVwRq8GHf3hseZuJb7/h35t/qK5NSltSNrz+kSJX+9p
AGWCcALyRbV7TTYtSN6ivDDDWNmWiCYoAmb9z1/qv3bN1hkPy/9hzkksJfqvAzqFsDk6LU6Drt5F
dnTYZMqlYA0oRYdRfEo55fAhsvShhsrREWAs1ue0liYh3Vjck/SIfjrO1/pQsJnQYju8EJalPXkv
+cprO/hnYNXw88Ri7FTWvMngP1yR6gSTVqfORsC3hezLJ2xdmk8SNt9TJa4o8Tfq2Vfgxc8f5WBj
gLqYIoKcICWujPW5DA03ZHkBXpc3tnjJ1u0OHG5Bx4A+BvtZNTa66i5vFDcETXzJoe1MPv6EskNx
Q2s5Z5FVEJ3bhor/ttUn7TjntSKlL7QIESa2YdL6HRldgtn1I3BdbSGMx1nYBzNd/bdzHX0jpCsS
M7AcYrWHnD7+gBvl6X4GdxUyJI2AZCkJPeqVQ6vq8MkKX0d/IHTnMBtv1omr3bVuIoPQ1pr2B7OJ
V0EZ7PuVuWZ2ly+hKoknI+XiSyPcSNmbR8R9cFoAtI8AuiByAD4bDSqsYhBtFsVDYzwfn1MH6lCt
pMDomCWnUhXG7lt/fxmKDigGvj5+rMkPXoPRbsssn9J1YRIj5DDjlq7pD0avly3v6NKr8WS7sPBw
xOSdCWHdnisRv6+eEeHOTSHAPS26wyZB3xeGcAMMcmrA6HO+FBaA64im/LKekl8fHx84MqHiu2yu
oO2yGuMAK3fUgG4AJw9Mv68qyovI3u3gdodf/G17h3TJ2rqUwD1Flw3PC7q6t8dv+Oqbt/KaUq3A
wxZBhTrmb+ZNOOS7dPMxg4csk28CAFoqh/MMY7TxutgIQKEVTnfAeWx+fqj5MG22jB3voGxsoPgt
5lEnUYujUFO+mwPHqNDaSrU6hzJZAFRCuASYmnh/1qb6emCKxPIrWDlmCe95e6PZmiXUhivYsfFc
V8/5FQIQGhA/onEXCbQKzQtBaaC4gIvPP6HUYZkZu7l7qScerZ5e/CC8PdiGLWwZOY5DFbDre1H4
9O2WEBxQT4v3p7IEYQGQ3Ui3B/514u9hpU8IchjhhmFFRbJsT9YTuJhYrJxe8U1t6/MjO4sjbdsz
2Zg4ePMOnCFAFkNUIMTRGVF1yyqcz6ewY6/WQFPMcJu9S3ARDymmzJ8+Pb/oYVAyqQQUHoazwtxt
IZyvCZOJ9vWXx9JQq/4W2jWzyMUSXaEYUMC5zGpZB62qViKLHGHgKLhzu+rK2tO0zb+3nNZmU3qW
yuUcBRQR6PiBofBhHoYy+exiHl3Z5LxoA5MdWFYqUBLJrScT/ughUQfG2lcc5dP88w8nYeOnHkxl
xeQ5jpOtt//zYpmedaQWzXW74UlGa/LgXFKidvTkhIMzCfU0vWfbYPTZc9TEAtlN669bGho+kkRi
vz/Yi/C33NrSuZ9fBVKV0py8mG5wbg8kAlsOmv4uZctwT5o2y8/jtMq+J0a6MG2X8TX/P04mRjRC
2zThDEzioIVm+7xJ9ZukLq0AXWCA6XFvSf+brU0EUAW/C/1p+pqkdACTVHpiZ/VhNkIC0n6WY11d
QrZwIXQwktWLow3MK3Nn56rMprbWZWNy/6pMhxTFSx+fpsVEs2315Rhr2nikXZMLrUmN7IPW9t3N
Hy37XwnWDPYtmuVUngreVKjEQtHx/oXDEPeX0h9cXobqvFiEWSNC/NWX51RLc28Z7g14AzjwZuz1
p8CmpuRaimptxudwtUFo2Ip8fpTpj7JtOhAbXOkIf7mZ1AV2YkR+R93b8ldKSkhSg+GCXwpp3Nd8
wQEzAJgIf1LHBX/mbc9egoV+FH7T6aWByQ5Ip7ipc0aUMlzaqutQ65E+ByR1DGNw/mDvOOsXuPUr
1W2ZJHMVmtv32+pV/0zaLW89fEAtMPcZLOznOZcxbDagCsuhn115utqf+W4jNXYmpwa9aLtwIyAw
0/Xjvr0pMLjPzhyupSFa4BVrpKPNGbiLUQTXe7it/IBOkZQSGYMt1HwI4BDUN5hPvCJGJzk/Z8ED
oGRgXYPITZWn6yT/v6gEk2+DEVepWBxtyi1hAFjOfnrgwr2UQ5Yf65DJwSs5nKOSkA6K7Lm2Le3T
Ys1fqSn2Ezdugmp+GAbCd2Q7z/WjZsV+yHHVvPzdBuuPLbEObsBqyTTJFjeGQWvcHJ0TGx+4TgtS
AT7gInHN+8xi21cRLrPeFHk/CY2YUylzY4TIfGGuWfoaX+NylPvnA+qDhcVbntGKOFHKP5B4NSVi
Z4zVJXX2PGJ0OTNel+Twd87tNDYpRtVS40Q6WIV7C0ILWvW6RZvkrqGQhmvnoysgu+M5kQXcI8fX
9xFvFkNuRQW0zBiR0qIq+AP75M3Ky4T25VMQ71Vl4AYVZJpSEiktEy+I6Yu5wcnoTX/YWGo+A9hM
+lVALpxX5D4UCdNg01QYErgdzNPPCFh3SuhfjzGRFiOmo0kI8TqWCxe8Zv7yiAYoIkn3/czkSd7V
XrmRECVmYGuSPp8bsEHqFlYpbYiQ5iIALX+2P9QS455bcNvsRX+lgbQ2dCmTFnGDpCx4NYo/LcJ9
aFfD40JfdB/huuAEEiaLourmvDIAnWi6GqE++ueIV55X9TIMQ8QOSTArPjoCQ7s6dMzG8gpN5AiI
e007oUHnqbTyCgOX+476mB2BpLQjZj+cR5UjGpD/5vqlZSntA/CpyOUOSY8rur6v15nJ5g7oZWPH
0NfQwOphHn/Nc1+C2ByT/OXBvb12/FnglF+O2xQ9maHJ6aC+eGnetiG7cxu9SD31auJSjlwq2+Ra
pe6XTbRLjPOlRmLi03WZ+zscF9q5GKDg4J6qbUPNeO57dgHzW2gMJ857dYmNh5qCrIurY1s57dZC
PeBzSAfKChKLgKbFBnxxdJByQKqezoBxMXVtdYDFYPzw5tuJhneI5Xnz5vUlCFQ2qsOz4i+K6ng6
vSkGQMRfVdjl8se7S/pOmYItny7ISv+UIjGEwZj+29YigA1qKduRTqGtyfNPiUzn27cSmqCVPsJq
HtV/pzJxHQETWRSo8oejKgOU8WDH6qU+Ztw294d64RsY8JqXigkm6TiojKG0JltCFnNpoNWPEFxy
Ls6Tw7NEZcfduuqDBzp9/NFOHhwvyuBPoDXXhQvicI+n6WGRqTlYbgBXoiyHTnTmbbYxzwhh3CBy
NUXWg+n3fj0mv/zSmMV1l5aDstNzQ8VelGlZ9WCIg1xwsRgfpg3klvabmraAWsyk+RuLEvewlQ/z
bMd4D6RXiBpu5jyzB/Th6p7h6Cx2DkuixgiiIXvecO6hwxk3gHrZAMAJG87Qg80rOhhx9xkqxyFU
ashVZXVzKlTuIbThonXoTs6O1lT2KaQ8rwbArDaVTS6grOZutupCIHskLKPSyH8If5cL9v5ppjqx
L9ApWPXh4nwzUtXYhnZFIUM/j/nPXFK4S2nui/nOJM24X1sJdaPcm6h0d9cQV8ihpNHTIbT/96Ls
D/eEEw9p2BJ3co6cZMiePPEEhgP06kOZi1G5iuEAkvwyCArUf9sO5ynRHxaCUoMB/ehu4jM9h9W6
B8Z/UhV8RP/5/5wLp6wh1afA1n0NMvCm5FPQvR20r0Kj+vVO8E8R5HQe/r16v1Zl6+HJOr9dbHgQ
Kg+wTQxuG9CILMzvexqD8I3wHXUyLpv6q0sd67onEn4mMmD3Q9dBIkfJawA8/AlvptMS+6o9QvTB
j4eM5yfE+jGZYtehcuqeIkh8pDiufe8yBbvCSiBl0KpdSiNwmgF9JykFA/Cyqy7loR9Y287LigFE
XC4L7lmjHSH20/LNVFDiPhbPVgwCaFzTmhxIq4n8+oG1PUL6Hbrw0/6Z2ISvDVQYLAEx44D43OXq
RUB/VlBnP29X25rf7gOtkyQ+KJ+p+zxuv9cLulnA0JWUj8QMVs4VwRTssmcOzaxSSWDNnguyAZfX
x4rKXalFhO9MBPoU05w1Sz1EcCngR04f1O/2mnLQN1ubqMjMmP2F9qr0af5fCRWYGPWQ0QO+gBA5
5CAQOJ2LX3J6JdViRgpcojofrk/RTTCviFS2RsluRFJleo4i6HUIK27y0ITuXmSAisuTHBn8JQvQ
ukb2vCncr3dUpzJtZDrchDwf27WnBHWLqjhubYzgUxyQjZmHCz392SY5stIXMGRcm1PPNpsz+N2c
GxXwTrUJi70sBAhhZHztT/yaZtxURAEZDo5XrVJ1UXKV+nf1trpollywZG7zVCkViKPrQP59eGLb
GZOqOIZvNmHDlAzPGcD4yRQVqinLCSWYWBr+MJ3LuXe1o0O+EjsDydVjCFmVmk+Oq5zM+8Op6FjC
ISV+eVyQXEezoG+RoiCeB+UD7AowLqJDQQRXY/b4FgQCo4+yn+10iJHoBPkCGBB8RlvDXIv9zLLb
oNXMqmGRmgpaOelsliXxmBrCuPOdP7izQUSn3YP+UZRcnrfNS+lgH86/4Gm96+i2NJlFSNUdBQF+
DgLnP/qUHalvRq+YGnx+u4dIc9bVZFu9uphNVGkM72XY7RIK8j9NTbqCHvMHbBpJipkOSKyIi4BK
DU/qthxMQZDJhWV+dNJGzh90PKokpnkuneeCpXo8dei2KcuDyo7khRHyvtz8bj+IyXvSrUilNKXQ
3TSElhzeCbQn1rFAbX2ma7SH4Z4W0xFKOk4qK15vkG8Gp0KudoepomGxjiaV5bG02uJ6a0o+05uX
BB0+sdE8071a0/ah/BMClOHHHP0M4AmECWhf0XBkLRbWdDYpmMWNDrJFlpEMVzmsc7Aluab+64MJ
rj1PO+5OSEg8MPLU0FB+pKPQgTohxFDaZCkCbnO9tcO3UdgwDQB98gKzWeMrpHWMkwVYlrKkIaup
zo/2O87Xr2wCgkT3fnjLqrO7hOPTHZWejgCyzvFV6yY61l1X9qhrZVMZ8nUm/NQ1mV/U+S30N7Uq
P9UU5MQgJQPOpH9LJBAhzbn29ZdolUtCwvLbz9zuFJIjvoIGs7XtpSznn3f2DtW1bF7G0APf+vy2
/lBdVw8nkbfmHWEyUU9zk2vNaHlRcwhMV623IqAHtIE46b8Z42QCyTtStIOX1fXeyB/kMEk7QJwA
ATIfFA6ygXzMPHJOHQNRM1AjCq+oEltWHG/oknoq+CVwuOG+PFYhePbaJhx6wbESJ2SHDLCXoF4a
anYRRmA3TFMHwe2bt/NYD4YnxQcO8lQ24/Cw7rNsOYmBshkD7K9DjBBfARC2ha92Rg4W6r3Mg0FG
u/A1yAHTk5WdoXLUqnajkonfK1XzXXc1G17VXj9IDw+Gvku1AU2j8Fr0jTeeMOgU6erGDlh3KrC1
odk2c0u45aTL+WwKso8emf/LiszwbKE/GArHChwOHmX3WP9DnH0mC+6ikaU09pfw9jMzykOUwV/m
DccqzbXDkvJJGvF3sl203tZnsnuJuLSXdGL0gzYxbHDJGfZB2nfMsH9hqDNjvWyjd8RH+cClnj9g
jARBVbb1BTkq/vkIgMLANb2J5duwGcTxhhqiQlEKbj9k9iYVEzOJQhRDdCcjN+IiQHelBRGp+Dqb
J914kCxiaKg6WRnVmsxtdYl3UKAGOnBJnMjV/FpLnspam+JjcleMWdAZXW18PJ+bLwZ3t6Yxifel
UWtq6SrNdTlEyQ/AAGbk1JanMcEE9BAbAB+Pf5xubwpYlqFXxU6gVgAnKvAGvOwj1RmRw7JUHvdk
1YQZAMEoU1PsYpdBlU+mQl7xNA/kwoilHol+8sBGSBZRCCVc24hb6wfZ6y3he0RTIXAK5AURVrfu
C+bElnP/ef62loF7LrLRLxEQ+C6Z4c8ZiHFg67ZtB60cI0O/HW6naGAtgepT0P7qPTDW15dcG4lI
EEBYIwn5nRt/VY0B0H86KFJd46W4VKf1bENB1Gg70TTR/FfEwtZSpPaTnjQe+Jbg48yMSna4b8PG
MtJRxWOOV1zmBpEhGRMkLCk5YEpac9oZ+Jb4Dwg2mLMHCOWiFb7ko9ZH9g74AfYlRlSMS7npk0/+
ijTZszdEB4JEbaichd2cFUh9Aroff/gCExf9oLAYIA/3h/GU+mcvyZKax12Vs05jH39i9wHJdc4p
OG4h/ttW8rEMRChIFDvanffP9o/JRKcgxKc3nlQImtmAXBUpP705VfPmEqtyoIODkPmG47oqbOP7
rD1iZGEFh95Tom0bE2N2MisH/NV1PJ15dpCj5TPXgkwysDsi29e5Jo9qm6nUbXH9XXWawEr3GnOU
Zhisit8pMZ4XhUBFhd0ArGFPBQhm/Wq+3zFeWxbmKk+kScmWhqyFaXRfRYwLqVGczn9Vn2eR4nkA
vCs+r/VCxJUjmM5ZXoEMdC8BFEDJ5QKAmIPvz6etU/Rkw9bgR3RsXrvlfqGlXnLQS+HXBpZy5vpW
ZtntVuu8uSTTw5CfettURHwNkwA/dkL8MHSWU1/SUGRWqO6qoKIAkILQO4+LsRuyFS1J6E8nmeqG
XoGY+JZ/3RbiwgNevmUS3qThtOc4goKDpAr5yU3ZpivA1fIby7O9+dvRyf162sUvTzC6jvLx2MWT
4u6pcX72qbfnp1doLg2KiZ7tLeAptm5I0VN0voGyaJGw/kIuLKmQeTQBfTDdGduVr8wbinvxf/+n
sBNcRh0tWov3lUAjT8FSlfCmGQmW1VFPTEeWUrdHpHA8kDqKmT/k+Kn9NtzP7M6UFF8yo8xD/7xA
J9Ux+BgoOsKuJlzBd6iVe7zKiU7QDiN71G6ux65Y2bNp7Ya8F8TOLMwlFhJ06hDf2eU9YmPn0thu
7eJ9aQTszf5mbUB/tsWkKWQI54zrMMOyDsg09UlQGNgJuR4qNxHYvID9sNUGTxkc7XecOoJxWVdL
z8sSNm2VszUj6SMkgRJe2ZO28PMuUrqJhaSy0M+6El6/pU80qYbaWc7zVBJt0xbDDw1iNXWHuCMY
eq2fHgYhtWFezZSAB+bSLbW/Wgiq9Z0dDprp+hcPp2058K4pWXnfod1CPXjwIP4mnfLB+2HJWuuN
Nb0eKAv52ai8khz6AMNbwnHigKOdqBSzgSRNHBnl/KYXeokov2HEsGJ4FC6q6UGCxYAgN1h1a2Dg
SuvtUOwpty3ucGG41rFtmxF1gbnErr09VG0VbB0eUA7eVkD6MZ360kpoP47T43rj1wfSeBHjc4L7
BxeiPr50ltydBWpp6laoSF8j3T6yMcA3rneYqW4BEUlwgmuiHsEfxaUc1Yda5zMdfJq0lJ/H2EYR
P7EUQfTYMctVJW8U6q0pE56MS9j40k76BjBGNh8GzQZ3HmRW6Lh7eGEWxtL/UPekKCgaZ7DsXVSW
LlhKb+DWVueZ4di7Xds5mKsaHwJnMSI1CQXM4zrB9l5Zz6IWUhba7UFvOnC6QMIp5gRUzFgV2A/L
C6lIObSnBfOLqt7eD7khPSF5a0XOO8fF4aGXERnnUsygyA088O+29JGYZ3vp16aohnu/cEfUL/o9
OO8GQs8cAxFjgpgnSZYfi1z9FZFgBoHQmPKTMZsNpXJXMW62UhgvAVMmoOX6yufpN8xxj0mNSAxB
k+MeBjDieYLBTcZC4GUvt5He8zx5P+0m00e+fEkgRDKZVRIjapXpmQB34n3cd/Ye3wHx7Kj/B4ta
TUiFvP65GJDBjX80Z9CgyAUa5UTLrXNbWt/AiJwmWygXBxSfhxlkVPv77wD5e9+axeQDTTOA1FCF
nZOQRLdSELq8sY5rt194uog6gBhorqhBeBFohY5gW9a4cYtXH+1AXBRVcaU6TCS/MTlDtu+9mQuC
bfq8v5l9Wnj0TjpjseypN0fpCzNDT521iGAZYTELdAfHuoaqcD82BG0I9EvswTBV7QktIilSynDI
utTbCcDqroNNrV2Kh6oIwvmqeslzS0tQufg0SfWPnM1HSbhYhCSgDHwyd7YG8s1UPgY0t4SCZ8nI
AvDQ5aojbLqM08FTUImW8jYR4akOtAuwjphnVkImbl/ykCytMa6rzbCcLJpFPB3+jPtaS5U8t34l
JiTwgSEUstouKH+YFTgMm5bNkLGh4K8IlwfxKNVk66610geHaheyW/jTA2wYxfuwB0Ssxi+1eaNd
2MONxR+BYRkF8bGg2J94evZg1DJfgreks01hpmfClU5M6EvygWctOD3yH9JzdwXSPHURI+3a7PaB
/KJMRjQBy078GSicl8VFoYPoFTiLAGK3Oeoak1qwrYX6pw9yrQoSr7HO9Nsb65+GXzs7A5Lytbv4
W2Rp17KTBhZyN4mOjm4UGziQAxq+xtij9FdI+6lLiAsb61hGMBqrn1tD3B9LTZ62VfyEeVPw8LSa
6S/OeFRRHfgUk+tVbai5qstCBYJpvO0qVZWlA575yMSgV76mQDxIYhwB0IXVqPEbFcOoTdJTcgsl
QhRxd/T5iWgPqxdD7MCHCRk/0wtELcV0bzHsCUCT9+FQ7JgxAtzDB7KnQmxmHaQdr2e9Bk4zUD+t
919qyhMGMNVRJCI3rvpxs58bDPUHJ2cujhauNWcnBYTDgeZAEHYNoWQYHySwMUP5AR/X6U5422UK
iB6IsSifl7tP+Wb6aZLMd0kM1NLjZ2O4OAAQzLWRnjOUjo3MlSZyHcy9/oNLrFt9B3y2rVCZbtaa
ui793GR0fbnUvvsVz3S3fTYZ9B9/xrNQjHBRhBp8F5ygbi7MP7u3f4z8MzNwYWhs/yXAiADOuOcD
mxhKqqRoWQ1KQMsEuGf3WNppLj9KSEdza/b1gYRLsLsHSzYM8p9sCBWy0+PBtu8DXFy0YUrRBifl
W1qu4U7AizyxLjmp+gFEHPR/3vSMKIjVdQvmaPXxOeusQ9pL01RdgGTZbeWZCW9W9QSUV2+o9h7d
N6tvyaHUIb56zmvPpeWL9IkYWm/WE9qTn5g9rd91cDQIji23cKmNE5G2nTcI8TLMvgO+vMfA+QAQ
XMQEQq6jw0inYEcx49pEhSC6rs4pABikWRsveUSkbyAgIPr8QDMgmHZcErsX5LY9vw7xvSn3Vroz
LWIdwAUcjYBIQ4lcFS2naNK4zuMvzrP9NB4+LGBuQUNtMtURMCl057fwUeddp/g3tRygq+YZcgmf
DiJae3DdKs7OLRJwBZLgvIgSs9wQK09AWL/nQ5VrWFbGcL6k9Ljo6QIfIpLhWZ3Zd7lu60HKQZp3
cH5Io/LGsmysbizT+AuGyFEARkeIym/FQcSVp+YXka461M4Gb/JA12l+RwrOYEUENJhadRqatbbV
6SPyvsbRn4Lk7i+uGKN3YafTFVUpb23iCw04jCpJFQ1zNg8ebZPom7f8SUo5tVMlOZb7ZGyEY2gl
2GkhSx4yvfarn6UXNrDLeWp4D4DKKuO1SFpq8YbrczLmbCOsMQvykaOipE6Yy7spHS0ra7ct/MIP
tl/ttvNcHK9T84m8nCFyV22gAdop0S3SVZsRsbogtrkhlz2IhIGfyfqFSwXdKEEc8Ld2IWICD3pn
jh2TArg3yZxsAIgkxQuik+Rog4+cAnU9hda9+LBvJjcRWAh+fWCvnWu6vW8yPHuRKsI06t6tIrBX
dqKKbJX8MSIOJAvEpn+Bb67n/qwAHJfZLGGLitUDEJGiqKzYjvggZgNpGz3oObXqs1OcatSFWAer
wEpsD5AvpKXP0tkoY8CUEIB5iMXtzvsRvKuYalJHPX1/04xCbuxNi55pKAIk6rNoaa8lHSDuSM13
w23e/HhVPs7AcB2x4S+6fDE8RB0b6DLHoxrD5etgh7/y+IKr2pJNtiaj4uuvVNaYRPDEWudF+fE0
SzNgN2pd8HIfVN6FWChGFt447eWVciNEENq3d1yTVYi/bPZPCgBqGrQVsijcBn1tVjgTHFg1Z6Ua
hGqUhrupbqw5PcVG0Y4NC+bD5R3XRuS1h6hOVyU1SpRspfVZLvtSDnedIqntyMHOctQg7nvAWhy0
pd2zkn9xEtiGMc8g1m687q3KMAAFah76s9Wg+P1kv6qYXT4HIFYW3DGESVs3dFq13lbO86ArwNK3
EDx4HsaR+0ecHVgApewr9NnU0wTxkPEJrvSmCQjplcmfmTSfZbZx/aIBrKN13Q9BLEi5kZ+zSqsi
OGkybogw1BMji5zt/OGKIvQW7N1jiQfArMOMFnvmLKLqtDufnsxc3TAwNKtTcIQIDCRWdWJWrod8
e7w2dOr5QiGVr1SxSs34egM/t0KaysCkTVd4O6Hspzawf93dyCvFsBDsysvMKDQBCfdGV1B+Wxw6
S+B7M2c7aXpzfevCxnbTzsIXfF3S0A0IXnIGecgRME2YTe2KNp77im46tDLY0PYgd3Jg+t8ICe09
FOgjE85HTsNNxaWVsyTEnwlM6yVM2XXz/fWp0/XdRlULS+DPhQcmkWizgVTKvrpdRmH60rGMz6Ea
BvgeAHvbOE6W8T5fHjTJSK7XcdtyF4wblOhmtsFmByJ25nyi7DUQGLExUx1SyZo5eAy4bvlFWyqQ
PF1RvM8v6OCmVrMQdwLibxEX7DhU+0hZqzWPx8ER51wJRuntfH/P0W276s41QSJyYMP+V0o6i1sG
vWlWB8NAOp+05jGXjq7fDY1tQhk7PZDKz6Nc17fEmo41Ua8zSFA/aQx0bUnO7npXoSZkUpRzCAiM
Nds9v1YrrmSpvDa6iz02UaoNS9Tsriq8hlRNoLBbE5A9FrNnJ9TP42l6IrX5l8GHok1qsWG1MA9a
8DxRIXTjehS8ukY/tQAEDmh0/ot7qinznbzsrseGMf0hKvP9mW7E31ofbBdY/QJvBh84TKTQkw4/
v5APYpxl4cQcUzfsvjvi7ZPhi073oGLwGqgoKrfeZRSYQ5WXjkyRai3DdshIxMLef4mtClTMFk2t
Y1A1oKcGFbraQ9VQy1HrB2kBhtBBL/v/lw0GVm7T1uZvDHy79nrQx3NlWNc0tzDfBiMapO9PJ7v/
Nc7W24WcWq0GFvEDGn/aVz6aQGEcT1IjlRpc/E9iRxpZycMll9TU4E9GzaFZgiqCBpRXoTmo/HgD
pkKMSjB2e1ceC65pIErSLcDPxaviVO/u/bF8Wo090jXpQH5V2Snst46G9KkkAS9ctBnjUZcbU7Hm
jNxDaDS6F3bn784jRWmgoBW2MAoaIOQ/JA9tbf/TICkkwc/3NVnUTHxU9r/6kt6ceZme7tuwsgUq
NwFukoKegMjNZAveyDFM3X59NhTRz6E2HnEFdF+Hh7vuniqpvDup0L4cOY7GPvicP2dSIJLkKUFc
IroSF8sh07YTaccRbH+Pq4Wxt5jnjzV8NND207OsOfm1RhUUjSe3NgEkOnSVIQScQVWck4M6S39z
fzUjLY8ZvWGq17hHy05PliI+mrqfSWp5VyC+71rJKdUQ8R2cscJn3wLtZ4M+pH751dnv2t9nprnk
r0aVW4HQ1mz0qhhf2cVIxRfOi1Xb1vujKDIS+ds1YugR5yUSOSBQnH9Z3C6TcNQj1hyc95Dm7MlE
wQgLP3XiR7I+rvSYpdEkbL8umcSI9bLf/tdfApZvuBhYbXB8kVADYmnmuJoHmwceuj/Jix5z0AlJ
I6HlGk50RyCx2F23inlMCbUns9HC9XKU4W361QV4UhjMSpefsz406lRH1fMXV0UpBoN01lMCZx2d
OjlnalTBIk+D1nySbPvkC4yuzHPx4rFHAR4sjG39Rq+fZ59w3lsCZx9XvmMWp87K/LiwypOjZ8aI
W+RFm3apQFYtzRTZc0D6qF16boKPm6Ga2Odw493eVE9S7ZWze+M/X+Cuvnv0AfJglzXu/8wekL29
hFC5bbuUCLzIU0vc4VYCKvwz7Qa1eT1DAyOAjZ0BJ4z4XsuFc6dwsU1LCzeFixI+IyIPwEIeDqfP
FVX3ltOe2i/MV/oSD8C/s7uuWEHBmqTi1xnzqZof4J6/kbbwIm01ze0RDyrW8zdotsTC+oqRFpXc
AOX+zXtV5CplfSt9c3cKYZcZQWAo9PoWJCySHWteIyvE7rB+dVdMzCRGNFr/NX0QNSUKO04db1+6
HeJWElyRsjJvCA7kj/r+G84wkEDE8EDUfQecRdfQ5kUxqJA0Y0XzCH792fma4WfVXwYBmt2OMnGP
99PfbqvAgW2UKeI+h8M0Y+S17squPqkiWx6jWqtqWGknp4LbeOEg5nyB4IVw7Am6PBr095HyOGVJ
dM5bFRCfj1vw4LfmVOT8GtoLDlaXm1NrFu+uH6FI/ER2Rq0QgC9TYW8ag1jMkhshhWUH+tZrnkOW
fC5iMstz6DHkpbeDNRq+UZcUj1B6Z8v1GF/CoBezgDxCz0sXs69Z6KDP6i+10a+KsK4r3hwuoXxi
E/k8CxEr7ZGkLcmZLlECeXWMSSQvnQdxQqpAK1MLuC+usp2o52Uo2hqJCFWe5nhZYygzEAhNkXCa
6ATSAU2JyBXN4i5PXFlxAaF75tnp3YM9HPOldIACAQCcvAeez6A8q9BSkOpGmAarjjmk8d3fZmvZ
zmWP+DmgzLxEOKSxt1N9Jcf+3eboYbNWV2toTsL46n5OZ8vIDkSkGKHoESZMEVdb1boylQQK/z1i
b7qlbGrLVk36IpDhcNKClTPAup93IfGEnwX54nPikU8RNihPYhDjNvwkhnL0/Et/eK/29K8cnpuK
RDfuWQojI+YOtpJuIcbu5B4tmRCCJGijN87YUKjEUw46XsoSl/rto/101i4NyLwujkqro/JKhouP
u47wsJQFIRv74HH71JD7+5v4Y5890QbXyppw5KE1Gm4+rwdFtrPha/MUin0rfU7ppcTzqCq3py0i
mWzprW7H7qVBHeVFHMuAn/8zwQQeDo9QVxv7ujbMwavjfEsL0gn8ILB7ju4KVVFYi6U2lRAkl2dP
atdK3f7yPOoTWOQ78om5AgwJ9yt9uErlB1PIhhLiwc+TuJmJ+RbmB2SrV0Mv3jlK//P8Z6/idT5G
L9AvAw5EW9u23xFlcJOa8DQJVkNxeEeiiusWCvrLJX6X26SNKsWBA/GvNhfKEBQgmGFgnq0I35yz
ULbgXQAAItwx36af8h9JfBFeo8h4JjYX56jHgNBoXK/huDTnCLeZWIBcld8YCU5Vkzye8+A6i9+9
twT0b+BlLm6c5Ui2OapR9ZP6rnzIiGeL07An30e7LX0dMffWfAeKk/bv8DqzsTT2Wl0aWW/QTPFM
nTCekxZHCLdzXzlR73G60uMce8EvU9YDGQDQgbeyeHJD6xln/f6XUPSV6CpDDv7ntbtk11HhG5Js
Q1LZdTGUHQ2Vy6iGDQrSQZKcES02ZLCmIJ7jUHoDbKhyPk60HOnDgrdlEsQvxYw418pbdZr5u0Eq
7s9wBJXVaZAwankj+jyI8GRFfYBOfBOXa2ELihM9V1d+70R0eHF7NW5iX9/NTIVb4OL/1H+vxTsZ
O7Rt8JJ0WoEsE1U98tD4NHjrIfreMqKqvLlgdKLE1gjvKWduhg7Y6umjsOOOKwJg44KumVQuxjr+
Hfkhe/ICf929qrZVG5vvUIZ5VzUtzpG8h6mmE1lgL0kY7Z2L4qfPvKeDOGjQXyhLNDBPZyne/m+/
nuaDym0fYD0AEsIvsLdB/ft5MU1DxZg8kNuAYamkWUekZQDE6YDS3PzsoZh92s2V+q7AbfwYPA2s
yly84wzRoUCdqZFhnFeZuJCO3CwGS7yCZmlFCFalvaSEgQI2YrR3uFIiOezAjOHG9QbgIm5wuybo
mchtFeazYo9asIMTNQ0ZGTc6tn0Whmv4ZOrehUABM+uuAdEVvibgelV2kFyg85NXQyM5Md8rpzF9
CMKl1rP1FtSGKjOSoAMMxmSNBbi/CJN4gdUBK7XwEahIQOkShghQhwxzYJ1lMzSvaKQN858vPD+0
dI/b1df87BlVeamyL6sErcP2IoMxa9Na5J8AS2mVqP+sl0IHckn74yW32Y1020ill8o2C6nnmcEU
QhSCLGgd1lKOZpIfHOZ/CakDb/WkxP1bXikoxmMX3yL34Idgvzh3QvHr8O6vKlONC6yJzddbQaaU
l9C1HOA12OOkulbyLWoUls+X9o0Fus5mjF3Ap17RDd8fyBvsNuSBmTMcYrvngk0s9sgXchqrRlK8
q+P4wyRQH9lfx6ylHTdxKbHDPaSde7aJJO7pJcHSJ31FTPtPw3HgRzInZgMRnhIcG+LoMspiPKvV
avhS/Qtexk49cbPC+NL8DFqaWx4wS9FaU5FSbAT0iYkmOWIoORaiQmadrrXpybriH4w6C2OcjB3U
ZPGjyveFdAE3BHXSflXXtQyYOeBAWvJ3UDKJzKKuLZDzi6ZI8q5ugbO7VTMST/CBpsmpTRhAN88Z
fvdUYcVEVF1c3keiutEHQfr0l241v8BNz5UN1tP8uhu5lnOBQeDnmnlKiN9YlSBvH8mT0fdkUFVv
O/ch60G+uA3Lf91x4HKglFgmXRkIlKYubHddP/cStG46j3+3WQY1swwldGT+ZDAj/jUr1b2lhp2Y
kQt6MEtfp4/AF/9Uri4uMgrSYSzNBm8N1Wfe9Qod0HNLfXCaarjHy7B8AB7uXEY2En18p7e6R7Un
W6aHYUe4hpu97yAN5TJEpVGK41xgkjyJRDNq0VZrTa9TQClxB89QZ2xjkiOf7CzkAWV4fKpCsMi1
EZVKxwOWcpYiG0RbX3vq11h6ULEyLRA7+7USobwqn3xhIt09XEuZtH6P+J5/V1shKvBUUL2gD5jc
u39JOtidgiT3J5VVUeA6K/soLIqUIE01lewMqbHsHKDrweclAESLDWCUGF5S0wtkTO+iA50Mlz8w
vfD/u0Zpc9UyHLxAAIzeMAypMTTEC2ziby6ms08gjcHjhk466CbFtt1V+f9+jPdgAQNi54q1xkzd
npThwpxiblCb9DXMyQbPu0FFVhSlFdVIbFA4IktjSGvYCZNUSkmtVWsqeS2XWDVn9fBvDERW5LRM
aT0DfQW23ouUFeCbVSxG37RYZ+mGRVCqItlkyTEHbO9NQDYC6aiBez/aTnZZsk3HQqP1WCS+ROm3
KOPF/167yNpRl41OLsDZAUxLq4oE3Xd5xJ97gvCDWnj09S7o5XKH93BlTXCUInkDGoDOdS2yYO4h
gyKQEACwU4Ke5x//gOyGszBvRaEOvcIJPbFzhJbo9rXomKF/f5Uv5EpKQ7KR9CK6NYhrZQ09gt+6
bRi3AbIzqyJBpmaqPxEYr37sMfxlSoKP3jjkgyKCjx+65XBV2INFmxk2cs6H9lL9bs5FXxRAgvWI
IUhy5HUOiO5LmFISrt389Nke2statmU39vnD3MXT5/CxUaqfc8rm0b76GcV0GkrSv9Gd+dzbQj3w
mcXVBlC5CsWfqjkOTR/ippsI2LxyZ73Y37914htBhYgItwAczZln1e09c0ZunrdwWdHk9OMPoJzI
P9eAcdmo9QuMVPn4BmF9mHoU7w7xAVUgjMqv1hYOnR2HijqO0NFfrErljzJ25bpM/cLPzjY2MWLX
2Xd6UfKcX+B1mUv+8yrC1YvSKs79qEEQzCPtqBcXV3WYp4En5f6sDL0qVROz8ckxikTseU66rps1
LDhL8ypFqh+2z+IVEQlrlZQGF0DMxXt1MZfGD2p/vnvcUJ9QNVZ+d32qj/ppJPjxTjzow86JlzDE
AmLwxvZi5fqjC7jcKcU5Pn5nhZv0/AgvZ5T8Slu2rceitPMV4zshcNxQFfsKEL3GiIUk5+mnbo9w
VeXwEp3b4OEl4nOm50HWOvARmUgD6s8j1bVBPJx9AFsV+HqcJS1ivcCBGor/PpQsTLwuTl6rsPzz
cRonLFZ1qXHStg8Sl704AB3YU/X2TtFkD8e9zJLbUuGqzMqjmWfGQKwo20A0NFZ3LNpPWUSjZTo5
ZUgLBNSB/iIgfmB2sO0ih83B7yw0vj7YQz5AlxMjBaQjKmAfKhFxmdh9FHJYO4/jXi+K1WNWRliX
Y0H68JF8RtP59DsOJ81sJD8biYs602jLWGAuICYeoGPA4iV5uurKbwRFj74k1sYMN8ikuxvYbaKZ
EBVyhEC7PGTq/AJ7cZewxA88dxdVAK5fxwdjJbHbp+thpdaTHqB6AdbywweHz4J28pGuE4/SnYJs
GK4YaYE/y/OXxHlX6awopSrki28X8HmqOpzZTG8h5qjzZTf6bmbs7HF1w+vDs6kzHQjh6VJcScEb
vkQ2DiY95dgsq/xQL0JGUV9KPhe+4RbEZMc1SA1vpVKBF3zbpFa5tYJ+FWyG67rqDVVxmQMQlack
8KpKmsNhOCQFeBB/CGA9N6R4a1eWKPOiKe2yLWL7I+bJdU1pheqaSgPlyHTx1pJqyDhidLhh5FV7
oxlsP13TAVaxNrKtDITAunnut5jJunD2oxiHyWcupZGc6bj/qSfjECMKWLK01T0RgUGcAvF5Yri6
+c+iCN9zSG+4cLZN0oeNgBGkSK8L1A87PiGVA0EeiwNaJ0n/N/M+f0Xd/EIf8Q1Nbmi8dH5wd1bb
Li8dUWFb6Lphk78g4tF5d/ej9EJS+z8gP5jjanlLQLizFsG56D9GD7tct3ppSr0Kdn19NibLRp72
nHLRRWcMiCgG/+oNsImSr1PylhnjpfwXi/TTSrrRmPPTW7thT9bDBuzcbczaXFAT7vXUQMcprH13
JxBBPLxUbnpvqBYfykCNBy+oGU1GlEbAIeJfdk9DAP9/S+JD9OPpOnVCfHTzGATC8HjvtmOXipsV
3HVT3vrlydyuzVoqwOs6NMz83RKo7t86mXO01A+YGJAXzhbf+7ryCeHEkKdTLErD/5m2GXixPYZ7
nxRw+Z2sWDaVRSzX74OrVDnKpRPdd0kT7wIk5owcQq5KCUJoe+oBUjJuDRZs5qPwC2nQYm362MZb
cUPHizD7QF1sJeI0Y9Yns1DwGIsCKQJT2Y58tyChntFsHqrFqUcl/eTLkK2jy0xYonGsAfdDeS61
cCmS1PpgTit4PIQ3t7oL/X2c5wCV8c8XZ1SZ5LXKE51Rhhbm0yFgZ7EhiuSyBYzNJM/9+423GCvr
Z2AN9X2a5jtHROjGqR+E2VCxxZrg3uxqS07zbRgOjvfMQixhZOBwS91D4NOf1+EE/x6WWbkn0Xuv
1jQ+V2r4wa0IWiZrvGe+ZIagtDZas6eivuGMzCUAYPBrm31LBwkN9N3y/huliWnex2AXoPvWRQMg
TlObR7QUwZMS4Fwk8Q7QpKkNAZxwLR2/McSJnPHVq5TWrKiljvxxOX1UhN6XYoPYza4jrEP6h+2F
aCdI+vQY57H5lQwZpa6VsqLMaQfq44wZv2s48RwB0MWf3/apRaZWt+Whb7CLd4BcdkN2PEjBtiKT
RHhJHrA8zp0EyzMIF0uzT3prSz/V72xtUEWSmz36AxnHoAbuJUQeX/6H484jsVDCPq97Gc7AJm8H
u1w/5rKofJ4V7AS874xZd8W0QhP/rKNnq7h3gptcFOf6q7MSgAN/c9RrQQVFU73A060KDVTGk+Ci
RPSDV0g3OYNbP52ZEQfort/RT5RLrKB/ToaOnec9L6CFjXV99cCjEKby0Ry+c/FjBgNrCkpBjr5+
kMkV7kAj/zkG9FoowMRTGqY+tSAVgtJFilxZqwnxPLvVseh8asO2UVszyR7utgY3Dnj41gaFHQGo
Y8vLiC/1JWfX5BJl4hnsYEa4GEf3PDmJdLv8Yj3MEf4bpEt/PlYWpFQr6RwTo+tGvkyIkoMagsFi
n3hbDkZy0yJf6rJSFil5i59bYLHeckiue4lOeNQi1BHuD1bx1Nx6DvkBkcbOUG1ITgsbiaZRjp4G
+fH5a7h2/SOi798JnmYgooslVHRn9BrXzdoMed6tvHngaLGtOGQ6WG3EIxUojOH4H4MxPO2vmcmk
v8bolg0NZTgbj1XiggzYuV7Pl/5Rrwr5iWHWKpa2e/wx8FiYE8nU1am4erAduxSWklWKCnDHM2Uq
WoIjaNF6q+I0Rkpp6InKCTZYFp9Z7fR+kCxMmvoOu18JtU/Xqq1K87Ujh12Q5PqKnYfz6wZttgR4
E9cLFLxSO+Yvp3wZ4ASPm6sjWBPa7GQN1bFN+rDCPgCZRz3xI3RTT9QXC7AJUjis/E2iv6Aoa5Nr
4VUoFmiewUmWerxgBsiQ8DVD6xsoEqVj9luO2F0qZWBT7dCHcLgggTazL2w7lw5bx2sN62VhtjFm
PtFTyuZoTCW/wjCz2gxYOHRS58EY7vd3bUZsW157uPFWuMHS76GQkBIahZfjXzxtP6awME6iyl+6
MbfmjyFjDYwlO9Ujl0DTXcxKesUYlTwtHleCv9Z2+97lXofqc3tBSUrF0ulPYfCZfPgcpRgPTFN/
LXzdfp0j9uLzWcd34e3dTS02JgTQjrTpa0oJb5yeIsEnixW/oSExYqktz4GWRvYZIC2z83IkaFxt
4FQtwk09ljatdeNImH9s175IhuP/i51czQqeNVK8owususEIHD+ibGRwlgRiK5Fwe0vQ+nblIxv1
M/zbCb5PlU+5Top84QiVSt1LoXsizME39xfIHOo/rk+Bodd/hmtYMN+vDPV3sjJ0dyT3bwEAFAkR
q2BtAJY7w+tD9MPDMly6D9Rrq7A8Gj4nc3hlafAGTPQtmnxCElv2zixiFQhljNh8wff5JOOwoXgs
+MlEriQ9UdC+XaDH0P05EXE9ami8nzHpUpHWk6LzIumeXYHDSjf2xTVAlfNKyco6nMARYbjir00c
VruzpnhCFqnIW18pkB3y8uPrX8AX84FkfKsost0+8MysFhiH3m2NXulMzt655CjHhzERJNGSETdj
plCXF3ugteb1/LSURPBvzfu0S9iHOgpwxwCtWDlfjx9FXk298u+kneh3tasKv2utjvWcOiwTbHFM
UGDsUONGd2Sn84MIo7b8APfGwqMQ4o1+hO0P65jGG6ABP/+O5Zt7mhRllsfMI+K7VbZXag/Mm9Td
jdOXKMzjh9Qb9Fe2KVyV6E7GbpjyifkGuFzrmamSqpCxNwTDK41IuBaoOSJ3rTRuEIPVL1Wrb+YN
/hvl/gh08PZQa8QwUG8ZrTGuB8QVoOioUWaCk2Eqnl5LeNraxW1SRSf/9uF/NBGE5Ixrx4USH4DC
q2LYdcW5b+LWAqPEHIQs9owR45/Kej4OkB36+JW3/C2pOqkDi2xeR/YsmO87vFCXmwaONrFbrpg8
LLBDPNWlNWLgqD8uxx5V/xKohxBuR93xN6PZs8eIiINiMu+tVaQjO4b5tJhOheVO4q8TAS2u7aH5
iYTCIMCMJUY7q6KY8wSu21RQeo9BJaP2rMWAL34aYP8Jbsxjfb6OjPNrzS2th3IcVDyMcpdmVuY/
vsq/0yxZQP70nTAbwOQADK6zujU2nGoQcVnoy0mpxNQ7x3w6WBzzIZXUfECmUlBzxa64BcRGUb2S
Oak8cmAg754yDFiCAlBKSRHRC3mSPKgjTtUhpYUzWrHF+cUSVLEdn4K/gmPPPW3W/95fmIucSCCK
0TqsUQ0NwkOG5k0iooJOMJT/uNmEsvZYtOf5UkoGlFUiPNCFsI8g9roT51ZeK2rm4QkApe/ewg4/
QPVrfamhZl5AG/oWml7udMfNbU1edzS+p1drF7bBX1IlEErnCdscVa4Sr2f8WFO6rK4xlqcXs9TD
huVzNBHNmGqksYYxr2yu8CQqY7zTO06yjaWAzXy7MCQWPByWvxHaMXBO8lBCA+4/SGHAsDVbsnUq
wdvIBs25waOTRFrzO4sWn3BJSPpWoRVlvTVhMCOew7spSJPSxZPezJxWgJ186UAcZff0PNsA6OPr
vM4aNffvBm40acbvOIn0Zi21EHMjj9D3+2XxfgQ4kpqpDiL6gmt3XileredHMSjff6il3duHRAWO
OZ6aejS+fkRE12xLsOFnERMtPc5xOIM8t+U7to8jrNzyMz1TXYR4UWQ1RACT7J5YLgU9JCyYGX2z
nIbPCDxPvWe9CtMijCZt/fAGHRQMddwrzMDCT6yqq4eBxlm6ehxd+6201V4JwySNsqal4Amc9Mbq
GXwd7BFZ6fgSmhPdx55mPnP0gX4PjMFw48Hx6oFjpy3IHhwU+YiKWLh6Q90yV9sGJyHwKC57+m2Y
mTZbHm/FmecPTDlGlwCxXAqLA4LdlgN1pgMf3Wa2I8N0lfXqYsRfenohkhW4eLdBK5+Bn+5dYLDF
BHNY3dZdbnQY6giCqgt+vipZkBzZNsRu/MH4vVLsdYF7iIZ91EumMZemypckvr3bhb3g6f7paoKv
RgzTcMDUTne/izvcezg5nh8ohxmYA0xt92nW8Y685ZFZOoj3qetufp3VBAj+Jbu0AGx45foMIFU2
C7YWGaWHkoMNtkwIYpXZDrDogUKJ48/2BZ6pBnsK0WVK+67Y2cwwtgYyBwsWMPnF2dLTxkq0PBkZ
jEBRWXtwzxJuTVNnKAp0PG/Y2odEz5URLn45dYMjvsVDJVtlLynkkXM3QX40PQUdNkkywtTSwqK2
oq8nFpom5KLempAYyGWh7FrZhCQQPpdLnLzEY5j9xBFw46jYwRTBTcNtzQ7jMdJSFsihxxuJrwzS
etQvDOgc5XRrPD+9uOLUJ98v1aiG2IYbtcKtoq5r/5HF+SlYrJa7qN5Cr0xjbOweKBGhvG2rIw6B
XHm91H2H7VBX10vvuTTyTexJRZdj2V+0FicQVjC271drLM66czJ4q5mTC6FkQ5Z0knbFzBBRcQdc
yZ6Cn5H72ga2kADaTzt23UeAK1cN+TPaj/tbq2BPLD8lg6VTKJFtR6US55v8EVDF0EMwYcHs13Q4
AsXBMMjnPOSYWY+vpVhMNLRE1nIH6xBYYA7dbwrtT+KdATLS9e/V9PQdPH/LocyKSXpqcnWQIgzd
MbOSDPtB2JR4/6/gl7lQXo9IoED0LAo+BaWnvdR/F4OOGN3O4RsNov1wdo5egbguNQVOMO+7YFdI
h6GyZIBUpj01qnjkV8i1wwLqFoLfamDj6EbjgqaON6xuxIdzWLmucGD35we7Xo8ijMpJNTKzUXJo
pYKnIa8F8tPXcEFICTuG+6/zUtuuzhlsHz2O+M+/zxxSZ4JhWBekkjRYNbV2ttkf+rk+0+Q5kKxa
Xr/IkQ/Xpgy1kxHSKzJJzlhLFYzHmNhotMbFBK7p1u0TT4wqfudfpn9vxyBU6AOfavmk7KrHvUhz
XgrY+SlOvxKjeQtHIaDXt9qDMyXI5n67TIy1QiTzCND5F3OX2W/3z2tYaNNPE6CT88uwwNmGYMxc
sSe1eyfhxQ2867YXv2vX+8u/CWF3eprho8NXO2EOlVmB+cFbXX1Ru+uJSmTh8gK4g44Rjublmo2H
Z3Lv2hxrEnndCSjmopiIKW9tDIEmjRza/Lc22B6BL9hfuiAe535ok5OBIqRSsflEnBkwSiEOvp2f
OhMph3+ll33OgQWHeY8Y2b0Ylke72uC4hjt8NtnEE45qLlonMWWlA4CPyqlM34khqXI4PKc6ErPz
K25zcJsdSQVCNW4AfmZB+tNh7qbNWGarsOTYef4MNKMeBgvc1rHoSKPsAcqrnvvjvk+Tj0NzBBf6
C82hXJy7xCB+gkxR9jcfZ1I1Ts0XRemMeU+lfBcAVv5he7G15ibfA/ZSKr3CDctG/hjyf8Bpd1KN
VRexgGgyplPcOxF/55JxhsD23WE1zjGMUOmNDTR8wENbhyEaNgS0P+ItmdsiNYLGg58Ia+QRiZ8C
75YTWz66BgJObCfk72nz5qjBGo2kNLJk8EZSCteeDcgAoMFSt/mXOvK5LJuJoXohJOp8mX9vwDpj
21wWxLSg3E9wE4MxVu2aZKUF7zEqeZ2AiPutmHJ4g50/0H8+5MaRbcTkG+36xByZVORDDXDFaBQh
E1QYt9Nm9N8nFdwhpg/Kg9KkNBwzLGlSJPTUwjQQHwu1fcoD4oluO5sGfRE1BYTbqevAZ4H8+La3
h1h+mqJHqh5ry/jxRWyVl6Sc5F75ks7OfZq8/GVRqsFOpPj00/+slmVrNfYj58T2LAqPdIf39s/N
gfqTxjTUJ+p+eM3cMOpvZ15da/cgPIpv20/vz85YBCFtpAU1j/iJdVCRLxgYY2yKO02mIW9/CObG
uls7Y6iSsUd2fMonHzLmptkaJ4g+5lH7MGGBPVbG6zPOkSyp5dWNMeYPLdDEOa1i0rQ2woUsvX7e
CNr1HI4zCoEo/YfaQVmkmaOMRPvfxdDb/AjrpU8kzWIqhlH3HAUQMUV8L6yIHMfTC8GKznHHAKiQ
frafCL5F+IZop/bVzN+Jl04HPH1QnaT9ALMAuvCEUwOeTBCOxRpvgDiOlAe7Yrw+BdfhObcngAn7
m9XMycMx4HDsxms/lnLzg725a7s4aQ0aSxO7KuR0RShIum+TvflXsT7vF36kmlY2TihsnQ3o0H1Z
deNBRmCp5s4ScR9jVuZe2ahtMjzSpIdvStcGE+Mr7RrQWIGpRpjSJsjGAOWf0PkPvfge71yKeXcT
zxRIp8v91Uhrnq0UE3u0GSZLh2cv8s9ZVlfYSPA96+jr3zOmAq87TWykq0RtaS2YqdEMngB9Od0D
K3L9XSHD8aDLwd3OrrB1ZXlClA5XPqwHvLApdLAT9xV7B36EhX4u5UdrAQLs2IRDbpnlVV++10yK
4l0XRwU9QxdxLKqjRu3++kqc44/Wluta+s4rH/DsNtihryPpXtW2UHYHFcPzvV5+xZ744n02rp/8
QuOlET5/oNm5kHNFt86lwbJmdoYxAWPNIRUCDT9YCnDxgvuLVr1HfI/RsOAE/QZuj5FOL7Dh9FW7
yItyE5rJC5b9GBlEE6FHog6316nVMmM3GL7+3C51vJdKxzVRgM2jCrPg2IFFJ7RQy5cyvjIzhJIU
4QUwoME/xlyKj/1KjMuVnhvf0nK2G2Yqn5HoThdZXwcmAu80Chq/nW5HjCNy3a9UjbCQlaLt0tWk
boD/wE8ZfIXwynNDpessDwRoP1nVKL7LyKMyiW+n24z5r1JxvbaBGliJcUmRq77nPCoVIs+ugM2K
OOj0/h3BcnQIeMIk9dql32E3rEmTlq4gmK/g/4eBCo1Pn/heYZrDEl1E4T+KCQdTYJ3y6qj6+F1G
CpbVhVaPNTSy8ixteBH137hiiJvmZhpBfGD7wU41x7LXZ+r3Ye0iSxRwiZfEsxOA6bhfjo0NwPPP
DZSvXElzN0+Z1uNPAv3dt+ZCeii/PPmwruuo9xMpdKth/5+YfrG4Ix795ejVF9DpWckoT00voOK7
sZmpmDBe4bcp8jAu1rezJWE5P0bffvLjzsbiqDbPlbRXc6YMldj80LhI5F3rLZx0N7zGeesuQfZK
2S+P5FjRbXAhPQJVOwT1+Lnrn+6WXfslNIUnqMTktRFzqkc7lU9/3IG2gaQOtbSsE3edY94luyB3
HqbCx2UaBJHI23PQp55Cm4jAfK8beLgKcr9e2UEaW92zNFrbRRI6VTpa1d6iL1KJtbpSSwsLA149
+4U0KzO52VMR0i156JIVYa7Ya294if5VuQQPNUqGm8YIFi9M8eJ7Pw+mQW2P0VRmiXCKdy0B2aw1
3Gr76RTPapNlhP+uJd3MoppiJcfWsbPxsI2QJFlzIbipJBbFrQ0WechED2Z0M23eUHNCngDKvv/X
WDMlejCYYt+/5EEad+yBFRxIxXi4dZcsPME0vX3v7ATeacdpHS1VmPxEuajXiRQR7cixamd0d/8o
Dx+sgQxPFzvXr/Rq51ddAGG3rlObNy+3fFgmHl/7sl9R9LaJN0HeJExpliIDvN3PplqzhumT4975
ZgSe/enDvXTy2/esF+UXCPYbZMqX/eeSj0LsPadSezXYEgdaJrxtKGGAwN6ECmv/uQKthYHFPFIb
OmWs0ldcZfdpiL5V/oMW/qqWpDWJzQ7rDhoGpr8qjMqc4HK+towzITbYvmDZdr9haZ980s/5i5RD
xnR9vIXKrQECqYIGncG1G9ArLgkFHiiCol690ai0TlLEqqtcZoueEr0ZMUt9XPfPgGZ5godxh5um
9dCsOut+X9RsA5w8Kz7tsj04OLV205zUyKcWh6se1Judep7ZJnbIU2EojRBrl0yGFeKzkhtahO7r
trFkCBZlMvdLZAofa8DrZiV55mIX8xszdaUlUUhI08/T9pN3KQoNVJH0WIfgwe126gQ07x5gx7eV
rJ2JJTSEQsLHPuup++7w0aGNJogblVyGwDB45qXswd/VwE365fEmzbNilI0RQsMubMCRZ0Dwahhs
n3IjYgsYK3Yr2tTEKMC+CbGNoNvvUyeVnHDXX/CkDF2ndIvugprhlGXO3n5SE241VN/39ieYTVI9
mUdpPmGAtTd0A2qCkoWMnkxvdNXUnwwQ+UfE/hXrjWWWcaBrc11qUKP0vGTTZrqLP5+Pzrb4PM0Y
imPXg/fg6skcsBtXUmr+71aqy/47iVo01WZKBsXmFpVAWRoYuJjcscW26oBqcuAwW8BkHJNDGcyV
Wcvm0Bwnu/T/cgH0jelsFxRFS4Q1jedFCJvdJzfLlp5sK5/r2KalHVGIX5VYDbjMUCVKiDQVZ+wS
6XjxRv/q37+nfcJPD7kDRY/ZrK8UczdYxFurtzN1/JRceYgbNCMQv+GRXXP2xlZ5kzzMu5VAUgNI
jmAg2W7KmpoevQ5bqc9DvCNHegbP3csfETAzy9AzuNCDl7z1/VB52QiJRfxmGUcrBOqS7mPrxsyH
1wwa4Y+iK4ZN4Ty1DgPbxAY1Kh56EbravA2kAv8DOc7pi8DQpRBaopaFM1uLfIkDQOlse285p5ae
qNywVDEaFlqMNffs30JpaOLwaoyxmv48ox7+s8sfNEt0StnsZmUrqBB2ONwiw40ebP+ZA34LYJAO
Kl9XqTAkyC4CbEDrtMGBtdCR/TPrxvS1LaO0w6GCSm7jOxhFT6ddppmflgrvw6oA6+x06a1XC+aC
pnCUjQHgCr2I49VqBlJr5GyAUvXHHB8HKY1uV+u9gPgm+HMRQ4x+5IC2d/92ynGFxXLca52Y6ku1
fjmmvWmxIgP0k3U5nEjT+IahA0UCp6wy7+Cu9Zc5m6n88FOZsiLBovbqlSrXA0BRDqkKKPaUZaf5
VFjdHFBujIpxntI65ksH71B7yrNuOS8kuponaJMiOx3TaJEzeziIAHoIaogyumP1NkkKk4ogpvni
bRJ/I+2Vj/hZoEHtSC7LS8UmDPiMj7mvpzdUPHF2kJQzWQ4Wsks2fSoOebSbvaXShloU0bNLr9i5
ut/NCMBANaYJ7CyvJidXw0RI5UqTCMSoGzkPhoJETGPpz+t1tSE6c+/ynNAhweRnwk+0xpGgPO/d
Ycj+jB4xKV0QtR6ixdGV+dgtAhjoOkVmhtlBfXQIvAtBuXtOfgtfJg4wM71gPd+y+yP8i+6vwMNR
PIi4bWuA9V/KTyJS2JL+2WYXcmD6A4JoqC8w+WD4FetDAN/2hVb78NIg02U/Rnuozj+ViqASAZFa
rnwhdpWJRqAmJ6+NpkAb06+0DjQ8VxewnwhwlhR9y6eDckXL7q7JKCnFTMMeWxn1u21m5EDhDzAQ
16sFWYF/XdjokaDXDGqEjG2GPHakCFNFuvDAu0CVKxEghy2w60MkYFDPsnLv9HaRpqzp1PXdY8Ny
r5ZymBGtMbOvufeDngrIEvZu9fnQrS66RiQcni5d+7AtrHAsEODFG7SO3gfIS2EHpeZ3YKO4ZeAO
x7eBqgt6s4TmR/8xTSjgoZzcdWFcEL70PVzXqn3dmvVELeHrm9M1hv2gLAqKVviBScFdI0h45DtK
8g5ltCpJwN32/+Q7FIGX5jMj2iOkN7OhV1kI666c6uRqAafhj1aSPnu7lLfJbgV2Cb4GLWjUwjm7
HhW3wMalLjEMk4nwFuyyUoqJC7CvmBJLAD6cVc12OAPjBQalB04Rx15FYB6hW0oPSEQ7KpEv4//Z
V/FcGb9P+FMxJFbvDtaf1mv5tROrTGjoPAHhMlVhL9naTQ0EC3+VA5b8ONwOzOLpm/jmTfIgb9qx
ZUXz5v7Vy7cE7dfj+CoUUpE+r77tkk+1TCiHZAm0WXK8SQTul/P8K0Vey2raS48mre1O30o5GbjP
sv6XHTVn0gBTDZLWKc0qCGe1XZsflWlMfrNiHzdpgdT5iJbhkReyTDmN2t8EC8e4uf8+NII7cBKD
nkBHJngvQPbbnEM28zANSYiX/KT94Z+ft8mDpSGxk7ptXGeYxwx9dFqm3smoinLjxeLpmQ7ZNDoU
plgiaVMiOhHxfIwsvGKLWxogQqWaEafulDWYdpI6J9Wcnp65KdclQwyHf0Fdx8zLaL2vcV6bPTYw
e5O7oe1xV3W3UEEoHtoFVm9ExRmoSMtEZHchStt8ne/yCFJLuEfJ8UhBQeHzqVG12zZSXKNZQZFK
fhVnEkFu1CgEzLFD5DMKpSPvLKsE/bUyBTgCvogewzzecnS7von5D//k7NUba8MC1+NmyJ/+r+HA
LSh0myRJnv29RlNcHQVZKIil3epSVwKMTG7g5AAp8w02muWfi58MHVBLj6/L3lBsnc5FUBt8zPjY
S2xeMU/Lj4/H2r3E5BpB/Ik8CqzFLHXof3HpGxsOt7KEBPmqKDxoJbSgpJbVSamtRe5xZNtK4Med
O0LNApekHx41rMRbbyTq8pwEoaUHi4y7siB5/Bw/q8pw6ZbfPDCXbWza9gLfyLJB/t2uHHK9n5PO
nGcV00Y4W+O44keWB+OfZGTpp/3Th4RuFHVADJejZ5tU/nb4E9XnWQ/vwOJlBkPNbAjaeu9DqvY+
HTxbhTnB+S5fdqBkBVXFNvpF7TguKK9hK5jYtH5XlBSK0N2o3y9pNuGUCWuFr7vKP9I8b5iuh+HJ
OFkwxJ59VCSyB/kVL14TcQfE2BM+bvfGQeWLLYxqZiHBQuOKCQbHb05R4DkVBJ3JmPtU9UzSdmCF
fkUU6pi2AxPSfe69Mu8GxrCQOIi9nt4gq66Fc5r+XEhrBIeblvWRb83ud0lMlU7sj2LKuOMevrEM
TWtC4Vppn9948dVOjOOBbLy+mPdXSQAPxLuszlvruV4u/Xcp1LMhqRl1LILVRYbhnhY5L5JHKLl7
xMhA0n5wb1ae+GKTqqALdye13ij2RBYT/7s9DreMuFP9UDgMi/uKr2Y9h4gTZP3KqwmmiIfD24Rd
3+7ooEt7UOyp48Z8/YweqLA5ujllL97w+QNs29nXOq3C8oMeAXmm1b2qjK1mhOZufZf/p3ew9bQK
i4EBhqFaenu2cXsNfTicgKr/aEDOqMjJHhdtwpnj+OYCVAW9bhBTcZoleIsEHqt/mlD0+Xa9ZhMV
1pjlCa96G341rZkIAmTi5GPL99/RzZ5d3kk5tAaljeVmhFuxhRbOBHEmHYlRdDfes7fMM+a9UWZF
X/PN8biZCven4bMmOxNq3I20kxiV+3pfRdIVYZcHvzse+qneXq0BXq/SgP1rWkGxihZbf1gYv0mJ
AobHoU7b1fbfXrRfaGTUplySx7De6Oa4T0qorCYe5BAFHZdfsAvOK66/7y+MfOQeaQLbcPsSv5pc
JyoeVErayhmBYkSdmFlPUbGgZjOL1VjmtGyNZVs8lFDyUVqDxzB6GBwte+/PAuTuJ0Un986wnhwu
tkVluMp32gQJEaN3VDkhGGssKOouqZJ08L4yfpNKZBwP6UBwdVrH5ycW6K44RBpNFaN8im6zSSgC
3GvHc6/PA6EkhddfScLaWz+dbwaRyx899CBItnN58uVn+/jYqugidE3pqgqtGbnJwsoP4p115s0n
ArcRgHZ/sMhHmyBgIl+WZtDEyg0dm92agLvpUsw7nmm01vMUyf8jxhe+/FC5cAmwfihw50EVYTB5
wzQD4jrQFrkl322RDgbL0U9SsE6CAjSu1pmMqB/kpbCGRFAK4v+UB8bV6zXymz3sk4TXyStrPsLa
ZZmoxf/K6woLjDOvKLhedqJ65vRPeOZuNPmjgufG41PgzQS4UQD3p5FXd1p+xMZkUJLAnhGHBv5b
m5Ay0oG/aop4m4YYspxEqMgzS3gMUxF3dkk23HHZo+lsO9UuxjDV/wDUK6P46JWzBQmrprOWwDIE
SJ0hZ4KVC+usp3ssQ/xyvau1R5HhVkoLvftxadTlAbXxQdJghwlSpVqzNWdb8CqIxygwdDZuD+wj
6w57xSvc2UV7MyecyRkn9qrm86xDS+BT2N6ApSuMa25v72x0zN2093HYDUA1FbzPR1i7xBfhRGgZ
UJfuagcdQoJFaVtQf9DhnOO9gLFg2CqkmZ6sPv0SZtz9tBjkor4eQw5KiBVl1ts3kp1aRmiMafTr
nA4xXbilE63HimipNXUHHHV6lLyJEN6NxTXUvR1uD0ACsuz0FDHhLPzOH9lTXhXjl2YPkc4Hh+/g
RK7ItpNd1trxRQl0VoOm2IWHtG64KhcOrnZJcMpgRPY4Jxjy38/EZfnqxd7CDSuAhrLvLt3iAqdA
yYmP012X7zgvsHi/zy1kcNpo5mMWyC+//avrRprQBHR5TkU0vK7l6RwrieUGoADRVA/B1LAUTzRy
83JX7KJI2GWBfl7JPrXeupPc6ODvdUpIcWusVQ8pBkBKTdcSLdKGKos0W0JosfLPWjDqOH4or6s7
z7UGTFaxKo0USq4LMGoZMiW3fmUuhmaVV+y79sNxVLJBNFDm7HoF0BD0hXfnNmD1Jj7Wf5XCDVfr
Fsme7W1pwUuXKlOEuwZBGQ1A0xB6PlTlg4GcOg/75uJXb82TyWI5JeDUjEm/703eDy+F3ZCHItrd
DlMZj7fWpT50UaNIOhDhBXdyk3A39yYkT4wNyAD+ZhxTFS4y9eOmH5AeNn+ybpXu7xTEUhcLwjgD
M2PrIeKtD0wiDPdhjdDA+GC8nJaCvy0dXg3DjMmZbXZI4eg5zwTBDckd3SojpubcKcYGHluSRuSX
DOGee5p1S8QA2hNL1ysB8lDEeJqjihMXeLwFPWmdgWYEPtDvpnnfnbnfKtPxuGaOOQkZlzqm0UtD
6euKpz2DCvL/2GKhQZ3zBG0rlIpBdMgLwXFspOcZ+rXaf28i/Km0JO51vWHr3E7WM3L0ABgzfZu5
hYcH7o8hvfFNVJF/XgoAlO0jA+r+QMPR8l53KOXJI31SuUfqTV7AcM1dHHlZFQB+5CEG1PrUCnrk
bzfalmK5wlqAv6+vMjc+K/0YXOLsUDm06AO2Tve1uKt6RNsJ49P2F+/8wWy1zO7DBZ50qww+9vVK
Y4aknwCTDg0/t2chGoekGXKp12VIziYtHly6Dt7rsSskQVZYzkIABcPTw11EvvL9JN9cAbF86gNB
hYmLb0/vF0QFB9al65BNyVhBiChqmebW74TLoWY0s+zGbBLSFxpjizDFAYe7SBMpycaiNpfo5DBU
NAk7KItHsdoULVCinGgNoBQY0mH+0OBkIBYi7AmKl8qcEydz4dOez4mrE0aUh+JjISSr/4RRzKq1
E3RxGYzZ89YIMLJhLiIAy1UjhZKSyh+2vwfmYjLfKmSxRPQYiWvcCjyrPf+lJVZPx7obUeI7AD3A
1ZdNOws03WP6t3gabXZJDS6GkKfCsvPxaDzP5Qv0LYN0XKvITmZhN98kiOh1VmeZRKExafe85cuU
SYZKgqnJJFZseKEoWiFhK9T/s+gsMmWU2PesnoKeKiy+yThq0mDZ5b51pdwb4WOpnowcYCfrvjmL
UVQ9Sil5DT6DnayyKPGbVXU+sgWLDksGuvDFPpM2j59cVL7RaI8NmCUPfNA4BYtqU+A4aR4WiNyX
l9hE7lCFM8RIZFhbHyqt2ARUs1jQgOydq4g+XA7ydNxJXNaImc5oyhUNv09MqrgD5xyfXjg3bPMa
yQoGGBmM/zzTYLVJ3tsJ0fUyMfKg3P3WvHqbc42zWqFR0pQAn2FwehJon4DWbrqjFhOTrtpANnaE
EuavMS1Kkz+0te8e8WbMPx1ilcT8lEgfHnJHvHwhyiMW54rWpsjtKzEf8cKxTdFv/XvSKo9CcsTB
GD6XUWLD7zUCsvAr49se226qqTR+HcD3eD/zmhQB469WxF222sDtjHaL2TcM83qBGByrPNYhkOq0
3ksVLALyskeTSfzaLWhHchyE6IKuQSsuafcac0W18tQFz76HjM1RHcTIqhAr/mMBb6Y44JBuPPyf
56h9eOH9HFkRd5Bm9k5LVKvKuU1ro3Kc50smD6G8VV0HjDcTAhDWk5VBGYGa/k09Xwtj/Iv2gWNX
oVfVdr1/EKAEpeJmDs8YSaTiZghXIsKMs9iOjAqD6WZsDILtGnrE7/dnkSpA79/tGu/DBeUMr3Ha
BrmEoenU/f85S/t3hQHaL5UcMWxNUS75t91rBe4Hv5iP2Dri7jlbYkRrjIuZB0HjTjezmGUmJOjL
NqXp99nrmUxPA2GuMME1UfdtlfzR+4Y/5Gg8N7rqUzqYZWL57JaZgbzcdRGknUE6/ZLbC5XYHo3c
XqHZorLFxy+ZvWnl6F1hasKTavdzw9H2rj+SPu77dP8nr0qE/1pJpM2MXYLwiT2Xk3sRQnsHVvlY
vqmGqlAA3uj9Eho0G6+nNUlRrz6107h9sIFfxWH/6/C37YqubLUt/IQaJ3KCBhXM4Vaupdbt8u3T
CNfX9/VaFQZ4J5yOLVsvSyeIM/DvMs3lUxCl1WyPnujXoeiogwlzAKddfJsym9xfPYztM8uwe0Dg
3WiR0xW9oTSOJ9z1NImCHvMsnDbdqg+of/g/p5sD+gW1Fz+MqwUaDSPiqFSm28CBIVGqDJbh1jmZ
I/4HFBRzkMvtOBvLFs+xVRphA7b0Qi3TNvusMEfnXT8lg2XckZz6Jfwhp05qREC+v4I/jYSJprPW
e5BB4H673vcosNummH+Nsf0B2/gzDz6PffTQmBzY/l1dLJQZYDnsnmslbOsdUfkAwHwxeuV9pSJd
FfxBYfBPaD/STK50VfAHHn361qVbR3mBqu/lGqO8NjbbbmO7260Uen3LgrUYhWxNFJnIPiCQN1cg
kwxpKlQJEbnB7KwKtLb2Kjj5X3/CHYJMs7x/FwnzLuNV8fR/LejfXbGwECR+fuTCEa32JXZLcSHb
gCSDSsrnrbCtgfpv1fwTPY6w8IdQsiVxA1E2QgE8IDXaDgglo3NPl8s8kDiDaPUXonrSYRINSust
tZ8T3eBiKWbA+tmR4w9m0dQ//UG8gYOqE+1/eAytTLv0jH3uxdhgOT/KzWMSmzCMkptpNIhOekZi
d1pCSK2h3f9Ae2fQoWs/flZUvZIdlp1KJC8iKgG7ZS/LjJwxB/Yr/Kx/ZzzNtfMgBd+mGO27cRbS
AecWewcvs2qLwsQi4+xGyflD/nX3R01XDun2tuoJTXQwd5pSfU4b2fyEzDydAT9u38vz8Ao1GR/w
rhE8L2GzyVOBwD4qokGCF8wlZhaHw1ZLyyyp2amtP3xeyYgX9mPDcHLXnlIT7WcMQSkcYPxCn6d2
T3nJ53uXHFkaJq418GNCbXbZYpiysP6igjIpams/Vse10tAHtNl5EwSXmTb9bgtjtm2Qn67WUpfr
Y79xgQXrkZJM4yCpXzrAzN94ZDy6o8lzMY71WHQDLVAiaJhcSAbmVdhIGlNHTc5iWBBXsmp80PbE
//lFGsAwcM7CkKLQUDHkidWRGUzNM6wABFUO1FP23zciD7OMuUc6thkd+TC01y3J9tlq/CBSpKw0
LsnfTnfxDUgKObp4zMcsREy/Md5W9aIPtNNqb5UyoPxRHOWIfNZrrLwKPrbOEPPhZMv24FS3FE6D
lJyxQPDi0EWUD30kbLDYfCM00lU7mhtBrjCNtjbU8k55BVBBTr7i9SMSqfDR1Em2zJj5vqFHl7Fj
HysJizke5b6WeIOY97V+BpV9pV1/jUn0MATXEq4thQK2CM7fqGxwU9cDgjCnBRCpoA9ttJqR/gpW
+KAGoH+chgR839/x5+CJI+ma9MTee68QRI3hUOOorb10h+IReAegTCsyw2vnQx5UibkshKCmblY4
WMQ2TJ9NristUL5Wz0/2oYaNpe6oRz3GETvaiWvFNiwxog48vW46MgEOVeJbeQy5WMCb3lDGg3aT
oAZ7xjfsaWTYVnjtAr0IFdvzA/na337LNNgdKcp0aJ0rFmiqOEEVzxfeNJZ9WkKWEwpwpcEU+kNy
t9+/GnAbPziZ8lFfGByNj9dZ6Vg5F+is+29XB71iEQMjHNOXLriH2m5wFfT+AvWZsh2jROpkMuPd
Gsk3l38kyIQRyGaD8hRaek3Odj6Xhc91yI2v2xICKIzM8DCqGcvHtYmHjCGfxlvkYRfCxM96ehk9
v/s7AFiCfkOYiZpIVNkDPNbzgBDMhc6cjKqfuiYsnNPoAP7S37PA1JsSdTD8r+a6+xZYM+t++IFI
6ukCBFPclZLgPgbre4WmUdGInOZlTn+7LxS2dm7b4lbsc6xhX7+Z0n1eBXMeuVDjE8s2RwvBBSiA
JBzP/v03d/HfVZrRdLjIP2jmTnJIVpwOVGX0JkRuL4Vj9P+dbc2X2Gi4m1ES1xcXCxqzrRZfDVmw
Ke+OITlIsfUJ+OwEt7M36ItMpPMqOylkWqIPetlti4DmyoiPvlMFHiGtjTe1w0Y/qyMqP79tEdvo
s9LX9D+N5b0P+VOXhStBQVUXsR9lyqwHt9zX5WWwyJApfgMw3CvfroV5o/KQCI+moHOV7uXRLcY/
GI7pOvPf22+su+g6ONL0Iw425/AdpVOFN+nS2euVCL2uctBRde7WCjH8WIykEQK9jqqyYl1c3TfS
iTGHMl0KMBKhzL1mtyFeH6MNRA0fKWYvQ7nF12wg20N80n+MYSN3M961s6tYe/5aw0Fh1DLkbnIa
OyvOR2exnMsEuN6YSpSFjBC8f7PH4S8M4mGvxgfiDFykyeWzunCdwrOkb//Ak/nHKJySju/R9lzK
cBl7fp3ZCtVLrrGKjIHBnyXPwDH8+kuAkKYzsBQtsKfmlARxQQO1Tq7ot/A00H86kUABNvvikZ08
mWgNyM29uYn0RDn4LnFq9SJ2xA142+f7JQ4qJLMCeT9qngQWbj5ozfE9U/7oPilfSaxmlM5dcthb
U64M6b5YZB6FteT61MSiomFBvQHFyN6ZlMmcyZ7PppgUC/6CsSiDW/Zu9hLWZkyxrptHbVBWxwsx
9kW2O3oc+GnMsOVfKGZ2GoxQEMHi7Bhbxqtuv4I1gbp4RsV46PLSmIvRs7a9FR4If8c4iltpCcPk
rMPpZOWskLbYJd82+hx43YRuRDtRqfLEgsvAqTBwupYy7uGPlEVwZ7gmdlwX2PYGoJbEsNZ+E6d7
3Nh+WqB5XOLkjdGqmdAyg7UQUJJftgaDQB7roRU74Ggk15lhsAc3uTm5mp+39ESwGXurniHDvFTI
jTd31fFe07flw7bVY57NTM+GRLR914iKFGTArXIm0k2M3ou1m3B/dgQObWQcIRoIFf3n1/lENyTU
+ohsSYJlnuNBLR0x95xtxvh65SdYRJjKZGJOl3R2F8oKTpdguJSOR/ooPd6otyvTLS+aD5MULuhh
GCbn+PS9vVciQ/Ut2SPHs7WlA9UOxJayQpJg1dSiN/8xds/WqIIOniX7Viy2J7Gu4ssEKBBW+mYo
hpGqfj0SzTruIe7CvASG/axd8T6+NsJCN1bV7k4imZvYl1ab2E8jRnVQk7rdl2VebS2gyAj7yNEi
ufB5k5sjex/iESsLmO4Q1WAEtE7d5srXct4yCqTX4SMD1Y48W3aBW2cIw6emGR8d34wY70xkMsgj
G6dKC1r8eSmNvwGKIGYPQoRJI1I942LhI2beFao/kyxrbr7FDYOk/3iQA5R2rCES6vdCKOSQ9u0E
TnAru/jA8sLT0xYOFz+IzzVrDb+ZTChEuIjgCK1JMMBVPZt8JjMf34QrSXF2aGPMIA+pK23oXW1k
XvalVV3oP2gux351L0b5OeoSxcHmH/z2Mk79+/7C2ROwyquZ9835zuAU4hYjyXTL8Ck6BUtKnqL1
bugMU+0JlTzdoZveVp2B7gFrUYKuwv8PAxaf62KDuNDeuR0RgY0yU+oEjhZTpVWamP4Qc5XsYy7s
VISicgaQqJYirjpgw38o98kEAzJglrE8ybDJJnYSF1xl42ZuVZb2bmmmsXfaQgPpSM7NBHyN7hpy
EcJXR0xEr9GLBQ6E/wh+mVRdPFQPzoHY8J9eMSc/uZm7u7ErucBGZxipKPhao91ayVF0rhM2ggbS
2hxsS2meH9Y6FIK73tg0+i2c+s4WShvumvheyE6T1388q3dFjdZzFvpSskrf6QuQBhGXuAA/OdH5
TP9fAf02XkKyWkZAL52M34s4K6e+QuU9wrTNveBHSZ7snJ+Wm4y5O9AN7fnW1yKnTWdOFuc3LNTu
MB3UPVi7+rN0iCH+4L4jlpk0Hek9EogwCzMOLLG7tTq32YX1uYjw19o+re6UNimyK+j+A5jzYC1I
VAdFJBqTxRQeJeycVssQe05Pl2vQOer05U+5CX5pOHaU0l4zm6XSqTU7ge22j6WGeN03c5v9mdze
9ZJN7D9Tjkm1JO4E+t+yGWnx1lkeeYKwYkHON6VEr3Kta5vGVnKsBeKr5xpI7yjiCNmk5f5C/wHJ
49EXei2RdDgf4/vRL/e9AY4mwXfG66ixCuHwhRJzBUrKrFQ0Pg2wMn74wvSrKvSx1DUbYqWei/7K
9Ilsiyx7gFKxAg9HlRxoS/BKGcEXO3wGS+Sgy82YYoiW6+trqlkkVykiOYixfT96SXofwCfAqWUj
SPeCg7nUywVKdujunUA1Xvowh+eRGn+8SUp8Rjlv28iJpDaiJESv0LXg0Zrok5ImvQpIKZs5q/X/
j0OXlsYsbdzVXiVpJsvJbeTCMJystLtJNfi6rO68J/WnGFcGfezqZoR/aEXw6i/Bfmk6dhdSVh1L
RmtP/4hZfeOa+TSwvthFBTjNIQ80qOJCGXbARCNMtjXZ47n0HGgFLWv+1mgsVogimVP3U8rdihyU
AyxhF4bDSBphlMAgjGMsqQ+dSKxCe04ESnMAEbZ8TvDAwDNydZwqPpcvkVb8wSE2oiy//5ps1kn3
bMHfRWCT12cQMZIDvZfoG3mR8+C5ur6uFJQLNVsKSZtZ/LSefbDOGgUokeMhwc/7PB2FEaUAy5q4
Qiw416Tg+xNQO/tofHgr/5kXdbR8A1gCAm9nPC8APU6eS5Yiyi6M665Hj3Ij49d4BMtw0TUlnhTZ
gzfJru9x6XqWoW7hasmQIx14KuSoDrCwnq/PMRXBBHTQ4b5kptTX63CBQm6iIxdb2lpS4AT19TaH
JS8kLRZLPNvMnvq5CbKXVmFFm23DyLVilzlLY11yzTI0UYpqZbEVk6O9aluak7LWW6QLdNKOJKE0
Sa3Kawn9KOCwoQhp/7oDgdx6tB9TqkKupCwtuEiKIFqtrIv/Xf9MouD74+RXYfm0Zu4iX8hO4fwR
yMKP48z1Ye3YQDFsG6Y4d/tEMje7XMM9b2qKzcOrsT7ni/7/BmpKYY4E7NUyYyFYaZz2Mb7K4PeK
GH/6SYuI6WuRIn2FkQKsLaaOsIvxqaUUpwh7azi6XdIbeMTg27RYpLkrX59Qo4jQXkiPXnryhu8q
Z4OA8PcGc6Tc9ul9Br82cVjFq3+f/pnbd1ZFJak88p9u5PiTqcMCbxlzhmgZoMfrfJ+mpYLUJpFw
fEwUjCbvvpz//R1tur3lzYMKGm8/TqY9/OFFXYjR5DD0gN47frnBm4CTYvsg5rEoBS/Fu3STkCle
0AGo6IDBf97lmYm1UheRVnl+ntMpHMwWLj+3iVGqUv86/Qw/Ib6yXGDCxlgjVdx1Tv9DoeCkBNc/
gyuCQLd+5EENju1EN8rZ4eGtZLL5ziESynIUnZswUy7Leaqy+AaluKyGZmsoqdRIirsWuIQfgSVq
BpQgvRyTmKqxvVxTTbhwIfWwSb0qH3YEsWTDujIZwt4mfIPzpeoXtHe0UYwf0Ans8Ovq6Gg+v5R7
DATpWpUoFHz3bsz1avB5m7c8LpeiBrskXIHbY6DtOvLYNz9DyZOdknxZzD7i5m+TaUgssPpKup5b
MerVsiL2kE76rD3ESjKl44j3tYCiDsOAa/noCRT4/1rXqrEdYcKZjFHo0g7FCRF0CDnD36zcDLFX
7VqgNoIS7sViqC0dLL9QvnaxFdFFwQ2FiczdjDsxtnDedR5Lm8OHhhGgSknI+ZE5cH6Pc7hSuY1N
uix+U8L3GTsuTKydyugoctQAOv8AEY1CNh5/3TOUt2it5MLtzaxftuiwHj0ahzYUUBjWloc33sag
2EO7aDAXYuW5Xe3/ARrK2pTOde9G/LSjdgpNtBwOSZBZ+APlCApEdK4AEpdGZC91/AiZ7R0pCRuE
+IxHrHsMh58Kf/KNQ1kQ4JQFNgFew1wkKJufm5G72tiaLgvympXQdaBlqpaSqODJZ63raJsePjls
iYZt7hZHu2ZCjB/5da93m4C36ET1vYD2nkICsZgtORUKpELAXRfWN7wP9NTbnMi7ALDcRLEelKzU
FpW+MDUzF7tlOtajQZ+qxB8KaMLocwmcwStkhJlPO7JVtcqDZ+T+3UzI1ZmhP7hBDMw3xrQsw+h1
vFgAc7LufLtbJcZsDHxdoYoeKEhuXnZUhgTealphVMO+9Chlft4pYK2QNveOUcFH1aGjQ/FLcZO1
7CCL2OoEvCQitPo31Y0AkodTSG+etUifnrRjxEjPD9HHH5BMcFoPL85+IYEYkFRBDpFyNbJ5JTBz
xRUTGWgPqQJnBruMQjBPKs6ZD6Aj1Ud9IEbZVJ9HCiUx7VVcxUddvY6IrwAGsrvVmeGgB4MLJFR6
F9sVrnnfrdq7EEFW2PV+rlTAopUO9ajHql2KXtbo0sCVWPi4LmoWrc5pvX21BoiXoFUhbw89iVNJ
OE2H2EnWw1NrOqDdm5pexqAmcNMibajJ5LuNX5qgYK752wCJYgOgG5zuXKl785Myo0FwUI4ACq+k
/6aUFwKFnatY35SUx13K3MrlwwuH05Wq3gcWIo1KZr7kgADVN5k9awHHAU5KluG+SE6hbwDGwg2K
yGhxZlmswamFJFu7MLH5HUFNWG5sJ59NHTSVtlce014MZj9vZeih+eg/WP+oAEIhHgNIaCgO8/T8
kZOVcgtYF3Vgw4nM0y78XiAEG8CZvx+1JxG66ILgFQc6nZdyTk4786Y3d31JeRdj3WYVvr2k6tSn
vKmSc/eGzoo5jlbS4bi2B2dbcO0kywb0jmBaE6IJge/EboCbmXPSRhyOJAH/44HViOT78KOgwx1Y
lz/rxRVWEP/StwOMDL6xXK60B+0aQ0olzQy7gsO9nUnHUqRsPK5XjAQ18KrSiRlTymTieWAXnKWu
6IrzKvqrb7eOGvW9bsLdiSFRVzRor3O7YUUI9vGaEHHtSiu+lC1omxws037FLSOBfm8zoonT1zNe
ierQi2rZXHv2v0NPnUnNKmtAf0xD+mo8Zzdxl34F5wq5miFOYdnEhzmvDVZlYXs+0thomICm7FTn
J3yfq3/vNJqcFnBCUOJ7/tdgU5WL24STJ/De7s2r1oTgbt1GQ2gaWNTMtqjGc8pXyHD7YSWkVb7B
I4JouYSVgT28eGTC/qGO9GFxw21fEf+hX4DyFdn/UKuBKnL1gF1M1cy1ITiWFs2lkT6mKT4LBK7m
OCbLl4Vb9+JjYpEPQjzu8N0bWDDBRbDbajPYjzkPp9CHbYPttd5pf7+Q8dogX7fAdpo9pPM1t40C
8ZfutZqyrQv6SDbRiZLh1eKQO7fuyDYnOGl0jDkygQpDSKZeyGwxznWvyjDH1GsDgJD39NbGXgG6
yiuQdQLz65poDoShotBB2bw3BfnclFHFCehMjUWVqm+zBvvpw3OXh7qMtvb4NadIVHp6xxtkh2oz
qzDqT8nBfDfUPC47+tFKKthfySMF5SqJNPqJ2m0c6VybxEnOvpDlhqt18Okbo0IAQjXUeJMUj2z0
0Y7AnuU/Og/3efVw2Gux+CLpziC61GqpsKieFLyirig32K7weigDJjXzpi5N0WFaxjuQCtqPseT5
KpxcVJlYttG+QEKJsnUpro0b7CMqiYy+w7i0nsc2y8VFKaYBQ7IZ01Gyzm3qQ3npXnxepvxcbrUx
rs4bJDl7728LAY9+LeQPT7MvmAVmjocQIRfzrvN4CaHf/C+tcoUcBjqrM0bxzo03cnQ0J6V01VKy
8xrtxBYBZvuRVqfCB1lR4VWAc7JA5LrHt/VJURuXu14y1NDLS03siOmZzmttKwmu3wfmrMi/9xwV
w6/aOxxyqFAbSZfdbVPCx17FD12mWbseZgLc7k8Jvl4OmwwcWpGuY6GR1eN8k5VEYMIjPza9TeGe
R32/+0zQShMirvMKgHXNet7HpxFqOocmchoQDebGTrvRVENukJeqTvMFrLIp9h1yMlksztq6ZLJw
hT98/YxXufRUJK8qc/zMWxJ4cbE/9q8JKG0+0Y7thPM7bi5KGL2F4hk6ycZMheJMik03ocxfPsqU
Kg6e4bAaGbRw7BOZVUy2+oqbxk7ibeFTe+yOsA59HuL/29wn+JUrkGsQ0Oxk+jCrcWObKUOl9pJF
TmgGFSFkXsMaNMMoXHzeAvIhDlCCOB9rfc09h9V12cjsL9aiiyqRgIPtlEIYtYUCVNNSmwnVMLSj
cVpTjvVPvnDlFjt9LwfbmGvjkbHTdl+SggrDz+hBDrY+myRXDz11BtAJOIcXc14JJv3jvHkwg9ZP
HjJr1GMubjhUSRQ9ZgNFqvkhsCwfwWxATHI+ETw4h/5vJjrL6MsR/6WbWqM3llT1Jf1XjbJvNilF
u0OSyJfVzN4CRABEaG4QAMo3LdMB7/5m2ZPURSjlpoVJyiNOp8nW47AxcIDn8DkDPb8hiYbkLMWn
BapDShgzZxp3dvHYKMxaCmt3Jr/vvALFOAHQwCWqF8m2usA0x9FPrtsMTJRBbHyUsuAkpIFsvc3L
qzJJaHyPQkCjwu8oZqL5b64mEh4L9r4eU97V/EFokOXt31qgcyWOEbre+iAkYP3IFQqHZZ1/JLLE
yHh1XKKDOFvVlMWrp31JgyrQNcg1m3r1D4NxGJWoLkuzf4mIYO0xAHTQzoNeJ47KZotI/dhYK4v0
V8Us1DCE+RVbzveW1rTglulth7GGqdOzgoOVd/35j0xz01Z0toegjMOVk9YpVmkmZ/3OmxcLNsof
uilQQxNyQ4qf+abIi7CUsD5u85d/rhglGutshJlUcfY/CwmzDpCakqaOo2zaLReDyBVVhGlUvBmS
nNHSuUS7p/WgXR/nYCJYojnXfefRKvBad/C398LsA6gGz5g0jwdBAiQAA877Eis27umViEHT33Dr
aNZ3+r3t6o9sZLBHDwQFe2eQ/AdzCXd4U6C4YJZHqU+kduhzWX9d/eTyIHs5mlP7jnhI4WZUyY+4
iqNcySC5yVoxBIrkv4EFbVq4XVDMsbDeCS+vwwDgTvanGr6CKuEJFi9wGjBqlKMFvpFWzSHwDnaB
K0ldwL9+U6Iz/P95gADuw7a8z12ko9Zv4QBB2yijGtd0mlrzvD0I8ajT3tZVgaEaCZPk/OuHbkPf
mM7yoVWDwFeqBw5K1JypClr9JgMuvl/EwGKTeNENlfrPtBSGHaSN3ApB0e0FqpWbJ4lMD6ZBwlRl
jSk70U2vDcKXRe8gL+M/M5A1ZBUEIOl/xmYrcg4Epk+IE8Rg48g/t/IqDGYgJxjZQQKHH9mxW7VF
JdaD5dLIcK8t2pNEY4V/qZZ8nqgVG2ypxaQ5WXDHGe1HnG3uRlCctTLgeyvP1ZvLCQyZOXtzrgNt
bsBcsqtKhMahNuOvVCy1XDnmnyEXgtiS1XJ4cfJIiA4NGivUqBMZI54toxywYWYiGs3/fPVf7Tw9
BmQaotm5cc113LSxZrZG8va7rAKRqZLxDDKIc+W3VfEM9dSInMkLvMYaDdJb/3twhEYqC5t7UrUN
Z3qZ8ZdyIhbNCWaKy8Z875tvXxHhw0nOpsfpjJyZz5q/yvLHtEQqpgrPG7bZnwjUi97OCMEDe3V1
EeV9bZFlDB/CarF+b139uovzn8gekjthMOUObq44+KeP8RLSw0qUvcpaJweIl6nfaZbrK+NMkyct
U3HJl6YkN8Vng8daxH4xC8T2x+Y7eRj1y18p7I74f4Xi3Fkwt9iTFUqj/PGIcD+Af/ak0Nb4cXhy
oSNJbRZhO557RwjDVt/NVuu6qorQgISgNzyvrFY2Xy3Zs67yRYbJb3WmKlw5F5rUpIJACJSx/Rtd
3TPBQTymDRavq7Z3PjRJ2H4cei4vdYjbi6Dm3olA6Daq1NVhpCOf1G61p/Ev7VjdE4L30GeQK6Hk
5diQVqKF+kuFR8CodfCw6dXxK5/J0orDWuZD7UHQdW9zBaZsIuSebXS8zx5O4flN+RRqERz0VbU+
9ePDkrTfFPZjC/W1thZbTYYPCV22wse8eDVHbWQ5ebA9O802hGg2KqpwDgwUlBKYfsIcxfP1jLJh
3ttNb2O6H1pAFg7VIGLxmSh5WKXvKl6PDTX1h6IgUNnrtExSADcwtcYT/j4yv8Gh+PbetO54rguD
/rVLD51WKxJgBfGz+iE0e7oKPLQvJM12Wkn7yWtVn6NCGf/aQlWqLrN5+nzVTW+tKIZpI/b0uC7z
+NvMWimGXMeaEbaiLr/hiU6cfLnnvh2mi3Q1R6OE7UoQ5wzO1wqKdywMNRhuonrgg7VtwjqCEGAb
ydqckmTTDJ1iyq9hcNv/hlrIrkTOkL4zEoIxawsHLg6imO9Y0MQvMsWQCIBhkCcIZ/nQIyTx7mTk
uPXuZYvoXso0bt4S9/2ANtvkPrWQhEobrHcgi0ZBmeHq3qnuZ4lE6Gt4TH5VdCihuUiD8FnOj5pz
qoqcrw3z69Weoe3/EsDwcpuPLVro2s8ggkec6/9eUK0etAhMPLobDRev7lGQ9HsdcE1dV+kEzVU/
fXLBZZus1xeG5J7Gzkw5RWFEm7Pq9Bo1DoDhbeocf9XuzHthoRKKRs3k0ifmqwlP67zsJroNTU0q
Lhmufcm8oEodUQn+OyAR+Q5hs/0nJYIyd1JJ9J3g8Xh3UYMOg+gG1heS0HnK/dEfMgBHRi5/YEFD
ocfU2L8SLCMeGZ683inxAwnYRD+2SL+eQ4s4GKJ6+D8uPm0n+g3tzGTTDO4+/QXz5q7yrgduijiw
0HWUfnYJ0Cie5pGjAZhnalPNs5iLOH47j0Nt5EAt91v0Pp7+gS6d9mHhZ4O4z20INJ1fbwaOUiHS
L1Clv9diFTAAURftScBGrRJtFeMDEXLYLSmaD9nhb3Tt7ThC5YEo6an3b8v4gWx3JOxAISvnZunE
9S75ojo10zWFWEepH7VTP3Fkcwn+J0TZ2qqJzD0yZVJ5t2481zB4X+pkBQL4vgGgzHh6DL2zkiSD
ZjBbzm5Pm+Lsr9KU2n3OjBxtwbzHXxbFrB4TgGM3bhTOUtJt3/y5dM3SNaOLU+bImSu6AZVWTEbU
atmuk+saL1D1/9ZmB50+7SXrIDEIDFq0ktV1KOaSSoEQrr2QGV3aPgqKYwFc18H7gdwXj0K639MK
PNJiyzSOoIPPBq7lm3bAfBO0dIG3LmGWkx5eCao8H9z1ta1ioJc8TBYyzM0IjrPIm3U5H1jxovuO
qHSHCf+bXxwZj9YWx2HyEq3jglXtOvemIAZBv1rMUbKO84HVt65bxVVq2z312+TU7pDykbXD2Cfl
+31j0/tPj9Ivx034vqLxapv7+KGWtlb+47IgLukf8Xfd1UJJ7u//nmpkmCLnlasf3i/D/fANxeSU
+kmUMThrIsPS8yIrTdw+zoBZy+ZqBH1/NaeEQxdOQahjGeso3weHzp96SUtSMRdCY5e0Zijk2E3Q
+EJfTwzXPTEkAHZzjv0rCzNKAhAt7R0P0in6tt+shCHhQSt5uCnJ8qHS6u8IBAi88A5DXsukWdqv
K05Bxv/kpSoKsxWkmNNOvlbBTelSOkuJKoh7kaRAvH9llfWTwJ+9t29mm4PwEHTEaQpKE8rsEcY6
77iS+pEbA6SrUohu9yrX9s3e8nkH7T7oSyJbOwfcEbhRU1Iqpi52jSDWKq6YXEqwVFPsRs2CRj3G
3JLCzzdookEIljAOSbCrhjlmtmsOKcALmgBrVUy2l5OxF6BQHLhMuU+oLDJVdeqdz0gBTNDpvWNe
NHYIAca/BAf5Dxv98KjI60jJFojEGoupb7csSF4vE/qXjRWbKKKkPSZivjCrYklkf7Apux/UP+tk
cegFsyi1Ow4AMyB8th5TvdVNM+BwR3fhLPDVRhj8d+o6zLEsSmIK+Y65IbISxhikCGmuKrXaURyh
x0bw9dN+kCMq0KyR9k5lIC+Mjoc2PKN/Ks/Nlslqn7TmjjBhkEMuo/L6i/peIosXWbC2U3rHCkB9
L9aePA8usslvT2QRQhB8PtZ637puFFtJ038fMllVbKXoyVBK6OZTx1LCs4FIaoo50cuxPvEVq/Ot
v9sH8Qg+CB8uqn8M124/Opl44kXplJJWpV7sdhcocSQxpiLfAGIaWLszdsKxZiCbSh1VJABZJ2Bh
kroX6N0MZR57a1kLXAqZhjpIcOg7QWDqbj/ZZf+mStBXMo0qpvXTKMJ5+dddJVJtUNlzvzF5GclY
ByO+8aWWqRzDrHNnxq8cq0OW9Pej+Hx5W4x4UXS4qLvVHLcgLuN6Hs0jj1A+37TWYcPZN1TloXov
HsDL/RyTnzwx5+cY2RoZLBIvA6aMkH7WT5KFXZ9kQmEo3jipPo7djTW/ggkgkbbtWUa4KIjQS0to
RQdj/F9pQelG96Ryjq0EPOJOJkcC4iqGjHzRuna6eS8P5pjxZNdGHANsax4VWYXI+i2FGTVwvDi7
ccOgaW2wRUlszxNnEbkc4jiD2FrOSBlFJaiTKgIuM+ztSW8+dOwmodAOn/ioMIfqqM/UdLiUUQnT
Bq71G9yt1SI88lfwMvUFecx/6yUNufBb8OzI4dZ0VELQr9PLCbNjpY2xOyHAQ0ZfWkUMtA0rsOzr
hUfjKzDdIbt+vfTLY/YotDGOx7xvGMOf5ouct2VJiT9W/uYbQ8JAXW6mwYQovy12NdjELvYFJT2i
BuvqJ9fEY6z1S+duGLqlZZu1CU6Hc09jOlzKBd3xQo/gPIlYwYPO+jQ/IgyxIDLggIoe+gSn4NAi
d3NSWvFzsZzNwLVlcAOxDqUD5ou3lISiF5RyoFpeZy28iSCUoX0esaGAOfm2rC9We1kZzNC9qLN/
ugwdnMIleWzNuVGdX3KPnVQnBh64XfmxCdVBMKa/6IHDIxmbC31a1RLdNASHWKloorKPoqY+08fp
j6CqqHAoXgzv9ah32bPujtYA+GO62x/iqkJKUZb1hAdPZI2xoae0Q7bt3CJLFHQue8vR1Qh24uUb
JHatEr113SzfKTLcGZ0uX2FHg3OPxykqCPoFxJlDSZ2Uzz4V5EUgLXcp2WmGtToalCYMKSSKCNCF
rileED0xsG6VP/mfv4Ftl7F4S1imhHOD9FaXUhnZa4rNKEu6FqjbX6/6DHkR1OKl7YgLloiRwV3F
ITXxk/XuyMaEYnIcF3+9S524hd1h+PSFNjCZS4AlxwAaqoKdT1alrPrQcFUhz28pkVfzVz5cD32p
138zXxBxPUWhYPzyhl52Z7NIVm+9lEyCCfiATdt5ENqeIWxBz8od3BC0fEIsKDQ094ADePXv/mFb
aUgLwqT6veLIgfKmRwR+SiyaHjAFgOmlo/yYDD2Bc/3LMUQ3nB6BcACtW847nzr32h8BtA2Txn66
yXRgEdoZLaprUv89uCCL19WruyGMHleqRZcYZVVFzxHEd4p07+RqFGo9NEHNjjIHLW1X3NO6xi4m
SjYRBdBPOkf45KKk3rA0OqPlay9fy2aAwGys0nJheUM9Qmfcue5AQ1c2R+wbA5Se1lEHbgLx+amq
qNmv0s0Us+tmRNZ3lSIF6CCi5A85eao379jknTsUhBVmXwEnXjXeQ3PnVMIctcES3RPDdyAe2bjH
z8BJ+KJHrebOtviaNTZK200rGXL7yS4LaEhpa4gpPZirTI3Ox7WaoeSphFEIelB2kY/2QZS9SQ64
qdgji3zIeIp+Yq+XVxvnVAbEbqvHvXvTLZ8sIr70oY+liir2hA66YyuLq12eWAsLVOd27OmPWChK
crcpx/DNW3DI9M45LoIiU47yoa9EIAUZR2392JuajboQebSdYknmM80AjPlq9jj8nQNnsNh/67KH
oD9Kc+f6u2qvA2AyFynMaK18sh0ink3bh4MrxiT0nx7lGgIdLg447SWHbyLUmPQf1k4r5LNwoepr
IXoenM6Tzg27JTepH16fFAaT2GdgBAjcUbmhvgNT97UTnYp2HHPV4PGEqvFwD/AcNpZxjMJsxpu7
pSRuWLRaHketjBD84aNxUJTQvqFrJE+OSzjzM+pc2Wu5tg1RwHK0vxMU1p+EsGccK4taDpfO19W7
1g1/EqVNfbdERh6O4LOB/4YtzQIwHkh5y5A4AwuSYaRmGU8n4Odfcxo603vQs9kMBpecpdv6XhfY
70FmaUOg4z1/A6erqXnXPK5MgyhGuM7jJjCx1qjFMqJA7G9jDpfCevqupcMPGdD/u2VyOKxR+FIw
RKwL4shGwXxtyWG3WmE6uyLMKyDzC/Ps0SJgoe8Ho/1zMEZPb/mM+zCBdynIhE9XZGrei/iS6UQF
i/U90qmjh6pnQji6taF0Sg28/m41afnLokMB5YwFJfVt7v13VHoSm8VXDmUcQ4TyQj7dPh2ELYwY
uh+DLz9u76cmjBHtMgWTGWHVW0/lWrN4ofPRvRqA2YchXepH96yvoHHgmwYEU6KVLXsMTOI1uDrE
uWxFjRpBstIosXpVns71u1mDuGRc9B7a9bxM0HL+oZjRAI5+hpfuumX1klizqAFkev5PG+l99eU5
F41h7mEBLDiq3q7MxijDGHSPDj24NBgdtfkntZTSroFe9iSNZzxUF5PUJ787oGy6NkZuSKSqa1pz
6SWcLU4aqCRfN56axlynkLqk44WkWJACGMlwJCTkmLTSj53oMAi3FHbv0g37bKN0XXxtURl7wYPw
3okvUiTjrqrNrjJdvFu0otZm/UlHSK8VltqDH+Dp0VA/JDlObp4D7+uRJm2WvJAC6Zyziw1zJ/Mk
0nHTFb6A7MREHL4q3O9eHaZofMc46iBXKN4RCqHIf3eUxXMEVRuWWNwNsnYIeE7waeE1DOzNguai
xKTkemQ7ZUqqGWLdmNDWpTXdBV+zyQf30MEPcmywbNUJJV2GsfvavtHBsy6xu0KX+AlmaYFX/e9R
J+V9AlwBzde+IA391wpt6I5yvzgKobiIG6fUPFPnFxL7A1g5GxsLu2BOfzPwV0T5ILUtF96oTHDk
REoJwLtveU6CGKja5UUoOkse/hYgR+Rg8dlRGMGXRhp/6tNLrg1CAzzIS7J3+/tzEshZOh8MW0zq
YtXXZlgWyoYlqiWySaq/f32gf7V+5Ucj952oyibKMG93jCTC9f2roG9LHVnPX/UEl+B2lOO7+rX9
iVssOQ4zWXCMD4KFILBnshL6M+QjNCWOS3XZ75onnDcUNqnOi5Ue+8LuT8IKbJPz6IKvb4ErouWu
lI7U9H8tn0P1Kis1FG4Chn+IOtNh5SyRzEhn4evtD/mCYG+ODleDDXHuRQx1HglhM+EKMBcM4F0g
cY/sJ6zcga7ChHu1YjS7m/ldNBs9jz5HV9BQmp/CutxK+tIGk7llaAsNR9E2U+LdDoT1tqFDAKyv
73wuK8Efv3vED3E/AMucXPVdI2xTkvOIRa7gXw3KZQanIwTfAUvB8Oc2onF/ZdRH1Q+WGs3FKlf0
hwGnbDtN9YNqRxgOMyiXxkB9HB+yV3+FX49sKA1jhSEU7SXDeh/jTWd6I7SsBqes4vzftr0q1KsW
2oJFKMzvgwKlTrxSdZIj+wCGBf4WDRPb7gZ3Tr2t+m7zm/tLt8VOhX5FfVwHC0gCReH9bPdLPHRO
S1fLbcEMat+A3sjiYF2iVxwuz49AxQVjO3RWZdt5H2NrEPmZJ5JQ+iNN8AMnPSsi6aAILHXOwyuK
NaAk4LJzZVF7FyRZgiBtZPwEi3VwpziV0PhbtrCQbrnn3cuKfYYGKG2KXqFP/2wkcHwRs4tikqVa
mqy28wBlZoQ150lo6p54UZlZyR/Bx6w0QUK5vZUulZsh1/cjfW4QH+aijIHm+O//1fgI4i1nPPeQ
l04x/abyd45MNNWuJ3lPxHciTU/DBE9ci4JGwRPIgpDlztcP55aLOVcSgfBv5kERaYzv0YJDkWf+
tvW4yi+V1rGd2a8zK9cZuCtRLeq1pvktxuEI1gJRWaAvDm+BNWedZsKs1vPTC9fqBcfJ2f+Mdu72
rg4Q2XDyj0JM/RUllXKJrVlPmJJAabIbXZpmx1XjttzLDClOqyzVdCFXoNTRvPTWkRvt5aHUExB+
LV5qLymWQhkTa8zpA/OTYQpkGQPOdSJEImaskd6KjnngVx+QzuwpxgrCvh70g1Aw172plDM0X5v9
lTSu8TiuxEmTcD1vrIIaPg1h7RXvxSlcwNPJBQhndPFYWRJ3y7kFfa2m0O4Uhtxvlbh7Pev35ZnP
VzxWmuro3Tok/10g0S+cPgI0EV3HIfZm12Bkvi/DhVWSsgL1CJ75uEkzuScVifQHloI7rZa6kF0K
DCT1ftbwLYQULwDUuj1ME7E5wbINFjnA7/tMWxjFre8RCGI5xRiCNN9vWVcxyUXhBh/0jZE5bPmu
bphnXyL5ZiFc59aFnHi7sZDQiVUqM9WVF1FtIQ3SbLEZM8eBM3RCw7H5IrBMfk0DBqduHhAOm8Wn
0W/HuymltKJ1mdszJ6I2OpzLUBJQkAw4MmjajFphU+/oywjiHaKWDgvI9bRkwWbPI7x7LPLxEZyB
KAM9IsYwFYRLRxbbVVfZtfBOnodmb6IMc2DLLFqEEA9KuRCaj9Kau95aF8kanuY1SVKGS6rdVYwh
VxKPymVznvlSEv4//eNyolJBm9xLPjA05vG2gM6BnOzwkrRsdM4/XTUBBi9hXLTv1Dzp/MQGq7pO
g9tGFUL+bjgX11SGW8jqIhgBnlCticvqk8SwapVLy9gHFCOHmPq0Y1SUaeO6DYbwc94UbRj+44hr
6QDZwPKAISD9YT/qTxRBZApLPOV9obmrS+19c38HsfKg9LXu7YsPsWEyBO75J6YGfJ1/Y6KeUyqt
BKBhASyC5DbdzeXrYkKpt5JedTRnnjRmesoTFE57/a5/GORgTrUb/F29b/f2W4tWQJeCvOG8S4+n
/HI6zAUMEAH6H7LybL9s3fGsxWeEnRPqHtJgQ2Nn0hoUFXfa8TMjHOVa55Y11DHfezSpTdrzPAL7
ja9RwBmnKNlMcWeHKGuxJjFg/5HD0ypIAFwPcvRAPc0G9b6Adw68G1BO3f1KcWnidpT07vNx3Cka
hUk5APBvv2EZRJljbCVJ2BThfTGAjnV1PXdlcWPYuRg4YpiykHjWiePOEuDgxXDXF97QQoFolnvT
3aENIgTQsj3Nu7fiHW880SFIog7xgFLxPh5T15kpOvFfwW1ciB5zNctcAXcg/BRePLiBDRJxAroy
RseVW3f8yDCsHxHw1P7yRYcsBm4U7cRjfjvuwfAbToXACk2/c2v724xxraCAqsxX4YP3xSGrHtVd
4l/a6UE0zG8BY68qUCYSJZo6bhC2qujWouAa+NpPwu6n9DgO3BOK+ztIFd855y/WY09xiotejpCV
OOjN9rHceixAaWN+PRKcI6U8vL0kI1iDQVTVmXf1zCnbidgVoDceXiMeWi/8QVX38B4vB23MrOUa
AAK0sMu2J9e0LbCJxi/k5/tiPtg47UaDBS+3ml7q6Ueki+o97xo3YSWxnMJkmFoxMq5tQgjeeeSv
y5yzcObsovhY8VVlHd5P1vYREOU9Bba+gELi307FWlOqLxJMCpuH9eivvm9eofCYXgWctB/lF/Af
qs3O9DU+YHMnOe7XWPzolT5a2CCgBF/jtKU6b5dvidKk8thBk0pNcS/RSlzSe9ec5RB1gzUzt+dd
kdmhOmuoYpad2bF4w7/f6gRdY8KcmKYHq9VorXiYXQOFCJyzhNjwjmJvOky3wZbc1IlUrEJPGTcc
HrzHZCqA/1nctuNvzy9DqkyHXvPf3nW327PZ1aFmCoA8Sq/MlhfM/OVVjlWqGzFj1wNSZebz+2wk
II8LRAHYt9wkfx9HLRqzBKLgvEyyJKTYL3YUMhFodkea+O6Drl7nYThKfvOZOjkxjtbJPEDPb/+P
g6AHHWBwZQAmM8IsIC3CbZ+g8snbB1mrC0POM/R3Zvm33J4uXaxoX0TCWqzgjpYS4u01WGAncvEp
7z/axWKjjx3WyXf1xoE/tBbvx4qsrRjJlzxuz33EWJTndVs2pAD8WqDsU/E8dk0LS3GipnEkMqI2
vqWIkqwC9/LdyfzJns/Axs8DrEOYE/CRTiG/j3q5Moq1fg9GZ4IFY3NPZ1hto0ehh9rM7d0mr/Zd
9e+HM+x3EeA1os0IatTFqSUvKB2tfFbIuRFzgEPYG02GpiQ91X6gLnLBuUhnBX0XVjbDT728KVPG
k3qkjn3NgK7XXIGe5AggMKKXCdha0WvrIzabw43pWonDjp6OPc6iVbleli9FlsYuk40l5x9Y1jaV
5ckMpAtFS0mr98Mw1WGfxkKt7ncwFiBhDoDCKvLf7xclS/oK/7vzIB3uSw958Qcz11EOhiTjYesB
TtswkWGXggf3YVBNV9uorS8Xyz2+N2r6//l5euVaGCKrGzxS+WJjAi9qHIG5W6SVWYadEs364E0M
3GjqiaPMWP3JgwQZvAdvS8/wPvTAq7BvVcCmO6Fxj3x5k6XZ5xpGr5dZ6JdUubYzBx93K7iw2HVq
op79MAW2pkJK3AYfZo+hdHRW34aUwGsxQOAg5OYMnomG9f2IJe8tQ4pAV1nfojVaZOHENeI8b9oe
HxxL+s5v7N4ve0VBmA7m9ecs6LVBDfgpBeBuQlcMreMNBRqDg2LWOARVRPCuVFQbuVu9DD0070wE
3b4RM+FfJSD96MuOSIvLvmX/A9oQy/xSfcCcAtBmx1qUK00v1oS6LzYiZs2SBf/NW55RF0X5lPAC
Sjg/aAMrSWrIU4y43Vv5ikNu1nDLhhnEPBoBCa5hmR8lUlVXyeapuZcL1Uxuj4NxwdYiGyb6LDl/
5GakmYOMeYFaulLMzBzIBg6OpfBs+8KHYJoqafGsAgBCG4quOHkGroZ1/MwFv6uIbxiIT6RS7cwP
JQkUOpO9bmi/LdmqQaBjzbKawv7MSNm6Ik7rY5W8PlAFok0HhnK5OQnwaLzjv+tEpWKKJcPsUpiV
/7jXPOXU6pOToF+oZH16T2pTogfb2DRU1/6qwjT9siuqHP1cjum5myeSARzamHuKRPh413OWRf8+
LZ5R/BbnXjjH0nwGlNc7EhepYq+bb48Gsvas4dCpgjpN4dSvgy/vrkDgtbcL3ezDQI6CU2ddYxYc
jWNcRhDMVJbsFK1/TZTxZ2vlUrhzfeCrKOLpXnRMtfAjiNdgUhB2lwNOijWdhmBR6nJdjPO7VKux
TXjE5lzzsZU2Q+k24qgQRzFhYOJDMwaqfXxAM95P6yNNMPmi6BNWRjFShK8IlyGcT6iruKELtoXd
uirdi5r4g+Manizj8oUT/xnClXE1gzj7eB5sSWBQ304GaFFQI42zP8u3mbjxoCrIesaumHauVi48
fwtOZVYVhXRtgZxhEbqhtSxTvkAj7x++GntmNbTidfblomEmFhI4UNrK9lLmiBXVjLgRt/fhIbDB
BjFW6/xBrXs0tmKT644JDPPDt2pWSjyLsQF2jJ9h2jYPLslLBLhd3hOjlawZMMnve8jCoCBh6bMW
V9DWIUClpyzwV3PkNC+0nnYRayQUZLe8uxfjEjFahLcui0rJdBv4YfrTP04hpi5OSIpIP+5QMsag
GcEZkEsS9IwWakdyhyMHJ+rUCF/b/Qn5y2rulyLClPLtkLYEgggAOZJKzsgnN11pqEgw7/haD2q3
fM4wFVMhUP5YG88F5M5WWSNDnP60T/PDXOhfuw+FU6wpwa3PCcY7O/u3VhGdLgwVLNGf4ZqacYva
v/SPSQXlyY/Ca1AgfbDHZsYQcAsfV6/EJq1wzROmDaTQcTYumy1hk90o2xv5jdRJ6e7eOd6SS+6/
YulR/jcbpFwBKjLmtgS/fq5QZ9k15MWiF6DgQsnowN4yb9xp8NX0ZEodHBHCbQFxfYWWId6F2iUG
lcd+gz0cK3itE0rclSp+qukuDPVAtKFjsPtpC8q/BGY7owKqxBNbqAZ1Q2sg/gSAON/e/kOH7YXM
lZSA1GKTjFIRfedcBUDKvf02/ZF1sTpcke6DtGGqn/hRjZe994I22WQGWqfgXcyqx/PdFPTVR+ea
RoQqVoUPb2mkC45qw9LiMhFkcFXs8IFlAwuotbjjJG6NlHQibTL64B/n45u/TEJ524Fzr1X/ZoQ7
K/wb6WVr+WzA/Gm7NqS6kUc9JPvNHYH+pmPiw5ell4xwo15rWvr6X3dUqtIzmzekCtp+u843VbwT
Gk1B/1/l/KVkuBG4iVlCyBgfdES8fyqWUNEY9IYx0HG3OP7AWgQ0ct2y0lT+wj8wJ5vQyf8OHdfx
ur2CA7ZTs7YawekUrEyJUvc9ShliiCTbXzJeUeZppuy44m3HsGIGUCpJbdzf2Qu11rniXwP4OgDl
4J2FJ0AY29pQ9z8MOEJ30Z6/X59Wx0FuTrQcsBGzb9ePixSrovJ4/+RTtJTHcOQvt1eKk5jCkdIm
1PsakwE/fTjX5JK4emyXvx2tcAQ+PNRsq9GHog1Px+flFCkI5EeHGJAsfs1p8A7umjISis4zbRpU
A3P/x86JPBM9l1cgiy5Zu46Kmecf6hJVgBBSHLfcLWiCbwokd9lsiNEXmbpWA5LlOz6cUr5mr9/G
BqAmaxViFt8lp8597sxL2sXrmFjzk4Dg4CAyETV96JoNjmP713FpDedX8PVBCDtTPUXZQ+jxabuo
a/96MMXKVvIiXFWF5XWWtxdqO2qyn+Zk1kkC6Vc8nCLZguu2KhXU9hSykK0nKelHQsUsuygztoni
yMWVP8Gc+u7E+o8Tayr4drjs1MsS/nkOTFOQYuiaUEqpkw0Y6f2PS7yxGPqGnU9LGnJhyoK4+FEV
pVeRK+BUl06mHKTTveNOBX9bZJzZe8+vhTcleiqEufD12dH9qh4JxpecnItoWUd46goPXE0ionsl
UhbUaa7Efwycy0b/EdPdk7kHAPzXQLetmvH9QnmzwPfJapm9npKoIT5oAxrNJVh0E+DBaW3kVgcN
UVU5q4rKWi7IlpOHDc9NNX+WLT11QXIX7KYsx8JBYyYDibD1mbKCPXQ/KqUeRuInbMoUSbt7shTP
UEU/waZBFRca1kVft6nEqwhgIwC4QXyxoPBQk+NVcarkpY1rmBgMK0DDKkY9lDiV3YrWf0MgfqqB
CvUy7TENJX9Ead7Pk7g75yS4SOjFCK+wNlNSNM2GWBRtSbrK/IxQCpV1ujilFUYZ2W/UP+nBOZ3n
w4Pm4nSsEX8R/4n3ZDVHojZXnoa8ETjZNH7BELBxo5+d38PSF2puS/zV8wg4nhR4exdyM/n8uyzb
zqMa3Y9uOShoS7QE/AZZuL6/AtjFO41tHtg6lGp9PePH9TEek0wFx+WHNDJZO+DEPDEWdRd3e4vE
3reMaJeTBPQd4U04QIUV63KD8sPGCwHyc0yhFiM6MrjD+Zsc1HgZZDpn+wkJPnmbom/vom2yOBpv
5FWQFNX8QuJ6QvZdnw4q0ACaSmdju3B4wwit3Bzmbb9yXH3cynkpc75uM7RriPhMv7iqfhIBYC92
yz1rZrOZIA1LEQeJDfFrh0KspHvZ47V8ZtwVqoNJVqx2OO7FfZ+CKUi1nQtQiCg3znXo0harJEfK
8UvW1won6dkdCEwJBdmcQEAgh6cbjeYvIWb3352ZyNcQ682mfiQ0jXv8HvEPv9hASYgDLCGiA4A9
jOt7bWGUXzI3ac8WC63tuWTQi/vpL0DaimMvqiuVkNCtWSueAmBWjk1Nbs2P9bedv64kXQbMQRZm
IOvuhi+xIgAIYDKrBdQ62n4Q6qi5eK5qWjAYGZ7tTMKZYclGPjGSa1j6h0ffoaDJwQy8B2Z0yyC/
hZpvbIRW5edhJL7ox9zG+lA1W1BqyTq4ckVokX1Ny/h+Y+iWC5uNQTQmwO+OxgvSJ7vFGGBzs0SM
UPlZVbRrQ255TJNgtQRdNAFxyO2bFfMq0X2N0/qMYDs/pHPeRM3K9SSRXLstAu6hayDDZVmu1+cr
TnTj9ANz9NGMWIzf4sMfpDT6E/ornmGY7YR1CA2hQSfX+hmr3T5mgbVagLhaNAnWKp8hfMORY6i5
wIudoG+GZcTblH8w8zUFxa1DDuELZHtrdXmMFzmkm2AxowwOJ1f7ZPes4rpW2Ui+Qrs/WP+tVmli
4KpL0FIDd9v2XRONO+cUCMBqlOAcpIlv0IMmIa9SK7KA2NRGtpKPWOsmmbyMQi2NPyNSxa6G63vo
55y53R9LoQm+2HAx6Y+QpsRHAZZBDQ/FSIPxEt8nqhtPppjnqKg9WmhrVG+MZUhY16xoZWjsu9dw
0aRGRRFacodQoWorAMXOnDuiqRZpGKl6su5WXMduRDvbDm3nWjJFpQ6ouIsk5IZlddDVIICN1Zkr
S6Z63GyfPhNYTNqfPmksQObyKqrgG1Prv31DKP88h480GIbTMXoEw0O12DTX5rQe2FvNyPjyhU71
W+v0MNAme4RobxRdTjcD27h+yYJifZ2+jEwPlqMGmDYJ8GFu/z703wuOzLw+/tr++LKsIOzqasgn
zAFE/uLEovb4kTmXYsAXNnB+GNoRrzYHnttWz/T/gc3VrliUCPxi54k+O5OemYQfufpUN6q1m789
PQ2xFTN63v1+iZiwpcuVzKKOjQQIa0YPhXcYJ6wcDyuh3o6LB4iUIq4Ornmkg5lIsr85yKvUmJ2B
ODQkRCrsPAVuIH0Sdb0Qt0p26eWzlyEAgQ0EdaHUzxJLPYV14jhBasvbdxsmQwOoxHsW1QVDSYzH
7anrx1Px4eCPokIXcBbgzk4zF3X+edPgJXXL9Fff4khfHrPtuWtDa5fMyGY8fnI3H6HIHV0r+rHQ
mBdZsj2PMKf/n3Rb933PAUJOja3ZIQJZ4gnX5XF0xzDZ/8C1r+jz+5SMGXoOSwui71VSGCc2cDB0
mO62bc5nO+dzRGbuHgC4jYAhq51/nS0QZHBfM8WoQPP2znPrK34anEn/ZIisxIrezRwhi3xlYkRU
tSrSWqbzxf3sO2iaP6PWExmJSFdkAD1BswcqRzk6C5sw86cq+h5VgufnlR9ZCzieSrEaJFsDmEe3
1PR6biLMrJaiHyRUXh+6Mk186zdJOQY6ZLjbH98MfCMQx2oec9o1VWKaaAyx399nPl/emt0HYXFU
/MieMMy/pfK5C9s5wrZFzJOtiX7iN4a8YSNcnl64G2JFg0LrZK3oVEkUovfMSbzVQ7OFQqHvpgLF
J+0tUfVtGG8DTmFbHMey40vegMNq1DBVeLqi4S06/7+WG0aOEZqFRaU61Kc1YC6zXjGgsovmdwe/
l/LkrcN83ZOPmrTYEIyyj7eIyTykhJhdclxKgnWlkr25GsN60HOoZZvaoGQf4puFWw43YG+X0upI
M5sI59cIZV/FE/2HQ3LJUyzSi0iXfRCzPxHxxETIH4GyNzHRH9E7i4X8EnCewAcZa4Sf8BZslTXV
Z/577K1nB/zyMFRvj8pjfpY6LoQEirfzReDhODV3mgM5SWBtORVO7Y8zZmtMYi/g0bQnPVVDneLy
ELzZXzTrqs5/NSPfdeRKMfUca6H9GxmbgjPOj7xUzvbTjeyfVloFDlFBBLFXaoDDR7EWoOj9QZ9H
NJEX6Z+VZUAJbs3CAwYH1ErNM9hCSUavT6bKgg+V74rQ/VnmHT+JtK74YrCuatZX7s0wg/o0zznE
3w9XLtLwizpUmncxNjzHpS1FVcovLPH+16kFq6BWhDfJJHtpmPK77DwWt5HnntgZ815JplXsSja4
xBeqlRq1HBC0H9HM7CNZbBwF8b6mffROOTxlRqRLLqM7xMeIt0Nbil24HjgEn3T+Cy+DMr3qts6b
n6xsjxXxjFPPqvR+3ZaiYpn6zXOY7vu0UGFP3dWlYZ8JvTRw/3ue+RqUnbx7ONxIq2GttZLj0ACU
wTJBy/89qy26gATxL5GpKu6M4xwkKpb+ozYtYCMwWFk5fjPWTtctm5t13AAhrV/H3R4wY7tHHTWn
C2/TUND5P54FC2ufHwAfRrkktlulzTAlgzzFNmgU7g27oByNoHF2ZahoksFMtX34WNdLzBrKi+Wj
FRMjUR/JE9IYvtQ/p9ZkyRY1TaT8dLy0o7Yer5TUBqhNboA62IxJYc+jKbv+qEKuH59gEkrTVmwW
VbPK17uAa3f6UrErXbI7cDnNkTzfS0mPW4sYQeDd54bUNXaiyy4C7kp49Utu2CiI1Qxdp9gv4nex
RcprsmeIjehVYsldRh7mK+QXPELXVsIPeVcSmHLuVaUlnDPeqsDaWKBVKOI1114OdL2lx8Gq9KqW
lZ8kAx+XT4kPOJ+aXPuPfPGJxcnuwN/ZxzZXM7t3kALY42PICRRnASuXNUG5NK60L5/NprBDM9SZ
iznzLKH7WVh6p45zVnmUJvl8ayfhHlugsbGTsD88IaU3G9z4nOSV16nWegRQcWDqWxnaGKK6fpKG
252njXHfEsq17dHxg63YRQ3kFhuzN5o3qiOcBJmB1kMjeSyRLQ9Q/UBVM5fXviNKWMKsrC1uAIwL
cKtyhSVquFaNm5FyDRfkq+SY3cWz9RxdC2YEQAULurw7LFhqi9dhkeIluKjwM9ckVegJ+XWWDjiM
11SyH8RUacCnzo+tyjIMdybfdTiPlYLUYzw3qY35ull2evCxeHXfn6C9bXKuVpqspNQqXsDvWe24
7Geym1VTxuaVnUkdxNWIgWlWJBFQ4bIdbSHpmOzWoJ5lnzF+I0dV07laE+7cvPfV//YSqWsI5Dt7
1N4d/i1oqT6XkLWwwYHp6B5ZbLcb0MpxZZ04gp3vqd4LI9+0orkFzy7YlaC/QqJVlHq2G9cPQsOy
+TM38gQZubCBrJkmKeUtx3pefN2lKOnAjfepFEMIubVzuGyGaCdpG7mshaZ7X2/1zTURdDDAlnsb
fFUduWGzbFQONCzWUZ8fbEHdWA1Nfl5fWbZIQ5irPRM6EDoFFZmlKeL69MbR1aljOwR3VINY+fj8
hcCE9OXDb+R2N7V0PHAny1flUbp9cMzDTX2n0rEOdI9oLQ0hLt05FRpE//nFz/hX7IkEaaq8fa8C
29ehF2g02m19SsNoL8qPsOEAJaTtEQX59As/m7f9YJU8WtTMG1jpPyUD4pry9l+Q/BPrfUEIv2Yx
nICkrRIfuQAhBEir8IUW0PQalLBFHfLUQvsV7yVDduc8bpnVKBBbyEP7ucoLKzDEvNTZBHlWp/MN
tlpCxtu51V35iSjNrGNw+1aYG+3C3M37tyyuZYPZNKbeKY1/K1Nq200YK3ixRDomD3hntZMohDhS
saeOP3JzYTF0D8IHy31NfYo3jLuvevFRMzTVgH+f5rWH/aRdbl+5wmgtE7dZyN/UcaMUt6hyykNT
DO1J910PyztQ+XZqNIznia7EGspCrzs2qOxaZcaMPeMCcA2IV9NcZ4IV06W/LNHXIIAqbDgYajQR
yPIQCTkeJDpJSOwTbu5I3RWGP9LCnTGJ5gjHWfWYn70VKhoOqzXPvVsymls/Otw64ecOOPBKfVu9
zxqkVh4cBYlfNNS/h3kJxvcG8Xah7+oxQKZ1/eFd3its2PI78c6yylwjVqeGaWNk5L06LA8ZYc+f
LdpI0+AnxtoqmXdVxxSjAsmRErM/pvq0kIa6i8DuCq0Zs78GZiCzsTzhnhAnZGwxv/dMsNQB9TAm
F9dMy+uWFuUe4FcrjSLEYNpKkNj1zU9gk2VWATBzFsEw3gGlSaBoKwX8u+zc6cNxEbaztedMPwuW
yu5K4F0rJ+DbuCXzkdW6JfX80tcw6YEg1dRRe9z0tRISSRs31R8Ct8LRAXEDICRQlhOGSOxJl0mi
/UNrJQX0cWqZzY5Yj7UwFNvPmHVk3QMOeTW5rIrSHODV+IndR4Z796atmn5jPnwfzolbf3npc8cW
PhhSsmEnjQwpzxTIKmD2f+Hbv/kUcIqgPKEnFRG78KpziE9K7Dc2Jyx6dxC4zTBmHuHZDxxnnxgG
B6XNGtUO7uUu93G+kqOLDqaoOYFczAq3AbbLOx+yv8i9NPIWsHROVJDdhvjDrqFdAtqEew4mfnMV
k+m2fRJBemSEaK5+HExmka4IdQSohdI1XRnwoEl4QAuxjGUAu9SP8v3BiYDvxgbtSkNHfvtghHks
aOtQrhTRuIAjaEGfXIo67paF7/ExKsWosEwVXuymWjEr7BetAROM6aIaMMmgtdnqhvH7SGqWkxXu
qomOCNZoC8PIeTEERsMCJvcD7IsrCF1fIQViIwrFKlZ/tzz9CAnkyloGhDJNoJdCCg7vOWavE0yP
f0SdHoyIbmqFI27m+GDCZv244eTzcz82c1XF70LiFtSn3LDYsYu7DmpIliaFivUogioSHBlzx89W
IahMRhpS5fe8rSwNQY+Ifr820El1/iPrBHyoQ1u7DQgWQ1pgXjbOmAe1fpDLy2NziJXHYtywSafg
rpTuQmkHwGmKwyS0AJfEm6Q3RVo2Tavfc04328YP2q6bL6OMbCl2juuMpcf5pPQAKJBXI5fDkZyd
nIlg+Nzb7O499knbeLWu2UQqEVgtZ43Zrd9SxWV2pnkSPSImvgAzRKyrturEFwwYPtQNJF4gmEyw
xzHudToxeIlLMHvev8FPu1X4l2K9XBk43NT/2q66R5KAHZvfWjpSHqk3CVPIK5V+dBXd6Br2N1vM
Gpz7H4voVo+YvYWxOpLghyp/oTdPUssDy+KW/m0vqaaLLSEbX+8I8r2W0+F1XINq0H7TLy4Qoo/f
CDn2NPWq5VxwYLbHa5UoTQxN4/ra2dby6/Sv7mqnI/1RDKmmX7erCn7CfOyqWGd8WqSwBAYRuP53
m6OsILyKNjyacWNS1jnKOiISeEv0CQHDP4jGg9nnurmmglfzIDKdzmPM8nnTBs5M5djwNyrPEf5i
rW08oT+qJ1i/pB+s+bg4S9qw06vQEMrv7abrIoqT9hmCk9wYMfYA9WfLhqixY0R0z8Hxczvw/qj8
jKSfEJngOvHC6p+1+i70iT5q+LjfopGQsFyFI2cxorE280bK4YndlN6eqQm3joESKPWKnZLE6SQ8
CV4KpEAPN5PfZz2qTb4kVDiO3mle6cjZWPqcFGil1d+Al9jiZ1ITz2SVJRmiZfzvlBp4KU1i7yBF
1r36KZyicJIZkHVtUoKSPx/JlhMQB6mRYalqb/mOn5aCKv4clvZljCFMHsg/zfWc1qjsW2bWmaoq
pq9yAvhEeHscM184kTPrpYTzzRo8YtLntQwluRJ6INWb2rreamXJNkOEgo0FPWqOZt6vUqwOn7ix
+Fpkidta/H395YT/xL3O6Yof3OpTF8AOWbH98dHJxNrxDWByoHPM8nPfY1ryI/pzKc2QK5mLmPdQ
tCJNIDv2hVkE+MOWJ+j10QXKjlvJ2KnAz6fMsTkZq3oK90FMxWZmbhMO5kzaH74jH9GcChqyLEHF
sfV2x9ehgyJINfbw2aB0T1LWUBjv5iFDZqa3w5w8Zb52n8GEnujq0pbmRiO0C9GzWuRxM2KfSggu
DuiZfThFHWOKAVZCDic/NRwb9z93J0ZliQMZbqTGOEPUCQjJzRrrb7A/smWL5fsKy/AaG7KKAJde
hxM9j3XywN3OosmBEMNbMO53SJdV0hwrPq1tSvt2tTDbHtF+1LIHuzHWVu5yv1iynsq2o5Vj9z8y
rQWgkqQ22/Oy2s0o81hQ/C6abkvi+OT8yDejvcp3JXX8Gv4gY3lAybh/gl4HIoCQXmhyTT4wo6/j
pZZIvSRBDSv3aE7o8ycvMMK+HnxgJNiLwF7WTlK0hSTz59zA+05W/6Sqnx8AWyQJOWq8KDbzPvNp
o8MW35m4cTKStNJcDk+mmTvXhXPzIjdvtZQhNygJ03Z1r7ByoHgrUUR7sgD/m1un5KDM3zaxu4Xw
QTH3qfOFm7JeAJBCEaNqWZxJlzl6cRvpFivmew7KP4zhuP8JZtSUrym+grrTPFBsB/wEcx1YM+Hx
1jJmFZboyeE9EUkcTfPUsUHfAmV+d7+zleqW+V7bpHvbypaAq9m3QJoKyGlg08dho5Zh5yleq1Y6
JA313GKvy9ctUNofNBkbusaKoc2fhnA8gFK53GCF6fc60WCHtBC6oiuRvWJwzoH7FuDqghDptgMG
v+hlfvXZjdlO1Fno60Azimuyy/bcUjDQCzy/LrSBHw5kXsCV0tBXV5KPTuqJyWK8DFxsWxd8LW91
D7Ix2ZF52YNPP88H7ZsCxeoyo1HfGw9yL8B1UKlIMr5gCXyQ3Ev0UoXTqefIl0/jbQ752Qx9qTes
tKCcCg6c3ffYvp1iD740OlNyIcEuBENH678h6WctoiqgzIyICSM9JhYFxaJDs8yg50Ioc2bdOAp4
qaaloXfP65Hgo5ll06lyRQzHgpaM7WT7NQNXzFgVBoiZ4TemwEy55yAoKMDwxQXHENupXY8EQFFu
ueG8Fsu6DtmoeUivgwEvZH2J8i/uthYVB6qy2IWc8q128tSM4w86afbzQo2bx3W1jifiepixiFke
iIJ1n35422Cgoj3EbzdOr5QmTLfO1I/8clVFCW1gbWK3Z2Jq/yJx/Bygn+cFzrTQeNq2f9Wf6Xu/
mEkfwBityxpjBSkQtkKPM3onDq3MENRMfBak9rAeWDi5RFJX6y0Wv8J6MPTjty8Y/mC/4DgF3XfS
B0w9MbgJthRCN0FpzzLcyvku+wz0VCrflPJFJ1c7IqHJCB+FdZdPT+eSzeoJDE6NwQ6RIGIvJH6D
F3huBzhSHQ+TJUH1RFnSMUJ+kDb+YgfcJOkxOvtsjejs0v71NnSB8p09sfmw6B5gq5ur1b/4Xk8S
KLNUv3ZCLjM1oSmWIVNlImOODHUOVNVy8sugrLh8SG46ghZ9rK33Y3e752MFBIs9lpnFVaEXk9cX
ewGQ2WPV3dttYjDUkP8NMO26U1eyOjmk3K6EQjvwp9Gj/bluZQ5oGWk5+FDRD/peC0xEEnsF1wJJ
B+5w80xcCxwKuCQd/Go39kt0OaAbKZ+NKdvm9Wndhvag5JT0T2Bh/bUnF2YZDkC0wW8i4VpoO48J
uvtqGF0NpUg8uZE2cjQ7/MiaP75kUudj96ins7NwXJ1JXABmlrN1bG/Zmjj9IEIgYqM0dEXCTaVX
ksVtO5XzG1/Mg7lk32JY0Fi2LcuvFKYYBq4qcbChQ/Spdnv+MlyIHZHnikrP3l9OMW8UkaaRiV1z
sriu3SX38LN+nAHrXwHpenocfhwHBY0i3c6QsNnDB/xAWQaphJccuxkZ/1Yv2QviKR39yeU9Dghy
uaMePVQEVtWw3WWPUQc4ADiBr+hOl0pSSZDROlR2KkidtEMORjy0edxz8mIAl+zakgKgaJPbYE+V
+TMWjWd/dxG6/Ry4mv150Vc2LVRPBG8Nq56w697GXaLHBcEXa+JDMJKnbaFv5WEE6owmMRJoNPPS
ysNctGVkhpbg/kChq7qJ144ubJhb19rqamsmxHJrOYurFrkjLO7XcnuRfwIqFLNQxIbbaUr1/Joo
qrjrUIQC/BNgAOZLMKPCt4vtniz/XmSTZxgDRqacK3RnBDy26F4oZ2WGaTxmWKUU8ebI0s/brH23
SMHQJ1EfDyS01Q5VgSGtPaHoUGCBhE6mIrPhuLC+OCWvgAk8SSUTH46lAy9RxUrKS/u4q453UtP1
ij0FgsiiGDQVHKLaHV9euXPLD1zihqqFyVb9VS8qORNXgUeU84vfT11VrylvYp6sPvfHOjpnoQRo
GA9BfbPggw6IVesPPEkV0e/QY8+kREVtSgoAEc3u11/79e607cRrUvoxvZGU/6MPauIbO4aKZ0cO
gQRIeVJ2t1KZJ702GXXEFFjWpOJfsxCShAJMC1qWeYLpWXLQ6KhH7ZJ4TtMnSPya3NtJBR3xgZAI
QYEt5nymQJRWH3h3EM7li8rQm01sbBIF7lOgivfVxXXBZnzIpkyhwZ51P/i3GmahV08DDWxqbORu
m2neNUEIgRaFk5+PXJ6CrwremDR2zrdTdOmz3t96VCgTFROeVRoVu4DzfQcVRqwv56EPZl8a2F8U
HfWgyIZjHxARhNfHlKHD6KTA81ljbdDQQnhqdPttGgnTQrU76BbZOyidL/Z7TrL8ov3eaaBAcRKn
B6TYV1V6gENqryk1PUpDX9ntONBJXE40LP5PleGbCxCht64R+tIQVo0DX3YLhHAzT+qkUAmuLBUm
/OTIrrbza6RzuucktcHs2OhdCKFjnbTVi6RaGSTx1JUkCXPoBqcbDRtENptoJ0YA69x6O1qQZhoL
B277nHiGdX7B2ii8mDANTM2zJP7X4otYJ1J0qzy9gu8ZGYrSXy0OG5jcNMhqyMqnnheerQoxlfma
ttTqeJ6OsMIEvc6GrxWuXGCg/mcIgtqdVv2d+H9mHEn6s9U9hdrHEw6kzMbSSf/PBJjmm2sY54Px
Dw2G7jo9l89hgoyLGeylMFdal2AoMtbf7Ha3HKkbQm9/gj3cj2ITcDgtUp6s12RJp2l/JNn/8m4w
5yQA/Jnzwz9gY/kzQBMQyv0lSWEEkMTPJcrBYpd3dufcewmI7DRieJfdAuIJDLBw5bbX+38oQd4R
PRayc6lW9TQg6rZQKY8rvzOzlI0/8VuOgUmfVpB1MMBhZJgTDBOYTYq6+3xTpoVXRSG6jk+70gPq
pad8r7ABWdgP4ZfhjRufYDOWmVDnV09yH8Fs2C3+HiIGze8RCsLjnpTSofGORtwu68fItDFc0DuE
T7TwJR+db9a3rBoENzi5poArihtS5q49aa0ZTZdvAdq8OqQLwdZyw8h2eq9NjkZMDzMbc4TLtNHv
6FQ9Rzhq2KDHsIS6k4qW9YT6nayITbELg83qPfN/N64bgG4xAImtWbqxHhAf6QPr4XlGqmkX2JBf
pV3bP3SZz1qwbJ31g7LwDYZYrIGP8VLzOcFqgYFxhFR+wwNgthoUSIwddwc2WwZP52RAvY5SKB9c
BJAGjjR4dwrHiyUQlWKtpP3EfLDoXZfK4LEH4NNQyNw0cUQq1nIO3oJNkXHyEPpLc+fMqtJPy/IX
2ILf+Zv0gFadi4qM3PJqW/oGJ3yU0UTjboijaDsTor+Er23y0wUDR5hsDZDiAzuHat2lWuGZH44m
78khiWIKoJFvk1NOG475CQFt8qfaaB9r9zo5T+992TF2ktXmfurqKkvrTfHR4ITBICPK9NVNw2ph
k4df7SnHe9BKFOJZzH8egGYogvhjUQWszmbia8eHVCvHNuP3AiAOqidiwOk+TjgoHq7qCUD4Gkld
RruIp191yJfZ9bko+gk99+MsMlcT4aHxpuyLc0cCaURwMCCQy4G1w9D3td1Z6+K8sE4xyunkieOL
6R+xM2J9sEUw+HnrwnxCJcYWwTad7mK2n079aEn9bcTcse3mKfu8txdaIiuq+pljv7Z684R1SACc
05+XzFXxmpQ1mQhkROFGIDdogW85QutSRGqFvD1bzLOSHGdszkznRLwlZ8BPpdodQpZjeOt22tEB
3kOvKe62K1iltYeB+osnbnKypPboq66kUNYwdOcx6yvZYOKfFk8QmVnD94sXoPGrA5i0sWoY4EgV
2R0m3qaIezV2jaurN6uL9ctKV8wcuZHY1DzRET9KCFuaf4rtytsk87ql0P7XQJxZvv8KX886+2hV
xcsJW/S2TczXbD/MNdirfVkER6+W34wH1oa6Xf0RKAontPvlkf5hBoOBMLmAZD+7pJbmQuD9sn0s
yFyUSGwk6Cjzp0dwUFB6OEwGYk1Gahy3Crk+F40uAvTQodsS0n3ogOqgqMmw10drsGxpggGgi6BF
d5Ev5+yfMBTGBgyZICiUiqd8hdKjJD2I8jz13Ub7OpbKj3Dij8V+RR3enoOiqDdE7ee8KaxI/rj0
brdWzizuxtKmMFyuUKZDVo1RxBKtr+wgICSdh4tx/3o/Gt4cgFvqMhVuooEpexKEGxYy6eYYKiwK
Lyo//EgqE8rYsvr+5MGjkkub2c7DKS5lQPPYIMD7h2+qa9CciKxFmDrl/x9S1sGJI8dpljRofsnE
8TPjYCiB3+81hxjQJC606zkcOux5Z8+YFWJOI0J9iSDJuHfnQswQnQmL9NxtasAu0L5FdNHcrc/K
hjA2ay02MecnHfZZiGEXXzeFjf+CdoO/X5fjZoJWL0avGBZ+tV49qDYLGL09+QSikD3uf7iPz7EY
Lpvwt5GU/uFGJYbVioYSlIbimWGTCcpzlmHJf6uIpcyRPAOJXXf7rcgEUUs/64AusPoNwEVA+AK8
HeYRoKc2sAqQOpugHrYepoNx2g63rnnY7IrkN6oLIuYTupUdruifuoGw/nriFzVrNcHDG8OOjkpK
vKfZbfABRtEEkEoBXBbJ1akv9NZa8PRx5rA97EyE84YWSYWo80NNDuYMdGIcWYN2UL7wCT+4jCx3
kV4jh280LhC6ziIfX7hb/3Mf7r/6p2RH6O70WJohxq/oeFAzWJzdDm7aVnPbfSJRVq0cTOpLTchi
0VplLq6C/m+rqLrri2ufYLz6Vcn+6H5Qy/dnhLZiIJC0NKbUZfFMTVwajVQLb4FTSqR4cvG7zHdj
/MN2irfxGXhzD4U/9VSBsOEJAJgsssYzgKaJUBIE6hufRtgYZF4WOIK+x2E4V+JmYJAL5hLtVZjU
afqbjOXtVxwkCQKMloL4BKVzwIiHEXmJqLseUvlCp8b4NGDA4hbY9diZfPokuB2xGtkR2WdcFtSk
1+e1LXERnL1Bjw39dGtpagPWMG8XJd3y155Hts8Fi2kbNtXyl0E7GhbnkvdQUbL7g0nNUjzz88vX
KT4kmY0cUJMZiwD2AR5HJFPkhbHKHjXNkXvIo86rhvFdYelLIYOxic54I767cTy4WLAUxdU1GNZA
ZUZRbXkYXm7uU6ud6nX9WjNSU8G3BMJR0rqcmClxNgH7f710FNQj7dM0fEhh+5YS76op2F/XVCC/
YOD4pXBJ0A2HlzdguRkq22nUtOuO4u7SBItCOIFym9Bm3w9zlSJ8vcUh8zbuvDsz/K3JCjB6tr4m
q+YInSvZOztcL2aQF79QqnWjHT4i/YGvPS0aRXlKh1Vqg2IwX/7WCMbG//ZsXZsPoVi5qRWGYsJ9
ngcqGXEvpQ0QQkZ4IIH2NGZDIY0/AoCNFF9erRbJXkKcnqp7PUOktPY2iGN3Je7AknVIDURiNkUi
ronAuOcKT5eNuq1c1Yjpy5mOLqSfjx5wOMgUiBorl0UA2Fbklzv19M9vqZ+SgF+6qq7GCsTHingc
Tp436XvMWq+bmgxRYB3RavzhN7kmA3pFSVgJcY4NhmwkJWn9Wwg7dF88Zu4xLy7poJ951AMvZ/Ao
eYKOEGCafDfFV/TJ7WzKtRz/U2qqpbksb6QHXtx7sYLx3MumpinAp0r3v9K/dbtb7MsrW/lXE5vB
vjWQVVG40xyVez5zqBYYPuy/9xcqPeNUhJX0VCXllJgDf/UpbMZKq4m8w/a9q1NlIz945gaogCQU
o8Mi5ZYA0hoSuU/sYAE1hNvGEbYY8yIapJJvbqVSzE3oqoYNIXKNKvKc6aIufCi0LW4ogq/bUV4y
UdvuUi3RKPcv2cknu3AMh80wviMSq14qcQuhLGkEKElx2evmZ3UKb8jJbmSbTTA6r7dJBXBNQDfD
SMRkFxsaX5HqKTjHfqeypAzcUkSfgGl/Ek2Lf+McOtCUbzXoGqmGWwRhQ/zvHj3pxEr1T+nEaVhO
mYxVdF1G763LUTdgEuOw8RahHgnXf9I/EG2+XJ8Cfk16kfPaS7gQq0ewAEa9CGqqbmiGiIKbzjR+
pxfoEv/A7KnEeFHEI0XlanL8agmepjYbsynG6eJj/s3VzWFwyDF1f/aefuEklKfKq64Ma2L32lN6
qV0oYysIszi0yeYsrZ0Biogwc/c7Ws1AQmK3hld6Po6AS2vf7tue6hw9CdqL0f/X8rmzd9t0OXPg
61UefWxvH/afOS8df8X1sidvK9hfsvsUhaaDMSrK7rCAVnu5jnd2xmdJzTtVHo/kHVFruAEbiRbC
nwl880Y16nK+WycTo12JYFDkNJAUE/dFLgB6IymyXxnv03HXtx0tVyKtVvIw++GOmTPX8vET/pHT
ec3DXqijRGbcIYoT0hDToc8PMnxSdsyN9fwqieofnsGArr3Ha4QEM4K85/2uAq2l4za8GWTdj4+0
iF//9xJyy3j7DkWC4zjUC1lzOYBPOYknps6mi84AiM+pl/IwfC2BvEfrKq4W5omK9yw05jXHBoCv
dCaXfRlok7sa+GKejHWltSjzFeXJIVZPbSvwH1sxD0LH3k8L3O9sAtj/rkAG61eX7mosl3a9RsN7
9YVUxLd1djeKTHPfRLs2HItBCKhbKQX+iDJybOM65NMSY6w/2o9YHyuZmNR9Ky72FzD7VW9m82fR
e3FsyZDZdeNK2yRYbj9k8NAqC+fKNKrOl3fKYd///ngkY0lTj19F/ASMF2DZSOqo23xuATKIdcGK
tO2pn9MjYySaQxY8bBTEfLSTXE45cYl2xthsDfcftAXT/86lLG7l/TdAZUUyx+0J+TFg35/Q1EPg
CXhHwDuChGqKwnyxnJsupxcsAhLqh2o9LjtXfMtRaKKmlfThFOi2w6tbNHNPu/8Bn8Zhs5WC5P5X
+I/cX690tpb+ec6xAE4L15Nu/2y9+RlONp8FpF5vme4yKh8pG3XfatshMwx3+qV7jxgNZn8OqkL2
jcNAqTCkmHL3h20eLRVaoTh3ovbc1/8tahILlxt0EX2trJ/EO+F9eQQLqCeM1va43BBo4695fSkV
x0FCoLVDyUKNZZSQfoj3POMm/GbFpVo1xAdma5Oc5EfeVcbkykcF2uwv0FNI0Eygsq23LLmhAIV6
DGLOlhPCVoCuYU24ds/3VG12PLTpuTZ5b5ZuYeQemFiQMNo5WfEQUbAJzAE9bRTyaeKWosJOFNoK
bcYveFU+LDvKVEC7qEuCyzv8RI76VTOXd5nzXviqcPCBLRambWnmVcB1RZdpj7PkR29s4JSs9PfQ
D1c3XUHZ3OilcAKzGIw1NQ0Vo6J7lBvw74EdI8NI5lmFsGKwlDfTQf6Ws7msqZbL4dGuuk7JTRZd
w9muyI3k2PAYBzu13Xz7aDf+n0vC0zCwwa4JKrITLvMfrd6DX5b1BmhCo7H94jh0GXbv4+Fj6zFq
f0OrlaSG+pjhdSQyckaOpJm3eRoXleD2P0YFpFBxJjOAetgWuY8SXq56qa98Z4QsnJOLW5P+zTRo
jUjbfgoAJGDdCOBQAKFkHfsOWhBkNkqx3Dc+v8RHZUOgokPkWyGFbqDt//rqUgDap9v65jdelwi9
QL2jyXg2PsMVFZ5sJGZ0ifHttWkZljFqWG0tE2zHQNAIxzrLpMpZfiHNZsDA98ePOgaI+BEh1Sru
zFISL1OEmbp6tjoPJlB2TjHmysmhNsh7H7JRtpIz8Q2Wo4Bq2SgrVHrimJwoBVQlq9aMpCCrzTIe
M2Rg0AyyzwO9gBKS6XxHRb/WGerFjLvrkkcRpqxXb9VhVhz40ggjfT76XBY4h5L5bqExBBIfkOJ0
cfvx/+ZUCyF/NExd4GYCIutnUua+bpND8cvsq24Y6ZmqznTGkorUewpSAyYyi3HT4+j7bS1SgcL7
xo9ibiQWKA5TjNCrA+uWMlt/xwOv96jt6+U4MI5jH48mklqeFajsGE8QAqVLCsID/YxXlBjGQ89M
wM2LylNQSCcV1nKbGylUq+koJbkfpKHEgp1uRJli65ojao/6s8lvRKFgFerpaLEdVjbfRQY+vKgK
nvnVO/BUujuUjXjX8YetVEU0fxP8zFVXWa4ADVeHul29vLNjx4vMXhFPrMWecGr+ztdf7W63ofK7
vhzcKnRVo1FoPj20LkPJ2Ln3KLU/0ubESmkimUyPD2Fd4hqGM1Eea+NyhBVhidd7mcTM5z6btKql
HYlQt9F8v6owqJ6gRE64/lcycc/yQmPnD2Vh1QI6aTWxRjSPDDeh2ylE99Rbybc0APouifWj1yk9
tpUbWGIthVHTvE+YseVJE8C1ODkTdFElcT++lHcRDZP9LobtpOyhj9c/11tFOFNr6Sdrf1pby/EW
Tbbfw7ms0lPhwXWHn/g0ZY0u4sObD9nfyot+0Xjk2ka9MjNEsoy83oE3/VHl/HyDrXuDRckL2s65
PGHhOj3AW21IL5bJtG5kzR/+fWivAdV73CZeh68YSHP18xPnqEgnJGJNjyxurz8fDlO5/W5KV4DW
JAYmwgkj4LI4sPjyjAWN/wrb+ZuSGvmHdvir1EnIIW0xvkRiw2/E92cJIC4c4wvnEhntIObATb6q
KkskQIpQQNEYhyF+oGKcIWibGpYRe3qczMpLohWdCar9V6Ke1ger29faTF1tq07emYTzUrmBohJa
gzlT3HGY3RqrgqDbYTVu1LkFrNPwZdpp4A03tDOBAiOTBBMso8FFiNRg2fuNCqQ3WZ17BluxQ6JI
3oVYXcs7UQy92itOL2ZgOifx3ktE6aIqeCuGCAigBwKZPFnyiLNs+jfvXoXCHO+os5W1NcAZdJAf
V9QQ6XrFgfYu1PTuKKBhWssMJuApQOpHfwlWj6TrJcL1fcQ0F4F05n4ew8ln4CS2MWvrbyjVnR5Q
fqN5WzGjr6vMRZAFwsYLxlxfeo+NTBW+aPcDPbSZIW3f3DwEj1vdkdH2u0+XcPBRYm8DxybuqW28
BATVE0RG439Xul/kBYzjvTOCLQVxaqsFYmkmJRRHM4TBZjNvTia5netTWDzkahzw/ByE1wvVm/UE
Xpo7aF3HuYBlOnluplg0WnJlVL9HS+Ul7OtXmzVADIYHBc1tm2PddblXyaC3p+dwu8S3x6HhNMDd
liUF6Yg3uiB40VBN8jpaymmJJMDHMA4hN84jQ3Yonvwxq8OUHicESeOcwwahKT2durFZN7HeZUrt
QyEu+dP2IvGWXmCWZaI71Wn4fZ0vffPhb4GOllQ0y3ip7q27ajhZy4V/74dD6kGF4fsGKJcSJr46
5m9dhofI4d+sRx9NROTsHxGC9dsshCLLZ5ZDRcC/dunsA+nqVo26s67R5CvRpwIHXNl+uZCc6yZd
kirQ2yHW4JM1FpTjQCo0+bguiCmYMtTUcsaJZ+yb8ie9i9GsvLm0yYi6F5eviyUkQgZ/j+/F1s/w
jfl3yuO6aIqJ1z93J44EIg0i4yA+99vjs8kFq7MYY9J/U+6V+nNmyEVwmO1eHcuXzLv7XsxAD22q
XKWQsiy8XWa05z2HGVz0X/j/NgXuLZ7h5DCV5qayaw3cqmcR+OP1kgXbRMkuav3e0Db8OSD9DblJ
ZF23BmmDM8HLcy6NrATSWoPAIT2ZFTMZ7O4O6uQdGKSlPkxI3tZUmsBfvk+1HsxCGnhFTw29I2kA
vPyzm93dBBy50IQ++Gpsfj3DWYFyhI9wSQHbvLCO1m6SuYnJhW7lZ7Au1zZ0lZ7YHjLxOhkYhNgP
1hnZspJhCqIfh7no78CLlkMnNdVA5FuDo0kPhVjG6MYlgDK+8sZbVRAzHAvBPDajCmuwbdeTvLv2
xfYU8mB1vtCw7A0887u0HKr99vBFreoH+ij3k4zGmalbSm2g+Kwg+nyolAU7cJ183Uyh0DrVMZL4
kgbgYjxea0tKOoGA0G7BMm2gjOG4gCL/BL4kEQzJ2PvA8mys1k2yBd0K15qvhqI35IhEj9ou3PUf
d3srKfhOOo9Al1rbMRFXJKJCaXv02vZbOUTqYtJKCQn2s638GXAdOcVGyHZx9298a+3Qd875Bao1
U/mHJNLqjO8vEbCjTuuEsKFehNxTNjnT5WNq4g0AF1kSoWerypGfg0pwd5R244M5XJwpMbZYe/Nl
TP1fu8LZdiEkkz14Wc9bhYIPutKI9GAT/vYxwCRO9xZYdeR3yot5u7Uk7i+ZbhGjKfCI+sk6oM/5
bEK8AjXwrpJpXaDiRjK9h4jSl09Nc0dvtRofnDUYW4FDkz+qOvX0DkyG0LnnzSUjLqtHcmkt0YLK
ctudpK8OyGD2uNtH4rzwHjj3eBRsKPeNVBlf+qN2G739Wxrc7eRRbOeMBlrXTkmPzRZGgJMGmVEK
HL6YgKVXBUc4MWAlGWeRqsIIclLi/tSpPjyd7ux8+YRfxzmhOhdeeqpaCcaBYs/O2LevDNFCx9l2
0lHQiM//ADHhyI+u+9a0L0xIb2171S3sbH+UCp7mFVAiyqucpoXkmhbf9awJjgLPAVMYcXkG4PbH
djdvu//7Yw4aFlDq7KAyE5B0A1bBAaCe5b7J4498aeZbUi56icpgSQxhMoEuI7OIR5Tl6vP0nQay
Glvw3wdfLqpJp1RJjPLeGieyBGWFwkndVY/Uo3bw+SbBH5aGXikkonhmezO4YIwe6IIZcI5jXz94
p9ghhCgxa5hVgX9tSku47qsUWN8GdHg5daGUdqAh8ytCyGX2Wl3nR5vVb2JQTU1H8+RXFlvOe4dM
0SngInWL5eaF/AcRmp1YGjwhgmnndN5/qe1/kVxzyZvJ+yuXHQTvNLnzLNeqqfReXSneYujlTGti
71lZYlBx1YyTScuQfklSp4bN5JOjSjtER+X7sMWG0EpYbhzKUi+IIOaKb+4iffI9K4ZhKu+qxQS3
8ilMNFndFz7Pv89oeAsG4nNnzQsSwIbWjBkOmHJjWCjww5HiNqNY+/sO+KN/dnVAxkmuU/AY0b/1
2t21M9oHO15FrFo9TDAo0Qxsj3cgdSQUcVpOAtp8jPyBQ630soNFvkEVwGOZysH5KWhHpHGbDhZ5
qWnaxyq/hxoQoZgAbWgtkXOlQb7RG0/E3tw7A4BDc9cANQ+uiGXs/vjGVEwMUAJ5QhXWpZsPxcrK
wLCgnkNbuUhkoHVHHlq/Aq48ycuTnUo5D2eEYHvGpo1wuBMNW3FxwUPiS4mB9LFQSSECnBuJbJC+
GdvGUd6Crvx3jiKAuhYpgoNVVTLUFPpmIhXq5y8l4b0am0wEvKV1X9JxD1JpO4RU+QOHVndqdWeQ
q4JTB4nvvBa8lr3kK0Suwfe5mC2ZwHtaBMmF+mm0gD0MG5vtnBknglCLOYgytvhJa6BnjBvxRR6r
GLpoCKAiEpPL+wEV9ccOOiM7/hyCwrQjr1g9QyXEDASUzTapMPe7EkUPBSIjp7NSEJKJuTHW1mCV
WptUZ/9ZooM72r1IINgTSEDmCu88TcgtisPzLmQhevi4lg/HFSSQ56fGMd+paBLKU09f9jiiIhYQ
aLfJo9FURrmnQJC+6QXbuB5JBszhRmSohoEDe7/H3UtCLE+FtFyP5MDVhjb188PG0Ben6Rc4eREv
a3IotC70gSzgFLbhK+w6gCJksKC0eqTZVI3GKHnoqqFlc2JuMNF4qhdBl+lSQdHR7jv5+a7xveA2
/u+aKQyx62zInohVuYOXOGKEq0Dv7bwsBBWNHG8unph2leDBdZtQKBwXqgpSALVP107+He/Yi7PT
W0JsxAgKlefWqfko821SJ6lN0tWjiCDHvT3UnQCQkhlgFf5/97pLUaxm4jSNDojevRpzwrHBwPFE
oPVSwlUMN58aE0sq6TucWMxvopcuqDarNmoJq6nbgqwel4Q/3ge6Gvtn47ua3nmpdaK0UQbstW4V
dYAtqopHZQ4yd9ZC1K83FIA0zZbghVPAIVnzZSxQf2qXs9cAtRddACbtsFMlbDP/auH+OVK9Tmq7
erwjo+Q0zMArv6wE7v//tF6ArbQszia/iVet2BhyMQSaGSQWRiolgl3xg923VKXiltzsWSddVQYC
LFf7tVFzf2WFgUkMMSi8dtXWixAFeAyK08INxf9eKMAjygfcE2ocy+ZAgLDZooS5lJPnsXDhiTNI
/YDUC0DK0tAB1AFBowQdMEzHVc0BddGG0hjo82Tx+APO1hleZBzIqA+vEukl9FZX4Eh5sxZtQJZQ
f+mM10X52DcPNTsKD2prXPCDJEhhRu/nMXUh2Ar2di/SSxYIuYL562IWhYO84ECHr9tpokj4bj4r
uydY2iURGeQGJ3C4Dk/We0iXP7UMcaX1E/aHTn+yrMs8v8qRTwsM2ZanwbUXmAS4qy3Aijuw+kl6
IJcomQ8cPKeYY7oWyluHbyWaKs6g4vfYW+PHR8VG5STHJ4Mlas3R0gVvV6KD9c/1xiIGFD+Za7gg
zaPFDEYw7e/xKfoJ2r4l//hzS7obQ2pNKlsLwAT+H38lgKbThPVXcE6bIez/IBXVGgOxbKzqnXv+
FWme8p7xiwgJs6qDwJaBNA+YYYOmj3hXhmj1TfqvQDqzBZdNNWHpYPdpXhydnml7JqgzHtXCgaeb
PuNg9ENwzLaUwKaQ8wOvQMaPQUt+G5/XeFYN4WlL2T7GNxj4AVKDZA0yoyP3glLt0hZEidftWI+F
YlHLcG9RxYhOBbCDDfF8u9QqNYjyb/l4U/vp+5hv7X4fUva9JtADSOr2UUTgB0RUh9pvI5uIydIT
I0j5lVhsK9Kxg07r3CI7AWcgmiCzBarPquTwUffi0JTYOhuYqOxEeGZSXBiH+XWlOCTnNhviLI42
q9lkWJxSNMjhLtP4D31i51rKG2cjq3mcVxIQ41xjE1+gvDGNFZ/D5C0Md4q85LHZ4u54sgeNjUhO
UcWcrzQNrRD3LaLXw0BWp+l7sPG0MHLAdWjOERpKLnCSY+hQkR7YgIDpqprRFJ1z/0MLYAg0umS1
naSVfcYBmMBLbPZqnkFrlDI0P0GzbJOCBh2Gmplp0l0V0OHGxvQLIbaKGsmjhtRQsrCG/9h4rN5D
9BkRNZaswQ+TeeeIjpv71UdnKXNGckjasC6Xh8STuooSdGlwpmYth/ZBGX5cu2auk353Bb0cB+29
eT1SUi+/KEKQr08RS7mWz6AODchXcS6izG5cLKdDXmrqJsYkVYn5sqVOHLB8qYAjsBBeilEyhf3d
f3y+tTiJMzaRPkUo4zgG6dgLPWtcSnQ3mLXnxYG15mXGgYpwWSbaWChk0uBcUq+R6ySAq+iMh9fF
ryB7+gpbxc9P09NOTk26MoD/I5Dv3lhnJsZLJvV9JxLANnneWt78mXDCSlXZ0IwEgpGOL3DBK5fc
9bqeg23ivneUDZDnoSIaKdfj69NlTnOzVF0niEfoLahNM8BwIwZ+qE8rXlrkdyrMS8XmnnQHzquN
PvLLNeYhBvd18GQz0a6al2l+KV8FoUUVtoIcyHx3LtXligTDKXLCgk8Gy2pi4bTqk/f4o4olAb1R
qeTGqw6i98TmOVG+S7JbB+TauiUCj78gN4JauTItZzXCv7lz7D4oNDsmTxruIGnqYfEGFz/parxS
nw//sCH1PFt8RrFXt39ncqqXYcSdm2FWharUR8+Xd8NPi+kwGxfcpgStfTgZupWvPn8YlCKn9Gap
zq8ZRapUNfTjfPnIMI1F0A+/yBviBLdcHr74d33F+JAx1+V+sD4/yGP1lznfpyHZyqYmapsiCOeW
YvWlo2aD/XZdOxMAwR96i0T3noPaicv0c8EW6EvYKiqhb+XfM0PZsazNPIPKs9awga8cNQIxTbd1
NieexcFOzE8LswS0QTm7ts30wQ5dD71kbdmD5aXTKh6xnIEPsVaud4zGyDosHrrrAj4pvjNADwq/
gDbH0DJ/lROw1Qv/b1KjNh1Ed48U/PcUT29ephIFz97RpdDxRK7ssDH6yrFUzHyeMni689th4/Go
4AwbGt7foKVAxRGucYy6aM6P+MI6CYxyvz3JLFYI1z+3twz8wUvRrZSw6tFXKq1qgPDQtNYMFH+Y
xDt138gbRpdMrjFg4KiDk6e0yxAsFrXZ6ty41TTmms/AydD/VbMffXRYY1gt1K1ZkMCVukz8pJ6e
WmvIl5Kv9Xm5yYwRgYo6h4R0Ri/nO9mWTTp0sorEZqnnV4qN9P3ZblpIuBAETxgtXIMhV6qb4C66
ceIj0HEja/byyDzRYZQecMbTirrRKPQX4GcjAavafMqtC5XB0FKhymTOho7rGn69X5k9Gav+XwbP
2BMzwnF1RAPkV0X039U5Bt7dbYkhd7rvCiLvA/3Ut/alILyAGVctzE0HYlSuG5BvxTKJq9xOjPgi
Qf7JE6GhPfYPcRuV4ZYyDv1VTnSbaHYWUFd4n9HpEjpudrW5HQULn+ePGGtEPbRUOb8plhBJi8Af
ThnFn/E4XfQI9ZXdOKRVIgd2YWuSoaSpOlVF6n1jC1D4x3KinHNuCDDDVtN9WcUQyA2eW4T5cmNf
vMb/EVnk1WC+ZZ6JWK+ubKLjLfWR7Kyml3BHwQHPGzxWjul+HaWydkXyrBKePoBoWUeNqxx4mRHk
txjWRK2qWBSiHNsqEtx1QW/xq9/wv8oSL/Of7lyI0BBxQXkLHWrESnsuRqOEuExJgAQe+d6dyMJm
x1WID0rau3F/e+d7+Gz5T/jDOO5krFPEM6HGdb1JSLIP7vYg+MqLkIuHv1LgO/Gx3OpmsEbB4QrZ
AAHiwGccehqKoZem8J1ThxSNdMFVuOD74aHE5Jee1FuN13bc4ZFuEMBLY6n6FpaMqBRMAmXP0Bho
chgrvQhKDxFrforlfXx19eFKoxMIxP/wHCUAyeGtpbDkizjcFmLRWSLK9GTf6EJjSgHIDQ8CMQlR
107gzXiWxK2jWltY7VSZn8BZVLieHnUc0FBlp2IqgxoNvATImflHNGzYxJs7jCKBSK0lc/MPig++
BaSqxsq4CBJSvy/ZNu50BHuMlvUgjPLnDijiUajgSNU9P9ctubSTCHXbE/iArbxZKQuDxe1GSK2S
8eRlT5MebzxwmSJsn3Y/uo2Cxh4jpaYqI0PqswW2LmRtWLQrQfACrRiv9byzbz0seNl+gsrCLn8G
XOQqYzPoG/CA5N8oA2/zB+gxF2cratVRhSvu+/pNFFSxoCpACa6h/WI1T2RVuO4Agor6oVf0qj+Y
ZxXuKmr3HjotSAqt3zaK8hLrP79vchbiJCg+xAtrsyPupcuRjsrVyQzcKw71sPXG1YdZsLgvU+Vb
1RV4KVFuWQBDghlGMi4hoLxYV+SUhNiUiJcxtJvfL+qJZKNCK9MpLSywJChHF28+n8ZYyTWg01Mb
51XLRAF85J7R8KMI9Ohzle2q8QGJ1RmHIAu+Y5Nw/Pq2LBM1Qo6Bas5sEyujsCZ0ohiTweQcR80K
Uy47NQafvNXE/+dgPwPP8+affOLiX/rAHBxTEA+y9/sP85giYzg9srXGqDrKXYFAc6HuoDCRq0d7
ZfNqw81Q/7bd9kcMH9Xc0MSiupC1/F3mhTYEpz9Z0H2d+hhFKrX1ZKKbvu1CHiH0wt2hEp5NfJ5N
DYYiSLIxcsiQ5ut2IbX76xOcrMxsbRjE5hbQwHdzjS/3QKeDBb7CSp3TRw8Un8EDj5/R56wWEJO2
DioxXBVa19ou0IDUs/Bou717PaaZdqpbHdVEqU3uf/wr31tcCEMem13O2cs3FcsRgTPTdh63ajPA
ag2O26XAMC0LIHndkKqmeabRMqsk9D7Jnn0fT4ndKdE+lY03XLWhnUzkH6HOxwDAh0ahl6rpEKBV
xiZqDUqQCelV3w8O3PfNnMhOnfmZEKlmxBJNKAnYOh5p3v/skdIjung7UEyl2CF8xGot6ht/QMCp
0m/0Th1koSnidOiFE3FgDeOdjYpuEgnT/R8BAVJRhfh4682hI/9BTizVLugovlMKpoaA0irCEFrQ
YRDJdH/e6eNLedIVBr3B1sVfYU695/jdN9BiVmJ//pek0E8FkKmtWF9Fq0YeAGPp09U5cWTknKW9
Io5ySVl3EeacvZqxvAc41TTA7rSSxHxJVu6QggSx1bWDJKfI9CinRq2rWi5TVPu5Se5C59PCDCV3
N5Ahh35eOlB3i0UxGEBIgOhTU3xNxYz+J7aVULEEVC16MRYDzFEzRmRAiaxDmhzmVK0FMB6T/QYX
7J7VzkIOjznSjGpT3hSsFknlt4EG3dG7ZBLoUDfLXWAyR0eXRkLhUy5RSbmKjxGbPHgI18Q47V8U
G4/vCdWM+RZSLRB3CGj2Y6+0tzlyGSp58MlOwGmCZrC/YO8xC0QsKQtsF9tNBq5gcymh/OTQIHm7
f+88dojv1eDxbS3wh5gcHptc0Giz3ZP7Am+0pxaJLCVTR8GTS4bqOgCkbIZSRp4umMpyJuuDpF+k
t9iK+spa1p4F78krOA8XbPSUFAhBQ7OJaKYo7gKdQA/HgZrzum6DG1UBIUMqjnfVvoy9VLgieH0D
0FexlyM/AaYqU6RaCrSkV2sMUSDr6iQyLhsy82tlGBGyJChyJk7YxoFqg7TEDDsHcPDO70tXmPY7
enjT4za5NMzFkNzGnEO1ihSBtVdeRZ3Z7gaXUnd75cY5GH+tKtu6B7vjlsXAC7Axd89t1kcsCjof
dNOZddzqRKyiqPht64yBvbnTZ9lJwbroYGejj/U9m8D3KytmesWYQL1GISq1GH6qJ5zA44AtkS/P
rZyOrcVHgspXlMLycjvFEmjtNc4KEieTxmoNxbcVVsngU0a1roPeTAdpFO+e7eqMWAN5bsagyEu5
c8zRouXApqApNuXUhhayUGlS4JnDnsiX3p+4HTLWOiXwOD0XzkEbMs/au5bAFiqn+LAa5wF4FY7S
HQ/DZYLcjjNpCr3Xc2jVEWCv/ubM45T3lSrMGQmzemSorB/2uz7zrdig9SifKJQdhD+D834CTPE6
lOhAN7+tVBSGc8M7ecqfvNFyOQdDllNcUZgeTulUyOipLnQyfE+LH1dHndkxJ4xKUWsL+/zg1fPK
qbKz33mgEMQkTD8lojLevCSQ81ld+77E2+mTY+/684olpMSqLaEPzTZbVsNEe0ZGKEqQLxYTAoud
qsgTgso9mDf3l5FmGbykEfXz23geHrhIvQP/892wxChl+I/ONt2BdbgJFpnYX4IWEhu3RaWMc/o1
eUopAr/+VD1C0y+FpFDyK8WI4qRJu6nS+vcPPj4TdS4+0hX3Um13YbJWV5By4zM7VCsx+Y7dCFB+
Gjqee1lC6sY59LiaQZJmJZn7zQ21usYIo7YaDLBoAVfRFflyhtSJ4GXfpXWo0Bz+b3hHFKDL2/w1
7sWjmNCD63HUQzRmMRYm1RceqLP5IaJCiGs+KS6o0wmv3J3JIts8jS/On8xWG02WXuS2K6bELqyb
RjicKJYghpRrVuGrOFE7F+6BWnmXCUaxWSgbnOlpUDjvOaeZLWUacoDEoi3639Xxg+KFq6lZkWN9
pQIX8yvXRGeVK+m8SVjf+ivbIUbtU1CHW/teo67di5hsFsfNdsY3s21CfkfT0ot7z2fvfMqZeOB1
EFaa+6wnX2UMpPkcOHzItW7OLWtF5G0mQFXZj5IhL+nmuJPzBfRwXeCdx1C6ELy5l8YmId5q8RG1
dX9zlUvGToT4VU7G3QlejjE4xA9WqN7KNAyrTXZ/SxCyJPn1IdEKH2HUjJ2+dl4JALkeRL9NrtMW
9STzI+xs5+FXxetws6/gnQ3YwcBxFmcbBGj1ww2DvkTuVagO7ezJfmFcPXfoip5EODN/SkJ9rNmG
Hz5xUdXZaEfFvNGPbkvEQEW4NmLlqVxnutKy+KZ65M67YwDX6D7SBVogItKHnDMnSSE+a4PKNa71
BF2w+DU+zwwW/z9d0dT4pI+CX0meiICbUK12X2QgY/opLtKu+yAH7bucu1yceqNLO/KmkZDfECn3
9qmgehhOOtoFH5ytH2lPb130W47YXmSrjG72O3vRFA4fi3iAzDpeBpE1mGQSku1OEIU18U9JccUe
KuFvaolF94mYkHXMFnzeJy/lwd60256eMxFHGIP/V5VI13uEARiTMozcboepIDKCzGkt3m2bMkeE
6WwGClHRWVpYdjUzSc9uDlm4Z81d7cfIFcR3pl/XxNkME0oZUGP7EPYHC7bngT6nLrZhHiv6KQqw
MrWqRK/EHw0cNTav5pumeAyQVDgq/yY4Mb5Q3H1Vv4w1ABP4d0duB/cdcbS8fOC9TUJpg66XNJXr
zRokm8IiVVx8Luh+lzbU9mXyoD9OKeSCVg7ydNBBUxU7dERH0Z+CR8UqhPlUasHZAQCQyROUdoJb
RVPJ31sn4HJcd1Siv06M7fDq7ToXTrNJRzK/EPyIOlU0CZl/obdzm7cGaKaM00sFULE+fIvkT8CF
ML4XP/XkPtRjDzOniZURuVA/59rorEkCMsc74YMuEbE4QpthHv+9DA2zf1k2MNiMHrkP1EAO1I6f
ysG+NPW2mSHdLbk/JtTcZ8TpnhzPF8aUcpiuGRpmJSt4V7Qxob7bPzWDYqlXqCGsITftM6has9vW
b9DMX0zdoowpoXHmsPVQAExqON94tLWOIdaqvMVm4QtNtRURbpCD5f/pp55X/BZwqvaiNzi0DbyK
/7PrZBpfVUjcVb9fJdqLbuO8FhuImAeKwFZgVqDHTB+RK63L3N4hkIMM50/9chThuXN86u/fZJkX
l2tV4JmN71nItxbhgWqMJwqjbjGPRN0x9li4a4ey8icTFnFEJwUIuEU1uSRWxHWzfVRbxJXHiZOn
UlL3hIbNZM53JZf9bvV5JBZPktGVY5VyO7lInEr4yT4hdFnjFawJd93dFYEvHgj2snZ5TERrmCzG
I+4Xlo+7kDluV1x2NoG6E8CeETgLGCkHRt3+DBcW2rWw96ZU6G2wLNyOKdlS5VAAaQ0mpcO6Ouji
J1JQwryMoi7F2VE+kfpWwMoG3Mm9ip+wt755SxC0Lpkn1iOLcZsE4UcNeeYq8fQF3Uj7pu/a9UPO
8DOJqMqSUUmTpmxlCg5mBBjqKPv855r0qtZs3/CJA7HTmJmtZZMKlbR5bzYZsdMEBQrrO5JJX8u1
7otV50IQUIGnR+d6EEDvhcHBoBu/yeziqgN6OLBDflbYuiByhEOUsP7DUM64ElQ7VfJ2JQzMxKvq
OQs4V1qgthWvYrlEDUFCeaisLR8iPWTInIPMRm/Oyk7W1hufWFkL9GOifoQUmgw7YT/tEamo3+Jk
++cf4dM+aBGsyEUGvnoe3W7lYzpPUHuKpsicsPAK/rWEPxlUyXS/3PTkH0UkyRqaabTSlCFK1s/x
5kI1zslRFkeD6XNCksSbpaTimUOqbjLov4dazwA85KXFV6tdWYGPmIKKSs+kvlecdvGm0Vq/I/aD
uR1yOgeu5TMw/jrexcZx/SITlyT+WZ294PdnnCqkt84SoRVSy8TqMp7eIdviUeceveyJRFG6LNcX
GipgwvRp+O4SeEhrJaCYEg1BX7ZIdPBeaP7bp2uEqVHLECLLSnuzb17GN+XkNsgoO3QzBvnT4aUh
nIjehH0O0ztm8F8uOtFWBVZqB/UEi9vbw6K+2O7jLgHvhQmmlmXL3b32DP5gz8hVsP5VmBdfZlcV
3mm8+13CZomrLUMdMVd/QOxD4u8eCcXuHV/AXDM26mK26rRNeErHI601ctB+xIHeCOA1orPyZWD8
W23ZopRMRuBLFFFUxrG0q8zIY3KX9t+E7Qhks5H8LRBe3/N5SU6USLROX9O8h7irp/x2dDBQ5HD9
qiLbOl/k8bj9C9sgAOIu+v8Tvid3b22d/bCi6gXSwlmCiXjFEBoN9qy5l51eK0kq+Xq5PuybvZps
fNslUIds9SrzoALTGvKEwHmFd0zYSqtytlnyDtZeDDbGShJ73f35R6+SNu7sbCAxbMi13Ob1U5Qj
UImyVuuQPJXJRvJh40mbekwwNaeGT9BsaTaxE+IfBJjI0IDgU9vH2UFjLbdVbCatgJoptUoqq9fV
urmRG56ao6xpdHPKPmF0M0LYpJMvjXfyjs9KCZnN0GX7F+Xhd5hntUdkDdeFFZ9xdozvJW5HUvwB
oxrMz8deyQDh5S3XYSBX/6AZY+kpyqQutJtVUkoH2T1nS7qS7p0Rnp8eGjxR9kdoQmp/kPo+1yGW
dj6vt/mbqhpyhdxiBD0jdJOs33FZPbhJHWmERxSHu944Oc3DU+tTBs316yYETIwGTtSIaAQCPtRh
mRbT2Uj9Gmagw9aON6juKMlkcOBEMGdVPUYjswdWr6ecRu2L61JpB2a+1B/uC1m0LpA0O9M4V0fq
YLCR5qWHyxQ9d1+SdXZHNYialBKZmT8obx+aZ8w0e/+HGG3AqLCYaUdywkZLcZ0erJ7hyI4EHn8p
iFGO7ogMpdsLtHCsKaGBy1urulxSahlr2dn25BJN4ppSOKJ9m5IpDhafqdpjUcsnfm+ftvl0aonL
z+oR/EcBTRg1J9wI47dlaDInrABc1Gx2J+YEvzbB8zDOkNzEOLlIbozRbRNst99neW0tkFTPujy4
juxG9t9FtPz1vQg9hAFl9sm7gPH2jytu+YstBz3VimkjaMteEYhpbAfvj5sNuWHHdS8gtymATuYY
9BZ+GGqkcQCzVMMAl2k3ePpcvYEj5lSWP9xh2pNqD2rrkwlez6oCFp/rXAxpVhreEh3AZgMLMLFo
PbqaE+PixFjsDbrd3jXOYqLpHrxZVFVfLlw7mnH34bdQxfQRoR6WKEk2x88E0W3BhEgiyun4h0ic
UxRK/XlGwEJ8grKeGLZ6hTtYntrUFo57xiVQxlykCyFdwo9noyZQQaq2DLoUROZTtAy5kff5uwMG
mcGPHNATMWZ/Wq8a/bJ0B8Ak1Gij4NEnbzjJB1zJt6gc+atMAh8nTKO/0xviu/YDPXj1o5D74GSn
HVXDcxnl5WJl5G5VDDhUTz+VN5pqeqoM0t/SdemQ4B2b2u3PcqtwA43afUeYCJrfgoAVQG8doVGM
snySN6PHv6RPMNhFupenLtpF+JOBf5d1ZtApUhtoF20+cOIC6qtFFcoXbtcOSawFQ1FIo9NyYUBD
ZexG0q5fzhMttB8xPwwr3l6T/3hXadjZzELBeWVoA7j8JH5k82hZTvDEUZOwkRh6o0/8tsS7idja
qMz3oqpoQSANhyrEEIWofNdiW02zh9PVrJQ2IbUxDGaOEwatrU3U6gvrhc5Vn5Zg+U4VoXseZNbP
BuGyWAnc94LbXteQiIE87ieeG8I0ErS/bNyH7i1d0I+vrMjxkSR3tnRx61+znvwkwzfxBE2LsdYT
t7SJjdjBnM28fp3+kDtsFs4WS9gE8TAqIiW7Lqcon4neWfSxMiA0qTxr2dQUDTuZCmjcXtXp3M9r
Hfmvmp1hgQnig1bONtU/1GV8rb+/QdMkvieTLEWai8EeOt22QPTwrcHxumVkH2wWNQ/JesFEDF0q
FNvf+YgGeYzqlH9LjoPL/6QUSJgwexnh4mqLl1OSD5hbIosaJ07KMI0W/+bhLbiSwz1P1inK5OWW
OQlmbGdp/KkkDi84IYZwq529IMAzDYZ+7V1M37ITFbTSCax8oqstDPRKTMUaTzyS1dWNqc/ZTDoh
HYQAYrZj0jPSMp8NDZUA9zcioVGrCqvi82mOZntFxcWGL+ix74IFyiFHCKhOIWSyCNH+jOVaU3mJ
e2nUgQiMsUoYg6pynebske6wI5UTGl11notWGNtrYE3Rpfn6B6TmYIRES1PU+5gnqDvNoSI2HpGn
eh4wA7RWZpvp73TbVeo5d8e7QUfeUs7kQAIafcH8wA1h/6V+FG4T6t72/BeQ/yqYRToPRmvOb6Qt
UzBwIj1/dxrSD1kjeuR8DbJnZSP9cVyk66QOqXeHlhzg6f2a2K5XmbYNK3wkG4KoPRDVXdHWJJuz
DFEd1DAikR784qikUQOhSNFWAI0f87JHG9Ho9Me02nEuUuskAi+yJCXChZdsy/gBS1CnJdXEXkkc
oULjH/AUwSjZsuqriQIpA7LEJTFdO9zO9mCYEYrQ0VAvBhCDr+otePZyWxwCjxRl4GyyBW6/9y8C
XGV3ZeiMSRPnZN3V/J1M8j2at3OXsg+3gBz3NZagAQrBRcAP4sgvbR14eZcQ7cHy+Ha3/SS663xc
+UrVFkcZkiRfhKyol0UMzVO97KNEVrolyi9xwHggZquJARuA/Wm3E+0osXY/Pb5j6lh+PCG1B1Aw
BV49k530eltSLxxMBLRPFnVG0850n5vAYXIgXSymELEs1Te62nFqlnwbDg2m8vMDUw7rfAnKzgIL
2N2/Q4uXzkHqG0Yu+VmhJ4+wxMxlsZo1Cxv8g8EIXEUj2fFN/SAaz5u79gGWHYxFE8BodkhoFPH1
Bl2s/FCBInVJnaJ7KecIS67S0/uVw9ShejJBFjOde2y/Tc/hwdcXGHHQmm8skiHf5doQZbquNdMe
q1mL6rkcL6RoJ3A/iacXeAw0qzsWNSTqfvpeN5i3Rk5n+B8flb636QbhcLOd0k459J0Lifs3OEMU
k7R/qUgfpPl54lG4MBTgPHQBV1fHtiv456me/M5gvI8VWK2hI6jpoJm2bg4S38voIpPE2unRyyed
o7E5JZHZWBLLLjrgc378d5JVdHXsnFAI7NeP785ZUdQPs9NQU1dEV82DBjo+B+pTMUiUoL6+wsFZ
mjCbcZ90THH/8nVN0/AcmxpR9BS2TZkWgG/k9F5aSZBy/U2TvHrz5Tlfmjwku9r3iPqssMhwuTjX
83ZYnDVIrFadBHxaLFeMGuC9zOjRJ5dwHdzAvPEjqirty2TfZOx4mPAIDC1Dj9qtOzVV3Xtyj4Nb
tScAtqhCgF2HRCaw4FMv6Ahr62Vd3XtdoOPMxsMFF7b91DYj3F03bUsnjRHa7Lb5pd564Zucy5ha
OPa//waP00h4TM8ZQoy6Naz1CwTSRS8kmS8rK6bjdXhgI19OozN1qVvv+enp8W4DIKyVVosiEnqK
FUPXLRRWQzLD+tUvVX6kaVOV0fZE9ybSpaldwC+2ebRudadBHQ71wBY8U9ee1rGCyjSBDppu2u9h
jej1eUfiODixKFOqm1KGl6idNj47XTjHfgQMy4Kodq5guNeO3H7EpXpvzWM=
`protect end_protected
