-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NClGvze8GAxNzj9WBdGy9GVT4hKGXAr4fGL5W3EGOPzhbMBhA2gKLBSqn98BFD2Q0fvhv0NhtkM+
53Bn/UrW4eK3TGS9R7RXzj4Bvw2G/9DKhseMGNgE/j+Q7tx8iYxl7OGaKeezsODhVC+gUI8iR5MR
FvVOApuDjjsQ+VbmZcIaY2ZHn1foMoGsTBb881Jyun8v8Gt1GcaT7TfdhpbND4/WtmFoROKJ7BWv
m2myI8bNOZeICIZEplrMS/qWU+Tngk+SLiPSmoyYYVH/iAuKFOAp7puhXWSLkug4vnZhxc+wDizT
Y+L/Qfums3azDK/a1w06SA/MKbWC5uHG1H43rA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
CsBzpAMEfHiw+Z5oNM/jZIL9qkvs/lS5WCMqAOy7z/5u1W4PXBI0UbXon0tg6ztnw/MRi1nKe0ie
IIN3mZj0excXB5Yy0eF2KBu2tb4mr9PwEfzi5nKQFD2gX1JYkbFQ+653CaxHr5Ep4L+8s4nKj0cM
UYcgs3Tonb92ilL4spLVJSU7OgWwdK+bA7AimJd25zjuzHh3N6tW4CIzOv/SiZy7qNZw/Wl/8x2D
hDiJp4N1A3fvlxJ4pPuTXN5oifc+w8wBZIq3ZL0joC46FE99ukELzATyysqYDSeDGpEEDD/RYqS2
7iNO1Bm7ypG2iaGunnSxvGfYRodalpmy9lI9ZWiBgw3iA13+Xayk3TWv/7Uax9m88lSEw6assTUA
E7ioaE8bLCpAtx15HInyw1vD2ozPNGKbDpwKLFxwdrIfc9FoX9JsftHnHLbaYxsvwZiHu75xNb33
ZzYhklVLEur/uEpGgm/R6NyRfoRHPu/ROKWxw/jA7xt8xWJ4xUAuEoJ6nI8rOBqRT6SajABxvcvB
38aZ7lmLzrfoVOtWrfJXZQ1wRxiRYnoP83GCQFycdehErGd7rLst/1ejN1Zp35poTYQSR32SNIz5
rg4BgTCeFNGb9PftavIr6v6JJgeFeou17pBq2BveeWrYLTOIsy734H2q6rpZ3cHQmRCkYF9aaZVW
MNzlmxcYFNIeijJqYWyHi50m831wMf+ffsSP2S82KVURo6OA/7PNawJhqvzAXZIeX7xF8TRoffVB
1AKUdGUZzzUnhMgShcAhfVP+u0kDyHx7ZvOfHBzUDKrBv32/Dl3STxCZh/wGPS9gi6VtpKe8iqWh
axs+bWDRAmTExRvQkc268aIQOtqe9tDgCn9Ud00CT3zPiHTay90Qi31CYiQZrGsWIgln3XGyEtHi
tMOJO/YbsWrEmJVcDvZ9i6JhypyEc+YTwkv3402U51KCz5sv+ts5vwQOd3RQ8HbI/XIB2v+8RE+w
dGRT8copvnYIleoeifCy1y61m+nEcTPm+bi0mztOzpz5luiz0l0gtCcdo5gDPr3oyRuNGbaICbaw
uEiAiU7wuXOB7PQ3BJiLG8wmbJz63tY/mNM+5EJauYwVz6M5jwWzoJj8KmJps027m0Lohj6UstU/
boIs+zm6u+GMMDw8KlyAuipA5RQAKvr4d3RxOjtZE3BS/HBOjWzXzpY4TNDTPWpUzDajwqMiqrVE
vW3p647UApbJnT2TxeMlOCaJ0/DOiezMrWgSWZIS4mC1etph9n3alcC02qo56/qEy3uLGSld102V
PMAfrzlN8WQytXyU/wJrRAL+bMetVBfU5vNZBhVzbtA/P0EEaGLMLHYDdAaxVyCZbijlGhiDfTkV
9C+Eb6PcLerShfsHiUhTAleMU6ZcT8evVEQ8Is9AeueTrluUQgvmJcSSBe/tIit3F9pf8KZ1kNtf
h4AOsSz6d7nJr756komHYCa5Is9u606X35E668z52SSsrLvQKoi2Nv4cq6SSMS2bJ+QxjgQTr9Ij
ztvePqAYEtqJIQnc7UvUX04X4nZzT3NUIWNmJCH4eRb62XbZOY47US5XD1/TK9c8gQaxOZQH1Qt9
Oi9bnqC3U0AQDw4aaJWGLS80y5KuDeJJbaOQhvr484atQEuJ/zc4RCSvWWKa30zfa9kqimGi7OtM
2lMtatCyEp+h4jmulTWpTn/muS0xTGVvyLVcXbhdrwME6aDhUYj6OLzNkEBsAIqOOOPiT8H+tc0l
CPswQWfUkvf0nYWoruRapwZdMWIWnUVCdqr+lxcmScCkYpXnB/i3iT743a5DnDY6BrmG+Vdm3hVM
GV6/DQm/DlsHgWYck2ejnoie9lwojXW1w+cnW2uZokDeYUFMJbH62S8BnYAcFmGfa/9fHpr26dQ8
XGt6Z0i3Gd24TTsI7yR6yyEQBJqtr5LoMz6vub4ZEaJIO0NVSiFGdWJ2VR0ti7/8px9Xao5fLmP6
d47rYewB2zndImaQDeiJ5s4oYBJywA2c0Co3dTVffVKpMrhDDKuOkQYD6qXt3+A0F/wgwKrQ/8Fq
Bk8KtlWNmkTCXunlO5iZEHHT7Yul/aCOByeXxTwSmCPWNQMyHTstYltdIPZO9UJQeCYbaSIZ0lj8
bl533TnmNTHe01p9cIg8A9Fnfo7tXOiNWNVamfVw5msTJcImNoZPQhMKeph8/oi9qPgk2oMj2oWS
4sJ8DrjMwGQN2Q8O03M+KAI92rNTQUEoD2IYIZkJK9UvGO/WpO4jz0WzLBg7Z+1NOodSpjrZZZiY
H6PVFCFPjTkUhEBEjyadCeIfPZmb3fizd1GxW3DP6Rf9kH6+A7JaLvcQLdkzfdhzxlaBMw9FlIOw
ANO2asCyoe/ECIm5nygsFSY3Dn5OdC5cR2amXJjM2bOKiB34Dfc0OZhrQToIRd//vMPKZvQVDdei
TynNPP7e0aarrI7la0425vVWGwannPFo8s4BUp1KY22fkXt5GLwaODl63RGhUk1ae3e/+e8kyalY
dqVYGsXUfwDUomxBTrimA7oVhiOPnX3Qt6rjJQ9BgR+mUwTIdtlbrVSJxgd7rOpGbG3jE5y+mLO6
vowChmL3lvC/ts18YQR2pdxw/6ZVofughfGWo6sgq6CvQ2p8y23SCtt6RwtUD7Y/mjtbx2tLKEIA
SPMT0fFA38VboVUrED4j7fLrnKYF+Mz3hxBsiS22v9610se1x16VwFUSQjlUh994VoGS9Vo5rkVh
7rF6tt8WlUWUS0UsO1H0L0Tcjn3g05TQbLiXZlUyrpg/q3WhIU+ADm28H5y0DghXzM39EY3WQusg
nVOgFMEblnoJDRuo7g9Ygt9oDX4/66emuE8k489EoJou7R7koxPTBSyiWpn3gNlzqcVRJe2xndWw
dyWRMmMKBNqztkEJGKgNXRdORYCLLPgg0Bkbg8oqTnnPLR4Q/9AKqV1dHrQ88ZFrGW6sgb7+DDN2
iK5e4PL8DWyTitqE7kLoqctMrZRUlm+Vz8Ze4QP3ncMLt7JFhOqmxXlFfPIwUic2ejVJHGsZkI6P
1E3TfebK0OLpTYG/oqphkjThwnW+3e+AsZcveWlM1fFmWsqfsE/7mGa+lYwZsDl2eVqKcoF5CGif
ATYc549xmFw5/PjO27HRAfryd6OkgQh/Aln06fbq8OQJzBvJR1D7kjdf4j581TTtdV2s3tXKk5MT
R+P6PdunzzWouR/57/Cgg2A/fA/E7fwPfmZ5kC4MxFCeETV7fnwMnv1HTEX+3sQ2PJb1t1KdH5Qg
XbetkijD0WDfownA5oY2xSGFpDkg0ZcP9Z1esUxSX4iGtmYAZOFcEnTH6cOCCja6yU8n2UMY93sZ
yzxFmJDb3OVN8x6i0WTWpz15dZyBGLRG0YbulyERyqgcU53NMi1+xaildCp5F5P3bTD5AU8Z+8oX
+oj8TMLvvP1RcoOSFnhngv1Mzk6C+9VKAkWvX4hs+y49dZXlENyWxBDCXSDv/qc0b6gGRtrGO0PV
0JJ7WmaSM55DcQyd3Oepi10iLPyS/mC5sSi4vLHA08fS1vm/UTm2fMv334nFO9WFsK7MQ5vlnwYG
Gj6vnlQAye4Q5HUqjXZu4P2oxjcbeC5ynAI+dMqbfluAzQUmw0LNwj0zvxwBPRFFsR3/kZaTRZca
A5U05WjF9hpksTGm1oXtzAMKDsGndRa0ZO+GHuwwB2wsbDM9srFaaUceqIVLt7ZFlvAZPYyIocQM
QLxOE/V5QxpuxkAhoekXtZb8jNt5I4FG7EX51RuEny744+MWt4EcIAJy+XGh0gM/BRs9SoKfLn6n
t7xQCBXJfAdAqXctxtSnBpYb3uX4Rkg3UcvUAmsqrP+RRyTzcW2QbArkq5IrJLqbE5324r+oYiG3
zpK3BK5zNo9ULhVHUsQlpUTeXRwCVbcrPO/jG2TlSgbPDtbWh+RUQfNaymvfcXCWV1v/zNUV2/G+
LvQdVGytkJRUcn2lBKLlg2yXyLg+le5d4gUSX0Mw5H3tFrYik3hMx4w7LxBhCOUKiDgd0hF/3HGK
OcUN6iBr4jpiheXyw6iSTwF7GPl9AygkOz3tL5e/+nnEioaJ3vgW7w4FAov+tsuyvE8sCdbJbsy6
tpqh52O3Rz6sDBSnG/IvZuQSue8mNLxrEk547fn6MB7mNWy8y/6lNWY5/XsKJ7GdTa4kjMqNkGUM
SgXP7VL7919NsDYQt3UKQa6n8/U7gHp0jF1D89rM8t0ka0q8AT/gw113N7jXRWH7ljBXQiD5EdZk
Xgi/u4O80WU9pgoffZcNoxCYUui31ATxeCLZMooSj3Qdpfez9p4i3/onbTgjgf7XGJNWM5YAZe9U
/ZSGu3Uzd9+85aRw/UaJPk96+czrbX/t8QbMOZURvS3EAerSV8C14rbMRr3SNFKUzZXATmiAY53v
Tdjn61eJtk3tqSjzFKpJVtJL0HCtgBk88fBzaihw+/Aqt2R1k3FumOFm+mQ0sagRuefszBG42+0m
M6jaHPaxJ43XLinFDiOHLXb29cdbCD1k4ShcaCNg08nfoOhl4WjYR01vhvSu/aKKjJrW5Od1Gn95
tsKFWK6yoOGRZwRTBGKvqHdxq7nCyuOvP7i1afm3yL/AgJbvv0y/9zsjw/wrnS3rL8PBlOuvMk5E
mpiuuUu3YWTo1eeQpCVZnREAoagVUIAFY1Xnz7E2/jI+Rvbu1AnMCKa2j7fA2jKxLzXsCecftILp
cbodCyE58RD3fbaDDPzI7ietzolSArF30AsajDc006h3SfmrnySA+pZ05n06FQvOzxO/f/dw7t4b
BqK9Nt9Pe1ss2Nz/ld2O2ogKND9m2YI4Owur33PItYAlOX/IhxY8/TZhpxWk1F2VBrloBMnm+GTu
0rAbkkq/sf3ssAmV+EvRMbL/MF0Nma3TnqlNvJJFpVlvqu6ZgbABqiNjho2D9H+hetZy4e7Cj5W5
KwaLlVF9Q9YUC0SPxP1vg4FT18hnS1Zo5bnOejTBuRoMFkZ6aDyGz2oxOfYV4OymjSEjodCmHrVc
DfQTrXAkDpfra6U7sDhcFRkxmJe6JFR688sY+u8Nwe+feFdh1g+mdgH8+lAM241qfZ11M5eaoYFX
ErMdmXgOD2EK2JZLTMECToj4qjZSRXcFBGwSWgZgL+wBiXqPhzwjjiZYn0cJtLSPwGZV7q/jhprN
2vR1Q4hxrl+HUcNaHVzeTitzfIuiNlREvUOeDTVligvcEn1L8zDzVkrZsyolzYSwvUc2PsaqbCcL
PQZwk6dRn69ZMXtdfZXNoBvRyjDpMlhB2tSIegiKDAPWmLmbdxq8ZMbtM7PoeOjUrelJI8Zf4ite
/KL4Mwerx84Y/aDI+sl/eO8iByJ3VVbvnu80MWH/ueVMX/V97wXNOf2a8m7NNb+cgYwlkoenVnEN
tiuoljF/vs7DChCr+MuYhSYG1zqTj2EfKAAV9SZQCkr3LMtVW96mPhcLxSqh+A4QU7ig21Jqodgi
wiV/5UPSu7o4e3vWLfBdTO9kSD8/1rlaW4J22Pn9yTRp9nS5QK37ByQtCoSBasl1Er9mXs3P8ldv
qcfLfqkaEQWHKDNTGEc0qrO+eF2Rm3Dwr3pg6cMmlfycruZEb4XQtZs/YFNaNGJ04b9PhqD7f6b6
C4q2UQZi1hlHRTd4gLPF8B65sbYcRiF63p3aPKvuXGoE7k1g2aTtc0KhMmMW0xCFaln6yrlC3GHy
8gHccMMoiTX6xvXje3J5lHkImJ0H1kJ14b5WLMIWpkKGaxkOyrD+rEw+aN2rheJ2cmO/hAAwNnf3
GeoMAygyJswUpBFdWVOH2DQ0atIY9p59Q7lPKrrjqCwSXXMr6lPS77ljQO5plECFpsoBzq/LJn9f
rgog0XYzCsgYm54EK6KbGWhdbTdmPecpZhtmmo3s/tR6gsZUeq1ieEy0ye6kL3sUbiNyf8SnKDu4
7g32AjtuVePjsBbh07BsmI+BZWlsBK17Cm1cgzRivzhmsciu9k+s2HGBtMOIuFY6yDQeF8wGWhMI
hrLbwqYBdB8Y2VdwWGvbNV9Yr+/K4qTi/26RVyhTRzbjuiq2FqFZv6rssSukW1aMvCarscyAPWkn
rcLzod40AESIj7gQ2V1ZL3M9OpOL8Pl6XQl7E7Wmw+kNfJHuxAusnwcgUKwdIqrDbq0wihvuPn24
IYEF63TwDKTQ+q/Yw0ujMq8iYGWGTibH5c5CDbOhdazVaTaraxu4B5vhjsG395akyKGfdF/VH02D
hHouovXixLft07UzvMMD1n8fSHnnR9lT4ZSGA3NIcY291/u2PGO0FqTkU5Hveb578b12DwotjK4U
riuL1E/hBbAMTCgmq9kXAmmvBY65kxHK0jbMySQoO21QsKcIX9EAGhMe4x4IkO36FdlbhHd/Z61y
Ju0tahEm59J5nkt9QtWy3SKT9X09nLg3pDiPiI+Jj3zlyZU+yMSrfKTkEtW3DnIUCKP54F2SBSol
IDM0gi8vh6KCbaVDz2VkwTL2b43p3UMbr9EfS461eMHHLG/Dh8XOjXYk5s/I4fUvLip3diDNokgA
pWJPyqZGPD2ettFXvzd4uyrZNlXoCWIpIlA2ktsDCB4lYf/0iitdDTo6yi58h+EPKS/39o7zoA8z
jCIRJzt887pf50xEz9awUWkgCvu4gfU26iv3uCG/1r2GQ/9HjjfCZA/J8jMQ1TDyM7d8AUp1iNk2
vTnj1ceJmArIxp5mh5qWRv9BmPKRSlFHtuZOj1ZQT8Y+LCBBxDBba1Fg0RpbLBw30GwI9S1a7Lsc
2xmZ2Wj52wOD0RhuYSv34F6jyoBLSpz7TA0Crve2O5Y+6K1YCbBHlu6HUWCe5xrB5DflkYz4IZrs
njEMsEky8h8OggIW2oABsWY9e7YQ+drrDwW9RDT4vhFzE+yIFJjhCitP7N8pL+R6SXui+ZnGIsvN
Z9A+f5Kh/ORKNFwOyIYa8WNQnEx2Sp0y4XdkHLu713MnYMEchpn/WmpzqEBDUneWGT7ZV0gFBjRK
XMAjtJ+DNailWt07Mu2iLWk+w8lbeENgJmbPW8ztyBZlQ9JFjsUfUdwDWd5af1CBlQ3Hq0qggj+l
y33OgmzAqnvwsAwY20KW0/bNKwuJpAK2L8ICSsQL0hksP+FC3obe6PJJ37aPYFMssQjRhJIhqJqS
QIL9zw6Clnl1qDRhMR17WrpGqIZPaFlz0rxMNaXz5wx4lfwjgN2Ccojx5qWl4dixcFulZKEYAGSb
lRQWbdHdHo/tg+ORZUVsuLjY90VNfatqS0UutuwQi2Qld4iUHoiKcB0zHL3Lifqp1sFw+my0vjnl
gbs2AEP23qSt0Zf8e7MWbOCud1Y484TVNY3D6WAn3RALxF8SFxqBjrtE339Ik/LWPBVJAIuJdUzP
s8Yd+xmlDqShrBRyemtSTl+l9zfgF3Tb4eEp+LVvFn3w5CTHM7rwMDh8ja92jdBKgYBVcFTwVeZj
6luXffe0f73W8IIttNfxYjMr9B8zQUSPg40wlBW0lh6R6SBS1pj0/Ev8VledDQT/fsYtqlFcjTGc
kB1PydEs+LdvVTFSeqjNvyAf3yVY/BnVlLET5VwpLvx58hzi8owWUU1cwKoGDT3nGF99cKteW2kG
YW2KWeRKXV9sW7OCU8Bxp+4Yjy7Z56K13047/Gfmg9IrYsqbcBXETn39vAkznw5kp6gdGBGsby/t
BaW9iTrijGF0lPGxWQ0cmio8x5mlSehcdyPdx260Y17noRvvxXRNK6eEl21lB9Pk7nKVVOS8HzyU
gihDTGntnuPoto1jap4IkbX+1TqVjz/yLzjOfNfLX7kYH2jXq0JYlNTFAnSTW0LSGVqwCH0AxR7O
YJxAVOB+ubbPjSwrvUcnmnpqoH+Lqm0/d/XEe69QvWSEkfDyu7yE0gaDCEaZFJLhRpeO8p41cbIM
xwTZ1/dsr9GYPRZxlOtBKXINYlwtOCiCPd33XnpFkcStFvNriEd6k+RRa4oN7W+RGznq554OCaMK
0CQTovf11Mwcku3tWZlueIR7dG3Ake2cf9SzNeyB5i7Jx88OwJ0YL9LrGSJ7plLJT2WAhiwd7y5v
i+ki2OVk529YlULd9LFWP1/TfnrDSz9Xx7Kvux3gyzbOZJHO3wsFdKftttYz2vLPpoVCRdwqgJaw
v/WaOS4iKGBgkpHJZ5CIxcGL2T+/mKVh/+6DxBdw/vkfvwgwhRxD/WX64YL9Bzn2hGGaMMf3a4WH
YJEUPRxWGmcB1SpwY0Z9Rn5t1FCgapRVkWq3OpIgOX/R0CSuIyhAaKNNzRArbGVJh59wxsNRLhdE
NHSg1Hq+lmho7cxDS4cgcw7zR4t7fc/QGdHqHa0rsW9X8zi/gPuyfuEBUyC7ymx4FK9P6sNPri9U
01ysE4ICSaOjXiOaw9/hAwqqO3+VYb179yhrw3aHWwDYhS+VtYs75cVbSyh5uS2tu2Q0oWdVHs8e
xbJQYkZKTPSH2/Sdc39JPaNKdYdE9mwr/GW/eC5tdg/QHLbje9peS9PiVl/BPPOXAPXSScaCUJhW
puifkFrWSThzNOgahQaZEjKo72xEWnNOKqplGXyRpEoE/Gfwhzrx28t/vSYKIxHRvf/1Ub2dROdx
LwmfDMyQrRhKQNjv9pM0PDgSlCafTjT9L8/rYC8fR1SdTiDVKNYVHgzplrPiHxs+qx/ZpJ6o+r7B
gJE7I2mN/2zEcc6E6i8kUXl+m2NONM6EiAk3WUrDCzo0gMjnt9jF2ClfeylAzashl0w2UEqlawLy
UFKAPW9LHlUWxN4nFSnZpQGyM8/2VS1sanD6X0EgYC9y+OSeVQKxwJjnKYn0XW6FgrOzR/IhlxWg
Dp1LNkMzUgdqx1MbMDkj+iiT/xHXj9BdCuDluO/AIt9X6cKTx+JvonprUQyzwzbuFUuqL95nj3d4
OXdXT5r7Jrss9ioOjKs6RU56Hv55mIFJwiOrEjrDa7CIvXz7UZAyg16C3nxPk0XCZQTG5wUo5X94
owB6I2n90rMKTYdbaqJtZ0PwuOpVmBI3xRiadUW/24IUcY50nYEWV670MCst7qIowGEw9B96Kivp
w622sLWDsR8A7C+L73zOD1Zpqj+ZXySb+QygfpT8qYKFZImHLYC90Ec9YNzw9yWsOqY0ILA/6qwh
fwc3mZM8iyoOrJNeiwGDVlW1qHZgEXXMAdCfHeDXo48JxUwRuUzGKzkElPAo+AMvNM8crumLoqXg
nQ+oIw2eOm4wyRu19ZdofZ8a4cx90yJ/Dcw7Gay4TiNkuywgJkeQrKrhg4RDYLHhikoskP78QLZh
m2yFfW6rVusmXxqlumDlXi8vsFaQGScK7C8gC/g3oEdQfnrOtdbS8O6BWVY1tzrJytsEcfH3rONo
WrcjBcJ6NqbtabPXx0eY7ESnSKN0oIOKkuCwVIK8Yu/T0MpwVxCHtgSX4ngUw9O/7R4aL7iqlxVZ
Q/+NJ1jepeQppLX7QJWQUSxCR3d8U4iH4wpMf1sfCWeV/3jg1Fa9UJrKv1nhfcrV1PdN04hNx/k2
qOCaBaQ9hGoURWeia9MgxoBnmgmB/UUcSxc7JwzRbFKGiHBQFmyk7XHPuxf/olo+30s50JhBR9e0
4oasv79FRoTdCEbPxF2MvqynRNIviCxA6FS4BkGOtJViv0QaRPpGz4EcRwKBpfdHwNqbHIapc0vX
74fte/ayXQPrXZa8eWMPsMQcH2YJmNN36qkKcaQf3/zdAP7w8jyfQzuvq3nu/f+OxPzd4s3XfmHs
3ZoLxJH/1/abWga1DtyjW4vYVn6D6KNz2SvLGfhSbMlgWr7C9ZzMIjJdoMHgOrGwj6sxz3QP/wxI
OIxXrFTQSUTH6QsWz1Jk9k2FXqAC/bSTctqIR/D+YJ45Ud2v+Kuf+lh8oXaNFqZPmsFTDYEvXBm+
6qRPlsJWR97eInHu91TV0EoCgKpx3yXCfkfF8BVTMIC2j2LCbXAuv5x+Tb+cWmp98UZ89QVyseaa
CLCr85/B5G6i/67ykWDNAxqZSYjEMBiTaIjLTfLuHz55zGVxr95TLP3YZrGh00FhWQIMAXSHF9Xx
jKN3w/OBdYYvWrDkdTRvNv0GZyU09EpwPFVuNKTGfpENUV/hzi8sLZG22Zyp2aBbk5qyhB+ypPS1
YdYQR8lO7Qpr6z0TGHL1QKNl2uhkeUqD7AW85GtYoFYrKNz7zg/RUGrXELSOVklD4sVIoOsUhB/9
m31KxR/37cPadLL9jXSPGCDNzjDOvpWLs4iGagVe/G7Irar25sqDe6y8QfjfeTlDyz9yBm9M/qTX
3X0yWICV+mDY8xQgUZl+XAXXz8J2upw+4CqKMXGATgHTWatq/qGpmxjSp9qq1eObiJgxKmRjXI4h
Q2IUHYXE8hHLHSEfalONB+uXEeLxD4lCWlq3KKapM7N8Wr3oJXPF1d9SCdHwTQIzrVIpU6+b24w1
p15KoIMcphYo2zIMDaFS7DG2qrjzNPTN4GD1jl/Z/Szm8FFYj9r1rTQq26Y27IsHcdAwTCVBB/El
X5z2thQOkebKjsM5olqlgciz8VrSB94gLx7WbrBn89psPYf9cTJsymRir4/qko0AemIDN1y1HZV7
Epo5VtxBw4HsmRJ/6MKrHXNO2VtEPeLyXfS6n5804YvBp3hC4/GYqOVIYin9xW8muL7khRETUmhP
lDRWlvM2p/UBG1ReXG4JjvwdLd6/MJ4ryP3QG4XksYeesASy//SU7RQUaj2ZDEtz6DhtVBdXT3FU
akh4rRZ4tY4OOiM0gVsK6Eu7Qi1ogyPYRvyzVpAtlPoCWHLIRGiCT1led2NbhMpPxx4OW7wrunQL
B9s27CRF0XgSYXXYvjOo9Gdc3vZTiFPMRd/G7uh+T5BvTZE5rd1FKUVBuCz5n/2OlUuZziO2lQPf
taRBSB45hBxlhSluKXCLSvR2BwHmtTjVF8yN0JwXdt6xCtZeXPOcVjrNyU0zljyIC9eCRcSOGagB
FaiyaYQ7L0bMM3QY150XmaUcyBTLNxOsVYwMs0Bk1sN32IIwg7WlRhEpO80tDlTAY0GSNsg3Ut25
vSN0M61EmcT6F3+TWJa5G44pcBtL5LKIOpujMcXS8uhMaurHEUbOHF7zbF/BUYYIACPiD8nAbSj7
U/T1JyA3vrBB0Mt2XPnInzE3GSh+jLSQaNulH5Gbz7T5Yw9cuBMPwNgoCa6Vfpf4coUCEZqAXfW9
4ecHBXHnHgcb1PGol5Ig3Km82Wc259E07kPw6mqvKJoY/F+4GSGVHqaydw5cJnvyXLoBr6MU3F2Y
nL1u3/Ck/kAUzn7QQTjHJUWSQhf1pN2Vhbn3xJo0YDthDnwfRuLGKyyEU9KzR/AxZ8DEaxHI3nhC
wtZ0HZOTpKr/sm1xJi1TGQtQoME3POf0umGB/8BW48MbtkMbT9KajV2VLN5TjzaWKt0sTnXPH8Op
AHgnRvxMem4pRKZusgBZiD8mzIxRZQcBxn5ZPu9ruxqwv9Fey9KU3l495QzLTPMCsGlSOFwVETNM
LSyTq6Ufi01hXh//J3PNUxUKYbBKyMdDKNTsEA2AJroqQfCim4aiMd+EPHkEHrr3NMgnMYHQIPON
M+BBBkM9bY34TKPf2rjpFBmMmeF15ReSETSax7qbbc5IjGeMQ6tW6bd+SxjeJRpho8rAQPZL1GA1
uN9qcr9Wdwq95ss8MfZ8QEK/+3TwHyqrH+x2lUf84IA6M+yXULzMhFtlG23eqZw0jDlQD8qE545F
g1SZN0w9grbijRsp8XOWESUIE+liU7ydFsBkGjfBvMq4Kb4+Q/IWOxKMR9AWm9ZNZUIsQxoM6yNL
CWSCm5Mm5tB4ucV/9p4KtNQQxO4P+4uPFa41Ibt3TnSU2a1W/xGHCwFjPfSEAPM9wGagtbUaXjso
KOzbkojjAfnhSUPZHxmLKaebF3nOJlZYW8QRfzQ7OstJ1ddL8lpsXGyeQWNnbMNAiA1e/3CU4MQU
Jltoz5+tlDcywjXtTwVBHpyDNmJF+2RvsW0pDUdRj/0EVpLVTAq7NPdKLV3BQW5KR+kA7Dam8gmN
DGQstk48Kryy7KNMnvyZmvJu01p5GClX8XPrvvxXaksIOWvB3v31kWaG+KXozoxGISUurdQfBdkf
HfeZBZXaI8Cg99PgPuJF4f9MO1MC08sofx6YRwjN0NhzwwVsLi5qGC7uub4sQfjMDVJ8jqmyNq+T
jP+mcMK6Hb72odpIqc4TcbxFD2m3p7nKW/MU6aOWVl1AwWT99JzWe8BWlCLi9CqDiJzQ9+hq8DGG
WUHT9XKD3gti7+hs4V0A/DtX1q7B1hIIw3TnOtadJmAg7nJaWjOHvKX7xJk5TISopujFblmfPiNX
/+bJE2Vr3fvoLxUc3vyqXhOrI8rohFY2NL5VqEEhDsGXqgmp2Tbqi0B6qyXQlvBCyQmSQ6hJiiTp
OBCK38xt9tCzt9tK6/HN19yrcBChKhEfbCKY7B7DZ6erqVNcxcg1tWawBXblCi7FhqdG9YviQwIZ
kGefKGsHCyc297gvBJ2kcmCqPkmdagGzcDcPrW0rzwlPuBtXCVAXs8zXARu9jZgnfuMAJu5bgjZs
VkiswZsaE3V69dBUvH0tjhSKL3RKJq3kTZngOwT1tq7aGxUmmrsiUJ6DOr0X8B0rmXMp2Z8t+MFM
mnYbT2I3JNksxgIxeyFlB/Ei3WGCpJKhIZJDQMxqlRH+mkg9xRFfWAT6SlXlzOzWhoUxNyhiduI6
u4g0KfbG5OaZp/KT576StypKivk1hpMKLFGp0suFc0TVQOUBIDVcu3HFGAHsriAIlCRn3840SNho
+BKsmnk9xcOf9UbcM+ExjRHprqwKMFp+Tv3UW6L1GzriQC0zSt82+CuIu7xusQfpDa4T9SnkWqfy
MaGWtBxm7/2otPHEM1VYzxcyTpVKJRzaz6vi6UgqdCbOtkwsc42CAeKziOfjbfOg6QBHWs1rVApS
fY/ueefxVs8ZTEUG9lBzHtebpH3ot6KM13qH1xrQaCttGewahVgFXVMMX95ZGzY57yEsm5O7hhmc
jjxC7fpFg5mabjxWzKFgaRO8OTiahOZH5TeQr8LD1Nmjeg70MT6zJmiggheRTlCPv0pZ4zw8O52+
5YTP19uL1WGQ4aYKzTkEy530XP3F7CmtITwShwuqkKr4z0v5M6uSpi44kDrbixYJb6E5Ldx4sO54
XfRNii9S2gv2gB6wot/P3O7xrsX/TMkWM+MEI1tOGn5vNtSRP0DTz5PTs4eE2hFL7QDkWGCaWZxF
JpxfjXDqKClB7+xmRgSBFstnkTGeNDKY4jtLKXUnJX3W79FsaEFXl0+KDnP1zjqOdzhiQA45176S
uC8udBIzezhv/VpsEeboPEV2btWRTS5nxARmqM5ykGaQMLmTu96sfL31sMxbuCn0/gLurFQ9vKtr
fYBpZ7e7JruzwAgkOEU7hPGRriPgmaBohp3I8OLo88Ub9mgRhWDPCnJ6MX7HRlGHaxWPauvYXvi2
0X9luYoYUj6AH4FyKSls1DrkjESWi57W+u6LogGPbqxIvInRvGnqYpnPcJcKpnZe4sZ4mHu9jj+5
gAv6ngUumEywdd9P+dCQW16mqNWLA4zaHk+M7HF6HUrQpfFcs0V3fdXxjvzICSZ7ANrMP0zfotvx
AYCQP2b8CG0JWMkICXsql28t1AEO3TXNUohOhkCJm+eF3vf9zGepr11ci4XXgD7wBF3HISYk4Nwi
q10M3Da+Ns5C1JdeUETUbH7OU8fFKo6mpE1siNsi9OmzxKdnqSBzkOAMqAo+DNhwnmrQZyrp5dWP
VKGEE3gOyHlX/xd3bUiP8eVc0C0wOTdmW4X5+WARoN/KoqmA9kkYEvngo2ir8mKyzNOmeoWY1e7v
zNHuZoYjMOr4w9g40VytcKWEntUM8NW3InyxGthIKMnKsg4geD/GG/L1T6Msd9ZN9VLTXzDhKiMB
qenYz8LyIMZCIfF4kyk/JMflr+Roy/ivhRBhcUzhAZ4D8HTE8SOV18p+X4klQmpFN4zaLzu3Wt3x
nZ/RnbCwpzdjO8InIOwfYgPHj2UXVAB+CTjXumCNJBrIXdkwlaB3HpeAsplJX3Q/WL1aO8+tTvtB
qPIL1KxQTl2MMa8TUKppIYSIw1ZoNeF4stkBJY/oTeUqikKqAJBiltiaC5tmQRM60Foegex3+qzm
Z/r/AmssYyq0SrLCkSMuCNYNWV8aNMMvHhoXMCkABDQqr2qGxWY5nThf6C46QoeWRBUiCLTU1SYi
s6EIGb1ozgtsmbt1MW6NEd0CRfMNu+sH2tQGDMONXXOH2JSkq3I/ZxnDtu7qx2xS+meb9jI1PDbR
gHTbAfKdlCb2I1GzUFzi2d9yjN2XVBNkjnGyInMSF6ir8Sz3rXIGZC+JBWk4DlJlt6EisJdh4ARg
lvk6pnHKhiBtXTMd+/Yw7ZobEgUijdnl38goKV4uIS3+mHikil4yaz/utdR+JHpqWM0noKKz81wn
S37Dcz2ZCdcZH63sh46YFBO+DSER3gvt4S8oBRm7XG4Z5scYPa+EHnLvL0RAdBXWCdMp9zO+wcdu
txszw73FqLfNDsCqCWrz47s5Y0gYIDA6G2IYjLB/04v+NmuGySpq4leEMOSWofme4u+zivvhYiA/
cuzfGW7XN16ES7D2WS1/opsxn+gdsJn/e9q9RVX7QyyaWpyLvuPj3kYTROnAAzJAxntRdWMW5JZG
9nsEVGRcERPwBTAaJZFQDORGA2DfXNyjyetc1NBR3pBxx12sX6HgN5PuFQ9/6hJ97X9Uxxu21b5m
EUF4u0R071FzSUKPBbK8FgyvpUtWsn306wP1d6EA2ZOr0OToaUxk+HZttKQXKHRYCJhLLvF+UEXb
fB59RR7IkKvyTUl3CaMHukEZgDTBwvWn8e5sr2b0dDzENvbAzYzzMGxI4IG451x8nI/8OEYbkox6
BL+WmHMyvvrFueFUZRoFrjm443rVBTJuE0kB3Ozu173NhWqwswnJzfRENvmQxd/ioDLMiQ6nwL0J
9sQ9EEo0rsFX2+lYLd6Y+oo03KFIY6ei6BLOaLLekDGiq4fhX74p0TNPxPYaeIQi7V9sZ0ZfoyQE
bQ9y82F1+tD2nyjJ4OAd5lX6XVD6AGIIhUT1TigF7v6np5QrnxfJPkAD31PWgPENyeM6l0TLKX+l
y7h+Ztrl1oCH1pKCRXpggDtVKvDgE4J1dnQ+75HrU9pdLE5IhTOifq/c/yozIiMDl7svfTOmmhpC
a9VkZC62268gPfu9I77r/6AlwHKm4/KT/CJd14wuAz/Kuqzoq2risl1+dfWYvFPSrl4HAtZW/qHr
EIqkFT2IsgdIlKHxyLIZmOYgVHUxD580wbIhaA8zu+2OergKK1Q/Mfvvp3FnSeO4eecThZU8nqUe
yUzckM6OjyYaGvjnOuINZJZLldYTTpZ65KarKpL1xdBpHncJ2OU0/QdEjgN1Cg+IUDqGGz5+tJDj
e8RFXxcxXMr1NOVW4eoLi6WU6cTzv63W+Q+OBvZ1hGJrrS01bV/GZPL1vOtZukv38K87WECv6lr8
Dzdb8eSyyftsbkIEFPxJUMPYHZF9L+vTr482P6hwoGGrwM1GcUfVa9xoMnQiNhHBiLGpZ7qCvza6
Up8uicpf7+sTmXq3bdD/9CkXybGNtlhb2xeYm+oPMQ5FXXmP9/bKvNiAMD2fDs3lemUOB22Kl1K1
zhm+JzDyGXYzmS9zYrHf5i47JJ72YyGzHbvR3xdq7qsaVQBw+Zijoo2rEr0f5/PKryTdA95g/Z/m
grfVqPVZjrF6OFXPSpNHBrA/PIA9saRI8VZ4QfZ3jvCIbCu6KiqJX9ANtJ/Am6IwPQOKVPfHG1vg
sPVJLvtLxBIItUElHEkiEMThGUuE4RZVw+UCIbzx7GFyN5ZDh5P7f7n0irVIsgH5wka7nsjjvFY4
9iZX+/qG3/Uk9C9hWq5x0GoJ/JhoXU16wTO1RtvwonWCkS3zYNJ4wSFNY0Kw4tlceJkaGfolnDRU
4CWa1ACHVkqL8yqPE7enFfLrS3CuOJtoiUO426kTeaIkRVvaq9/vaHXLPA2d622RHrJEFabZtYiG
OCl8QCc/J/FTEO4m1Es8+6AW50hD6NOoG2sH9D/KpwtyyF25n5tZIKsEdU5PAO4Jv4pIS877FSUr
jjRr2Rt0ubCdVR1wKVi/JdB9fvDA7thm/vpARMeL6Z6EmV4Oiufsr4AgOZ6WLvBwAckI9L2wxRCV
kGtDopTUvzTx0x0LU0A9UdOYD8Zj29XEZK9mX6qrnRaYu1WTbC2zRWKl4at1ZkJhzJ9p42ktPeLV
d7Q3faBK4Ug5CJjaKP+z5HYMDSRD3wl9btpalIciwmhu3tfAAlQrnAYpwbUTtnXNbvFBMFCICOG6
y+EWOVwenicuD5m50XRM79zUVFVtHT6wbOWYDMjA9/7p0m0h9/uBV/IPtgUM+2Ys05qQVIHO5csc
jvQMU6bDR+60H26ihBHDTrCjLpO+i+nDoZk0NFW+ayPvpRuJtNLCuYzOCuYT4uC1YgXgyeHO5deq
0mmY/UuvLsVXqTqhpk3s7jnjhHSHGpW33ZDwjZ08Mv8EfLA7COXks3/eviSVND12eMbOsUK9wG6d
v5EVFrgYp1jSPYQiWwMy2WnLzDCHj+8t/tLP2eLiUksXavpH0Kbr6Jhc0+YAdXCpKuwqnQhznd7z
KcqGuZDmQUA09WOzG/wCXjRDCmnIgpYHP8m9RlJbtVWQtaZ1jntrDEiUG1OA5NTNb6zAyfi4lr8/
Cm7doJ/urNnRKXUbfRPeq3fmagPKVqOheNn0gllJ7G5lum6J9ec8gtjXL9JaWWaaKus3YYo0/y+G
GFHKf2KffKBbyCsKdpb0q2iKA5/2mJVV01zAUnxUS7hLVcF8RIZmZaewupjjZGyVHvwmK21MT/wb
c+4FtTD389ibVcWa+Lv68w1t1VQElKufl9iES77u1Fcr1p6sk/M6yGO9mNigyhfIMEG43ysxn7EY
1UR4RPSeO+WflfNo4WDIXEMYks3mvpYv56dtXE1PPDN0Qt7X/9JY8dExQlJqgKh74H/S5d3u0Cf4
+PnmuwbHiHFH4M9HcBaJofLcfCtjOImVZ5D59tCAX3dFQtiFSx9HVs2cYWlMvRPwOYUSDc+63AhG
SjYT2WTtkcl+WProk1uqSsnDmTvIaNfPI533BdvEQfoX96kKVotZ+M/5sXZ8eByuYCzfNOggvemA
YpDhzYtbNh+l2Lnekd5ppoU6w46Wy1ty2Mhs9wIVj2Vnkm+q6UlMdQ9TTMcmd/04n6ctI23TWOaH
LW1CxDxFinGIkfG+V4FznZvxbfbVWvs4MBnt3CbEd878pmSyawWLmbep6mpLThErnablJly+N/cv
3yjOx7FdTfNu95SHwG41xFX0lUtSgVbg00ikzFaHsCpNNioJ3Z2irCMIgDS67RAkplvJoNAjZo+b
kQe+GeBLOQRWcjcPVFs+yXZE7aa1666KfV3Hq7TB0vsmIGoKB1xfqUgeec6TM5iKO5rFnnnGzLPH
c7retR06d8OZkMNi6WLRPXQHQ6mWJcRD9iAi55mNfM8KvTqT0m8rj3fDh3F/vDeEmXmzlXIY4TYy
I8Yxnt3u1Chqr3lzXYCMjFULPPOprziRS+nvosyRS2Rk8FVydvBYlmpQqTBY4eAf6us3VcJYqNSF
58g90UzGwVR11HfbmKTbJIy/WKv1UEojt+S2gj7z68sKh35GMj3cJ9oiKXTLN3LyyvfcREQVwm2J
sqCEMLmcQm4PcSyRhgGrZ4PpTJW/bg+FcGLFMlEha4ODaYwtTnyl3siVOIi93JI1ZAuEMTXPIm60
ndYKWzw2DDDVBv+s6obsYyi2RaqN78DkAbrgo3p8ey77upmCNIve8yhuhoeo6R4mG2OdAIpYmCUl
SNrWxej9+z8rryfHwNZ7ocEF7wxZNkWHMwvVyquPUsILU73pkuQlwxpSdvFJNYQ+3EJ/qk/A9GRj
zv/+/YFyPpUi+aeUqClBL7/Ik788KeXgqcMQ+x29f0O5Qt5TgXo4fGLTF2/KnNpdVhsqnjmELXyL
kdPglvrSASOTIx719w7IhNWck+16icRlR2SRROM5FFQizenSnvwJx215iGKgmK5CNJovmoCYMTlH
gTcpJDUQ5rQSahN7gnAehTgO7aZUP5VXawyvdLO8gYbXOOCMWdKdonh6fXrWfhkTlnpCHVx9mWpR
fmxEHSFGP1kildLzPl7xxJfedcI+/5tEqTsih1nYYWsda2N1vO+fNMBirCmcnO+fLpIL3GWoxBmN
rmtcpdYHnQn3YI2iaKTUTMqZ5trGZZo58tsPxYZV6YGkmjZ2wWhwRScuMEobVvJpXxHv3zPYGO5+
D8RYF6mRvc0j1v7/ngO4mYB6pAYjhCmi//cdsVF3zcbmFCPAxmfrWWtTUWIGshKH5d2J6anmfM3x
htDKaRp8l9xNu8W18JF4Op5LhqKPEIGrXwFdWGwq0z4fS0q3faRZc/HqB7ZFyMuQViIXj8gm6r+T
8vqjRGLYj/vJu2HqQNf4fNFPkCXuTc+brnMdA2EMsAPS1ehU4cQEt5taGs5Nx0lZJTSnBxgOJ7Sr
mh6M/rC+QWbfrEK0WupEGuy0r5sfMBl4fPAu+ab1NSJhzrl4SVoSYh1i0ruCldQo2xaMWNr6dLcC
KKuLKrT1MfUe7/r2TpyQkLGZ1G+dQyjU0WdBDb8P8qHJlnK0/A3x3Dta3meFBMEaE1LJE/DqVRU5
3I3Y2umnWtLqJpT4MNI5adz0ereBN6zvMXl5DRQKM9+4AbV2VqKPHfQQPib6qV6g3dWoh/2tcSqB
dj54F2rHc8XJZIWbLU+ujp9Ezt8VIG16r6toxkVhHWidrOjCNx1ky0Odtr8O06r6nqpJ/zPHrk2N
brlDAS5MbiAE0b+5sHU8nqGSX4dbqapT6Pisa5Q7leuRtqCXO6hWWm0MWBj3tA5o3Itr2ssjCTiK
K6z/SLKP+49EK6fg2wNYyWGuvBjyX9E1A2bs1d0HCr8oIUvUVNycXMS9nhN7By2f5KlFlO4vWbph
mtZIHStEsOpJT2TnaAGs8OGiXjBhHsZlp8T1/TY2o/ACY8sFjoKMmR7nNWNyBZNnEoWkLLX9q5Gq
hFOtyqnzUsEEqbFIJvAaWrUrqfX0JQnO3ox6UP6FaRJO8PyIV5IoZwDY2ZG9E8DgMLePDwysLWPo
6ed0DTeMa65OY6X/+ghPFiWX7S7/aDPqrRttsIrITYu3qgTSdo60ybh0vS8a7SaoDWquaIIvwIk+
3JIezaXblEX1qp6ZZABpT4pAV7RKRVs2vQVtI6voHdNHdgpWf5dgxQs385HvFy0GhbyJLrSUC284
8M30mbAJXa0DvK5PJyixpicXjw06gIpFASkraDsMYtX7qP4S4LTI2VjAbRp3hZCxV7VOfLzI2aO3
4xakDsnN1sL8elADfFTrMuB4rSARsqh4qGqHOupN2VIo2EoSNxWl0fVSOmXLvR8jvNoi1rMToAmL
6WtNYU7PLN0g+WTbn8uu5VhsXOk1uubpUjirHzQ/sCMnJZeqP9E1wRNk/LWxZZL9bZC0C89R0a74
SM70hdhYf+bOm2+rIpke1cUqkqPP1iOu3NTmghI4fawKUGH/nHhCv/7Jh9fBfRHVc1AP5y36QeCn
xJ3wskAokmkGsdRejCF7eUMj3dEPfMx9byopMKnwFCMlikABdLegr9mSwvl8ptF3fZynVOeWXBhp
3tAWKWdJx5+XqlmHpkV7cuWqVFPvgpmoLos+/LrEpHKwNBAmtriMzcS2a/5MBJfFB/hSIQrCsXDe
/LKtc49CeUjq/psABtQQ0ZMp3DgMW23fxvUTkDHGorpGkpnpNLmsptA0CUOCYitallRH6BtiA3jI
4oY2CmmuvbYQRdbQW+n3cBt6wsipG+jdLdonkQNDwXnjGYp2b0ay1YAHueoJ8kvSp3exosMX38YD
DTyjEXivEQ2wDKUBtVVF9X38zIjWLfeSOywUwM6ZOnHdhSStc34dkyv2AlZrL7KgiLmDmWELpMfW
HXuI9d35gdyqyqAx7SxpzlArFcg5KVo62rK0wmtF2S184BbZY6aJOuPqh/kPjFCGQaGwPvDjYU3+
Fxx814+8qfXWrJYDGv8U/e7odIMqFM1mBGbblVrlwXFQx+Y04qlpWcR3Uj5FSJIc5Fnq5S93EFE1
DafFJG5sEHT/Ws3EGrUoBLCiuONz77DYTafqiZ7Akpeh2vPY7b7RiDEa+YtZQQpD++cWSiBNsPEk
UW4HPg4csRLfa9TMMuQ8SESM8lZJ8scT/6zliZ+XYGHr8CiUkd2w6jYn7qKkfRGDU2jDHGwMMJtm
yGRf5Yh7bpmp3a+56GURMQvlGKHiQE/yAFO7pqnKiDw+LDaHw+//oiVnkajHu8wfBQcJtBLTFc9r
rpA+xNLeSrTOQaSGrQUVA60dEtxJIb+QBfRhaaDCYLY3yVwm2eM7WIiVDwq5AIeJNpGnGTe4/0ht
J/FBsOo+On+aisgw3Z1jripFrXcvXHpEQdE6YaYCliYfxo9O8YI0qTtxCScu5luiSN55xK8iJWOx
94nKM/8nu3YdzhQvz7r/EBNLPkc2ipG3IgVpdhhEbnZ5xviHB/l+Lyhwy6iR/I0DDdCgXqjramxT
7O2d9x9kl3jxWeCnBiphKP/2y4NsfkVCq8N0ch7WM9K/LvUumXqlpkn3MN96KgWv7/A8P6+H2QQ2
lH7xEzrS7ED/dwdenzhWcXk+d4sbCA7emVPQhP9ormlOF+epjeVE9w4T5lljFoqTRXcUcDbEzYHc
KSD/Uy8SBxyS48uCeU8RsX5v75sAy4qiqWAX1yI7ZYfgXS8O2DoAUiV43LYKILfDF0bOe58KkF9V
bPTb4BGESOsdNRuYlkrZumu/AaMLHoWNlsuol/AIpzI53unOQmYme/9iumSD2ru/sxwGa56LYcb+
BmYAOeXV3PBADgqGFuufwsprQZedTCSc9G/2GcCAYMo+80VTlo7/r0iECi40Aw9thdfX8YsOLt/p
hKflfyTakO3hDa5oHDMQBwNT5MqNzS9pDIhBrYNdfltnHqLO7ArKgMno1y8TWoG2QupCW9xpjWAg
CtnXLEfthpbdAvum7guw6SOmtMA8jRlKj+fQ8/I3q+HzNIvddwvOg06+DhXiOYc2dYqypitm4+qK
Lk8+MvWTp1hCEFfqKpXk7i82q1tT6bFl4z0MLZVWi6XHDPMOmLmiJu7UoXxeCdPvET27LxhoYfYZ
9unhJG3ZJGf3rinXhJzqU7jbvJ1VWVQX4zzG6JNXe3fobk4dHuIdJoO67klnPH6H81zvHoOrlxzo
Z+svHV3EfkuJKe4+U5+XaadCKFafKUCW388stAsgGJ4yvB6//Tn5nYngoFxJpkgyAlNsISqZAaRz
OlyPE4qyn00L2/fHXqme6hle/QY/YwlOWkhPTCKbNIDty17MbkNxegv+B4yWm6j6Q+pDrSbWLq4s
zWNe0jCsXLTdQtxMbFEMnGLaEkMFQdEzx25KXfVPoSpb2X3D6xkWN+0qEJVwOMhMmpxZKKV7BgJN
7zScvXnnXl25SDsTQt/6U6PDz1qkEMg1AdAr0ta5ESYH7Us2OE2/iTOSvTzP/Qq4mRH7BX7WIcOz
eDw9k8Jee1i1WpeIgKPWdEPOtimfZNJde7THy++4BS8Vdv3TblBUnH5ArY/d2F/FT7fnH1md86GL
kLIqFj5jTN+zqZ1qKWa8pVR42hnfjUDPBrV1OTS2tT1bfIovH7ctrvhYlbnXcoBtKjklcqKE7jij
FRxTDhnrZGPin/fqPLmn5wzeR8xrfDJRHE+ofxXxFmUgnqHkSJnp5eJUVetk+knEDPevGITMeIpI
5Jtrv1inBCsCmFnUsZyqF3VSO9Zgxp7mDXFWY7W5YvL+OiHq91ZuTk9oa6N/g/9rubv5u3FycGBT
T6bO9elZPylQP++HLwgC01y2nEUiHfJj3CPheY+bYh7uUKX15jWW574F4jBFFrsts7UsNzl3ny4V
0jfYIdH0rfPXLosQOhILaQ4U/p6EjO7LhzGFaXOOqtS0xotOT1IYp462lZowJ1pHW1SEi2XHJTbr
PLv5LKvHoxFUGo9nobJuD1rSZMvqmc32TRRrqsYAt2ivFK0XnJHcJGXghCjeOtxhoWVAzUYp9Kqq
SOBBLa87XEaKwSFWUpSXEUduev8n7kgQ3LJLE6tsIR8aTnnMfFXp7cO8FrbZiFlvZvXxL1SHDPE9
zxaPR2rBx9HXwuRw38NL0h/Pss8U5e7MyI+cIyl028BEBIcvBA6cGS/AseH7pu90WyfQwo1e0+4V
WdGo3eYgD6vcLBGy/NfKCDZQ5M+m3v+EG6MNG8s+mrvXC6cZPk1ahhh+fbQ6yLsJ1aT+dl6D425m
/PS5RUJmmbOBUXE5O3dUA8ZGz5TlxKKH6ZwwoyheRNzEzgfzQH7/fPPWGhJ8FAV/jpGbxmuTYRMn
TVbDRb6xBeEYx19kdHI3ucB7fc8HWf2U1eTxRtGmWHkgoktg7sbZ9f+aWqA8OseVKP12RMRAp45x
ivrqO5rNfQVN3NUm75eJniIUBgRNFZsLmcsFHVozujTR9z8xxgMV2Ao3CxKysFYq8V1VzG8HgeIM
F235jcthWMudbPAJQrlTE/iYibbcZDF4wOZUiSb+T98JtkjPBuTOdROE7xoXxNCJ7EGqHOM6S8aa
lxGm9PihOX8fDRCla8gcYR/ASnKZSVnZuXl4/LRcm4G8GdD8/i7CnBLGTHf+CSOzur57sWgrlFzc
tIVY4IXHWYtyK3UKPnFNcqFxKK2qo/SWjYCMMHkzKfKLPJg8GoloFjKFYaQbGJ91oHRKEvirK1b2
Te4a524y9hQ4Gujcfxr2Ka2U0CbNeUvrEqPwM+PpazQY2dfDjyqbliDH71F4Z9NLbBsFXtu5kIoJ
3GHFt6wjuH5jpWcqfEStmNWmHvT0Uml24P6+nIJX+gwSRjaxgnRcIufWhKstL+ZenTRlBUbb0RNr
etHjqryF6jgIEm+u5SV8L6kgUrSJBO1Fuf511AnZdRIg68d75Q6t9LP/x3XIsc5P4ssaTtobDnBq
mz08LRwPBM+yIzYOvABVQI8Pq4+NTESsr5jRkyVKU1tk3RsjSuHmYqC2clTy/AcwRybOwHwmJwbr
YLXw+v4HFxLOJnehQU1fyo7gzFeMaR18pXtJMmAcq5rs39asoRAAgwi0lWGGcoiTuTw3wzNI+qIu
BpDfgqgWn9vvgFQTkE/2TxmCdy3l2cPO7VL4UlF93w5Ufko0eEhWjndqV0FnV2QlPUxS8GARSVbS
w1K9CTPqjVRn0Rjz9o0lnGVF2mll6FKcTGLfMcywHz94o/Q6XY8/2hkcvsBw/ZISgTe5b/YGqxKs
ZmDPiHfWojesMZ0GQP9QTidBLvwz68xT5t8goLrtVLU2AmdaaPyop4msGMYgBwxIeLJ36CDlPeNJ
jwv3INuvLC4autvualIszZDbeAuha7sYSpjS+jaKnWt+qkrqbGNe8Pivgi/JQtTTTyH499274XsM
u8v/klf9CiXkdIiLpAwGl0v5xeeOy2kKWkjeYgJQ7rSdlQoDR6+jw6paaaxjkNfvPNItO0NFfhpz
whHZAyDwScSydFWB98lLPDluHhAnDkV3yugKlHgC9PYP1wzuaNIiMk+7wXrNz1D55B290ZJ6fHZU
An0aXLnDDHbwc/JWlnLBEKo8iYdOwKwEcPasempalPuA4py9Gyv8mZWBQUET4uFtkGku/18y1TVJ
Zmq7GFNtW0UdfAOrjpOKTI65XxTPTu35CltqfvCkn6r2cefXmDfzIrvsH7yBjs5111nM4BDEbQiI
Or7I1hJ3fvkHXm/kmwc1/AKUPspF+utMh/XV7TksY0ELfL4YuYqGEFCWvFJG7Y3pSXwcPmtJl/zU
YJB7RqJi6KOE7LWfVv9maKLSXNGuWTUMgz918HbNSyP+SxSEIohbw/mx+ANzYqiVPZIdW90JYkDF
rK3/B/3+58rczzv1T90XQgkw/57MeU0x2zdWVd36Z73r7Vq69ZdXmzXknAoNw4sv/2ft4PjUHP5e
u+Si0DTT+EVwWT94kZ9pZhz31QYGnwtTrZqWZgYW/zaRrrrO9OSDsPqOhEsP1VqY/e+XG/xAZAJR
mKmT2Kcb1RYBCzZnN/UcApMOc70XCWyq4M+dqfKD2Tt6TWvEYNHlgFF1YzAu/mCeATCr2rqTQSTm
WPwZ1jpLCEtSoBcNuQoPCzQOdEgY+r7Zq06Bd6jo6stJ99GITEv9VtOi2lbjFoLvX6DcIUHx9CaV
mio7OlPUneYB/HRUGDHo9e0NOhfIyjgKWG8FTKwfFIx7BVCtpp7kBYplOXfieeQzsMVU7DSWWOgH
V4Bw62UHA8/T6ppYS1IWFz9e/xAcsNWY/vV4nEMRDfJ16d3/RDHWtYkpOijjV8GVogz7ciXaLut1
Jk+PrF1NH5eN0jYzhW2N5oGVfWLhVzMteGe3hx63TJ7PGDhBzRqjXgH51cMMCGBjNBkhZN2ZXb2D
GUDvnSlBcQzX2iR7zOgsqUbT9YDfD5XIM24YXOq68YPm1YoFu3lZyEx7OwpwkJodf3zMdjDLdIfl
H1KM0svfyrIJfaG2rd6BYX5QkzYVSb2+Ia/ZzuhxMuS86cnEZh2Q9zaj0ZOOOb+u1caEx6lUWGY7
hLRfEneYH6kkyDb7oI9KtfGxF/T+dyHaVNxAkE91dizKuROlogW7JIcCMqeM/3a0QviqUYLZdPBn
53fp3KZ0MyBM2TOjBH3ZRl2KH+1+KSILs0jRn8DbGyWFolv+HulbbPKqHCsadvSv6bC9SVjeu7qX
bHqzG+YVoGUdJ7DGpZjw6+PoHW2xJFfupM5e9+++g5DHtXdLIAetlQZMbXllkAoM0DPLgJilZ10W
MsqlGT9rL+Q/9JTj3REN2vgJymLdxq9UNSnLdeqgArbj2XFMwXkZL+wGLeKRgAWwpzq5lBgF77wJ
Bfh3gFPN99O643nM4YMgguzpwQC73FSTXwNJDK6qgzKu8XrQd0y7IAVQhzrtlvjmiCO672E9jdpC
Nvn7iO0MshJv30DgGQBgQFaBTWo/rwCPvXpsFW6pnTvekzn0HZ2xWS3fAsUkxF+zzaBbegTBfb1A
cvuzspq+jrcCQPkQK7g8ODZtmC7Yvx0WRj13reMZNHiWUuEN6ySXdPyCEomkBCHGp24p9d9vITfI
eurPgPW2KHz27rG7FKRELcxIVJENI0ZBPAQRrbRs19a7APpNulUE222gZWnrHL8RW937VErhhi/2
znF4NZULQUmfD+8HIAatP/fjzbt+G4n5cx0oUesqnoSc7ntukTOknukH/gS4tDiU57SCnRGNskNu
iwgWap5UPLKDm0flMCXbtpXcCEdkU27NDnqTlxjJjIZXPcLALs3MEFLljVpZjCQohmHAo8pQBvUQ
v0kxJM2O6syHrw435htSaDL0wEh99uLs2Rjk/evAfgbshRdJFAW/FfwWj+Yw7MLxCqN/U+3V5XGw
9u/NUCsdePT7C44fVBJ64cfj5kdUNw912biSRNQsJI6kyM/fvIcVl4gu/bAt+sTywAIdLxYWzv/5
/1JkrYUKx15aFb6Bw48uI5Cq2HmRM+CjqQRZpycMu2yeDXVrbH69fRcE/KxydqG0enQA2m4EoCFs
tddoO2YUVJzFHOFJAcyuqYC175p1++ddQ+NdSwu7pw1tzlgMYNSFCd97dSROGEjSAse8Hvl2tWdJ
tjOcY/ZKnGT9G9spwGbam/ItZCvWwGIg1vzSd7/LO+ubPtExsVdo9p2q7lfid+C3fi+fpqoEsLkZ
098YyNONsUEZCAlfIXUNYNxGVOruLYu+EYgZgcfEwYZG7/dFMehuBLptuJXivgIGO4uxbrw9eIsN
2TpoCFVLq1To7TaKRL49IWs8fnb+y72pFVfDSVvrEiT9bj9m4AzAyPQC8/H3+IZEddpFPJU2NmUX
WWnPFG1Yo6Dktcf/9QSYpg+uLSwqSypcRApiZlgFiq5LdwdMRiH9MMOh01jvVGL9YvrsbxpfyIVi
H598OIxJe1q8iB+HeuN+pJ6hELxgQyx652MaT4oEDc0XyfIMq1hIS87xIWKZ1IUebN6cqdhox8J+
W8ZFJ6klrjLZpbsKYbF1Rq2bqvH6gfwggYzhe6reVJD3rnhPZ19HIJFQfdxLfil87rxNCqbsvEHU
A4r4MGKrXJLNo4YXEvrqvxV0yTRxuBB6UEIxupU0dbHy3Kocoa9EbkgV1gkFy9iaCEk1W3bT7fhl
1HN+2xksZwesR3JYwYUCAUXu1N/krQW+AblAsSw8pL/rudyvLu6X3r08a3QkC+hijh+fxUMvBgnn
0usKke+WG6ykU5yBBf3ZFbo8+/xk3IyK0TSpkEA243htJCaBNACcU4XAQFEpVJiozepnaw45JxkS
5jMmTMzeyCubdDtnhaehb8w8jVsa5Wi04ULdyfcr8ZJgBi9HWhEaBGIdY8QEtOKaz4Aak53nBP8u
bKgBLigSHDaOEb/W7tFzDPWmrkYr9WnchdA7/e1Ds2nhcTISCVYvs/ph26hGH1PSoWK3cLbOKWOB
3KJXGKjCpoYNBuYHlHY6CA721McDOuS3hn1EC1K5Op+34qvptKi2Vp4gj2dI4m1WFltpLLYfDF8v
UBjExXD3Z0IzzGXh5mLLBuMJacxld/GzpZU/Cwhpt5CSwGNj4fyTgwKSuOcLhF09Ki3BXNe+raG3
itCHs5s7ycXd21BsmkxDJm4l75VwL1d+Yhqiww+4JzhLnqR0X3dbZsQwnANcQLbp7VDMKptdZVaa
ic2HlEiept0Woq84uL5+nyccLDmxgBYzw/Q50siIpOTjG7O3uP71VT5UCW4zNKOgjMAkQDq8j4Qf
KS9i6bY00WRK+xcRyDJqGNnXAskLcovM7/vQC9wm4i58En9JgFqqYg5iL1HGbI+4cG6uR6NOQQUg
joB/90lgtlzr6xSv8b4bPg4H01CSfFmVYBbLjtDXIfRUj4VL9Xgigb1AhRz/sHOmSlMIl2YJDoQn
hbi8+8057wa9a5ZGw5iDPWFZ5/R2LEzbO3qI7xEe4nyNesq8glj91atKVBzpE85HEvA0k1irRzog
I3eKSEDidCOEWrA4peHW1MyZjPtbQT0yRRyx2VcY62eOm3FOM7WmgA0I0cz1RVvBYDOPh7Tmpn1R
oh10HanCZUrgzN9tPazxD62oBQ5yX0LEq1X1NIzXFL3c2hTzhCn/dl8DXadX3UiCFVhUeczCahOV
w+xflz7aw0P4AkWHupgUQoWbJC6/6tE/kF4PG7TiITxWYSzvVHBU96j95pe5RfuXSBONX/KwZKyx
BBLp0X/0SDRojumKQK158G8kgpqGqG+FnL/NM+FLzBiVB0oYdJ6fR/SOEmWzVnhxStBDhI6YkWDw
+YW+mCmQTjTOyQQOzuPLk2NLb+OPUqI0rgnvcMuQooT1cQ177TCFt+LRYo/dy88Csho85KwhVdt+
giTmy/78kXTvICt4x5t/riKVarRBn9+VDIOdrHdq4sLDAzx+oR+Co3YLQ/WJk75l9Y67ZUWYml/9
7gEVmy/pCZbvF6PimA2HBzeY7F6kkl6VIqkCUk0bRYG0e7G+pEca2L6tKed4XRI07aEmTlBX7R8k
cnAYkmP5RcSJXbzdgYQepreuWj2ZhSqIwZOTrueo0IsW8tCA7OOXX87SBqbdh2QJB4BvHvfTjIe5
AW6vTJnjQyDS8ZeS2AxwfMBDugTJLjtCCAcevhW7LsoyAlEZJYDzEbAtAlTRg5uEuvitEMQxazon
sRocV6d8trnFRrvwIabRYVloSER4Wn1v9T7bk237U/CPKkW8WrDZm0Pu2v9FAMKz3HNwMozMEfNV
UQRzcPvBkakk79WE7lwr26jB7bOYm+YGZ/4Hiy/UEWF7M94ueQBKj/+5MMHwQtzD/AKM8ftXlR8a
DsnSDX5kz7z0OmUSWNcKBZXyD1unYnDajBo/jZ32ltHmJ35wnOHpkgEds6XQFh6AV7Im8PVsAUJM
AmE/ltn69X6c66fLqfNlr5mPI5b7qlueXE9aExgVMC50jX9i2mNekSdo8n+EIj+inqwG1woFGnOL
xSV7HZSPqkQ+IQ3jkAkX245VWIN7YSx1xkuHU6pm5Yk7d+ROkG0mCAUA9gqMK0bMEORYcT6WLlLd
wW6xLfT5Iq1VPKQwIJObsG5j1o7Ts27LcdGB4ll+3bMU3SfQKhdKEj0fU/Q2mZWe7WNFUtnQT3jz
k4HoxV5guZZH4853Gk02Lv5tyAkAUUmcW8LF5VZvhC48wHI7Avt50KWu9yskZM1I2D+k+CGz+XnW
51Txx5xFlfrK+Gbqf3WAP6odEXVQ0aeUhqWJ3P8iP/vTBqAFtGjrU/0FTOyBdNXoTMRoN3vRHYnM
Zp4E9XX1w+lplMprr6dIRawoZC4YUfSUcKFA7I2EPyGfK/ONsMqPcP+ADa8+f410jP5yvOfqABYl
qg/YbEydFCLbBls0i1TWj3PuW5aebCwTRLdNAS9Pd44csQ27z3bGA+3Lez11Yksxt/0QFN1jTulV
NMnw9YKuymuOMb1xK5/V+MXQalFeP/BKamg4/aMBYrcP/SGWRJHVEHWK5DrJU6FD4bV4IUb73h3Z
ne4svzRTD4WjxT3l9yqRu5L7UsQhwrqU3CjG3CdD5wawycE+1mVDir9whEi0DMaWGw8fcs6m6v+q
ncvEr0C6YLlZdt5dKMdjIoAOXbpybgu14H7wbrAESkAKMzDYbS1zJ9rygdNCurmQ7XhEbbW7PSWl
IiIxlm1wqdPwjq5Dfl+p6tg+xTPZlhGQY1GHx7e8960IUndMvyViT9w7QPKWHVTzIp9k6krhpQSx
iDjg9pzAMKMz40Kd+HYrg0THL39EueejPLlSfFYid4V9E5mWg0gjrzf2Wkkp/aRAvpQheQGTn2mR
XsM1ERSWUc3gkX8gvRXkxeMVCdh7Yfx2csDx4B3l7NeJuo47hZAirRPwX2IDOLkqeUkx6mMtF6aJ
nMNcO1hBEA/2kJrLzYyvOtWHPko8n8R9/bD6Nm2OmOdGow9ffh+v1evpUTJ+QbQfUWaN5hI+ENF3
UyzLFaH7/oVi9oLJ2u5rDPEOWznhDWW9ZP3v9RyXDtTNBD9gbNDaJpT3NYZYzryhj8T+cMdgWYro
SX+6w/NxIc+nirKgZj73eetV1Kr6dkZQMqKIttJ1RaZcbiGU1t64ppwkaJ9HOUlN4OtUoruogVng
3sx/tiUfhzWM87lmh3i80KdYW4NpBlbRm+NKltGyMBOKymf7vrqqUjjs92FSANleNlLiILOQYUK8
PS6hTs1CDn07LjEwgbZHXFGJQg0etQynue82Qp+p+CJd6BeAwXMAqCweY5C+kT1cVliCz2tQllr7
XSG0YxmHC3UITPK2zCSaVsrOgtGCDljKahfRPRywrmpoyXZad1YfQExNXpPCJKNLLdwTU7RlZp08
0TCD04gvhyVXq56UJ77OcDdvyxpx9UfJxWDSs0WV2Z6fEA2COtKQrlWXvZWWIRtzUl1PQc6Q5H+f
FN1BI1spR1Di3JPXdul5dloKqict7L2in2QEIRy9GZtMN5ovgAzdFzfW6TSimK24REYMil5muW9O
hs27E4zRihE/Qtw9hskCbxMuJ/MKJxgObbd58nrW5L1AjdYGUReP/dkhD/+tzlL0X0hctrPwYjF2
/SLkiPVZY4xzfWtT6sZpjzhKPLqS74jWW+pYUsnhEQlJU4y3v2hk9emqk737o2JowY935wm/rrJh
9gz4V//WVXFG/eI9/jeiVFmRFzWVz6sMLYJo4asFsw95sF51heZYXtLx0Q9+sj6oIidbiHe7Alv+
DMMnlJUoWhw5s88ZYZTmxBibIMikGGZV91ZotTg/0sCIAkXTazROiD787PUZXjt+tnIL8jhstZr8
d40FTsxUJ3dQnL2TibtWChie280f9M6PdSZLk7Md1P/1SE8E/A9Ist6ZwdDXhiV8AUblzEIjDUij
sUXze6maiq0qbiHNHvPaSdwNuHmBrpuySUoBLWILDddrB414Cg535fz22qge6gMkyt4o+G92/P87
iqhFYC5KSvcTk5XIST4k+N6o4L2lmJ8RUcVdhVFubaO2ToCX7mlRPkWsFVHgPcalJ5125zH3FQNZ
JPN2jKY5yyj5X+TLO92VOXu1D3zpFpTbdLkeckhyVE0uSPHDGY0aGAHv0QnbJhDF4FXeVhgJNhST
YwkMi3nt6qowIJg35p553cXcgZ09CF9kFCYG2tXga8EsmPfywrarxmhibmKo9TwVTmQFX7RLUwcq
XU6cP24w82krOe2eaNUK4jZrXWAxIHl0skLFJff7NAdGjtb+7qvRhQfx2NeACJba/uXOsU4+7hZ+
OznrH1UnsURjsq1Ve0jR7dWEnSLKjB4TjAlKAW5H+AFKo36M+S0TDqQzkIfWc0Qw04OGgPoMSi2R
WzKTF0QMkbj72aaRU0WPj7x/N+xDp0WsZV1/rbUQHP6Dl0gvbXs6gZvXcIjTf49Z6kB4mIGZl0uH
xZRsvhixovakAe8+1nXIWWMqwywoOhdttYvtc4L72orqxn6ghC7mOeyYYKAFB5PTVrqe6rH9bu7e
fFUILXKOlxtzrvKPidXFChKRWZEHmGvcVTB8Yd2k0sH5EgxwEigigZyaT9B6hPcK0y+XFC1BpT+f
HUf3n+TXYUGgCjQ0jGCgeCuekGrkx9KhCEqOvy3sIQmVxZjk9v02AlFRRmdboS4K5Zz3ybw0Unuz
wpx5Oli0GAMD94lAs+3WmCPmZthczeqCOqJYedW6eBfQNZpF5whD3nAvYBz+wGzIQOm/0dOIrqtp
9k0muXkw61YGgwCAf9YZxVmbKqroz3Hi6C44H13OYzXY1h2oQ2yE8z7xiWx2tTTIwxmUPBESRdxK
goNd5FSlioq250gUKG/Fbo077BW5wglj0Y5M4I6S8CMI/oaKaYlNEt2kuLPPKYXAHyf/WATh4VMo
jOWgRWVDb8gGr2pGZ+vu60d4MkzsvqkXNFFJE+qnr8bzw3Faa4/kUU2EzFDkH7wVRSXamUoD2jQ1
qS8iWCKgBSIn6DkyuKpO1Wsia9o1TINIK4HbSV3hlFPUTfkWSsRhOOh6lm2XCYdMoL1ibGaq0vum
94mguv/PgeZKsbvxy59qSCAWdQh00GWu16RCsuwnwtfm2gePd7fC03KMLQt5McWKDkWDJwEDSPBN
ye9djFVx821qeOVELWeg7r+eEYm3uTPNsH9KJdapHRoOar74B6/qpTc67Ygpu7W4tPsZgdC8ePLh
aJ28/9dkVpSCOMPhplJ1l1pdPeF7B15BcI+weaHBiurkz2R7TO67lXfeaQqOo4IxhQjE6tp9Tnmt
Be+Ag0KgmFUjffcVx4LAc09v4uk0P9d9veC/3xRPqKcSyvmI2K8lua9HDE0HLFQcGDuzo2VfnAeI
i3pK6yOSp2fgZgQViK4DMbd9t5Ng+24+zsAMJUGA5mayXvuZsqccDO80ckSiwEqj963qijRuwc7T
RP+lcKaz2L1bECz/QIGyjmc4Ngx6985yU9DgwDzvJ+zkO5hmPJ+CqUMwSqOl6DYNz3DIp1Sfq2Lc
4nGkuKoKh89oof2Q15UhTvDy1EHY/ziiOzhFWOC8Cbuld907ayxBIhRF7MH0BFkb375F1EntvhgJ
A6zQRRxIT+9AQh+IMc3wmtpgF9R1Vp2D41Tw91xTRpYnZQ8+aPjTzz9qcRM1Qj2kRxX1gp2jeIt+
qS9XOWUucoTPRFt2mbfHn4Jr7bq+qiNM6X2/rZ2x7IMh9TobfXYancFNRSW8yrw1qRHivv/LfnkL
TUYa6BkA5n50z2SBi4TtIKqxMi8CFYrTrmuxLP16KxLFFfqmH7ngvqCZI4K/eLetx0nnCAXRxu9N
jhd+URFL9NiCGXaeYFOGZ3Ls71Og6v7Jr/jAADIiFiWSUE4haRWT/c/PEOvVoVNZRUEYlwjB7XRb
kJPBoWSarWwg9zFlfbTq+804hcqJsxzR03Y9vIbN2uvKBITGK3zoBbkq5/BlMHkrW2StS4YLCb/h
A+xynsC1adOQ6WtoRHKDKN6BWYIk7Y9OcZt6qMHvkEZ/zpgGi3P5x1imcujg0VoSOQxQj14s5kqN
gDtTirs2tjw5B6xznikZNQ8rd0/vTbZXWxuv44YbL6GLHt2L9QjKvB/vBOvt59Nx67LA9xZGpcA7
2kwkpO6V3ej5X7I3nJGDAZopH1XxDP3x+M6NQDZcQSyeLhVAGsRSUAM+ZSnCZmauFUJds50xDgXG
fVblnnuoKQ4CfdlD6I3e8xFLwGFoFhBTLyYz6yMhyYz7k99ULFNfj2vmf+KFviS+PiW0sFCkeP4l
w0DCmOtcoCiHMQdxgEylGAV72V2Rz4SWApPl2951kHEC+6cgcAzUtbnS7JH1ViorICL/W+YsFBOy
/TD0iASPqao1FWtjVYLZnGAHnK5eygOsajd2g1UGVMUUBCWZQQhacxQElvVd1mDp2BI4qhq34IGw
ji5dSdwt3l8HFMWfCJ7mlZIGKMpUceSr0ESIsyPA7xVcTJvZ8XfbIzGoKsouL1f/VfgQRUQuVSWB
Z7KCAr0xlucTeuhj4kAuURnf0EKMhoNAd4S0FtJheRCMO4KRvrNlVta8KawBMvTnKQBoaFnxTFE2
hJBvaPOEy+GAUTrmzLUYwSdA122mQqYuijjDdgLnooaMupPArXs+X1jpw5yMuUv2LcIj1sA7zhg5
XmXyOY4pGu2Qw4TNWjjTtPf+W2sQ9NJnWhp5Pqa9pYG25XnIbfld16bHEeey3Wo6uEKv5psCx600
bdg0aZpNXbzbe+EQ7TPa3croAlvMsYcnx62FA6ZybrqfP3kKFnsrw9JaH2v73b+ymVfZSrolDG+P
04yclJun5iHCGst71VBgZvvoytk4sX6L7XI7bkbViFpoTdt1oiQTslu18Kpd4L8g9sY6EM4trrg4
3uY2/nDKpaJksYrCVYXJntkwfs18HNyfG9dYms4d3COeotVAkzF0Xwh3HOpwNhk9LONu7yMWZtHp
VssdnCosdyY9isdSnzY4W7KgzyUbKI+nAKUNf6QXC+mhfTmfM8k9CYFKqsbg8wWYtKUpHgGI8tJ8
90mhsnRS3jxJA819rvcwzgBZ3wySyYmcqonU1b+qcYSvtzdmNmawpBNzaTg18sJCvlx7TBsJLQdX
zn/sWNbzFutUATK74ikcBpDeXCp0WiDk+aXjTdrCJbZw1+06cPFjKDB97WE4HqYdigmiWSyh6faO
1xVrvO2o4f55Z81iO2Uf2cWV0ssTJnUBA3DxSLqnz4F0ewz6Ai8b2v2tY13wpSd8vav/8yjhhVop
PisWYH1Z/Shw4EfuvMEyOOiglSyU69b10zAh2GsLZvHez9e7CSEboS2loRcbVXbOnJT8LolDGDjV
aHwnMnVxpv0q2/RzZLUSK1AUjqGoEyp2/qNYCDjYTgjB0NK3eekrAE+uQT7iUEQKz5kgkOJShhel
TX/5RrcPmjj7CzeGM+2BNWK3sQ96+YADh1PaaTnJyOdY5NQ8Nz1ufC7rjQ/KmXbeRHWX8U0phtFA
0Q7GomfMTKNiaJCJTGdKv0y5WguMJj9eQmoMSoeD/P1r+IQhh9Q33N2xak9Mr/IUp0tJy/C4sPQf
NLymykwrbwZqBg5xlwojZ/0TnCTCGM2/4zDa8SNh5mn+hhQl6h8g15FmmwuITGVtcZOk0AxfauK2
RLu5AgHrqFCTN1qHy3OpOaOK6PbFxbp07LCj6Vh53cp3dmzWgSR/qSNLX9mZ3JSqN8fJFabs3fhb
3KGN3LPg3lm1SPmcD8H3y6H1qjqcMhrw4zfXjlEYGH9DZgLgo5zUHpzLVMn5Ys3sYRARt6NFNVZ6
n9h/9GY1v1s9cFeaSWrl99YWnQ95WAM4P2t0SjPZoGgljL8Jip7NtDUhrUc0NmCa38ktjZtlWwh9
lrf0s/ODSpmOcyUNyAy1hY7sTWOSVeO0uYFeLWUCKxyQvQNSxo6xVfvdZTRkE0DwjY+Csei4y6RI
jJxRU1e9i6XNOe8PXBPKytKZ0Nz2itA+SKHaG5hDQrEYdTuheA72R5/nIh3W95vLlKZ3IsJ9+Wwd
Eth6Cnhuah4d04xRS0D9tF5vujFQrlDS9K9EdnZtJpQEPmwbHu0X0YMrQn4xdDRZPtGbUPv3Q5VD
G7ReJlDK5bbapjb3GqX3Ryq3rWpOT4qCgqKPolI34a1pNT7fua5lPApTYAL9Mcv5vIAHW2i8vgV6
uZPOjwkHJ4HgTChuCLHp5kRtG6JQxQX/47ZdH1jACFIVKFQC8MjijogUI8uCK4b6GVCGVc6/om9l
hgZaCLtgXjoZ1wR0BZNh0780PNlxKSxI5r+btjNGbhmz5J3syaSygW8FZXuI/kYaJQ3z7e0WRPSu
4WFeuIKjNZSQld97KLbYaLdbfeGQ0BYHu5TARip33vav+1kg11fkllM4hh00EgDOfPwWYbBvLpGJ
ek8r/3ffXukggW8QrwQiVa/DNLkxf8WdsF7mBv4xRKJ1CDC+DNbkfejAxRjcMhGBB9t70hZyCwUI
i5GeGKmHqV14i9oLyiVdq8NdqdaKnWs0zdOkj7TSIwTdiyZPiSQ2Lj0DHq2O0E8XRQjDT6yK1/wM
3+ADO0jL0eqH8BO2jnpnchjX17P0qxY9ZbJOc5hjkJ+6enHu3VtuOYqseJzCYqONNGHEncSAfYHz
rsrk0hP0B8GMqaj+qp53M1j4Q7CyPIYJmbWvbhVbdCaSAOm9xtLBC8lQ6aQHat93f7SpzIPs7pVB
c3IJ2AtBMzPZ2Mbw/ufOmKmX01baFlwd/A+8UKiH/KJPFClLJY/Uc1GMpwFEGjA5F8ds9zly1NNh
dISquC3AVc6kAP6JOL8wM0EyyQybrNmSJYqirCOxnPzqNW24kVjACQdl7Lcuc7GO5ciCrk63wIME
hvy7vtvp2GAVdSHkCoWriHxaiMYdlfiqDCR+2fFyp/Wh4SxuODjApFCaLyL4a+2Fl+9EZ78poZEm
7hZPbvJnMe8fBLjEsJZebY8vZ8DKL7duA/bgsLvcbpH0Ly3Ele6Z+6XSirE56I3wyocL72gEtRBb
tuz3nrKLmDHdZ6am1F8HrchuRj1pB1D2B5BhcuO7TRoMODzoZ2pPEUQJRIGmmuSVUX/U4/qldKXC
BHJrE+ycdTf672u6IMO65InKi3lxEpYRUVJFyr9yzWGspcghedhGjdRCHAHg3hCUu5VpguaTQXb0
1DkgywKzVt+e+xzn4YPtNfak9wv5GDQOxgmFSVzuGpb8H8NLi4ZZeYXlcB0zCnrpAJ+0E0jggSwW
Ux7WWVyCeS2sn1LLLsS/PKRo2AxNqoHo0o/0chJo0D+hdtFLKBe748oubSmyU52mNs/c2TfWvCg+
VNfWinGa8+hUf+e9pDCtwvt0UyxKtf4Df7KnjKYp2fylA24S9hweTVPrkhy9bkm8afVWC05biSWU
D9ffhervZkuoyXKEk444giJrUuQtIRPyDbRjMy/nWVeRJVRnTdpeomyOLr5TIEwq/kSJ4NHO3yac
X8JAiHX79kLxWbVc5d7/Cpnap3y/qg45cce5xMWFyHL4D0KYAFXsRd8pCZgEe78bXffO+qHRA/zi
7Yjb8tcYnEKwc63+VEtMLbFR49CjYnrag4O+LJ09dQytgpOR2dtXtL1IM5ZGuCsLzkDQtg5gaqUl
PhaeHxnnCyKvN58Bsg2uIZYzQJ4T6Sde/M52X3HnxIX/YyRbDcyJvzG6320KBvg7oesvESxRB2Lj
7kmhGpSIdSd8T06ZOQ2iqKFB5HbhC5cbxp6V2pnQkjwp/YLIuj+5IM0algYOMV+R/S0gPqomTJYC
6JfYQ3MUzzmBsI91MqPXE7EPu0HMn35h2TQlJpTORFoQeEJQKClrKF+mXtuPS7Qo5ZzhwbKMuH6u
3bYh2nFFAKF9Cg+kHVEJjsK4rlZKQzfYgCQYdF41EhWOtKVzzQn5ybThfCVGZS1IKttLSmuoOQGT
Y4aP3VCceB1gAjA3E5vQDpVr+vOTsVHN12h7EnVvvAPOhkl7I8WCE+Z2VBw35pln0XoVNXJM5qoL
/ouy9yKyDJ+Zc1rlNvHF140fWSVSbVqWpLa129TAUL1H4MvxafVnVEniFDO5EQF5YW/r5MLD/XOQ
TDh9PYcpYySZafL+jYurpCHH0KetKMGIiJI4zUoe6KT+PTgTnvH2OIDVpwyoaUTUWBDsJMBED7SQ
GhUsL65QFBF1qxEjgYV9rKbUq2tWA8KcItmB7pM0fLc82vF0WV5A9O2a3fouXcR1X5rUPFdr4xiu
u+zMdrPNOXJPw4whX1zfAcftU1G4WJJ/Fyrg+CRY4df4sN3vedwnIuENURgz/1btsiBqgxfj6WH1
YaUkaTsQu72IkFS3flarCWsKHZwwU+hvx+V+dr2bvmXRlZ41dnVfCD8a6PLoZ8jYwC0WguQBGFkP
Z7BalzU8N9Cf4MesARX/8ERfaKipOdbIz8+83GgYkQs/X5kEC7YZSvrlT29L8IPOP5elEjuP4K0z
OhdZhAnwh2eU7Cy08bSGVl91iTBMf76EQYk8HC5ysEFDFMey+GFqZmzuHZUpR9Mq/E/4K8DjOS/E
Z7nmKLfYMn2suDRnci/QDC3isl7IoQfLL9Y8njDcGdK6Aje7x9l8Lip6oBlH3ZWJnaBlHAOjHY+u
xJ/D77LJDZjj2/HvjE7c+MHrHECAFZTjS39N0HMvSgPhvnXF/2CMuL+m0wBxR9j0yAUcv4yx0EEX
WyO4W0xOAfowjD+COikbUtMeHQM4Lzd6OuSSNHQutSt/hdyEyHUEuJK/sMUAaPQgiAyFRGB/6KeQ
TcXabp5J6v1ah1xHiR6HmpcStyZsm4s7WD2+qCiAPF6fqP7CsPqNOUPNf8aTBscDso7D0cpio9MW
beirjD+reF86WXkIQL4G6h494yl+FtQjDKsuKqBVO/egpCdp5Nd6szfUj5xpGmWL5fUO+iGsqm4w
/TBcPcli06B3jw3n0thVzAYpZ7YSHE/4WNw2F4v0bWW6Li2CNmNWkyO3+gYXfKQWnET3U/mTaadT
7JbBIaPKkhuJJOylECOWTvG1sGtPEmrzcxy8TnMEIUdVJuuWgyc87fBp6sHHd+gdA4tQVla8zTap
qBAIN3DbjYeQrf8TdPxgqX4Xl3ssPRpvZouY0p+JtRudXS+g22DAeSe0F57gZAT6azvjsnJLpHrd
J5E7DIt4pF2uICgSa3F7g7O2OaHR11d4g2c9d8QRFLmbSJ0sILxP+aeIwZldNUYCjr85olM3idqM
4Wg3v6zmYxTuUxP+MQWmEVY1rKFCfu6MPiVS0MHJMsD4yFC+N/THXighwH9rPdf8Au5iJdhQBh7A
uRQ/icYfvfz+MyZ8WNw3c/9u4aqOz5k/bJerIiCFtr5f68ve0Vb9CvuUv68kHPTs3bUCn5mu6Gu4
+9LaT7i5+KoYs475xScGDr9lwtAJKitOOc0uHeU0moy27UiBi1/lS0Yq2EwRVRpxvujStZJ0znGj
zp5DXIle3NfjOmyhEXHC+U4W3OjdSkPnYpiB6JQjXgsBqy9U4b4zCLyg5DGNlzGIfacrbiSRZTZm
0vNKqj96nHpJQCQh6Lpc+HhHQ2QXuSxzXqCsjmZG/Tn5OPUjA7N9KaSzt3J3X0Hqn/u+1egn8ymH
H2lYV8n1Gipf2tLbBo40g3IDl7nAJsY5zQYwYGfUHMfhyMblVU2Tb3l3OiQwSwnfT0YbRRxoYrAx
HsW6qaM6yUtUZUgtu/qa3ijPaVEb+0A76l3FyHcbhX550/6NjqLKk2puxoTeR0wlmOqPOqj5r86f
PEMyhD8dJsj4OXSup1cYj4NfqmqiLjelTDWmW11USNZyGak8s017eXUj/u7s+dZuoL1oKbWrRnqy
bcf9Fe+1xrT4l7ot8zn2KHtOc14kxZg/RfABhnx7gb9Z4UsAjoNBgVboi1USZgZp1Oyx5swn0+vY
fJpDMZUHNtvCkl8T5uCw2obKaE8/UP7PZLzNtm5NnqDMA6lcw+hC/o63QXeovVz01AKgFTDUllsb
I8TaZotmF1d1hSznhwJGleoCEQqoirxaNfC3hkWqehRGtU2l5a039SSS/kLbTO6NZtkqaN49036a
jo/rpFqOXyeSeP/2W/ID7spcnn1rwdvUytED9paumbflHLt6zjgMcR/9dCvwQfS4zRJhP6Pzwjf9
rfzR0KyVJz0wNf2XFiAXkkZWbAFI3x5WnhzvRrq+MA19YzbK+Hy8phwbfFsTt/QBlIBxngjmT63b
aX0UjDHjl2fd3HZVag3I8WeKpP7GDrOMmoNlRfuAsVhRUtd9XZzgrbopQV/ouUYz9JbrlujMV9jF
frX0I5S0DUOdww2yoB6OUowYMwJHRM3hX0smpEiSLb5kku4sw/oFXF2MNWJp3eVSiyx3j2KcXlav
Vj2bNhK90+r5Q1wzI2GoPy4B/PgogT5Zdw+fVseHxxgtBv7z5lfa89ZB0gA0BBJ1ggxtMX4Qm46W
qNvqWSpPzl6eLHwrkGi/ZiV/Yh3tcSRYlwM/Slh+lDyLA+mK/1aE1jqOclp9XAINuMLg7QvpMita
rs6Lb8wzDzoxl5DZvY1i41okFiI03OiSQBtEnpdQkH33HQqmpNWEZnleSKMVEXSCqjYRqEr1bWm9
CKc9aJxz4s09ZGElaR3wF2eN80Q9B5ZGK8l48tVbVmgHNjyslUV+9gEN34i6WZUWDu2ON+5j+JZG
DLdpR1UvSRX8f0AX5qcOMu6+y8iHgrmtORBzd23SdW/pNeQm8waRNYcXmuuJ54JHzAs2Qf3ivvG0
rKsYL4GZ160duFeKFOdGnqKy/Y+6iK9poMkRC1y6g5A6uU+j1YohNR04+HKNYYK528ul9nutQR2a
/Nqg5W3Dc0kv5aTsJ2JbfNO/hIW7UUQymRVB7+Fhk9JgPwlrVGxT8NbvctPpJVfObhTXS4aMLvXG
QSQcrEYnZCvT8vBAV76ylOM6S5bDGOM4HfQxarz5NXthvx1mBnoJmIZsMt00uabv3tLfX+2L1Wlk
VyZDyZiEegUU3HUn+sI9TMdGrqo8vlulTIdN57M+2nDH5VDJQ+Q+1G1Anp2oBAGe8The96oFgUoS
iy/AjxoXs/OktXq5NRzrISpaq8Pe1hTrzYwywk5gUJPjppJtEy9vtfkmS4mfa4VcbUtl6wbSDQH/
yM9cQR+AYN8J1jepkFB68C9mwYJ8rrbjd+F8ujen/DGCVEiAgMpf5oD5XpQbAuF7b1fp1GxMTgSr
qOsELgkRC7I1r8J3IqEloXOdc5y2KxY4gek8Qxop7vk4WRruCVSWL32vPC5+V2f+ugJUZB8xQ0oG
xYsasLBCKaob2N6d482yb7EM/YVXmIzwik2JArMr7RCv01DCraEbPXY7/S2lf29TdChQdOb3NbDk
BcoQH33j2gz8vJo4mAchro0NIgLbLnemH5IVyOplg9rttKkIlAAGS88ppCMT4TAQLOBD9xyAHrb2
aiLsb+81HQ0qY5gIFDkpFDzW5UpT1jcP6RxdLmtx7rsZSM77x6+Ao4zrgO3hmuQViNb8Z1rUK26Y
jB9hKN+9GH9rxaX6lDB1H+oCuifosCyu/neKYVw8yLE7saBlC0ndzEuYKEjrHGj1vX+bFZTAOUPp
e6DMpsYFPxY8r6qgRjhPWFq0pKwX9a/s1OKH04lVkVKHR2+Wg6L7m7LBPvoJs2sXtfcC8M3qjWPH
7pZe5B11DNQDdcIXMOJzrnIlueGHS52mFG3H/N1+tjAx75di4l9EhMPp7OQ1NmyoYos2ZOiSnXL1
SwbSbRSgw5O1wyKHVezdBlK7zYmhP4PKeUNM/lTGTr7rWR7EJC+ZhyowogD6TpVGCpgLq5yqgGXA
HaUvpmVyqk54OCSjvwJImyQqDd4QkiKHhqjamcgz8mClfI2/RbP+jVpFw1CVyBEgC9VQ0n9zVnfT
QOLUZnQ/Yt9S6N88EVbsZ6eZn5AkXA5Ay5/THyE7rKA0sGXS1NyARH9GJcGdAUGiWqAt+46Gtpum
Sk0eCbndK5fyY7qYPqF1yNV5lrpuvBq75pHbi7lFCZR7LTEDqH80MUHuuLdHU20g7baAYO3HGa5t
sYd9Olf8Xk3D+05g0hHxMHnUj2BkRLTVKiOzud5Y3m20lVTskj/H3Tej0a/rrWV9u7mHAvHAJ8Hc
2Y5GMnOk7mbcRe8xQXuWmLJ1yuE6fUsbKG8XnOLYKya8eqyfr2XuSw/5jOkNS4geQcn1nEUTMbVI
qLNi5zzoagyjZbmsYz29OALc+N4Rw38DVqCjTref1ginVuvMU51FKLaSs3o+IamS1a0NclPrQWLQ
qdxPFgI6Vk0+CNtkOnbbjWP/fRxTa3Ccsyw63q2evKcbVKJZ1wasH/F829NdXmkV+I3A75wN8BIA
wYdLqFDwTyNdySM2fbjPSaoeXpvuzUJye9AbXMtgq1+hha3UJ+PX56rsh36dcGybw6shn3aLViSi
X1TIsl5QGiu24ZA1NJX/1hxaLuSW26s9P8k6VkJori2o5JJpOzkZKzcKJDzbmsVTzr+EDVnUtwfa
BciesdeL2XO2fxeN+/b7X7q0wfYJTizoiG6N/8OduRBLjNpxnb58/14Yaw1zWgbJhWTUu9X8e/pk
AG9TigoqukdyGnvVVMsIVHt/SZ1p0MfLTPsjEPYsCTSBwlICDbiEnbT7NFCbept4q5ECoZcfvIgN
pn8ODaCOjao4HKQnr11TeE8kdNccLacbvHfnQLn1dLjfUyYM3beO4y6dw9il0MmrjvpQw8Y6Bdo2
D4QCDWCrZlqqPY03cBDTw9DaxBw+c9IrJOdNnUDkYpq1hnKsHxzWDsIliD2/J7sAeS24VB/1+KrH
dZuafAy3K/fC+jokBKlXdrRdRZAzliIcZSL28IiOMF2yGZYtyrGQbixPRoJ9rYVqO5+pm3WmhzDY
j7isTgOzya33I5eNIM3ZLSDDCvehU/YSpatYKjg/LN1KE6T/P+MU6pZfTdazvqVWkJ/JN387bsdK
uxK/Y4YWEHlzs2dvolFL08GJiR9n1HsmMQWpdMyMPXOXbyvhn6b7NGiLMY83j3UxvDtz0XrMJIcI
D4Crn+VAwuB7CkHvS+mAr7jx6tjz0bmcCFKeFmaPBbH15EvjRFtwdNDs0TM4gfd+NIRX5McDgHXP
4gjhvEv1nJ4pN1UGEKBjb77wxWcSzlGKuBY3VQPU7BSltl5XEPIrUV3HWmeDVt7YhsDzN+vYzdMw
4T86oUj1IP2SaaL0ZTVQlSTRmdFfF2DsYMtO2begeXKymC79n40Yz8KX1XJblW95ZTrOnET1KQzT
5FywNe3U/4QgW6CTn2eZpgQAMC24haIr7CXEc0OxmxHpZxipcRQaWQPiuRmzNOkxSTDUusAY9wAF
moV/SlpMmUP9LUyzYkHs5aTnQ3CKm1h+chTdBiYUxlreA6Sn6p0wlUMjmjEMYC1gLkBB+1b79Ssq
DNamqTfIYNkdTgARGVYpqmPUcym+zCbevQ5ezsbPKM56V/r+meh5+Zsq0UsMcEIImG8rLdOA3+pz
6KuiYJXTr8IydKMp0ldKtnIuXXkWyVLI9tZymWlxWdwj5lTrS2IDTsSkTPQyTWM88FrPeRV1yjk/
BzzI+Vb+neu8yRUCJDE5yZvjbE09ckAT5UN3tNxhJBxJFuxEq7lZSy6JVdHnsqPWSkWnMyuXzKQj
po1Z35ZGNckfUx2uYdrrku0ov4jAe/xpKFh9Csvyqnp57jxHH2lIzKaZIvWUvuvsJAGOvAdfc9lA
RdJ+uEeybc3wWAO8TOj2hkR8Utl4OjB4M1bG5oIJ0s5uqXIHG8ZKEpx3xHdmBZUJ6VD4HNO3Mawr
t9HSxPA9beue01a4OB05QykAJ1D0HIz1vVYwvhn1gBVx/HDg3EDpATkBZ8GxMtrP+TNr9hYtr6qp
m0BbH4pr9YSEweFQFc7A9w14aNejbLSFaYQwg3UFWG9ac2HslOeSsqSEqcW5tkevC/yZvm1oQa7b
/Jm43bEAfQtJk6iTSd2eMxUela72Naa/YnRBsOq+jaApxSQPWfkTpvRAzURFo6cnI2G7G82J9PpB
zGcf+r0sc6AlHQ19jfZz/RlwNOWRrtUaf2S7Rh3godsTU1Ljk/RYsPO9RUa2cUGEAQB3/nyN15R2
JGWdmNNPij2kLvbNB4QrhY0KfGPNwz7/KzHLdVd1QbhgqIQuWYfx5SyCE7Yaw+zmRGsTOtUzWJHz
nyEwPZutcNSx4huDL8ZdylK6I2aCf4Jd2AGzbcA/bhDv0J+0U+Ry60d/RL34UpMlj8MB9B/1tUhm
Y8vIFyNuP5//OynfhhiyxU6M09Qb9u58jsVl8F6UNqzRcuTQdwl7PdztkWGkCV5459SQf26rk7Vd
rVg/mDp9Vln+54PKnqz+A0RTv1AHA6n0pM2my+lAxRLyw7+tTsaTwlBJETY3tYzTsRHL/7bicVD6
8+SfFxfw1iBKA701mK88jX9kMu5L4z3bjEH7ut8hWnfbbrSrPAwJhRqNuMvoBi/QCVCGzF7PuZ+N
y2Qpp2DmcKbiazHcauNfJakf5Wc+pgaEIni2/t8CiHBrtRT93jckt0i/aX/rQtys42o++8E/wg7J
RIgf+opgc36oWzc1o6/jDva17yCTJ7kMlvSAYeQjH9OdzqUsaA7Ks6nIuAj/mFHjBaRC7qIQsKgH
skpwjmfUp3opwbba1PHuBwt8oCCj2cRQpM/VM0qzU1DasoF6mK3TCVabqJMt9U44NtFSIWPacZow
lRMRWEKkHALVG9S1efi/ijOmMODGZq98YUXNRIpL0grIEWFnnAKZqnyC+A9uHByUHulqjCm2Bvgr
U+eig02jIQ8S3lP0EEVAZiJCdor5g8yOjNVulcn32X1lJSGz+ugwKRZW7RjJMvuK3NTYmxAwBGxK
o5X7b/347Wd8e39whTpGHP07mh2Mt2Apy1y9JnGDOyhMMsXEaNfc9paWmKQG2Im9DpAz5AKrD4Rt
lsKXeXP4Xri7dDI30Sl+ILBLsRaA5X9cdxQnsy2ANnZzi0K7DoxyqN/VPL3nJyTKR3k8igZyxia9
A7kFt3pFBYnsLa9u82O68TsLXCVBJSi+e2XowXenBiFd/G7GuuzfF08vF2iPeFfcQqj3jjNMX7TT
Kwwv1Jumhs8/4bEqkN+ZHd8vMDq9sa7CLlJ2czarPBZNAQPaTfOxnlx1yza488bTiAVjSVkvSIaE
AxIRho32LciAXwKiudadbb13LipPEMbRPqRODRA4WauFacNqBkhfaoFIK+Jss+XkIJJFOK/t/R+M
xB0A22fOUgUkjQocg60/dejDxiGdYKhP3F/ga2drfW8giomOovu2MxOWD2Ql4l9B4Zt7Soy4uv2j
/Ku3ul3maqUNwWh+4+ULXhJy47nMRKxMQkTpvwDA1/Xo4BSv8Rs2c7V3VU6bBaboJcAMnezG8zUh
SdzntgRr8spnUAsCA7Iu8Ia6isONjiLkv43HcAz8b9Z77WeejKZym7aMpVXK3HKRkF1Vz13RpdFp
dgzdDPXPB+lhcsQ9a3Hley+6K8B7ybJTVJxCxb9T1NtjPHzPLfCtwYE8lVjC27z6Y9YiQM/e9R/s
E/XsHVRG93luAFwUtlELYUkZ1yZVjk/pDM6g1ryuH/2Dul5TMwpBX7loL7W25K52PD5E+K/aWQDs
EmgASOnqjWGFVd4VGbUK9oJW02dQVGIVVBnYLCOX1jzjisSfTourYL+/A2SyLFfhHDMkPxTQrTNl
5jQhAKug6ea+JVDk+c4mpU1C7gOX1s47PCZaTXZ5YvFJjXUTHs1/qsFKopJuf4PRYFdsHQtvcqF4
fUoqKEnr4vvK7EYmC/S9g/vli1uNIetBLgXVHdGIW8mhDGaIJwQeiOl6y1NGUzDmxKIcKbnE18iz
pex4ogME0GUGwNxqb48KoJnF2vDztJVZ7QB6ElkGO4YdjIEdY5fhzcQaAz10Joe/NDsDmvbpLz/U
mTw2datJFuddK7u++qKAA/RS0nQbgoj6cVBSr9rR0lh9iWXglsVFjaq7gJHb0zqn4fhNjkOszJMQ
30dPdo9ubJjHr1mQ2VIdvlI6BzTJkhOWRN1dE2k0+aNOn+3mPk46ZePn4QYlxywJehaBFLsJG3hE
AQLAPJmV71myeTmpdaWGiSd+lZghV/JDgui+4d002pY0/7EJ1TQmCegpOzFLhejPxjsdKZB68b1R
KWcBKFBiiGJdjXM2gZZGJsTL3s5aP0jLn7L0ktKt17YWzsJRBxZ/WI6rsWGgkghDonCmnSJUPPJE
qBUTpStqsHJS73faQwHC25tPAP5JJOUykJ2EDtTlgh9bC/a2LaFxOBbQvYh5pLMqsCn8/me8ruKb
h7+/cd+nVxfXTGbXE8gAjpjybDMJxXVaK3/mi9DDIE2sccWr2mnEpv2+NuFKX7rQRIbjP7LtypSn
potyx2cyG7+4Q6OwD19VcuhZJmRJw/2LvVVN7VLdTLmZfRLrxCz2iwzTQqd1VRA5fumGybcDppXj
E6H4vuL5RqC+CuKUAV5S6sa88K0rbBc8X+5XqV9MGlNbmpy4JhkCOIjWDbohG/uvrJ1heJYezFqd
CpJtZcmXuppUwR7XSbAnhXW0KPhahLIPkHMK/JoxQCPYjo612BcZX9tF+/qlRz5j6M/++pMZxpAE
W2Ayyz3wsagUjnSEpt1PD0DIsjEeomyQshT3WF9UNKqV12m14lbrbnbHsEE+xtQ4+GtDkOAIjamP
iEznziH0lViEH+5CyER9+omthACSCr+3xfoHwEB+KCx69Zhe9BTYU2NxhoSJBfcxMudyqTW84ajT
FvBYNCIdFMjy7xGUDAnNQXrWXsJUA2RmpoZJioCtDkQ7Wd6tKsFuoPsQadwR6i8FDSJbqokJCNKG
ti4OZ8HSW4PBDg99Wu3DBOyWs4eI6LAnY0ZzSnQk4CEwy1Akvz3OmWzLCmYsnLUclkDjZC5xxHXz
MAAUyI3TWwYyXbhYIioPqUL5rlc1pchT239W7FIvX64erqQaiAeQWX0cYA9TTLZWJFYqc1HQ6x4T
cFhvLcuLC84p7VtHN7Kt8oP9U5A/6f/jIbMnGmCKOXPcPMRqhxy7vL5A2VnyQXtd/P3a0EECrrxA
Gk7UqGroQnkF5Sf/dl3PvHpbi4nb2aZindLwWN4ehzPlRqGwKMYgkyC3r4AlOnmLzGaDrac89Xkz
gFyuHQCJnJuYxWyqhjP86k0uxfn2JSgwM0yyYIeVVcfQbHbMdel2FKdaRr6hU4ieVPKHV23grJCA
6NqW6lcWn1IvfTfjsICZczVCJCqCJMMkwO9hb4RBj6B+UrQglytKg/xVVmdgBxRb0UjAwDu57nf8
Zu8CSwj0FLhGMwLzJoapeaYkaqCD3bI+US5GKnDOCBq+IRL0e6BiXTmPzjjwi2Ncj+laXYhDcHEN
pjseJYNYVjPVSxvyc6JCzYYkwVJgvlFrbPwY3fGchAeDKG3ao9AWin5ZK8u3cVcBjrxXhkVkAqsV
lA/WJ7TKDaMPT6rzz87Q3jr6koJ3Q9GvRMDUDPiNaI8z1eUbu5bEi2EYW59zErGd7hOJPNN9QsGy
xhhbsGKr1icuiw3shw84CFlIa/M7AsJNsp+Dg62GS73beKSi6vi8SFEm02/3+3HU5cxHGRJmN7Zw
HiuZasw/MTQgkP+XqBiSpiUeOMrNnBvDATDOkJGeVWUf+iaBBs9/9boGtzuYSvA351Cdgh6C8sZw
s4PtPj1/9YNOYOuaIOTtuGOiBCutUNQ3s3il8bgsZMkP//Aun37/a7xw7UFy/W3teVCQEm/t1pUS
7JLns7Ys4r5KpQI4Q1oxEJWEBtNP/yOviR/TjZWzEZUBLrkoUm1HHGnvtdAUEwtNOgCJEu4wRyoU
4YpMyew+mwSB21ai2jO2ca6f8rjiv8aiBYzjJAw19vdUGHLSe14zNeMURn4rZernH8YZhHVrqoLc
xMdwj8V3LQa14X/A6VQ9hpXm0orZ3cTkWxFeSg0sLwWC66U6E9L6Qhk9O0GlSTnkadkjP7RjE93S
QG5mtFoldGibNYCatamaxMo5zJFqP0plnWaniSr10giKfP6+AOOLcarZ/q04b7BBNrrr3yq6Sndj
VBzd0AHvhlKEvXWPYdGo2K3yroUrygPo7av7cd2u/bSbGcRPWoxQo29WxRTf1vnauGF2VHvOMcwt
jAsCzrqS08N93RXlEoCF0fwG7GngIfyEOP57w5jLXmNJSG12enU3YpFXUnu71dRshXeLUIdOZT7g
o40U74TUqidm5wZeIxBdcLltAwb98vgFkcsDDGk2+BORUjo0+c1xNcovVS34L608fxjhjMB+XzHk
t1VTeeK8gJIbafFx+WhdGSmRv8ITCTiitSdJ8Lc1cknkyK3Wee8EJmj2J2tVJiZngrUtNdYsQlwQ
3MxpQZGRVHDx1TAAD3Kij6t3IkfHgb7AgCGv0KE1MmZT8FhaOzNe4YF5irF7i9fduA71Dh5rEPvN
YjNIyHR6zhAOCxuXBmghLKU/94jeCKlTwF+6iIGeeCtloGh/3agXrYOPZpKAFgJIJ5/gGtypngGi
zR7cNQzEz/N3eusra0u9cmTh1niq/1P4gVuD3TwtakYaAm80f/2VLFZnPkj5naNgOsTZFPuIN8Lx
rTe4S80qNPzxOUdkRlr4WCMil9iK3DRMcU38hL/ILJL1ClCFvXrVVtSJOfIff6F2XtKsuY/Kh2DQ
jPA73r239KsqMoNXaye53bDzlPaUFoQahVDp0cjSUo7QJvQnIS3vj/fxzfCD/ZiQREjjbMYAkETR
kTpLdADCFhyv/Y2Lhqfbr7MLZsiRnTEMmI0RGWtVsgl1j68EW+zWCyZeplU+92+zwuDubIeINR9x
+6eTlfNdTuMY/SVsA9qGEOQ72PXBOobrXmW5dEkTeFjLDrEVzy1EthSvNQGGHsqboukQL8aXTZQx
kPdFPpCggk8QoebocZqPqfbAcP7EUQTqB1b2jrr04B0RvI4p/uHTzEg6Q+NC3NcktPxZGCwiXcBH
jub1P+ThXrVwFu7V+HyI8KJAG3hUKTyXGduMNGwSkmui9N5OfPnOp+YcF+RQr7hCdOz2s8DYpe+j
7VlODdFTCe+sEaMZdQOK5f+CeSx/NyJOKkn/1K/p7C7v26Or+gK573oGglb227t0xNL1tOsemX5f
Vm6tFpx1+rnbu7iM165xF33cJ9yMNzxAXxS0KZnja1V48WQmzYNApgwa89kWlxyyG2xUTKqdh7UF
imDm6dhyNvOL0B6jaP+UkUmRH0+h3oniyIsoTcRW+I5dW4m3nFHJy23Ir0lgZsx5hs5pyX0j6nUf
XDUVcAosRjqMvTZAU8/cIyDqvZpx4rGifursIT6qYTwMn7eV53bri2kfGwyoWOzEHjZLQgVlUL32
A+ojgJlQuHJlzYWHZq4sqxpqxRj6yXxEyvcQjbgCdrpAO+96oPPBKNNEfrJYFmRtMtAmAlV6y+Fw
ZzTANSJIDSAdVAmZ0y+Qeh9sLOAl5LFLpC4n146tU1yfGydFRpYhxRR+FEKSnfI51rSH3xrXMWI8
+zL93KX5HlhXceUsJwW5Ur1wYOaY4Z0jn0gp39gPVtikGRGyoGKjOHGCSwqEBNOvI0BLIIDaSyv3
mFNeWLr2+GAe119vx6h0sGX2Fc1vGwwKiZSgwRj6oLm/VTSxn0/YPyvbnN+5vCekIDDBS9wuTj60
NvLwtmYE0gUDdhbhV6lS0h5H+A1CVX4StpV9UsPgZOPEJRqFE3FQWXcNMTv1Rm8T/CTTYUV31MoU
FJCnc5RVHnf2kCfbupqC6i5KXVon6MGUlqPULcb/A67vmTL9DGVvj8rC6tAIqX3eyu3HaD4Y2Uty
ZIJ006lIDoUjPbtalM7V8IUCPvJRpYEk6jcuatC6JIFNrlbDoGoLvOC0ITSE7FQTCC3E6LF6U6yN
N6Vj/qDm9JnDVswF/nn9cUuycXCdPzxBWLO/dXE31MCiYkCcTdWWXkuMx6n9CYQHgcNJvpdFsTXd
5CwdSUzI7pfoe299X9isPKBf5KB05D8rga04Ug+lFkUjPTaUaxHNNiYxWNXI28BBgTIQgAmTqRcX
tFHBfED0qImZC/4y0q8Y4mq9+dcpBmGPAO8Lc5EEcccsUyWUKcnL8mOZzVAKce1UtPShbta6uglK
QkYLa1bi972zF29O7Etwp5zieKmesaGPUnOPOwmahl9UMxF0PZ/82y7MzoJGdEjG95rPLHF1x2X2
lqVhnBdJVtMgliTxbyqYCuc2a3XSCFT5Arz3D5MDyK98qme2bVmJPFEwaYnFn50VNrpcDuroOmZG
d6hpQsqZb1lkluHeL2Ru2AFUWgNYIVFt5XHMlC+ek4JKNnxGWdW0LV7dX9T+idSy5B/CxzL7pGa7
OlDOuw7axC7s6Y2PGH+mHLkJ1IRMx5Rv33JEN/+Mk+M+cEkMdhZ4FbtApH/Jmb3Ca05+BwIcqyYe
ItklQoyNA+loLu4+J02UI7Pmy7W9JTuxRxu8pr3bNg5YsqH01EXgygLjLb9UeN4dJI+v7Q+iDWuI
Uc+/FD89FwRRxXPmUC5RZww4TmlTJEuAr6vEX6Q5jMU/msdYjO7dhutLDxiuvxD7gkqV3yiJ517n
bpUPrbD4OUuCH3NCpAezYvCLYxk9fjLC6WNrzFh45qX9NKwYFmrkRldwsfvQyO67ZYMjr4QthTUb
nrKBaOf144iN4zjIWt1Mg8RehpAG77iOrpnZSf6I/XRw1WlbL7M0d+m35bizX2qzzm2Sdy8b0B45
y8HdGEudOcxV0Mvo2mbkTZXHqt/ZH6/FR0eAvMtZTQssL1tYoJi08WP6h3WHZzf6VgGW1Qt0qsPv
kLKn6JyAPNsJdnMS3J4iJSjNDtsdPKZyfOm0jBXjTsJQpEG3M5TggVckSm71H8dix1FwWPoCJ0XR
VZOMasZXO+b4MwMnre0MNg5SvT+09/UOtghN4xi7tzpZPxCjB9p5F+EUl+CEjg2/wpxjBdfrWHXO
s6UgAmNg5AJd/YVH09CPMrjnJqkQLvStXE/0s12+JZzO2ExRrxm+7sU+iss16dbFRvkifaORbXDY
/G3mAu4Mg5X+uDWEFudSu8eCTgDfmy/AmAiGQJZtjlapKW1c+CjAKqtg0/6tJj3imuwTCG6p4kqX
+gN3/bkBD54NlWIHmkRzs7wKY2J9Pq6X4aeu35wy3B0jL3mQ+1Bt3xScpwNOQhJ76HKkkoWSeZDE
BxFxH6YnEanR5uRrdml8vMEFLMVHmVO2NU04AZwNvajwd9xDNmYiIbawa16u/AvoBQQkI0ewZ1aT
vOUehcgOSosmSGssgSZCGMgddFWgbAGltsvv/4wS2+gFoKDkn+g41QTNAJ/tsU80+8UtbZPUKHV0
yA/ymNp/x8JPykxlG0WOmHtCBuKCGH2aNXItZCQEQjA2iWwEX5//HKGAXuFSNNl6/zEHVFJkIpFh
O7ceLyAUKMWMYVkm5YW0vfPzIODG5Zd9a4SWOimm0+Zo8bDyPD4tXrYjNic6qq6vFC1h9h407Sgw
3JfyRzFL7FU4uf42sJaaSTVa6jU2LzLe4Ux89LfwtgaLU86BQ5xrG6Uzjf0dkhPA6+yt+B7LmmjI
ET324NsGD6F1NWpRgKZJwOdB9q4U9XGPgsUpLDV6UFTWqAvfhpJ43T0C2KJVCpfx38BlMCiNBpoy
lqK5zYuPU+gyVQCT8aCBDcj8xvqTv6qUNm4ghT0NHGNTUnB7X2LIds+JQdrVYJ80DGNEKbqkXndy
5jyjrvGdRIuhoOTt4t1HmVXw6UwYRu0Hcs3DSteex54i/plZR7ibbfBxDiYs/ARXSEQWgZi1RCHM
OEU9SPqvovsx/kqEr4EjD3SHYcj7kbFzlcLuBHMkaaeRxRhkE7yg270xMhpH0a+v+hpIwjzh0Ggl
pC2DfqcQLePMAEyfZsKDKFtoFrb95DX7AgqP5zcXeeZpjZQ6HhewafrFi+MQJMjkLSOdKF/7ICdG
m0IQa68GjUxfezGcxxZ7hdPUCtPIyN8KpHHhH1ltLZopFyMn5ByMiEPiiKnaYFudAqebYIGGRQS5
tANpMrWvML9pDf8zq93c8X5qa+myf6TSpsfZF7BIMxK1crZ25izyKBQOWVK9Xs/PPj+XzosAOa2+
OvDPo3cnJj+G3nfIbdy5WHL7YniB+jtP1eVMM2Y4yS2aksDqa7+SAQbDGd/E/JQPCM7BV5AzftvF
9dE2cCdPHtvTd5Ds5V2o1u8e7QoIO7g0LuJz/4PBDU4z/YKkBbM16aiCel94+aeS6tjsCGb8Qs4O
wrkwBwkwChUmlgfQO7La2uokEH/OGpj0uU0F70LHR9RHdwsnXQlukLy7sGsLYs8HKKX5DRHN9QfW
xm83dUID5RVsz4SbNCB4tlHo12BcQ0RpTyZRM94z6KTLmInNj3dcXuCpB+UUF4llkFPgigqMKhk5
pNbhw8x2NMfA811xV4nHP6tyWfaze9o5Jugff4MZ5Ul9d+Qd+22hoqC72C9hlg+HiuWZfihSNlso
lgXg4VZoMZZpzJpz5vk7+X+PpDJC7C6LdfdWzy9S1db4czpgzkgMH9u5bSHuMvuvzft2hJI3jSKi
Bu0A04D1s/FXHF10ZUmLIu6Or+RxPCcFEU03X7NBe4xXXZ9I1wm7nP4O1ISqPcZZnuL4ewE9yrfr
F06C1mnbZp+bjNUwwqKCoUOHni4f2kFbKxQYFQis8yCQS1Afr/+uaUB5j2IUzuumsNnqWz7nTwrU
JIAfRHJghVx9JcMOt8acQEmc2mzHd4ICfPcULNnDU73vkEl/zPqDMlBKHWN4NuQEPEET77B1pI5g
tMCdyyrQtUGsGIYixCp7fbbwvUkArgDhSfHYqaUKkVVG10oIhGhs8uirZz/WOxVMN1vTby21sc44
HXJ405F7sK9RfMINOX9FnNAbRPS4IPkNWU6SaoYi6/GhfVwgKqikOKjweGh5vplln/xy8R3EVuuN
PkLojcXj1goq9zGDSK/8WXcOCv7dZisSbwnSyBj8kJ9FBQ/myrC8V0GAu6fxlQrIiRrH1/IFnzZN
D2dmZRcdsi4p3xt7TMogCZvDi6MN6ucE/SAQRMV/Hpgqneqh+BoPUxgGJ1wZxlVBFEGbHT61hME4
C7w7O4d1RCEPpgs88y8X1yxfu31yiy9NFpLVIqExqohMFVZbe+VcrZkJcBxnFXMVrfsIFxMDWTgQ
yY6e3qr4EIxcvKwfnrRNbnCxzJEaZmMMLnUAUmcnt8uhnPVEhr167u9qRG7IB5SuSFeCuRxpuMZf
g/XVklrgCPA+tP7Bn9SdBZBJhdc3QCf99VyRq7fKCc/A7nAwkl2RxlgyS6ygvQSBBig1BECjbmbG
44psAbjipb0TtZB8zxDsJ6iN/r3zWWKel3a9irdg/sx+efpJktI1sihtVJ4KbPTpYpfZ3Zqk+a5o
zVj2mfe9qEDQ44u+YaaDdAA+M2HeFn5NwcSDve7MxkNsEEX+zjgXHYED+xVP1E5Hm7DHEXQ4huP5
jAVZZn8JA6QyW0HD4QZqY5qXbUd1txTbe6fvDONNKU/QRMqwwxSOCCbzFQqOof9w03UQhOya10/6
GhstM3UFkvXNbbGgk2k4OOjehOm8+WhsXEUJE8xxRHO43xHOE1M4jBSuS3+YPlfsslSyZKHl4hPK
3UuVlo5DqF6go9so5ApM1IbJTujOCd3oSJxvJy3/Grf87WVpg3h7SfRTjEu1a7zc8DauLUA6QswI
qYOPKUB0kOR0AXBs04AVUYTx3c89sY+yuh/oXqgpE9MWvun9JmkaQU+cRVSv6r7EqBjGxxXwHKgw
+JTIkvYp4uSNPf65FYPEonX85Ii/M0x913nEKHGbV2eObobROQmrI0eOhuU/GhU3eklGESNwQAG/
PtZ5QZJIUeEoOA4SfCoJAcXuQHPs4LnCerB3PCAGPaYrHxZv5RtBw5RJLEgaKQGs0YiUmfMBH5RW
GhgE1ttYgSBFw3bLXIP9kbyhDPWsVPOKKnnwd7JtouLEkLcqoeOayqiPJub2lg+/CHgsTfXaJ5Kf
2rWYQRUe0daobnWQyrf/3fPIKhnVGTxs/LcOkfbqslFCmwJ7Y7UEVei1edgk9wrUwp6YHfQ85ZMr
8ZwtvbqiPhrLr0PV90uFE2podWqANMR2zFe3nMAfmrZ1B4CBn9cSQ6+2xYfN5JeFENqnQgAs0Fwi
rLluQ1wD+lTLHoTTYuOHuZiYWcb6DRFUOaQOA5qBrKdr1kC74q8dZcPb9rqfoSMZr3M4ZwWQUbQl
ktjlgHhEytXuC6WqYRVlBj3iWSX+zUosKjXkTHKjiJtrD8DWF15tXSRBfV5LPkcR04oJOadm+DRm
dWojEOOAr3CRSEpp2m84xFT0onSI+cjbC8gd2kzBEnOvkGUkFnY3q4zCRyVYDp6ug+HBjNRXDlqC
r5qXwDHIoTgGCIc5GgCdRChIYuzdlhSy90v/qsW5+s9Xr2SDV+SAmUF2rZ6wDwiBFXR7MWcLuv/E
2/caGc6CfG6IIVZgVWoXCuDnZqShJMvX1/jRPGbhE1hlnOaJYNHBqcUKEQHFW/RPkswEjkmBY5Qb
5jSxlbkc7Cxs95zgWf8m3kTHXi3I/oqM0jmfJGEn9ndFUU+YszHM/5knAK483sRbmbXSUASJSlia
GGFh7j75spd2kAqWMFWFBlzLIKfsiDWcyPwOzQizOX259xmQFVeqXbZI2X6dWyMbwdRzsJTSJTY9
EHKaW9hTbJNbYRZu3MUxVs5yRkkiLAl9ZQ2jpOQdSvx9rI4/xwS+wlncVpWtc+mEABf+oTJRDupQ
S7WywLjmzyQDGS7TTkcFKu5cwfmupIZfby07nENhSRmBBpIvkGlGht/iFfaC7QJOJp53dQH9FY+y
WOe4cu2VueqI9oKFLmUCUIZ1G4b5VAL7Cmc49meAavkToybRiPbK9a/QIleo9uqsrLJJdzqBkD34
0KBr4xeWWaUjK3AQCXG4dmcWQQhzlBWXIbLjHnsk7a+odR26Vp5qbIq+d+cWjv9++J1c/t8DbihD
WFZjHKYdiPKXI6X5DKngxD9eCmttGdUcRCEpq7oDVBJaYvuFd1mxmMsiPQD5bAc0i+H5m+D8Wal9
PdWgY3Ui+NqISS2h4Lx1WEm9i4piSuejxGaS2QNjeBbheC9ydkQ7nZumbFEWpyiUXB5iw7sCSD9J
TRaLeDzWIU+8S1zQAUPDZxm2dYTZDWr8C+rhe/HvgVWu1yKjNdULOrtN2RMAKSUuRvGSt+ZP7ETS
3hzvnf0r35jR5hkTeCRh1b+32kcsC0CbCEIyysyOdArV0iDHKbdW1j5IumBcUTRkC7xBu58PTd/9
VxJZugHv61De5S78lGASiR77XUxmPCQN+GECHB2u+DAENrJZ0a0pydohfCnCF18OCQvJMR1DGHQ7
GElXKZZf5+uw5R8BLDIymYmw7obfgPMfDM4pzhCIcYtEh+xnHsI/RBtwWRl7gKgTwI312rgH2OsV
7tS72ukIoIjt8AGS/FOUfKTKXdUFS8n1YeFdhNtS7+bEBhUbGSSTjkbrv5hFUdZbmZIbARpLVzVr
2oF+RuQngPV50cXl31mQqMMPIGHDcD7uPY5L2nyemqS+VRasRn/jBJY1DXpQK3UX2RLl7z3oBux/
2H4yoUZhhERTIY7msjAU4a0NHLsfz/gLl6+5d5RamFmIAUCZVzSQlfV8CDES3GCrttrQnDNa477x
1LMZtZlcLTiRSvmulMVFsH4YXfi2odslULT3hOSFOid1M5KJTeE3OS2ronMgaHpNdLTEG+za/Jhb
ZIS5+03foWiLeZqlrBm5ZursrEg9e4x0GkPpFR7KbuXgme/u0BUVJKV0riaBTiiTnfeZ91cwBvX0
/1YkqOvAV+cwwsY/eOOeFMF3AED6RMvFMJe8HeQK3CB8CDRQd3t8YdNRbW9cR7RvFGlzr2Oo9m9b
TgdA1fcJj+ksQJ2+11pUpO57huLoR8q3moA8Alkn8GASoT/8t0/TpaYWC8shS+9MjJMxxf8fGUtq
OXVj2GVWheWwzyqFLeFP9a1vf5E7trlLUkd6I5jqa/SGMfzYTu+uTEPXRXwUQq1sRdU2cdiFv2zQ
cg5bHl3udENvJ/8La4zExzTtsTbHJpFtY3sPfZRV6klPgnGW5GAiiYkSfMpUE1K48z7TpQKg6nfn
i62EWj+p+kNgTeWoGPgYbkmymWjfgbJZyumq0hARQsicLZo1Oiaq32QzE8jSh3yQfHHw0LdRdpuV
nsE9z7UojKcpLIvoPyMT9IO1nWeB68xOwpfb0Ew1QxGvYUC6QjlPfpBE9d3J/qvcF86HRKrqtRhR
lN7ghxj7EyMRDILr95XQpCitWGZrUmRgFDOen0lBd9l7EsyOGY+4vU9OErzeqmq836Hqmj1Z3YLr
x9CqFO8sOPLDiQNYhxlXNrpZlTIAEEMe+HmtTY0AlZ9pnZjvxEmPhRsT6MHk/2lHr0fc+oOKmQhe
TSd4l0yJi0KcbaEm6YTSnKbEKJSV3poZwrI1AFNqTQAbsjXLUWHJQVJcVuEMGpPYDlF391E4xYJd
JuDbDaMsQwB0y8ZzpWZlsmdlNTUZeoc8pZ1tGs5bHzSFTGlVMDM8gUl5EyS6dCzUJ1MQSTu+mPjq
uJHmcA6RdTxDCE8SAqT4KOx61EeCCibCaCX3090QkBrBWKhOebBDDye5FYhhWvr4TBLlruXbL/H1
NfpcJtcn1spoAlNgtklAVDZ6YIr3UjxdapWHlT0L8nAKiXEMq7Yyb4qFwkQ1FdwvM56TyArVlDwy
KkHUZo4EcnD+L2HG38uSpzQUY0UYXmt+ukfe6hLwg5p6c8HNGzjT3tdeyM9MNTToYus89gvbb+Uj
RgBHbFOP1C5iT45cZ6rpNieXWppuI6425ZrqLF6iJZIK7xqJIuutChJKqNIrnxGSvYNAPD0O8GwW
IUDOzOyIX0tSeYyzbjox5onzJpbMpRzWfzFlGG7blXRFY35xu4dcjh4UmDzX3l6O72EhADFFGmKM
Dyv/hxMQ0XtnmHc2klFAMP7gy/greF92yu+PNzB1O1y3rlHcpdw7Cp2/CaPnpg8Cqkdlonsb/Uqc
six2uGanHi5VSeBbINeqrMh6h36OKQYJ1FCzth9nDXmD/KqyuPr1XzcPSWPkGsQJEapuC60GrQZF
sZTZtkdBpBAX17O/V3ntJsAhhcY1Xn9AoM+rvOjTVGWKhcNDincFnfmzfUeEpS9dCeRAXXJUWgXQ
oeZCb5L7/JFgybhkP87ZS2Koq92r5fzmX4BlbV1XVPryn0smI+nMCd8Vo1+XvMXVMYZ2/dApgGib
lvB5ZFBVO+P8dwdItuXc7HoNVXswVkZLyuslp2JglvYwaJ5It9mBQCnHMJScYmubEY0s2p/BOuSk
W7VM7WslynijfAXAjrh+fMmbg7jfGGocBNmDEoLiEvAEGSpw8vZRGeqlFBMcPwt2tN5yYQX6CGKM
blfqfbL3nFOF/HaDXjawmxYQlPxkydHDu1cWwAATTVwJdtTOWf8+Bb6TkO2kpe8gpxbIY1MnpoE4
+ybkHdab4dY7lAg7IoYt5nuDFRxoCeaa9pYIxcRPxHN829wP5AXiq1yvCWxrtBMKIVEN2nLywcp1
+f8nMPFltBr5E1F/sG57g2yHrDuYljE3yZL2yLOpxfENYYszryxZGvf1y8RiA7ng/bQCQmg2IQM7
pGexHFaO4m9M4J5PXvD8pcm89Y16hI+mF5ZPxVZin/03S54BxaBTBihfbOJRPbflOFaSK7zEHDsP
xadnPOYiu0T1Xgth8+h4JfksoeNkwfwahhJFad/mvYvj6JGEYZThNAbl/rfj9lE2J8EzGMIJoliK
jagVGKsIrFUQ4tRzwoH/nOTSm78o831/35Fnv9EbJGm+Rc1U8wVSzRbryrJZea+ddc6sL59vp48R
RCzY4dkBCU+fdcMPgxbdcQ2FSpobE8o8jrODLmf2Cof/2eimKwAnzwkjmq9JVJQ5DLLOKmOLTxux
8DgVGS5EzEur+t8y/ItbwBLDZQ8SOjhMIHkFpkaIbO2jlNbkWr1ge21eUa22quu//js+N/6IV4Nz
nkyjAAmxQe+DitX1ea/JcrLDpqgIc5IcgmhEJS8/uHEa2pub8l3eK/QkR31YrNRPADXdUyx2bJ72
sUhDV0SGZtjeNIPoC6W1rTbcoRZVtPlHrHPzNH/bO0umdJV6ih/ZGN75BI/ET+v9xz4zEkiOiEAh
Gz0JLvMXk+9M9qZ3OIZfDgxmapOSP7tK9hZLYoplz2tSRtFMXPcNorHwj34N4YNLqKe9iXlzo6qR
LVnxQDX/DstHKvgIC6d22IlRU4bKYFlBL/vmpb/WHZRfo2ZUw7mkhSjcBMMO8qsT7Gueh/Y3djsz
1cPiXa1Afl/JWfM4NGq3oir6aY4wPlP2TsGqLDJffwNozeV34SAE6PWRMagS5uMr9IWVD4hlMsTG
Wr+9YLtc0nr68vzencl5kdG7PEwYDBtytqf+dlX557sp79RWxJ3MLqm9bICA2+IkDpO+aJo08yrT
NopAv2kUXpuudI17ypmlzGtxnqY6lzDNoyScTGAgaHSAeX2106HSOlCYMmbzu+/18j1BJtdP5Qy1
OOYp8tfe/GibQuZ2xnGRwlzng1KxDaodHHIBqxEzAR7sHYwcJPWzlhu+Mbuxg4HfV2dR5+4MHANx
GTg3RPyPEG6l68Arc1J0VfHhBdmklHzm4a739zVaWJOqnb/X41d+yJJOUfV+UOYwcEcr5nBRdg/s
O9VQaty1mTVXuE1riiU5PTkrNTjEWAUqegSA4TqPKCud2fOREBKuScuKaThcZif5po2fbJzLMlK7
Omh/zyGVjj2FY9IZptUf9GXUV78QANlqYd5jxwm0wtwX+P+8ZU2u0iVASsKWBzKFckA6Q6U+9G1p
sm+GX1wh1xFEkVBIRIMWBwi61JQIbnqYiA60YKki/XbAINowIplwombE5mS0R9dCrPKegQDXej+v
DMhRvWnG/IttT0E2DOaeRa9HkY1WBNtmQgvkXjPaZ43e+IF4qFtMIRL/HwoYvWd7cN6MtIBZiubA
nh796ViyV10wkCjkMqMDidorVFuu+su7tBstdT/D/51Ro/HNSIxM8Ij1fINLPGwLvUVHieWyytqk
M64FsXY0yqZjFnDbxbSO0pFMDzEKHVtentpsb76OykmRIC0H5MsbavqU0UBPd4AwS0Q0/SSa5+kv
rsZYfXrx96GsQNMPeZyjukpTGSkAHSNO08xJ7Bx1751FcRRuFcdxB4pbC+cUFFLoJr5DOlUlXj9D
2gWefojaEC0xqeE/TOGebcodV9aYnc/N+qZuRoQH6w39M3/QG9K7wGzOpMbzjre3wtJ2buuLE4Bx
8ze4YIsGfMMgiHTKDGrt1zFSbooZG/r4R/xdNHdry7XMfsR+bkiQxXz6+poTQinMWzd/Y2RXo8Yz
Rp2sJJGjS8R/8dB6Ae8+bu7ej4A8qBl4TTszOkKkiTAZ0mKMAOov75XVIXWG5r0WVxfP1znkP0Vg
3Z2e2HUc2NDfD+SkoQanbJ/sW0Z40p/73F5pDVCFe6xSRT7mNfc7hWK55yl103+wkKQuk8mSF+uZ
zvc08mv0vSgrIMU+DXLB0iQrobUso0ZWmxEsTKx2v1bkjCVqHFkL2nTmPIzn9W8Jrxg9lh0S1Cdw
hriYMkcsxC0c4g2Gp0q7spTeIeKSZZIGYZ83m8CCfgWVW5LtC1nGr1zYvE4SUTkf+CuOG3153JfK
uA5ikEXzQFgDsNnFBqfohqkrgC5ztbbasn0euS9zSap7TGgRCun7GDHDiop6AqmUJnYEAl4JW/hI
5pHjKl2qlV4Cn/kiPDsT1zFtJLuUmZUCOkXgqCWOtz7IR3zL5e0aemevPB8dJjkVI0tvSjeqif2T
MJ1Poy8ofBe5JmQngKdfB/1BhOEsItuxcEBho3tuSsi99Kd3bXnvyIaKrowpv0ZzfIay/jDJ5n+C
HniMf+HwXccyMrv0hJIJRDKAXv1eSbYBg75HeKF/CVczFykxm76zOhwV+qEBCHmFTMEROD5Z1rlX
evkfQ4EV+XVYlLwb6uDMlAR5X/II5Kh/ankxL9X8xMlvzbXJJFmncDI5OAtc9oocaHuvRh048EPm
LiDATeW3tT7E08bufmHYdMIZoZwZvv3PWF/ve0LiCcPUiwNGWGtLHsQmeGHyP/8nKO1JjvLJzH/F
TvNrucCB07PnnPglukrR7uYaO/gXOivoht7MahlrPlAia0humEWf4GX4h0N3nRfdM7f6dn8y/r9+
mgXtRrI5sGdAjNGLG8stN1rNZvmmNVtcW2HBbOGL/3vY/+Es8y+OAlYz0kIpk+4I2ykv4OGG5a4O
kNp3rqG+Epj60dbfIvDmDsPU75na8Pc0dht/jYmG8rB9lXawqEEkbdRx1G2P/Vt0DE49W28RwCeZ
7knQdla9RV8OZGg0LVtdW4jPX2lO8CzV4Ue/q036UOrKQyeBdEG0wByv2hXEnF8cfptHy4j3+BR8
5dUdLhRrRzKgczzM/IE65NZiyW2NblExqyqwxvXDlciWfPrqTDEk0yrKOQZx42XY8FN8Tu/FnuYJ
yt0IlhpFUJW2RkAID0jLQrOXJ8EignhvXEGeUoXgsMOKOT8CRGToc07DUVOMtVg3sftoieOwvqHR
v1ADV1nNgBm6nnzXb7CKAMqfenqPu+e0Efj4o1kIldH663Z7Sowkzj2OMPmAXLsc6GFsEQKpP9K0
rdrV97JV3xbuinn1Ti1iGfATgH54/rPQzI7TrG+NFbqOXhUCS/i97r/E0KTwBJKn59eOzqK0NVdZ
A0tkQxNkHC4y138dj9qTRZgSfQc6/k2TvBvn/NOqsFuQvlCgkyU5cPWF0NKB4pYsdOMvnp8HGI7Z
RvPdduBVjVHV1xtnuCg5Sx/wD9kY4kDnQF7ZQmt+3CpTcuXnKmxYyGmapDO9pM+SHQ2WbD+8UbfS
3duYp8klVEmcLIRtubcdwdmXkUD8oiyoMxT4nrv+umTOHPq/jr6YeLiyQKYHoggvSbDtjIK0SAvx
BY2jZAy24dTDgfeQAvBQpSaHbCqaPvLr8pNcNIKHvHsjDYqbCNmaQ7siltAgNi2JfENdckNhguL7
BPssWfdR1fGD00cVZi/jOgBhvacpTl+SOFBAnpoJWE/zW1nmVEmr2m7O0d9KbZyo80J2cERj8o9T
/ERDzOhWmxp3AC94qbRRg88JDCg9i5ZKqeG4Oid0yOJSJj/P8XTsFWmaiQskYXnEfLJnpqbZC44f
u7t/BS28ONrGqNgPo5V4wTyVAWw9lJYzJ4mpK4n5b1heQAc26TQGSk65IHVBDMWts5+FGZFhGZZN
o13c+5rxgkEIEtp2cV5JDSZqR7/7bAFnytCfZ4ajnOAeefXA493LjUFPZwX5wRLirXkf8mSq6aEz
SS4o5nlqsTRWM9aidnIq/O9vbL6PqdfM4PUsHGF4OOKIi7Fi8GZF5GN4FlB2zvwwEqhXKmh1Hg+6
iJHpS4ZJFc/Fu6f7rH4azW7C/ykdzC3TYkPPzdn2sFlnkHjlA4XxmVcXkQ9L5wZwxZKBSBMNZnEH
IlqpgT6r6DCoujsqDkYuAGjCKShxePYkuRmAL96hrwLGfCis9493Z9y2Ct5X9Kn8jzJNE1dmeJUh
tyEd4Wo9r+/fpMhslc/vaH7VJAu1iuq8giwmLNZJR/DWGK9S5eazo0RCjfHdM0Z7b5xJlifHMfhn
tRgwLknwyKcGE/fkHNsT0n+j3V5dkI4xEdiccVMrmpCtdhRLYoq+vO/xh1e0HouU8yjDLkO352ZP
XjDRQ8DHpkW/CxwxvzwG08Z0cKSmia31ZHDyZOegROfxLn7Yl7QgFPxtHD7f7KFoblLYYiDMKm9w
p2rLwhsyjGOw93sHIrycGAxIgzZriX4mKq0Sh6V2JEJeyYEM58LojzFYAMNnewU5APg74yB7ZPwz
M0QsiHONSHu03y2MGY1qmFVFJ/rp86Kq/ZxJxtmoXDpl/JC+N8KGKSSHnuIgcB3n34NZMn0fnoYR
jH2d/Nx62FokeQbMpLVvZRNEDduemEGLiq4IOXzASw7t9ZzK/1ZmRhXAq21zhRG3aiLqR5AwHsRo
yMwc0yN3OG/7VbdESVtuxOjNhrb2TH5o3syPPBNrlJjOO7N6b7NlkuNpf+pAQbqg6+0nTKMG62Ll
Ri5HZI+eD5oNqtQ589s4oKfoBL13buni/pgY5iBNxmy+UQXQhAfgy1LlTODn+vTvpHDgJ9bjJ+f4
4q4pz/bawhPS5Or4zQxHzAOWmpwJq/paV78XfeiLNUA1e84lKzPXV3by/2Yrjfet1zlBoBQ5cH3O
fGvqQ5FwhR2EXElMY4LpD0pjQqnNC6FsvieoYCwQRCJGaw7343Th6e+dveZORwbDu0RatK0ARLOp
YxEQ4ZbQsiWNcwx9ukyaY0IRd001F7Chsjk45k9iACyhAQAAELhXbh9shLCtz/P7gle/YmauwubK
JxdOaMWTH4+YrVUgzCuNo0XnMPi5c+PINw7k6BWQiAZwsG9UH7+twwXAedZbaWxgM7+8Jy/vS0Gk
f4wf3SUKtxr+F5/w6lWY0kW1agHTnlM5OuqzN7lXZUICd1w05wa0NEDzW7VdCyfIBPsqjuBvRv6J
UfyDVmQ/9xUwjerNO/c0I6EcJAKdY5E02t08UluAFd7nfHKZZ0LmVMybc8Aormq2yWEHwymspmrN
mxlXb7jflEywkJ90ONhDJy7vImYc/FtJIAu8dJ0RDARMp7BJpMKDXiND2iPM1c/DsFCbHiPJoIV6
hV9Qi2j3T7o+2geFnnxiXQGkQ7f9OJ3t7Lb4dFOFLbt1Qpqpny4wwwPqdlPq7DTrxJcqFY8hcdlr
SSyJKP2W3G9V8ByRNnNgYI6RpvBBXsw6B7F/tp7uYAbyV0r7hi78rd+me5RWA2foqQAe0QaCePJs
LIk9WQBnwW96N/MhKZoqX9NBsU73ucPnCqO1QISUeY2eWpaGhpgEJIW3J/7ETI2/YgOeb8J2vKo7
CMq78hsrIeIVsvS6CdHP2+SujGczFbizQwbiXcOj4CWHaV4D55Lf66FxRNaks1boSnLC8kOZqh7T
b4QwJtcjM5M3kdefLqvXWtPDeoqfE6G1oLJiM1Ncka5lfKGyaaWoE8ToJu7qYfZRhvjJa7uhnNzz
0azq0iQc/AEqinSA2TZ/Ivj39l7e4mSRPlNAITSNkIHb5ltxg5Wk2FvO2j3psqO5By8+1YHWlG5s
wVvlaAq5cAmCntoeBgJsMWYaCLI6IACTbqJGoHDRKUGJJ9iPd2VOqmofl1sBXa4391TIdl2DDOI7
zrNFC5u3pUu35FYJBdEgjKUBcIReA+/hEXAVUgG23ft0Cq7stP2fmECtXTRZ/Jki5EwkrHuJ8Fns
4UbCT/t2azh9iRqRBgO/HpCot/l5G1emU/Cm4OwJFDo0o0v1TLHZilJclvb4JMLn48WEsNNVxNKX
OI2kcOOKUyTd7bs1kGXbKvuSQoST+1ZC3VVesUXsub5yxTanyHHYrYZp397lN7gnvqYbatqGIn7s
u9BofxaQogL/e9zs8UGMI61qhTvKvmE+eyitX4EV9wxHN2egCW2nxgrbjsoHsphHgu0qO8ddnHrx
0Tvh5V/XAMmFCLH6FwcPAXzfqaFZ1C12LLjYiRp05c/OgpgsGaynh4/EFW52fPaIxvwEVfvjPYY+
R7+wYcL5SwecDVFJL1Hgnv2M8tIVohgzPCIvkBUVVRVSGpirxmhDeCYDsvd2ZVoh4fT/hk1wrY7F
ivpOD22ajIDYh8bSXYRXkjJd8L1VR1mNiCkOS6alKyPBYlZ0zrNAqpL48mobnJy5eYsncqfkE0Jr
0dulKNLGH0k/V1DAfIfGKGLKCzwzvr+c5sKr8Z92LaGXB8n7c6eH1FGwBwUT+640kVKCe1ENPbXZ
MnvPm0xVJDfexeN6w76Q4BALBTSi6iVA8ly9vdXBIKs/AIbFXZdlAkT5rFcsBuxsvCkO+AAgrTVB
3vFklqUpa3qmzO3CbiY9uBSr0gW7yUbewheZYEITyA09xCGeiMTDnnoao/OeAyHH8mjOFWZLzWvJ
CdSBnyrQO1QsYOT6zXzMs64+hizNcVKccFv0zQzJ/JjMS1ysajd7ywj6sPgcc7VN30oCfDtI2WQg
pXrnU1JfEaTARjytlntkLBSB3ZbXp4dUrA0ACNL2Of3h+xKYpSTHS2/M1qi1zAEQQFy4kP7V/86a
4sYW2lSEZrm6ePYzHt7EBXXymJjLQiYJnFCup22vRTAmrbcfcifpUKuyk8Fmr1TuYQCt2bhQ4K2p
XLwZNjej0mzjAQfajdXR5CcpWGeDnnj04086MkodKNpGvkMbWs3+yIMkmwRpqzrdEmNrEq5s65JB
zOWZdxxIshlu747JZR+7MZdOahcTFYAFtT+HGFB8dsintge/K8VtijYL7JrfBlgBfT8HHS2OXfLa
k7FxfQK96iis0iXqFOxL9/mh1QLAxi/0l43gczuQyKZJa0MW1FPrnB6hhLbsTzwD0dHzvkiMzQir
Jr3EYez9tjA7DG1IVcCTVrH5LbVtttw8teNRAxFA6fsHZtLughZ+2gg1WW1XYCAPDS4+qm9K0id9
LFnNq+E4NKIyeH+sCGXbC6A7BSE8IaYJJoj/RYQRm+lEPaTzFaWWTwFf9Wp2CpnR8RRjsTgQOAC8
/rFvpTwIcoYWQw1EAQ9fHsRWqBlsfuFYCGRzSWATrLh4NHnLza0lhCfdjBh5Kj+XUDk7pzZzPQQu
V545RVAdUbsGIMYJEVC8DoAvnZWFPMm1PN0NortBc3XgV2TzCIJHKk+K4VLgKHMdC/stAJG+L+RO
VIzH+a5SDVYMr/ndca7zpB7a5ugmA8Nv1zIHune4al5VEVKXC3g3QEY9WvLBRYeDRC9F9kmU8DsJ
BpCcfe1nunqLBXLfmjFidpr+SGgBH4OkBmQRrWaUZZuayTYz63j0zcB9FiQpy5lW0ekO19wbFAHw
iIpDjqupekRGZaOcQ0OEPGY/yCMJaUTqyy3V9Fc25U4l23PeFmItbK+uksa1gEiPpw9HVqAhiUjU
UWIDPV4+Phx/0Nt2CIrGHXu1p5spw+U88Cf56T9h8zruzzuWax7TN6ji2vKQAw/c0b86/kYJQIVT
jx2cKtHdTSpb9yDsy0ifx1FkZJ8NooFwXjXgDOWhMHMR0QFz64xpWqrf62UpIF8CjcKqqX9xOEzl
mdfZSeYVgDsNpoaa3n+o3rEAPMldTWIJD+U+Huj5opWwQXXaZDPYoX845+QxBJI4u4Bv//bbCXYx
lxYsjvoo3rCfFD5wq5vnZ4PA5VFro58zz06jVYPXw8EyjejtbCA+VsHaQEhSxALTP8yPihwWK9fQ
SwBv4/SXsj5e8laDc/I3C7o0ncpSgOPzHiL6WlI+bvUY8snXwZrqBeXWd7FNhesgoXwsmlkLH8TQ
YqTDbcfzMMvXpbfpjFpAMKYjP8zR6VSHi9XoEi0A43NeE0Xwkwbph6cCIREli2BN/JWL4IZ+KYKJ
VSb2WvAHBACtQABvgOx+ztK/8r6jOlGRKt8pkCndlPcG1Je7kiymSbKm8UjOH/la3lqaEyXMALtW
9YjITL5EoEC4V0eWSEgEpEU7vs4l+XnUpKlEjL8YBYxnh+PEn9zeGO0CvgLOz6EgkPeQXfLH7wDq
L/sk/78iF3+X51EN7vbTMl7uCo8zfKPWbGWCak/r2cJ7eaksyoNsT65lCbZu8nlAQn+t0E/19VY0
nFqC/H5OYMuLUkmtIGqwQ+xAtXCWc1ajqV3issdIhqfYFYVvq+nvAvObfT0+V1Rj8wxIFakVMpm1
88SCJ2JLkDwRJHCfsZf3KlH5PB9Vek9OQehZjyB8v8Nx0l4rx9SI3epnfiXi+xGQJ9Q3AQqzxO6t
iHsL9L4uV8shYkfAWtKT5wA0DgVBlNjzcw+puTWxIuOPEl60RXRrXJLOyE7bb4TAxK0XRQU2lv+b
Y8QUl9Dnd+1XjS27NsBIdx0sZLHRMQqOp0N4kqp6cB63L4ZcifEn9vUvvMrYky5LvfsMpPQ1WZAv
h5lab0qWchIgthqY2mJ/Yes6oeXBvaNXdpLleiazd1z3+TCasIvhd9JsWaDnZzFits+52us0duex
Zbt4ru0ob4JFf+jhA1TwyqfhzoAM1+Ctxrq28BcKcSsZATP7cZVNuHxiAFUBIgZjUoPE9f+vG/GD
9SpPAPhBCK1/d+ywzQHxmyg8VmTxMuriJL7MdXJPurv74MVOjzWmmIcqmq5uQGi7uOMRnhkuqk+u
b/T/V1sn4eLSYKi9Yt7GkDa0CGgTg9E7oj0BUzhGlflh08g61xt0z8dPv2zyM/Ep5mdviOOL2HCe
Lf5jErpheqK6deME9hUelQg8t+I69EsUK/ptT3MSKBLTZvFc28Tic8JIHqG1hyjNVasYz7l4iydY
8qJKyHTLTFJL+EhbgB+NtBvLfpkhhZFLotG7trqIvJfWmH2VkKtg98u6FV6y8Jsv00cZnOuI8G3U
Br6NEj479qGdzdbYeubCBqh6DqUAoTot73iKu5KBuVUGqBgq83LBcjzEaa2m+zl1pa/y1FRBdha5
uezsI6SJIkP/8tJHHlYPEl9EOsRQpcKx7TaNtY8j2GduIKd7302gUHkVHZbaFS1/JKo2IvdRX3X5
sJVJHjUXkGvP/1dk0zMw+oafyzfRJsZ6wDn/USW1tAclsjjbwoqyoNQ/HE68U8mf7xwbdPz8qQRH
eCaDK8OE6bZfXpbQ1qfwfbFMLoZX14bo+4MpgnIxFFtitkPX0agcvliWjCySX+YJpQ0/XJxQcV7z
aiTke1jHhhHT/lSC/NanCC/4NV8RN4iDUNMeJNNs0p6BN1MNgW+Oe0qAJImYqujkYjCw9OM4nPlK
tTLoARkipAkr12F7D/5PyWGygAf1ejWl2M2JZ1zs1vlD6CNk+z/t073FOz3hDXLn6lDI96pvRjub
DdD8ndYdPA2/9T4UW7ZA8fGPkGct4Cd4Td779CvENceW15E1I6bls0YT/Hbkiylr2OHAUON0DIBo
cWlsUVS41F1mmOCSZwGHeXwBjDp06fZNIaPxtyd238KHli+WEH3YoeaC/7teJu1W3KmMce+iXgyW
vR+8y0twvytJGD1HZCSgYxmebBK6oE26Y0vIHUby4sBIF+qboh13LP9daEnerIWQeJBmWGrIIRS9
mJ0H0D7W429I0cWYqE8XdbifFpUSxEgkzOxgD/aQOsbUmv6OMFqHbmk3YEe5wXTZkFEuUc4LGX+d
Ti/aJPaRCDu0TYS3Z9/pZ4fuhu5oOmlWh73CV+wm+N2oKzfVW46mrGH0FdattxTQzE2h3F327iMl
aI1uQsppCbyRrViZ8KKlWSS9hyOZkB3hqJHyXZreC9tenjwFh1EDiRVEBJLCTK4bllWwVyWmXOf/
Jjgi3QmvYhVUYhEsd3ELmVMZEQhbqHYKYZAmmC3Vpvy139VhCxZ3mwCdkHPhcwcuGIRsFWOm91nI
U8mPElXp12IRTZFVmXEIPbD4dfXqVqxjsw+W2AsOPg/voYVcKyocEw7VQ9kW/7pk0fST6NyEbav7
NYOSYRVxCmRxm7z8kG+5kfIKDvAYD75Cj6qkLbhDE4WzpXitbV7HjZCb8vDM42IOxEhxXFb3G6Kq
qM3CqNRaex5deDOJOhX6/uGNaVZi8KwotHeCH9/gQnYNBXm0w1eDuhPcgDK/MatzKqgDZO5hOE+G
ga7G194qDcg8DRjmGQy6TnRqdSzfs3wYKE7L2aGxg5iKEp1MTnmhkAf1Qfhv2knWsbNghiaUaGK8
Df7t6Q5LsIn8YL1ZJT2sCghV1MCIK35+aXsFNzP9b9iIrrcpeeMwLosm3yC8ElcLQTvOPhsAPQu9
oLwOrtGBL4Iti3UYQ5ZGeOsCURt6w1DGVPE8Rd8j9GTgZEwW8/tNb9NrRaEysFM1c150sNbhzcLn
JFBzpg3j8c7YIe0YFaMoeuhriPtcM/P4GWJv1kJMrrnY52OTyfVwzzKHSAc635N9waM7SXg4ChLl
VSMneTQOvmy0upCua7BOlQxqryYkOxu1YJeP7dcjtLyVuYWLZVneV4zhVa5eghZYvE/TroaCxIcO
YGFNwr0EPRf18Y8GgEG0ySurybjz5FshTkJWltGfRacaxzSZqwEvzeGCFRndaIEq7tuXO1bxVa9b
kv4NP0KZEJC3/IsHGho6KKgGOixzTnlceEdmymihKrhpRNy+A4H59YSUTSK9Fz48H4hPUATtU2GI
d0V+/Cn/tom2OeUr3lAi0tnS6aBtsrgiiW6FSOUspF6R4hzfR8LXJYWqs/0kDB2KB2Wt/4BTWm3g
2nsKsgP+4vLkBu/6lZU/WTbCV8DzXj+aveZSya0bQ2xbF2j0ckxrSHL/poSUNvQXhq1+AIH5qqNh
0lZUODAcY+t+jMwL0/ew2VXEUNCroum2jv+KpgGQp5zNR2ne8yshiHSktn+I8G9M++ZlinAWXBbE
4GlRBi6eTsS8+04AiqFM3c3k4y36xTiyGTX/8pMyen2e140WlIsL9v88lNZhRerCWld++HH0Wh+7
GcWdByCNkn0i7/OPdgISa94IQI/fi9D58JxsuiSJ4jZ2iR7uQLZaIlAgkqMhZX4tIVf9rOaawRqB
GKiHQjY6wDxPPcesV/JmWEaYQ3XyoStVErNz0FLk+EYkhXhS6PRp0TEC8b4SLOH21NZbF80wGnbX
Cv3ZGzrajS1jsEbkFD0eSnWldoC6FZzBlVzMLNhz3THKR4qyW8Ajbv/AP2+efkTb+wtOGmjWShvv
uxnOQATqx9U3GaAfa/mtlJHzKLoujPKrAj46b37V/jmszOeLqyL+5tMk4vUuSYFt7a+MJx7ef9gE
rrGvL9y1TEluD2EjzY0AWBqsID1GxEJpL2Dlay+c/iFlcOIKbtbBJPJLOlyycAfn34BZ+xbgikV5
28HUBSp0kLlIyq4qM8gRXfc5ftVDYTB6Q17FAuWQmO6iyfmwpS0L2/QRxenlfu99QwG16wvh9Z4L
mZ04RvgrFyUqWtvH493zH6uQQeQ3KTuk1Pz41T/x4NAQ3ZI9o7oPJ1V38j0MlsJu56MD6ioAG64z
isDBtnm1j3mXp+0/95nzCb9PVWmQoqlYDHzGcQ7mCvFWL5gxJ9979gv6hBx5SXM6yasrGxWH4/tD
h6JrfI61cksRDyMPWeyZWoyWiifl3/IJ9fDc5jJ5hP6TgyJvvLbh/4icq/Dwk3MjtafE6FkIzf2j
CCMdvZW18lkjSc3ld84/apSPu+gTJlRlFm3spXVcR3FH1rJnsv8fTb9JB+dwbUXTA9CAdYT+tafU
/RlikDg8QvJAbB33JkLwNJ++s+dUpthjTvQmwUBoSNpiO7mdIVmoHvCCC0YXLpCe7ngBwR6oEzQv
OybD72w0/EqS8tUGROuFDG1gcYeTUHnSfPbvVQCCeE2CCvqQmukI+wcSALiRj8BjGjGBQ0W9UZ5n
XUVr6HaOvFliTNJvek8gFS7lHv6+KCUPnesuJspG8ovU+F6PaKppJqhL0GAtmg2JjFH8RRfD8mYA
6MvrhlYdOlMvzd8I1ARj3AhMF+P6TIxLDu+6KiQEupya6U5+kxxKz7CDwnaDXzY0V9B5SH7h8FLM
xO0uhJTV9/uXoUN9BfD86k8F//41gpdND7VwzEXtfrlAJXfFyiIoGVgRvMDipq5FaW8N+3Ac+6bw
I2pMhf+9mRlGC3Ra0hOKwFLJEjH3qBhWE8YZzNcH4j3WMqpUe6WKxd/l6qcB1+agztPKSWYKnmek
6BAhfgi1VJbbCtypBKkIWy33sp01Uop4snjQCA2X8Jh7tYKLXn6qvLqR9hXW+aSTuYmUit5fEZaM
vLjFxGor1OWLqbVPJ/nI5bEnAG4+99/K1qvK4w8diRdjVrZPe2p7+Ls6HeV+K5saW4ecXlS1PZPu
PaPaIw0lUWysqQ9LbRlrTDH4Hz/AgPubUQUWY1kOL9HWFHqqLgBGggN379hvyWSnHfBbkgfeDN4P
E+FNbfMJhBSB0UXoUyjn6IIwmLhZd2nx+J0kbh7frCNqjgP9Q/2bMEQTVXtB073+kj1zkGOsWe7e
LOQ8FOMPY6tIO6eeqe3ebKlkk3mW10tgA0tdSVpfwlkG7QaKSEZKQTjHeDLQDZzhRQk99Eu1AaRN
Q2DFs2Nfxp5Pw/XeTi4+Lt/YLdXu4+OttkfVw42qSk2drY8sYiMqdWPZzV1+P3PY4n/B6EROx8Sv
XTGwp6Qxpd2/FOTv9RyuEczMCjhlj8rtIINllyvzex2wGhKU5riePnUf2TAugoW2kVabo+HrzAEu
B3QIgb3cK3JqOPBz0hnD9IKMOjEPoDvX+Tjm2hSBKPg66G+kB5SZEaZ1yNqhAT70nwO/dgMz2s4x
CQM4lsKB668a1YVrBb0BnHGHjEyRhDYzJgL1IZFaLTnQvAVAFO3T9Y/aZRGQ77kR41rHPT4b/kBf
lJuyrCCQEkpqfmy1TMsNNpPbT+fiZVWMfBqsn+2SWU3OJa5n/EA0wJZAyyjGlRx5InVHUxXYNLzE
x3Vq7t8lsGbQ6cJXWrgYJPAH4Ctrt+Kbvxoj9T25Y7zJqwICNwtM7XOl0FzBflXBNjCiCH54jVFz
w5YVIcz5PoOGaXuUkoBL3ZGLhsUSrCqTxGdRwQTTYNtrS9PwYQD4K05UjWqgH3d7G5yqjqW8Q8+u
BLTmGr7D30OGP+K2JNae99jlZREvD0TJw86hkpzMLDYMwOD+bDqbtfWVtJYgM3pXYQqJ7Vfeuo3D
G42I3ES6ykIkjP8O+vM26u3zDZNRyCZYupnfm0Qzzmq0oVZEV6kt8jQ2wQAwCWKjXpmdElktHLPS
8fCFsV4LzbwcofUIqCTGR6MyyUdndPOVoWiEkHHCHtBbnoKJ7Q805jt9tZEwq8GBDa8nQ8Q6SJ9x
vd/hVdJMqf0HObwAGony7g4hOqgCL9xgKQK9kKGS/bbXE5rCoU6TBw+H6R/DApnWKEWGiJ1FvoMt
tpFzQ2NzcAnMRjkTT37QDBwB4xn3CqEhcHyJT6ft58Jgo2YQoooJoA0RgR3vPxXsb/dP1rtoNnQu
gzYcaixHju2sQElGwEZdQvwFGX9gvfgqVneM8/+nbJF7II03toGx8FpNeVNOpQYegPUXDBfHuQOK
dAzBw8IDupx1tnpEjp7SfrpHW6QI/kR4V/SIEfqPaS2VBsmJh2g960pJjmSn9MISp8kLh3Ww2NtE
O7e6XgQTR0rVLWP7xtGtneCg09/yZazWMQUzkry6rzn7Z4bHLyjzjT4srtzpVyq+hag5aH+hYasC
GZW8br1tUTYyJ99I2yVbKAT2aBSBG4KpKX8msMgiWPsXNph/pAftrKUvMs7Jj16HgjDcSdw83a3C
dyOgkekcCQ7p5T1nZ6plzkrCiN7E/H1b/Rcex+Ve4uwqpCydB7xE80qNG6KEm92FyqROLvQK9Ela
PHZ2Kn59WUXI8S+QvVJ7J3F82PjumjBQF4AxwIARLlUaygbOFDZ7zm3Vth/D1n1ABQ2yekQqF2tZ
ZKEI7W47hzxOhgkY3zhoheny8rORfU1nrpIuzqaL7jTVhgvym1YTSyeQsZ4DrS/DCBixN9fBGPKX
oWAEH2U2nsBW4XrT0AG1jj81GqwYOKRjFNtS/JBx6qBOuU71b39lK5y6HIdCZ0AORcmBDxosv6ZB
pwW8GzKJgxeeI2fRdQU24DPiRAgWSYDskeffZ/AmHbi967IgqtWSHTGB3Q80UJ4YX3e2KOmJq0US
NVQA/XRAWeljSElyp+i8S386QhE5Z7WGRYziDM7Br9A7nmrh64zdduyFMAXuD0swcAj/5EJEPwx/
esAwJ0aWBXIfzFMwt7iYub22Oe2UD3f/NPe2NNA5jrfPrbHXvqjGJWPgWLF4B9pd4xQ/heZlkfLJ
4joplwxDgTLB1G4VxSZ7GlqWw+W+RmGVgge39RjDm4nseWhuTOLpizOsNChQTsam9Te9CeyQ2V5l
+/IsQ+Of4JngqvSe96GnYYFsWv3cBMFM7ZD9KeDFfltSiGvHBbPSTit/nwYhSlCiYin5805R0fkl
48aE/DQqC42nHbcY3H7XVlHRYZrj/fSZu3JY7dUXDoq/XUQXdNx5l9PnwePAnWqpHTGqDv5jlWth
P0ZP1KmpnLTrHyUiRK0vmlGN4Ga8HGVgPF5BYlVl4kpj1CfW4DrbTcVy0/kk7yfHoI8zsUYi5MC/
3kvQ2WBi1Lo4fYSanaKaVQUAaAXGwqXTHc+ZKw7a68Jr+PXwZF27DfnZ1li1ZPTu3E81NIv88wBG
MzeYvKAt3M+cn0/jUa9E2zchv3aQedwzNcvPOQPFOc1zXnvrxqnGFbeaPz8Oh0j60K0657ZEG4LQ
60ZFacsMvc4XPfQfpPPIwyB6h/bARaW5F1XJ9Wyc1IwsDz9C8SGSDcFeOoHNpZysqkgUx8IeFf93
nstxR2kw9l5VWPmpUUFlqAwe0/Ul+QAwriKHH5uJn2DTZJaIF6H27S0lrBxwY86emp22tSdnAU8l
G4PVLeIaoEssCeyBdn7HilzainaMonqoQ4PY+O62n7eY7gpKuDpg08r6/bLP73RrvRk+9d/vYx3O
xd0nRC/yrXDHg1SOwgejufDAUuD5DLAM002nwMvMs+x4P1WxFfLW8JsKQjZtZEZD76Zra23NuufJ
x+lDDHhVGKhd0uWwMC4Ip+QnPH7WMR99mcgEYZhE7Cb4L6kVWoRaOouoyZjonhGueTiwDIPbzwFa
f7CMWj3NVk6kzOEgnC+9Ar7RPIJFlcwhW9BO0RGPcGKyfmxAbvjUWexIdpGP/L2tc3kx/cISb7Pv
SY87wW716S1U7nYRAEU2pvrxuB17ORqzgx2wlM2U9v3CeQ4VV6wz8SxdHWXYOYSVzZqAnarOrvW4
X9lzrKUZ6V0lOzg4Z5U11XlIDqzuMOyq0WGxyAwy+ma47kD+dd6m+6FkCQmJjC8Ua2nm9ybi1K1U
zhQSwVb4FUVawcOQIykHlVQjQYZ00qYJOCUQUJAKYeC3Q+xW8jP8Qka0tFDEFjthmx2KWfQdJ9xI
fc0etw0eB+0wWdol/sSwaPhorkALT7bw8faz9Uzlk3h9eE2ILRgsfm+/dIHvI5PejlLIZIQjI1L6
q2TJKYdO4FlqAFrVynqmBsxef8x8SjYtznfBw2V5ONHjLP0B1fL/WPhNvzgE87gAfw98khzB0U8G
CyRey7ddLzAeD5zeju1I/4TJz3C8o46djtCZhZQZx9l8BrIY+RcTZE/hR++WoxriFc6txxtqzQsR
Envb8WQg3g4ZL25Jl6z1pxJVkTMZJ1cOEX72d2qpnuJro5ptr1tqWfUQ0gNSsrank0kED3BplasH
ZkjdUZ4En//N3DvmJ+GDKcqxf1dPVgXw0rNohLw160EzbVMQWiuCMVRHzlPi8Dp60jXBZPO1MyeR
oqdUK1213ZUtiQk51VEXJrsAxGta9yUOHVkkn30rUcFO+loAfqvZqSLaIsjHpWpY3Bu+W+swYoWs
YEqAoAEQs9Dl/5nW1PvAoqb24au+Wg/5HvlHd7hYX6HQ4i3OCjqAiW4V8+XQQ05DyuB8gI7eTR+8
JfaxIBGykSPIWOFaT/J5jlcdC8twWbSLmHuQxxg4gVAesGeFdBcVaOwa90iZQktI61IkZcbM2qtq
yF5pUOtK7+4ro5MahkbEILiYinylJgxTCX5nQ/54IbKXY18BMqhtRhAQD2RXz3eQJkTt8ozo3hSa
/eKtY2ZIVaJyyPDXn05DcDjtev6+hPNxdfrCNA0CoQvwF5RJEROeLCkLQ2VhkfpoRqEj4Pf89d+F
tCjVyoGMF6kkLRy31JepwvpuCVQTZWwY+HX8yyqVNdtLAXiIJa44LsVKWlS0C8OACkNdhTgwnL7f
vedOnZ3W0fQyME6t6Mg0RZDrOdJNz+gRAfgw3/8Ex3V0SPsCFFKX7BadaZU1R+GSWjXdx3VRckU3
8+TDP25dgesZxJp3v3do5a8NmRQ0K04+QrAWVRX2IPjE7eVsIwAYiK2j0HZxALMGZsuQE/mFEXI/
B8Zpre8N2dWaXKGHvhMUNGRWsM04Dn1JFCsOfk/a3CF4G5HyOqa7Ln6flhwYVmt0zvPD7rmcv/VD
vFZGYUNQNWmTE+iYvgjf+K9vKZOUpuZz3NDwfb0xNPHJTclyHzq92qcWVka22KEMQMQtPbY5X4dQ
r06YkBSolTurJOkAh9uO/Y/GysAJuvYr4bfFZCbPiYB1sAQ7ALPLI7u/nvQ+KByp2+GwKiP1RJzS
J9iaRouBrrQ5MXzgGJnbiZbVRDvITyBwJ/DkykEyXNUsNDMyqCS2iEqlBGEN6uGDIJe4bWUaFdv0
SRrxwe2g1oft1l6KSYyz5+wcwiLlLCKhbhRhZsm3tA9s+yOtYtbjrOnyfc69mnxTMSnf6X2M/SxT
x6s8Mx9QlA6jg668ENJ4n8v5D31/09FUPw57MbZmqZ9cZ3Q5vIiDygf7izJLRoXFm8aPEgAN4ONz
TCBMjklLNseUETN4Tf3z+k/uZhio11Hsp/BiaHKFWFPpd2Ol/w5fx0RC4AK6YxnTpOyB/6omdgh8
oUk/GrAb/aE3IOYRufcz9vQ+vWCcO/MOwkt3s33s68DWMNTpH+U3l5zJiuds68Iq9KxOAQkwGAaf
8Vz7PS+dxb3jRz2vmOI0Nuvp1l4gY6FOSvxCQXMZ2qDreA0s4xcNfwpWYiSypTuiwBkYRKYSAwJ+
6vBYr246TRqgzB7dA7NknkQ7oOdsZYwEY1ES/aZ5HfhO/NAna852ghGM7rdyasaCLkDOx/VTROkY
A/O3C3B56puT4KoX7LtI4fyrjq9uquUKDbpWaUpNN9XG1apRSKzKKZd5n3AbqblVnZsgbzUxZOY9
ZS5DdOeWBl8GlLQU+TgZ2LN+ymqGeDi0PYgDAIrF7Yk542DXzv4Fk3RrdwefBN+Fs2ZydlQ+z+ZF
forlAW3WwD/97Qb2nGGM8ILhBf70AQ6thD0ZVJxUo4fP77ojjrtulLZCYpwPwNhK6XLga3o6dDNX
XpwP0xkEQHxdx5TYR/ISbD2DhgbqaNcCFt8GblC5oLqhKle/YkZ653Ir2a4J2sOSImFE1W2knx4c
85e6dnlWQo9jr+govlt9gzGyMqh9xqNX7lyWKNuO5vlx3owLrgAAPU2RZAK2qKdvKgrgxHNgs++g
t9VsDw+scECips67e+uhnmwTG0qPUXmGk7sKkhcVM5r77gFRqRGKQb9aMT2sSm5gkMr+XxoDZA3Z
T3uvfQJWCgAukzL5ejK72rLsFuOR+KqSJD18E76I6NAtlPVxHw3vLwMOj1Ln2y3JhUfXfZPWN3aP
okzX3VINMg4IOvN6rgW+LPww3oAqrIxVaTjMM2q0MLt5JaFHSmj6xmHbuFjItsL2ZsKIRFiy4EQS
z74U+5873KfT21fV/GrIPZxw9PazD1KucRx5e4rSYQEPwYj3YsbSQ6cr2GiD+4dlTHkahRRThZ2b
kxx6+Su1RUMhKrw/fuF4ge+oFMWJzJrPR4zSSnnRrhfXsszwjOslrBCauJzDASE4qPW6ftr03BuC
rhIQlzvy4Jt3OWK4BaUEUfmHzzjhl1N6xpxX/XrcYe918kXVXwKN9PVKOQAnpFVFwVNKytkeTRGj
IruV3P0RFqoIGjvsG3gxJ7VGiq0cAR22yBX4l4XM85GqcMmKujr6p7vgAZkZtP/Oqy18SSgKGMwo
3QhC33cjYhkGACdWYEyG2T4Uw3JKcNXixOqpSZhdIug1rUvc5kh647iQ9iQnItr01lDHMkmzBEeW
cgZrweB9fgaNoLAV+FP/T7UX1NybiyUJkz9J+adRcI1ELy0iaQc1SFJzrDRQ7aFcl0eRqXnXfTlZ
juz4w/uW5/m/l9FWDQv33cAWN0IlEiKbk3Di1VK9W/ehtq7c7vo2/4uGgLPZg723xfig61ZpK7CA
8Vu2ZJX1w1ieoLkanwJXZztz+F9QhPwebNPX29Jv1zvCCkhBNVsgwAk7/t9zrABv82V/vWfjUxsk
qZONexVjJIaPjPHNSaTQmbaB/0kHDhlmjbbnnvFGwpf5JMcqfy/RDIdbZU3R7NsJHCRkhmvrSf0I
vUFtkAq8VCt2OZygOMOaQlX2mqmYO8jX23cWtxTvwFi2uf+cUKo4fhL/MeYHPXhR+Z6Xu3/5Xkso
D8RjW66iMxjhF9sstWkztAtjkfF0R+Wt6ZN4NVUcVdC32/tL/TxSDsAI92QWQjpt7zSv5DdFE2nn
ToJDmeb1g3GxVPxnL3j8p6ye8aszAUWM9EgHn4q+dUfnvi0+oSxTLnTPFFZNVkmIwQfEfqu7NVqv
6NTF6xmb2YAjaV9gmqtkJ/dDTEbwkxvCgKqxizEKtr8HO/XnWnO5AX6srSN03k6nNlGNqbd+BozB
KSf0oDuhztOoqIDiXTq6u2kLWPAfuBoQ5rahNwcEbArex8Fb/bOWAJ0BpNkdqVQzKBDbJdeibuh/
4ei1uA5N2RDrhrfhuzhhc9zf5oQ4v9kUvE56k6YM1/+vAiLV+DjUjqASsdyrQsJLo0UrjELXiNxv
wyvS0CbuocsVBkmLRvuE4Y1+/JWYxGfaopGqle+p1n+MBCAO9IFpF1INJ9gQSJaOau3ThTw4p73e
kEqfWFLQnyX8CzKVmmpzIYLinRXR0KNEJ3XAUOF0sYM49czgLUV7vn6vj0IkYEfqmNOBriHvFYI9
OfKqzw5L4AVq7jne5preM0skPk/v0ls1lVoNVDYKjvpamqt1U/8UBoxi+R8tDxtMCYT3+6MVPwGa
essgO27r/VQ/ByNGRteYE1S4SoN/McRIaT6vupdom7WP4N8lNOlFksc9F8Qg8qAOpOGNCts6K7Wd
ybvzW0vngRp7hfeaO1JzQ8PhHfloNcb4h7R4+Wz9l/ta5HRxFmBqojubfEaVpvkmvDzFgysVZzaD
Zv5/+Ewbbi46+3ZPnzZWHm/U7LNUMZ31bZE7A8HyzhAdvnOXP/cfWP8Iel1nKA8V1R/iKGGMBigx
dSOYEP/33HDMRHxbtKoTZj98xNKm6dXUSYP3E9snmL6egCFEptSsuDw66CORFWXaZzSqyqn7vvd2
BNjXnNRdAVMiQdkoR9oDE5LzvoeuH4TYfUm5N8MYGWRojgibO2A/toP1oJAWryanj8KkKIZ23K6c
Vh8j3fcnU10xN+mEcNTzZAuKTw7s122u1w8dY1Qt8wzSCD+fHrWpTny44W0uy0TcS548Z1MPZSY+
9vndA70Mckw3hBv6dccK/XWkYqwU1HF8I587sd8kyRyBrogIMi/CmYOar48Bs/xBQxTltRzm5Tcb
mGmduji0F2TI1lbdkV5Nt2w7/2BkOp5LCNFcmOc8e2FLeDKPhHT3fTIBAui3lrrIXvOykspbRNwy
V5UEO8Ps5eyqwLGLKaYrpKKLqmq6F7qLruaajLjIORyzGGoodZo5WYo6oGwJjbe9a/sGcrJyjRvh
k3C94PIfVEJ73J7NtHauZlWKXGJU0NpL3ld7yhshuwuvxziz/8ZHguYt0ijcGjQ64TfiBeNo5hHx
UKXh76JZyv/l3n3FjwpatP17/JqR32P3oIVCCX2UR03E0zydH7cfRzrugiXK353ulyhRb9EHDcya
6uB/drB0mdiZkJKgi3QsX6L6MQqhMQ2gRr4HO4JymrBtJsD7uUlVuOiTDPLrErCL+JVl685spVID
MXRmSTdLRojhDrx/5tjgdSdHDutNu+7cEOoAmVWFtHZEIWwHJzLJZ7J4gDdaYQoR4g+DZt4gVqGe
IsHsdTw5m+lPMz/p7MLrMTt9bYG72pT3TykFgHkeajrUdnfGS/cp9pTndOkpMblDXkOTWxXfrGRe
meJUv26HBvoD2WBn2oaScw2MTUoZMV0EJxRwPBPUOaOUFTApIqfGh7q3iL7mjUntBre8AgmNLPJ3
9/b7lAomnnMoYn9iG/yVb4pvw/WCESK2oVw28GM+vDsR0N028eT6lBpbDDLuNm0bZLkZSy5keXqF
gJHDB1jDQGd10lqbX5K1Fnw5fZazD8WfNA+IdyxHwDCEfD/hTC0wRDfoAIP5/uXj2jeiViTDbRJr
wcpOE93Iq8Q4go1xZrQC62dvpmabcB/pyloNzRLlH9nhwS1jP/vfKgS6k943BKO3ZF4GqvoQjv+A
hSap63FVkwAHRk8qpQXoFHYCvG5H54QZ+fpayYt6OLoQABzyF5C01xxj2aS4uuYoAEBvy7jpOrmM
JLjmpxLF2jxYLxhDkeWA3PRyQPL/DKQMNP5agLCEVQuXIE6KD0am+pqyLwEyiUFAtZ49teD6lWEM
5MMDOJeLXi0HzijR+bqJNn3vFeB927BFSnooPMSW5OK/eYF3GDXAsuH4DOu9Juwvt966B2vSjmAJ
B9W00U7KADdYaq0J1y0U4jOTa6BcNivR1bVYNOFXqDNNJVu7IYLYUOpptFBYGM01WK90bhMlNAlT
rWHB8y9x3KzjljjthGYDjFwo5XGI+EBS/euIUF6dHsxkKxvb4NKuD078RWc3nwOIQtRVm4/QisbP
16D782JWMM3VoAhLJsXq79/Ev1KoFbQ1ZRL41gk8YC/rZRu1x7AOuEmXY+zX4fTg1BfHdr+8CTnL
MmJdRW6Od+Po8aqPTuojb96edfE+DtN2Qo9kDDfGRIMXhiEe7RrtycSgXVozoOlB+KyquyL9ZXhn
kIZ6G9Q4umXPnYZz1886pJzfwhVexUvvK6fv2GM+O4t7/CJxq6+Gad6zXQTnGCP5Fcyc4EIyru9Q
FIBAUpT333mhWCUZRQi/VFHba8M9PDRdQV1spmz1t7XHsU3s0sXSFoqIlHWhq129EZbckthM1s3T
PLY1E7eMU3Y5u+68WtvysoevXd4QflfqmcYO7y4vDQXeeYLTIMHw5q4FKQSJGnUWghmUNonOSkrx
usF+NFGWoAtyq+7waUEmR7dbtXgQxWPuY9Vr1dFihXC+HTdWFOrWD0wfzpKc/Jwo+wq/ssk4fMle
NLjn4wpEtbtpA0kig7Z62VGrSm6uIfrLrr2Zj4CMWSsmdhnKyTAw8Bq5bSR1WiVJSjqrHUDho3bZ
DDXGMym6ni9v6hUQjlbUjfqVdFLF8KodTg9Ph0Lo5HUkL2seoH+kpfHOzNFCrjv/aoz5psxS1m4r
5I7tirBJIblwQ1INxTdh6JKkk4s39J7AZ47MiJzB/Nc+qykewtI+rLp2uyVi+rP13i2W7qxQHgqW
uAjcNRXuz6g02ajtCcbNNnsb/vXlBOtdGSvD9YsoKZinr4rWzIomT2rh0rcavVGEurF+i+V/xHZ3
iPvHSL8UI0n3g2DffgqOhYjLvsi7SXrubNzHsVmcUHd2VAwG3Bxth5wimDQn/M4WofniXmCSsjtj
ag5+T+LX0D0EO2/qaZQMD0YMxQEcOiDm4+YF9dmTojAYO5frXqr1gj2uvj8rbSzyaVDqzgk2vMNZ
8eWIsLnYw4pAjmwTLKoBg4t5xqh01brisVAZrz511fsg5uVdRZY3jCqRlX28fmyNcIhOaXJCrqKb
/eAO3BUtYwwpVQN1Lnxt+59fUuVFDbOCXvsbbf1fSZHAUtaQQqVtvnsSc9l3skYZ2VahH/fV0o7f
U1AyHuorcesSVZkCC+TiGRRoJYyZxI1AyZRHlNv5N6GTWvsNZu6q9bBw9uZXBPbVPLCpimr2+yTN
Oqfgz/dRHoog5WjQ3+WgZLf2UgR2qhjtx5qkEPs1OnL/MlrgUVrMvEfcCcis+p45rWiD6nZ/22H9
nd9smo74WBuUucXybtdT8rMMsQM3BehJfnBueZ5zR86KooZD5LlKCYgqakPUZfoA8Cuy86nEInHc
xBaFlZ5l+HiU9akeYLYxdZ3A2/etCoiuCULNYRe833M6FT1m62UqdmPe4MhteU+vq21JkbdLATdv
cE9o7uBl4nlGhgJ8IRxapniTtwLW+FdZV62oGt9pRxJ6vc3tWWP4ZOwQAxTWDMM6Bx838OJOwA0s
hkLuupJ0B3OoFLqKKvdQsSjNiBZqYtK8HC4mNQgoCvbC8w0bL3Xch4lEAPsLYpTvCQxLExvQveA2
aMarX0EkfzMHWv5R1YJvb6FS2d6aU/S2DkcVh0Lh6JQarYuQr5nrtujwNDvsCWxuIpLwWhVF1sRk
PvS2a62ZpsyxTcyRhe20R/uG7WB/GsU/25O8STWh/45paVKsOMa9Hd5/52II1ZVF1FrRpXzWzVUA
R6igYPGDEYoYgBrO3Wt8OBQ2ixcxjI/7wJ3ACHOSrD5tGMO14vjzzpKWMARu86vXjN+NUufrqTeZ
6cKKcFb9JDbJNstvtLIPo73FvtPWfL/Xty8RrPWG6muoZhNFi1s+esr3VGhzeRSAw5w9KKv4jWgP
uNCW1w1EZcYVBtGJqPPK6wHczIJ0/7tegfpgqbp1Zmo42RPdEnodyczFDwQTmXFNllDpZhS1acvp
7PXpv2zhfjL5pjJYOxaZ60hHvhZj1DBSMXhQJwL5+NcTN/k8IfcYfOPrQMXE8YENoH4tJFv9mtA2
0RnGuLYWnmyHVusu9WCLq2SIxpi44IA5Bh72OzzAvvoBlPwDyovO8npTJRmwCXdLD/DEApKAN+2U
BAZlmnwsAZOAUwFjayK4+Q6BPoLlK9BvyR7XdoSbBsUTVRhCmBY5nVyhiUiU/1orH4s4UmtqgBX8
SxKFoQ+k5gBz8BdJYW+z26fxbEwOxwlFYIAVqJp7RitxMq61LNumYYYoq/Uia1aYwUkUamwAHpQ7
abAfEofQtWScqFT3qHO+7Nnaxlemb0eBzufW/5F7RKAQupVS2ZDmhIIYwOaHOeTM56u4k+htZ69J
QaHHJ9S7Cdu7XnkWPIj4NZ4gWYcgf+3pva2dgNZ3wNx2FBsLk9fIbQ35j2HU68VlpJbcS/YI3Scb
gHaUwFJ9ZnzDYx7gk+WH3kS+/uCwsYE0ceDJXYxc6mncau9kh581AvHNe3ydO50wjoJMEJHj6AUD
hY4r1qr+wHv8+NXLrFP5JSl4kWyPHecQ+TC0JE+RFn7lDV7PuUbbOk6fQTYglQmpgw8u8pHSkpk/
fYon7wNcXIAWZlXG5aHeVHCTqn1TeNlJe+iAyBbKhCvHw5Tu0O6yy5cpnxCYsPYmYHaEroWL72F1
nD3fe6SH/zZCf1gJgSCtO8fbouhDzuIYg/P2wftyhXKFXlO0dP2ar7j+YDIE4BDg4q3wBoXkAgxX
OMoprgLzsKHa7kA8ytQDgD0Kpm+4HpVIZnqSYWMeYwRPi/kGmG5r+v86DqfKCd3WVGB9tLmaiF2V
Y7No6RPpQXKG2nOc3LLRa7xJDoBsNIDe32TeeRtkK2Pne5gV1PnNG7Th1j0OTjNUFWJ52Gc9Paxn
cVKhJMHVQBdCtQsFFqwaoGn8GG7520LIdf48SBGFVMrkL8ErHa7AnuqHXki6s5ZVu3YaIiK7YLV5
pt7KDLdqZu/X/agUli76WmJB73zIXncW9o30k8OFpbBat27NGIRDbIEU4JnlTssnb0hntCeWqGrG
EjThdbgoM1K0vFgkw0H70CvE427G5XUy+ONguFEVZZeQ8rHwfZP4fkLu5NuRrlKWWZ1qeMNQwDX6
hqzjPqfbqH1YfboSzb2oyWVeQFAUV3u43u3Mud3PXNBtlF5iXlxmsAqZKLqLXmK9gCqdl7A1Br9i
WpxB/YJi4AEmgwPF309hUofCPsQDka4vROEP178lB9ui13IFAzUDAPz2unvr8EwNAxCwM7Id3uuO
NWfrDFPySxxywTWkB5yKcXY9Bfj2IgUZqtndA53nNOBGvXkVnS5tfIg26RhAkO/kCi6rC0WB4I/2
+bKcivwNs4Lwod7tCZ9BFIPBAZdhVeVj6eZXnyo/ceHaI7Gr4Hgl4awf/via8Xlzq4XXNWlmNweS
i7EtH0emFJ3MBGW/HfWMBg9RdNbNQMBcoL+k0RQU2GgSWUsnMbbeSYDFvNnCf8fGZacZoZ7gXDOp
2UFVHgTiU9eEOsiFx0+LQF10xlyhyLvcG4I3ocdGaSC4h+Btr1n/aZ+7by8POND2zRW10MhC8VM+
79IKnCienfS/Nx4Ib7ggsSD1Q6tgdRi6y48Uz8IZfmN1+xjpbpN6DV62a8SL21gbXYiAZs1m8wTW
ooaeffmejtZZEwklvqvEZO5iDW8SJNhMoGvCIyYRVnIS5FUY+5tUAprxH67xXexBIBswK7ZDS4/p
wXIseLy5QSw240gklb3NVOnHee+u0MK+ONQUcbgSahmreWtcXnZBWvXPP5MavM8zwxIHRiZD23Rw
pgfqnct4HIEV0Oo3AEUTqzyXkFldbne2gf38i6cogW6WQz9KRAp95fvolfeqmBJK2GLUTObx+vSQ
ZcIC06op1H44syq82PbdJTiwLdjvXeLjZDFlSzH9dccqp68zT4R0R2qK/mIj6/7AeNG7AzjqsyKZ
p1AOYktKJxW46PBDfCnD9v3Djbfd/5LLHsstkBcAIM59i7Y/R4alnjnDHEJrpMhRDSy6zo+Be+7q
BMaUJhb46SDRPY/iF1mbprCVwyliWiXyaQLGlL1bFiO33MhqDY/ACpe2/OasZ3ADohwrRMNfnB9b
+In2Pv+Ftj9J9N7aGQ+OvBstPYlypqcNVe+Aqg9/2GUfJbU+/1c+owxNBmTH3pnPVGh+fn6ZWjo3
fyQH+iRy92BBbRYduJMPLLf7HKrrFJIzJAfHipOeSjrcnRY+3k7O1+4c/hq7EGxDDY+G4N/9bmFs
MCGvJAZQ5muHbmRSoyi3ebG3/W73/5oXvPnAua94ipf8ijHwqz/MPYsVxyEFsYC9U4ffsUNHjsy3
dw7RHSiG66i6SNZYumKdL1qzcV05mJtLCp5VrN19Q3dCw6pj7JPYyaLX5tg4cSGQz9veco9UpG72
rhGSGlaXc363pcL43xQ2tl2DQi7ajcZwqsageOZ2iphjp4XmusZya/1LXl6GT8Ln+sd1tnAdFq8T
wlyRs8Qh+CA76IaUvr8/7xFCd28js9dY5KaOhMUtq+lQ0ufzgIeSbqgYQkq1bb6/E5KnMBBaZfed
UT+wBPCkpnA00JCm4K97Xprsam/Mvf9QVyXXQP0UCDLSoRpS9gci76j08oGOjWFWLzhvyzwJcSRD
F2NSnoBaM131HPPpNMBxcb6CTmD80JcyXnoxjm6gP5+4U6uvEoMTOEMQ0CBIf2FEIUpO+XfWyhyb
jv2qpgDzlMqtkTawC0HseWYLC7M9dONhvyWIz7yVEpA24t6pIhTAok+8r0utz2qYrhK1bbw93Qak
BYfv4LUHg5LAuq3NvB9pxDeS4vbOAWSUgHcwgilS6J2k5WPcoLT9sPZm9iG1ECSsqNOD4bz49xRG
vBEbDPMl0IRbHqI1gzyFaB/vryzv4ekp7JH3jYfQpNhIXtpLmbz/UBgzjCAO6vCxRIgetNlbmd9c
A4ovwF7NlOhW7A6tvOaq3u2dbstIxBJ561c7VDwZ3hCmdYPOXVLkXC8mgm3JO7hR24Qu0ltPNUKV
N8YIoGSHtv1qr3w2BVHzo91ObyAu00EPp51Ib6L8A9GAxIx9Qjx8XJWtM1M+hw5+Yo7md/+2kx9I
x5sNs12VJV5KMdEydn7c9uLXb5PKtu1wq5Yrb7+jRnZa/y5r3IfaB0EPx3+ln+iZTUn3WlG2UDAx
r+k1llCQHSFiaXjGp98YN0GfcXkJF9Hf8e2Po3bsFF81SDlo6vLhIVEYcqHLihbQyVVAVb6MPZq6
Gaap0XEO7SVpAR6tmFKIgQUQtUGxfu0AAHsklt8KUuv/VZC8SfEu0K4EYJ8B1EOzrm92Lpyym/FX
nlgLMlWE3fpeSzPww/oBhSrw0INI2NnPWxsdMH5Fn7jO+5IJNyB4w/slBFRZCkNcdrHeXpcaBPjN
7MSTZ6lpAozddT1CHj307jFRzsJ4Y50BQFYOF8hnjFu6lMs03nph+Z083tPUKgyq/OH23uAO2iyX
2fGzBX8Lmhsa8OiESCTf/Rb5xzHIKrIgDBmVtyTcwOd69SvA9zEzqAwmIPePA+Sqex1Zs+f3W8SV
0IFJOouF1XhfaaiMlo8H1zmJAL0AhURd81qFxNXz1xEXJYmSs+kdCT8yqded7FtDRZohRCbhuXwA
fUxstDF5v0mGfDygwJVDCtkWmRONcuwDY1m6u3EKOHrOghF9obI55cyS1OndkhSN7P7ddD2mja+k
FTXDFW9bzy6y5r/DoRE9dHWOS0s3iAgoT2rUi23dkrXWFLwoQYG4nBbJhRS+QCfMTs37ecwNMIJO
PO/v15jvlGy0Ldi1n6xeUlS+2FNi7iBdT0KRf3SyCXLDO7kbLv8ESobCDticypTYJIWxOCu0VxMh
Jbx90rDEcx02iYe1kc6xT52SsY1GpvFPEd8eX91OooYaQUXwzZmnCekINJfnOp+Uxr8irE7c1pLw
rGJn6aWtdguoeBXVfaXnqKWEJa2lXd4MrANySDkSiBs3uXY8uV/iij+0depxlWD62BvxNuFadVDt
gU11GG74KvtpAuIcC8tQTMFgYqdoWVD3aVcyIg78+9zakMM88lfiYdiy9Q5ju+R0+y09yjx5rzNB
ZVc9Xc02znnSsj3agg7TNJeC4Gamr4jBlLSW4Wv/NC6JZU1YAMD9MV0mdVo3e7rimW3OlG0uNmZa
oqYClaG21otqTh3mBRYXCMIdxWUODtikPnRWRYnvkXTxRstDJDEA8TUFpkvUNc3+VT22fvRZsNkb
OwSXtvhtWQ+Ne/zZPpnaDbWRxi/T3xEm8//PFA15vnNHaZiYL5sSS0k0z1GQKoeapmR+fw7evh8i
VLyLa7NMX/n4rFAgrSIrdXPRAZD2NrB9ch/o7VslT6pvhqcEA3U28XnIntNoX8LzB4rg5uNsBR/G
a+y+0icSKrzFYu7o7d30/N//9uSiJ87S0SBdaCM8fG+jWL7wci8frY4C1E5NvHHhKx+qFPPlA9wI
5fNCUGS1WFQaGeYbLHRwZtrTJHTubtzCPup1feyHdpsYRE342v0cTaNmefCjK9V+wvScuCGfQKGj
bn0X9JVXOMlPNp25cGzjpxCjh5OXqKqO0Q4MS9G8ZBsN+59aIaNsvX18+i52bBw0pcscYKH2GdD9
R+2jDwZU72G0G/nvsfPkdTFTszJ8Xpd3cAHFMedwhgzh/Y2p7UAnNpkIJQVcaDV9JFwYb/flZadm
zgpuU5lcA1j7W0bVd+xwX/ZSGJF0tyltvdPhih4NAUHAS8a4eXrd2ch92WO+ilcoXcSTgHZZ4dA7
I4lzpd3rj//6ENoJ3H5aFI2OvcFsZJ+x4AwNRv04N2qP4Ic/nrxnPpLDWzEe5pSG0bg+r5IU3Un3
J7oM9rPKLH4Gx1Gchpm2SSlbpwpHNKAhoL2YwnpKwkUp0a0sdOlQIfjOSj1IPN5IhXt+lKKOZVGE
SJewuaEQ3DGvRte7hfA9syZT1nlkItRLb/wAB6LbsUubxlYF+tD/Zg7fhKgjnGOYwlPkrm8WC+jq
z1Bk6vPZfxITJfLftu08KmcjgD+bkATCQzQt0lDs/FT2GldqYfTMlak9zulPmX1wW5fWn8meYZdo
86+VYppqQEIh6kisjzGaKcgVyhzf67k1gWsEZbUXlHykmtwpMOHAzAKHDvqOgamNALGFDkqz0Y0F
IXE8lp32sx9pNkGoSO9c7iBn3Wh4fRdHiiYP+BkQLYTJRMOg8xuTR6vFzCXQ6LjGBqzMaaRUQtNB
1arruRK9jt3eBntqEVVL9IikUATd7IWT3br5Gpe6AHt5UoYLkZRJLttXfLRt+wXhPNROjIGHso18
jhg3zdvePM3WTkFOaneU8wMnWDsC6NOycquS8HxKW6aoA/0wPnu5xjWGZQpMjrlrUwkp977WYDll
u//Dl5LsdWIZ3og7Nk6UncdWqta7vBjfRu6Pcy892rj884fWHeWct8PRGHfLAkZkmcPcZ9obKe9H
QX7jOTRyW4yWU/LkhxvohLafRdGE14bEYgzE4MyibsG2t9D4cY9bXgMn92CxHyd2Vz7yDySieBA6
Ur6KMYqRVv2f/+0Gcedeh7W9y2jQrJ5CEU85oH/eVO9A3aLwKAF4dS9U+WeRjP/eSxHPCpCDA+GJ
H7NVQzFvP8mY0mlIa0Ea8Chnz7Mv41TD9HcevsoGIUaxtTeCFQ3GCwI/skCORoy/jt22ABD0MKKa
1d3fA1fZdVl7MkdZmEqLBHz7u03U5c5OTT9N7w0c+t7oQR1nt95jI+dfHKooCHXEOlw2Z4yAk9J5
ag4mhcCQJ7K2MUkqvV9rx20Q0s9M1RuqEoB8HWwbIqv8P4DdwPZ/kYZah4oWltZ6oopgn0pNsSQB
Dqmaio25IBFyYc1JcrkcIY+1QlEhGpoR2r/BOrVqn35ha5d/Ch7PG3Iiny9s3rdJF1qVY+aCYMSK
39mmO0tXbO2en+VVWerCGZGpMkvh5Cgwxpk2DyIcV80f8mZjkQfyXiNmun4Nd5q7jruoHUkNTt09
cv/G+AN8mnIYPDTf/qXaeDwvM1rUXBX1f+E9CF7ZCgYFa6ii4Y0dCPMXqpi+Jr+JcFrUT0wOpA09
4f86lAh5bexZVrTTjAOZUyuiXPUI+L3TiB5m5OYgekuhXmFtDtJzddPUnmToTFzbqr+1D/dbgJmZ
bMSK7lbfC6ryyyo0a+ZmZwXznw6lRY8F9Tkvc8DRBuNzIt1vN4M1ul9/N9mdPEcIdLDB4R/Gx2Fr
6xsnKFNVeytzZk+QaSymZcTWzLmwQ3RVAsd/S8KtrzVQTZJlwvhVnjRrsbGPyVw8fntyzd5WhEk+
CNlYQrmkjQdlj0k9unOMEbYkQRrT0ksdrhkt/hr1I+3IovH5uTZJBzGPt79n4YZEomsJ87i8F4Pk
kbCdmIvlfpWTUqYRN4bTseuc+F+yVKz99vPwPAO0YpRCF2QaWSirjnWU9YAlqA8ed2dxoMfSqXLq
12H/m0cwY4hV1zDaZ6lHRzwLEzRn6MIah3LRAh23zsoBJyNj45rPsxaYadrMODj9U/nEmvMuY3Hc
+iFJAXzHNY7etztzHGrifBlKvOqNR/bOb/SCZDoqYxjAIcqs8ntIFDIdd1lGmBpKcGIIPqDZd3jk
2bDxeZxAH1oBd88T56bSDOx9uihOQJ7ty/2ulLugm6O7gJ6o97byD2FY2vhEZ2dF6/3y9SaYd6Z9
nFlokqScpSC3R/Z2lFgiwi+KMO45V1jJ6BEGGtYcRQPDCh0gIaqrJe4eQKOpp7jCJv20d/GbHUeC
9cOKDvmmQoprc+hM/aQdLwk7eeKKVlP+GdnI8Lw7gkMuvcrwlQQudSRO9tbKykvdj/15y673NDBO
MObN9cBIvYfwew+wlx9w/2mfgKIRW7+zo19Y6kZZJrhOeftwKJvomp2Z6Uq7Z1X9gSUFvsxZaim3
C8KrPYexjFt2TmRP95VXe1EgHoDKF6KvceXUuVoSYYn87lLMCZAHga9srtH/S0yqw5/iUracaMXY
EspXYJcZ0eRO82/HF+p1Ya8uSZrNw8jHHQa/5jc7/GCC8el7BeMPG9gThEol2CTW4nA0ljcmV1KQ
8ZWMlcWjpjCkWKr392nlsZjXFY+Qik1zRQAtaGf8ugszS92ijRgkzMzSBz0gNzc/QWRFuEoz5Z6q
N1zvzkxx76SUIHyFZkwagFikX09OpbMqy6eJcngpy91I1xj+roBFpHBCihHHWl2SeEGe6jwuHnWF
1h+x9ZZzQNG/ga8mzUkJrqzHLqSlhsRhWlx+YCJfhrunaArJSiMPxg6UGh2znIh4SN1yu70ll5xo
/pQvc9U5xbVnFP86Da9qyfTxPfRSLiikX+yOrj9KM3Yta09j/UNLkuzF046tTBYBRroJVgICMmOJ
c84Fwt2kM5+kP1zvtQRssGKB41kGpQh2sUI47E/+86JgoJWQcKR2XRbsmWxErsiJWwIn+RfBPyhg
xVsBXrtHzOCz/U0NfpvdQ8PzlvA4jNV7DR9Y1+ox7YapIaFRAABXAHq6tl2WpzDrbUxcagKEtJvm
h9xw0PkBs7h2dlzoZWNWluxKSA9Bo1XoI3TBAf7WENvssiKVwBDMwMy6znZDGB1ynHPNWTVqN69I
rAbrfEm3lKsM4BFX7xA6alAqrJI2MS6adihos4Xd0ELy82+sGNl5YM7j/8i/C/pUIShobhm89WHJ
j5nPsLa9DGGsG3rJK8lZER36K0OOD+NJsYxF0vpabUGYRwvh5hSOSSoFyBIncpQKrjvGOUai9U0B
KXSDZTossoyT8iRXN7RdkJtRSZJnoziUX4nIcJ0oW2NRpxV6hAuhHj3pe9aawmHnNQKgqpFObDL/
7Rw/R2lXBaDjr7iLEZoSEM053BIHT5N2CrGCDr91N7/txIGKd34COu6mzjmY4jehMn5e8H1Fs1aG
j+uVSmFmzeZXIsyaE59/CZ6azCjU78JpqecKFgxNAq6AXKCaBhkFBL6pG8WEojs3zZblatH7xhec
oidT8F2Ut6BkiG653LfYD8c80um2QfRXx8hbTB/9U5MDmrIPJ9o9uXeISeNBaJXwh1iwo0JjwXgl
on0OQ9hAA2bEPnKe6WnJp5+Kyt9Dm7G/qt9EDQunJ3sdBitGXHi6qsOEFqEi9dmB3Q6sdhAxnIIw
t+jp/pnPKvySCpnHjGA4ozbnlixfYTMmDm0hijA21uRCgxeVpVo+A46Kllk6s20ZbNPkOAOXyIi1
FXL1xrK8ICMzwKwX4lcm4hqqQUqxfTd75HYkWCqseWl1Q1z0rtHd78Sur0+kz8zDBPqQM028jnCy
eYjLQTRv1ekGOPgtoCM1QbL6Nx1O8gyrHEVrm3Y6qvtg0KBAux8OJumNXMussGSk0w+55wG+/55x
HeaHAFzKELL9I9k0UrYMR+g/T+9t1g2JMGHsSSNb5JYbh2ePTPCyNb1yytLYTALVDAzQHFEkl4Qj
YwjBot2dJbO4e9g994QUHPosVdg480O+P4kjZJnYZw9NuhDY+Vzgz4R3wFUvAAG7k6No0JkZMych
A443itH9DV7D0XUkEmuijak5t1Q8L+vXg3wzbkbagi+taEkjZu9k2WVU405RsBNc/2NzD0opJ64u
i8oithuqkkN1xFnLpqY169F3rA/9McTZ9Iz6LsRw2vAGdyqXZpPOukbx3FhbLlhUjC6BLAMNrO0v
dZUUvOz2935JmKq/yieRtCd1an97eWWOFG0XdoRPuA4YwIrS8IuxwTnxACxh/cC9QMBYGYBJ9Nwe
0dzZzNz29o0pvVhjJrzt6PTIvPa0CvEZ7NLFrt8OA0DQtJnooAuoxhIujqQMzIs+BPdK25RRMuwp
Flp4q3wLjDzIbE4GPL+C4esev3dOZokO0gOj5JpIbtiK/clZvJ2mdA343jBmEDk2q5FN0TWqXIAe
8DwSIiU3Sx1cUeti9lH1rzJTzs3kc1B+rYcAWkbSrvy4ZXTxAjFkdoXbJST7utG0feDsTabmIemr
NS3FqvZ/Wdpp+i3MSgTo9HUeC/Q3z3kF1elTxmyhp7RWJs/i0iD7GfhcFXkqGzgqIVkSsmBJlwDT
kVl14ZOIha2pjT8pfKKr/0YtsgJyZE1N0a4LlfaxUy/nSy1hP1CYPjO5KkLl+MKd5a97iMmJcMTH
cJuU4F76sxpu7mzw7oKeBUTo7IgfbgtZU2ufn1yjGLFlRX6aHFNGsAkRn1ZpFiRJolTiFMqJWusb
7krX4GvwX6sbFUg6zrpBxy0bifUhb1V5aFnJh/VYLzirCoeTFC+uMLESEaoDARg/hcKIa2gCzoqV
cPc04qOdZwaBJt9TVFPtqberBrgyHqIG7IZLNPBKeOwHEMo8QQCVhf/y8BDtvwYM2A6+N8Kf59FC
UUceoYsv32dj21WCMcl9PdXdqV1Pjbh7Ni6sW1piScOOIm8LiFFwApRli6jjoj+qZRXDtL29mAmj
85wa0sMpCakMf/OjN0Wqb4y8Oy7moQf9PxVgsnDBpTeOKKgBLPB+1xqVjkFFhgcR2Sns13DpgwX7
d6oYKIYhJmimVhcG+9p1t/+TEhTQyTCfLyIf7RUHUB+DOw7fBSRIA/r+dQ+FNxnhUWPy5NgQQ1eg
rfswgTrY/hjOfAEhu6QR81pQokE/vGVbEqG5P7Hi6l32VixlMyr7fnr2dtPs4F6biv9nMxCLosox
GkuCZ3TRFnPaBzGJvUTcs2DZ5zyhjBHTqGGwYMjwnxSPAmMoq+ImK2RBjeKQ5ZBJ0K1mYRVutOek
wHoDXpyarp5GAh4kzAsRPkWaxaGc2mnUlQnHqDKBBkhzartA3sDCKBbdkUCTWQgn1QiZNSBZVgYj
TjcTBEl0SZccBWHZNZV5hlenX8U+AtRdYkZD1uEm5/pRBYw1ierWrWu/PBpYJIn+ZG/7rX1MNhFa
aKfYV5Pff1pukrNtXOkS+tEc0T/Bo7oMm8gnK4fT99SM9MhgWo/ee5YGzeJm3t2X0dnombCuZW/q
Gjlw+pVGvunBwvD9UBelymH1BlpfUmLJQ/7g6QYBBOyHQC1HxCZBmtu/0Bt+sAiFGTGBJgw8zko1
akkKuDAe3YF9riVOCG2yex7Ww3KP2NvbgXYx1Rnvrvdp3WFhdFR6HVWQ7JFnMMBjW6qRq3wsDFHP
xRB46ta0bpwHmyHIZapCLMfJ2UplLysxMwCb6qB6VV3pdzP2RWxDJbpum92oL+IPywVdDlln5q0/
vdq1vSgmvmbz+vQMBeHtqVTtqZlMgMxL5UBDYGa88hFXqigEp0blQ2GfCEdMdREKpPvNaaDulWLQ
o/BKDBaOPaIo0BPYYQL8TpA4TxytwiArBaD2z9sjqRwjPuyE6DupxtE9Njgc75QhZxPbqZIJE7nC
Wq9TXIRTPB/BD/Lmgenh63TYIxE5BgjBrR10SFoqpOJ79HrLcowoxu4Ge2aehAeOpfi7cs1Zktqq
iA1N0f5u5cX+7EX7HbRwKGFmGU5LaswrLYhoEDzmpwMUZTQiNOXFVFHiqL1E++hj/GTYZDpVRu0c
WaXVHrHIBveiR7Euwz146dJIBbDlV3nfzOTr5+5RlhX4KiWJkyvyimdUyR8dKDcXoZHadu2MtQFH
RxW4yAOCO2h+oKIpWKdh6misjH3DAOlJ7/BghWBpMYKCsN/fmlCfBfx7NZYit9gCNIuchs6yaVbh
mR8H3K3GiFNJCYy4kUbkO9DWJLsY4xeWMc8Sv94/ZXxjmH6wBXACxes0xILyjD6ttDyTyTvg1TS1
XSvWFTAQ8OCzL+knECCAH5rzq6/aWs6ZZgd8TZbGUTg3l4pc+pPdoQujTI76H9+G4zwa1WxYUDoB
4mJZgnNs/1pOjmfXelA4CyuzTdIF4WP5kULlDA3F1a/Uhz2byHc3kv5sHTbfkDhr6J9odRCmR4Dk
SJpA1X0Q4P3lmaVk3s69COs9QfHmmVoXNqsMkemK6zERAItR/sQ+3zU9wzw9EVEMxq8Q2do06G9h
QPShOf7ZCYWCIyn+JsxNx7g/rg8ylte+nhjPs8ZMUamMuezydA5uuUFZsqGIfI7AvB1ghu5MlGEC
7oXRtbxyLjuOJIUpf9PQYfnh1CpJ7mNwhFq/eQpXswClw6Cvt/ixde1jLGpbGxK/7MLnXClkP6H3
XeRx12OXk37dtkBOSf5LmHMeSTC0/UYWYs0/wFcuYTIMEfykw3STceG00biEhT3/lRadlLydt4qi
HOMO1ELm9/GwRy78EymqcVI0ZCurJMvbmT5xMHj+byST8gBrjkNIEe0DC39Hy6ZOBfqvLqeLUFu8
g8RpC8dSMLSZQxM+NktCFSyxoUDDDKMoJBTMxOIwADqBJYDOpierBcqND2fSp8RDj7KSzIeS2kA2
1+BR3clg/lldr+iazO/OGEW6b7RR8n8D+4BYs8n85in0jwocMJiQDiznYCeK27Na7dROZaqS8xEU
0SKpEnJQLHRU5/saJQYYfZMQgBIDAwPQ3bATANlr92lSVMg18dxy3cXKXSKQ/hnKhJs7vntj/tuh
QAjTOvVv+XE3SOrjREFhhoQLCboma5TfOamo3fmlgUkgjaNbNUSU55QW6NTszsdMqaxeVOTpyg11
I15v+LBhDVSixe2h7aHOA4ALQ7Ae9BV3pYl0n/cj9Nq5pKqbLBmklJ/81aRf5MjW+BcRjjQ9H/K0
PHD/HNKnlLinVVqYPzgtJzYu+biXVGmI4CEA3VuJZA+ctxXknWW53YTCpMY09g2v2GD51ewCDnxE
FGY6xlWCMZ5uLgXiYl6SWUkyp5qEmKasy0WK77kBIHjRvV1hYdNRemWuYLgEfVQMulaw1RCZMgSS
3ZesCVViqdAdpfdwzG4aBOn51g+tlzrS6PHXBcVyuvK7GWsfMiH5qOdiLRPps5Xi32aGsGekiW44
iuXM8rb45F+gOTgFs/loWTDAMuTkNifs8hlr68EJ7A/Hmvr1fNnJUcMmvlzAtC2+QvzJ/bqWpfgY
SySz19GeUWJpAU51/O57qU/iJkXUnUb83tEITvsON/2VmudsAEJ+c836gskpLYmvyg1X4D6RIhjy
kFIm1P7jl3yAUG57elrxGHpFcx9a1xYzfc6MiIBWcBLB7ZTMm5P3axg4EwWOTSaY4Je6Cl2RzwDF
qggtURSN3gCCVKbhsu5pmeC5PVkoFQqmTtihCkVdrlZhEjIS0fyYAiLIsFvF6E9bYd3tPQVyv1Mz
nNtSmyrLrDdYdWq9RxlKvn/smvLz+A5DktnuicVmXsagttLjlH8RFi3u0GzvpNhgT1CfNL35ElfW
mJavjEmTqcPdHDn64cv6kK2Ap+dT5/P1vbduaiIj5xGTcpTMp0EpTHMAnjwMPY4VSLeLssSU2ax/
swC/UGQcPsRvbIOYzuXS6FOxLSOBzgF+QQuzAJqQcxrQMgVmJYgGIMRNyAnxb2elo9mOUT8uA1rL
Mc373CngB766LrgaAG97abbIZXhU91iMMBaG5/uXSwG1M17pw58d5uAI8fbGzDHqiZ1TqUlfpAi3
oqnPgeLxgBADmTpk/gOAd6HuOlpigFK/VKXbFNVx7NWdG2vBfpSe0wJfVUeqeeN629+PxRayk0Us
ksKpGzXt8wEN96N3PtdzRKXINlLBKMXeD5uhB9WImS36YmWr3VuKqgGdgUEdwJVIp+HEWBvDPDJM
PU73AEIbehsXuML761ZfXB7wNxFuZsm7iQkBr8DBQyKZllD+YAngdLjOWBVa+BmPLafw+Yrvhr5J
9K9ynWQhVs6LiuiNCRHWcWhjrg5ceJJmIHUtjQs1R4hwFhjhB9UYywQqNWGEDsyZqoMvP0WXNgqk
wOuG/yxXAiv+1K5w1WgSI+lIQs4dwnOK/WGr37x7fJ9PMgfNF5z+iidS7j5OqpfAICFA7ys8AvVL
JR8NcBTz5hMXphfaBka8FmAu27/JnJ1mDdbk8hnUABX1bJG5KsshnDN/XEbc3zesQdpkKkilxqpz
IO+cgK6xUWzpaDulPrgHmkpZqXz7i1V432mTm+IIvgKvfwWRDS0Q/yaQbSbxKkTgI6/piy84KRK5
2a4xs0ORutYTtR0tMCaihCEEpw+IJHK7MXnuGSTGtcAp1HgzINdSiFQMe1BaUtBki9GmvYURa9YK
+OKt4QeSh/tx7qzOLtK1ffLUIlIPQYI6vqrToQ9rSCdMMcBtNXmOQr8j4s8vURAA+ogneigOkRCx
xBMRVbEOTGT1jkSt8Ky4gyueDGeY7mOZt4TCnwYCKgkJ7YmQj4CHGNl6K7fjEJbnpI0yvLQg2ff7
1q0HBdVFcrU5PAKq50mxGMP39HnAnUStKxCtGbIrs3TznD6RWwXUZGpBrUlFbmd+YiN3Hu6LpyOi
BzABeBiYny9nO7J7TAg9d1KereQ+BG1frXf4oqBqFA/iTC7nnd+0DthRy+2lOLOzDmpIPa3TfBU0
h40EfJ3ndcXOjHde+Lmmagm4SW8DPFxjY8loAsYUlNVStlMOL0HhAHnGUO4RWKUTZIfaakfIHq0j
i9PBdp0EAbBEGB/xzbpUg5OVp2k//cjEd5IORZVPq9PQpSqWvWWwpfza4CoAlMhbpSIHDYcf0dYY
pnLtmNNT9Dxn0Sev5EKOcZasH8mD7BgOS/k3F6RClSmbeJuamVHc70ptkvuhPsCpdZC3CBIhxf4v
IdL0N7bF/UFlpGOS0ecyUBJLQP44h3PDSS7WesyEXjSNx/XB9flewCxTtgZIMauofbcuDpg3NZaw
5s8IR0bnR1X3FtjtlX1wIo4HElXyAj0CIljBySpWcBU8XdE4w8dAW+viFC/CluWpsIgPxVfmZN4W
mJ2XR9ImvV7399FfoFCvxriQFs9wcpZvMaZodwvD1UrvUTw46bAa2Y6oyXOX8To7YnE0ylQzJCUD
0Z1GgBjN+hfjXLuFYi8G+sFjKfuhGhNEmzUSxM0MCC0WdzItNTLYiSK9AsJVLHqtcauJ05dwCJe7
A6AcxYSji12O+gvp8n9TWhJvUZqWjDYvU0x7MwM9iJIEIA2De3bbg2NqYOipo6FU2zc5Yf1+HY+y
eUo3KOLsYwjG0PLL2nxrTpvqJkZxJs2wwqZEIxoZcOSmTnbNgS5cue3c26yWNWmuHZtyBqOfJfYZ
nwuAEDgbpqiSLqNsdA/175evE4noZps4ijdK3VH6jG3ZWFru8mabhroLxSaEbYaPr/El1cVRww1B
L+QnPSj5ISk30UQ1/sIjZzXxmq03hG6y1YdUS5JRn3auEdBbhy+bLobfGsF2Ylzhvk9RNKbsBGRt
4FI41wqIcQoMPgNE9xEu2Nlzu2iWbYGxQ/4fH5IFZo1flFpVasOkGnbyL6J9gOOVtYNiyysrsq05
gEyPt3Q8XEY6Zov2ARRTyjSSZ5tad838PUd6V07w28QW5S+F3B4/4en0Ja+5eTHMHdfR5vWGCS8a
m9+kOdLGqRoZPt5LakWH8Uw0iv2aGlhlPgbMA1VoIXgM0HgS0REtIn8ZY4STVJUW7sSemzEM9AB5
OVyor9v5TCjgDZiZelX3bDnCjG4+O/qG1xhsG5c00qI/OGnMbeaxUyczZKEjmUSXa0Kzli1KUCTR
URn99W0Hn+xOs4TVp836QQH5mDt49ILU5CSdlKxILt/WYKBgYquPAAbSXoc+OJwTaPU/NuBt63Y2
ttusu8m/o8ARCGidG6Z2jZE7oYwgkG7LOdF5Rg0mI3yVvqWpLKB8iKDHfYaNGRe8t1qMY8PlI7EG
dPiMSqUzwTbYhKaFPcrhIPlhfuVRMATOg6mh/6dtFRdFBN6WZ3/erqxeI2tqcfZLpTGAmyhMjBQV
5CfJxUgA51ml/ePqRObJeG/9m3IIh0FgMwFimi966Nqd+lvAX+i3x7xlFzMmEFlMPXbLvbnFYNlP
2bNJcaLAMMhitK9vFe+vBzNcL73jbi4rxOND67zu/suOhG82fe+/CfJKAyQytVJVZ5XNBBi+o+FK
DBmp1JqF6xojc/7xV6FCT4YKESqWpgT45BGGTw7eFJlGWskWb82GYlaYW2dFnbF/pQ1KMspJoL+g
RqsEkyCFAcX9jazQRDV6bT3/7YbQ4n9yAb+cMTozP7qR2mAKuP9uyOcGW2dCrwvrhNHfm6aMS/qQ
3tFdyUrEfZC7vG7YsXlPh5N4ra4xIM6D4yr3qwtWSs5pfOIbo/9pT0B96GSJ8YZOt/BDEysRk5zT
fN348eFondDsAlJG/lguP4Znxf5mJ7EcLauUlwm6VH8CH7q3YNQqR1xHVTM+jn7BbIhSmDm1eXro
DF3rQIyHAM1gu3BfPdBYJ68jAi5qw9UjMhl1JPviGCUfN6R7tSeC1TVMVeNlk4hUQDlZNoIAOwzZ
a3wPT1c+ym2idaeEXhAYzOYIoCybP41lpFuSzUxzrrhN+b7FklhsM0mPHo3EjGdD/s4NWIvBGrhg
mBS7HZfHryGYZl9pWxBpVy5NJrbdw1pP3fLepKjsuXAG5ZaZDwNCXDW1YBpHrJMktlwc3Ecb5ExZ
woQQ4lwucAumSJ8paVFQc+wykme6ieSbDtdUiGVHj7sMX1Prkz825OT5rOPU1RO4IMZAQfNCl7hy
8I7CQIlsNbXqpOC7kyvPCqt028nTVGzgkT+tiEUozRkL89tJG1XgVOWpr9yLdCVnUS9IJ2Ss33U+
b/iUvzqYB9HYgDickU0nUFLAIiwVkbLzFU0eHz3x6nIVZhQmUtKZte7R2rPNJGGgKJmskkR33plG
4UpjnVvBUhOM4L0mka+9Fmy6W0A+y1PBJtmfvPdt+zoueOMolCllmBcsI/AStVkhTLybhwVTS5nU
tp+U2WgXtmO9NscKJOuFM2IqgQy2hZM4llgZDt68bCFoW1iB9/jUN+Qdxu85YYlCZRwEgkXtifUV
vSbd6XFZ0fRlW5stvMy4XqpY62tgbLYrrQCztU+jBX1epIZrk9LxyGIcckeY8y+YtNEBRg5qZERp
Wscc7AcN9pClATH8QapJCzmiN7s/Lfg4d8KqX4mWq5IBPxBn8ShDceF6275UdndpvTKUDLchS5Eq
Gm/GISdDa4Jnx2alMvSZlTzFq0OHKScFtoyX/b8Ae6LPLTJXnP+wqWZsoDW5g1WO9AmxsRVWN3Aq
4hoB+xx1HnDRnQcpR149PJjgXVXspb6MHUpyOb24mqscBBS62d7MWgL6zPhUGDWpBm8WIlz6lXzR
Hebs4C66vghkXx/UCzcTOY75VwNeaCcKSaXwOPNoM3M4lDYpxmRvicNhfRuB2tRCkmYlUMPLK+EC
9C6t5MPZCnVcVxvCjaO53v8oX8vMR+FPDFis6u7l7wsoJVb7bImt4P8jl2HBowY5u9xukgEOXr5s
rJorVl908AknRkiK7oyNDprwZSKHEb8Pn57ZEx2+fUjCTPoeOMucJ+jrSEvLfvin5rUpbv+1tzPF
rPMXpQWlsVjNUD+kMQDlf9fGWgLWzWtqarAl4TZ7Tdsrnwwf2zvhupzZbxWe8uANHZHtKH+72nt/
ItyKuQBFpm+k3H/hdKkJmCnlSGTbdL430rbufdlBa7GiYz+lFm4bIqRQrZ0ogIeVdelu4uENUja1
rxWweu7vJzsgVvLOjLJHIs+Ez1pfeqQ4ylawE5XKPRhViK0qlDwGJ+EjqVHo8hLVv1mXEH/cE8jJ
vyEHvUe8v0uBxPdUg73ucQWiNAvBvsy0TmQwtKP8/5fHe/tbPWeUDBM5bZvOtE0fUuPEGOM5/Mt+
P/i8n30RdESNMUyGHK1dpYDZ+n6xUNXWd6zLJjZ1h70EwapqcIsKSXmfI1Jz8i97bt/W7bA+gODy
7kJDwUQviuJ+K2zQvq7Ry5P4QYRMaOL8lrR46COlV+sDeQ+BD3M+g8S/rdJAyX8UyRBkv+yuORHS
HGDFjAjpLln4ASqpUgb1VBfMKfRjBDqRaFUVCgphKzqaZaR2UurjwZq/tTEBT0IDUP+YwrYfryl3
jvkStyWSz65nt75JgqZw3iXjxRI11CxiC5bfROyHJzG5QHxWEwLpvVuo6rxlQRXvNRKYWYJFgGUn
AJ9bXKHRc5y7KtG+CAMe0qCCdsGVbkyoicfglV7qV58OIxVZYGfNl8nBURYrwjMKpWloZAsIBhYG
HIewr5DNAiXpHR2YeenOcmvRcDWJOPsX93Rk8fZ9PyLBIvCwnSkJVMSiBXYs/5cD0KuwYZ6Wn2ZM
8DK5md7QBGPJCTSe7RhPQFllJasoHThxn+h/SpAY/4qNNYqZqGMsoa7zQ2io8BI7PQLONLP2VIzk
LU7kjF1zuiJ9NLkKAy9Qtfbu+4uJMeqQ8qs9mNEv3qZdBH8DFtYBQqGjtgEP4TVPF3Ovxvt+Js8E
cMzL/e4Y3ZHHyDACY4v566j7j7yIaakTkArl7GtXc49uwWU+/RX9qno9xysq+bzgseyJtm5t2jMx
eVhCAMjGNWN1FlA+kEQhsoQw2+WxWPiRj4HJsgd6fmAna5J2/NGS0LdFq2E4bWvm3eDxD2PmH9NS
BY1IfbyTfOobElAcq5b5fMPgdiLJlkylsftTuRuYXHvXa77rAg8DhFZ5ZMSIfzgs8Gu9h9enRxRe
r8u34NYCjwEXtQ4LRZATObMOfRdufi+cbKvDSzQ46QiixKH32ZuTdVVSkPgZCpQvP7hp55ZbB7FN
cGkqNPXFingvah3VFweBWCqtW0HTDHsVgDiG5WBuiW0++R1C3BAxmwV2WGtxjHGCNTj6ujun6kdm
XrmXTzoVG7VNozg9N58nKn2A9fPDgsTlNHOoJaIAhRL4fs3uKilLq0OK7TyD0Hs5HhDVsgLcBbOM
tfZ04cWrUbdyjjwrU5s82Jh8+MprIryFHepsT4SfLUrcmgrv8UUVXfQeLpCMS3E7Q0usGt1Qi5bh
xKcpfiV4vN/wHRPBNi6Tc0hqz/xHYIrXCFnOB+kmPYFWHDHMmAtl6KKf5VoK7FzPo8b0pR8kwEfM
hKtO9/M5QyGB7gNP7FWVkXQI6isR4amPsQuYli8vDp+vOPab6PDdYKKFwAbEx4LLfubyBH8tvCJ3
UBgFQtamHv0WaQ0jTILvpUS8SOHIT0S4wznDTM4VNocwH6TNvZ+W2kcMFMHd+Vh0gRZPV4cgHXma
1aDhtgjNrp4ibZdlc3Z+zkO+e417l5qT7BdSvcKDWP9TVR4adXff5IEyzx5WS+tqdR+UCJCbhr8u
rbTx5v0vNDWg8dpo3W0HJig90bBiCBZ+1Mb3208xl3a3olUFoo24a5UIId8OLNquilww362rZb1A
ny3at7JnMCKKgt3v7e8sKrLzn1J2t9DmJcKJy9BKJceV000A1HvaNI4zbOV+8kmK6oiORVcScfxT
S0pnHPOv21WWzgk1U6eiTwoVb7Vq0ZJW++zEeiaNUhkrWdatWe6KIbfC1Ca14BAzO5DfYb/8JdeL
qGNOWrjnD2vwZvqgndgMrlJENfpRUEHtADV62VpWlpkr+vHKSgRIjmulpOIoa0h3xTEq1x/5dJpW
XO/B7xxWgbMomvVKnWydvoY8rawaPeSLh6IY3mT1967sXineWG0MWFsNrrkr7PuqlusBeElyqxM9
d0Bgs/CPi4ncBhQTA0aU5V80j2TjAClC4gAZTEdkpTkotiCMaYSjLmoMrmjH0D1249if5FRNppmL
HbLATaaLUYrwZdsruZGGwsi8eOyKkUE+G+7tiv2/2cwLBMwzXigvj8lhWZFoLvPzSOCnbl2V9kyx
5bNf2HjZWHBv8BSN7ithRfwe8Aa20v9hq9Nn3R8HD1Aq8EWLz/F29Ci0dZmgWFsVibIWBUGMHhFN
cn2gc8SfL/z1LhmaTO0srR+FoAj7eQ/YcbXW8gjVxq4cHIKxnlbGJNmhDkbOZ9INLEVqVB50ofWK
96omZep52T4sVsaKYpTvWow9+euhErkQEB4IMOvb8dg/o3sqCa83qssnfgM6OE91pEAOwbC374af
jGpk0+RvRB4tsZjCjMnYcyrg+t6GGEd/2fKOqub1SdoRSyTZk1Xgx2vIawzJ6W9nO9OHRuvgthpJ
D0iLJOeV37nlljWhAKi70/UB7KtI/Rpce5QcLSg3qFIIsRyaR2ghfYf9vhKVj/9WwcY4QADk0eJn
TJn964Ezr8DDssja+DUeK1Rr//wUVDpsjg2nqAgE9LuOudq0YJvEOhYXZRtwpuAedjmWVoUmusrm
rFLlr7182AOMNPB/oBMe259vEaDWNa6xgUUIWw51v0qfC0ywFfq/WDWZvh+427HxtJhvqrta5sSq
nZpq4CEgzsKkthi6DZluGS89JBxvhVg3vNOqFeV473UrGhS6/cfrgOuh7mjw+ngEeFcAks4IEBv7
TYyQORvlZ4Prq9PUrPs11PTWuGSP1x4FTMQntEeatlhs/qdLrUP8XJdF93aIMsD2Qr/50jdsdgi+
89YbdrPUhRxg0VBSy/2zzPWBolpvo2gwLjtUWmtGTsk7PGId1pjjpYEyFpLXQ60cw4HSbGOQ9VMt
tYLZnAP01RJwhT+B2vE58LzUVvQqaiZdF28o1GDeJ6ZlIu3hPHd73AbCCAfiAdyFcdmg6nnLP28Z
zT+fQsMHEO9fHfuavzbTXY9Obs17ybZnlnxU9ZWTJYgU1OIGMNZMoYplYnpyac4mpwSsjJGoOvEN
YBwJl4CYe7Q6mmDRnvFLVwVNFST0jXRx4L+ptGo0ujjxSdpD0W5T4mIUoLd6cgfm+IjPeB0lvpKY
UsuhJHak53a1Lgvs+WZEMawxVvZNo6gz1QEa4IMU2akIkJen+I48YrqKlgU7SLarrICEe5j/+QDx
YUgtKqHquAU11IEv0Zle4JrG7nmWoCaGtXZVlSn47jS5GgeHgd2aod9L8liv/BSLI3i2ZWSnOI8F
EYIWb38SNziQxBoLz9/B16rM3iUf4TnArcBh8HQ6glrbxDggPMdqD9O3CG57d6sIyz7iJ9qBCupH
11gYt2phW/IcMmOi6uAV489rhXmVwvzSFxXPqaFCEaH6ykUmeCMnZgrw5Jlyy3n4rIgnh4/PkV4B
36gThFyM46WSQ6VM2YAhRNcpPLW5cFvHAye2zwl1RuPkXk9O9M2OVa9g/d00GdJb/tiWvGlfJCcb
DtnR9dPgwwCzAPNPZO0wAyCjtXEBTW3ILrk7F4DjzKYUOhcvNHVzM4xRW7F7rTjAY750VV+CMTtY
SCU8oGKr/EdAFlBf8m/jp1K8LG5CVih+Ty/qBWwDw8nGMq6NnFNBdequPfpRAhUZtcy2moBrO1d8
bMPs3j0nJNoHH3JKKGG5kZok1KOolejjmd5GjpYoEGHzEEUZhVz2MiIotUbG5MwjdmftLi4mZbhy
OCWebdcrUynmWcpO1KXW0qpFzz8jK944ZMtkhMyR6F7oqHCB3J1CONXcgCK7J/wSWeDbtmQV+hS0
alJHHzxD1pxwiRvJ/y00NP35gCuzB/8oyjtMd+BNN/2/o9rLcf8xbd1VNrZTfNrQBymCgY8zSBpm
B76LbZsid9dpfMnWxNsKAd1ZO867QahKyP/YC93s9IqsOyt/VUI7MWZYuCztkUJqzOwDBnEVF0Ol
OyaDVwFUpKEcvSPWPPw7myrJxTuEdK5lEY86KFeMzRRc1E7VFKujjN6GY/k/LKFYfEqErbu4Moq4
0ZW8xN9SyqNyWZi51+49SjxDNZKwZ7foeuMQ5Ns6rkfMw77pB+qpXGWDhvO1nEkV/oHEWZCHCWKX
kcLNNnyVEzPxIWNDtqTCXg5O49onRKDw9ODoCbwQv/9jtQq2ycz+lBV4ZBOeQPAr3ydCs1cPsqnE
IqbKADQs+mygRy38Rq+zNqyY6qnrBqk7X7na649lS5zIuSdziQj5B52w5piwyk5VtvLKd6IQlPfZ
dRJ5OJTOIG1YJ7MZq0//FCcmQdzGGXAo2liqJrneLVCUJVvW930wqUZCtkvMi50uT6e7PnHjFu0r
JOPk90PWIokgv6AVIeznQN7yw5nSZT3ykLlOFRdRv4jy9Pu/R375XQyy3F+wq0hxBH0+InS61g4l
l9subHJjDvp5y/2hJ4qbcDwI2kXvOpRPj+BBr52yeEa7JEOb26g3zZkOVtDmNzR12iBOMadeAXzb
BG6RSkEyBnC5cTQid7gIIGNiAjHDRoV46df2+bYXHqX021vKcfYCbMVZufMXWclUPq3p03UQWORQ
rr3hZv5afgzcWRSodiVTtdrRJirQi82SVskto7ehf6HUVqF6PcYXORpXIOsfCJiiHKHVM+74CqFo
8S+cMt0+C3msZKMuPxwmJpilaw1QlrfJl5kHOrFNn/7+EH+j6qiDmTqSfJNpLSPdsmpP8e0Vd/wR
mIxc4eJTEf0070osmdfk8pb8F0aRUDSEs+mJDJqhw6Z+/syXuA2Djlf7JFKrGBMPSmvzT1nRLRe6
fMpzFkiZQHgyGk76J4uIlBsUI0ZPu2vmgrTJcHVcXzsjF1fp5FFpMW3FXmG1u5ytTWInaPHc2/95
pTc7rAcDZ0rws1ZIlQDNCGCzIXFHd2Iwz/RMIIrB/yQVb76ON59107YqxvjqD5QubgVzQTQnLC1J
Ky0yTxVKo5+JeQJvSuAHVSeotGf67TKEn1+AauOw3WQchsHPBu3W+FO75qh5t/z4dpTv+f73Y7eI
PYi9ifRW4atYafaMgWE0+KRm7zLY/C5MdE308T0LvUJSQ1Wd2TRbpb9CpcZJIo0VB1xkYOy8uBiH
RnXXJxUVB89tIE61y6vmlx+Wp2nPQkHxL7jVtS4MCIaMsiV6yGJAoY9JxJMquBGsSBxAM331eKqI
+lOUxqwv7+wXWPk5XFfbhYHs8ixY9a1+DwXJOcSSZO27EJI7gpxsOf6bSvHQOCY4UMqlmyDUQlm9
QSH1Sjt9pWp3Vx3Ch3KHd2/EOKzDATIQyifQ0HpnKiUFC33Ria3Qmh61nYzH/SrZkn1GiKKwVhG9
SWVXZLLaWc1npWjBzC3W08zIF66pYdVp0EnuQyurT2Z/ZYIjW2TsguFINx0zs934JZ0RKpwhtXul
yooZnpsUvJdgXIQMk/p3Apx4Dh+3KKLnig0WbsHpA3FsYBhbEiR2xQZMMh92LpFcyR4F75IRoCPo
PegRRsb45X301tG3qywC+aNZEkNU8A8Osn6KgWz/a00w6Poha6eSlxKx7kAUTtZGYjk31uoDPnEe
8paeSFnfisBr4fKYLwuVYz3dt/JjrrNsXdUYHjO0rqa2FoG9jvUXU8hgnsYLe3NZ83pF4eddDNhM
Rx6Nl10BZWfgoNVcw92yzDA6NWnc/XBMg6f5DSvM12VP2o8q71DE/5IabhSqJQr68QbIVKGjMFU7
7VIDkaSeNJVRjKQQXXeB4PUlDVvFoc+yYGleoMZ3fz/J9JVvKOJVwjpXr/AQ34odP2TDFHrOZQ+L
86QKLpA5cyVXHIDOdLNcK2FeG5K908WtfmG+K4u7s5VlxRuF0PiCNsO0xzkTTo7w82Qzry8Tq9pB
SQ41BgxfcBVK/gydJgFLaq0r5T5cR/1KYkBnBSGeqN758HOfEI9KngxsfdV7nW4RxMbiQmvKiktC
w+yun9d9rHpYhWrufJrSHGe+SOthb/5kf2FqiVcITtaBnnKgAh/cqBMk78Gxn7FVNvhYUl5UdVOv
EodjP8CkBV7Kd1/geyYhStlJhyfiN/PyNntkTlJGuwEFSRW1pex+6IVOilqWBh+dvT0J8wr+Pdlb
CPYY5bBz/PO1JDCTIpiIeu6DX9qtz3BRuSbapkOeYSc3e3ohd7qxvhWFY+gYrN54msHY96143bpQ
UrHDylYaX6omV70xAHtIZkRXw2d9klBzNhYNp2mHiyx9IGWmMSj/rmjT2FUEHlk9l/bwt1CHlzct
DyxIU3r0jgpOsvCQwS7FyZAHSqp4rO0B3Dxe3wMxHz6SYjSbUcl+CS6qmc5tGu8p0hnI3F4Tmawc
rXK9nRs5gLkV9xq/JrjSM1dF+B7yg7JZ5koP6Z5k8uzPhDjOCd2eEzFM+deWRdozG0pOZGIUDTIu
uL+S0eKSQLDszi7PRbG3sQpJpnDz6df0q/3k0J+heHYSWwbUtrvEdC/ydM6bZJ/WIcYKNHprM4Zg
LyTMIxY8KXiz55okTLUd3dxi8LvnVHUPbEg2ES55PlQNq0K+N06WaPLYPNyeBiox5KUQoPse/9qR
EerrzrBtAhI4V3vo+oibe9Z8wRXMwXTOUwFnBwO0C+srSXNTaVpKYcOPu2uX8EmU2FYLp4oIvD8x
bJNjUCMMLht426o2W0LCpMIvdivJLL08UNxTbvzJlhObn0l7UPkUjrGW+JMlv7PpZWCy79gRLv0S
Ce4PjHcUrQjknA8Aq33boumbljtfnBq5ve+4QIKhmd/FCtHFvrpJoqKR4Zdc7uufzEXHApRXBBLe
iy/q86MXtiaPF3dwexodZDCMQ33eKxJYnDMnSSM+3t2eAeoPlHflBEv6xWnLsxpVSHewUBQGoF5W
VbuRpn0NOLtKRHfvSd6ffTdNr/ilADIA8J3C5KKSQqgieMjTH1k9k4qFS2cAvTJYD+YSzZwxraYw
ooSA4JPA+cTsc00jHdRPfLDF45iVC2T8WoAtDmOnCE4DRtg1XMGx3bwkqtf/hh18a40RmOr5uvfc
+2+ZZ0LxFQVjEFYtNBUZTdQ7HoYToRbXZ6JJEp5DEZKNegQwLIhr5eOgnnrwwBAwtz+knF9IhzDO
APSeETpjkeXS9PG0vTMLWv8JA5x27z5XorFhnF6MZd/xOFQ4utdNXLB4l/ZG7ie+xrHs5ptYzFzw
cJ7hDTSytH63mX5cKMRGeeCj63gnff7V512MkobjsVuEJ8nXBpCrMReATqmUG6Z1vxhS5NpSGLAM
UNRjqQOupq9/jG762N50R9qy9XbDWzHLpwHO0ue70Ls/b0B61ISyP2wyPeD5vX2ccbU2qMaLncJS
TmP8m559UI/lU2Ch30Qi/O0dz/aNUDWpRbLzWKTpbWxQg5htS0vZWp7jjxMlWae5/GoBmVeIeweD
ERrkxw4Yeo/dXUyvxWow5j8Zv4gQaxCziRE/SEkP/LTxzauxmPBw/d8XEyuFm63+JMZuu9fP8iJN
Yza6SQ2aBSQnR4kfj+sTEOp4mfWAwRb3Bp28laa+sAU2mYpdxxD+HO4PORONzJvbOxMRryN7cF4u
ubYR1lDT6uVenMUCMa3YZEkJjhkQfo9wHDRGXnjr/2xBm1mNY8NBGsnKCn275fWW12k7V7ITynLS
V6bbNqAQMkRKO+SzgNKOC2VBYSpWi/kCIkVUdo02cGSOqO1ufRlMkNaTjfBDvOfBbDLf9hTG5npu
l6wuW+uiOiTurIcT4bSXKlRxc6XTkYGzw60L45w9jFzjSGdlgcAFn6I7S6qvpwyyqfhhHAaLTqxK
rRKdPmGwq6bVI6v/OTKmyOYB7GVRA/yP5dQeRVQSK3e+NnzcbTQvHRcEWExSQh8LKdq1Nl6bEa3a
fHIBjOQFzXqxsL2P4LNGdo0YLTl9gOWCdIRgzbLI5XLPDsxIfPRUJ1EiA3izld+fm3pdbtkY30fl
EyD7MTaYvZzh9JORtDyP8V0Ax0KiEJ5fiSzaHspoLQAGpwiPCHS8fkmr5Bb74Q+eEtevBvHcc5iW
dOU/ESQKQemAoiuPfn2vYQXlt7/Nlw76pYek7vEmaPK3BPOGmtgTcMXcDRznuW7R9KYSGfSmm3jW
wgTD2Gw1vqPnashjn5zXvlo7pz6qyYWJ+TDOR8NzRbDyCTotoTzDFcpvxqsXGWm+aQOdXQBQQawV
TqbzDG5mJ6MtI1oEtHzx+axe0buIOpweJ7s8xkZgNSiw4Z0fyZ27KI8fpvqQmw9a7gWrcmbfJ1wT
fUW5/RB7JgkARpFMIKsdKSu4p+5UfpmShxZb4QQf+WoGUlE7nlEtuwSCZs/pcPCK/Yqhxr8ppEL2
lgPvakqq01O8wOPUIn5vkGFTkRLvGYg5yjVY0CcNi+IOGzWVjhq3m7p12N8lZCC80HWwjzh/vWWr
dEImd8UGxD0DxG4ujDhSZjBM5W/6R3RqZfmeFG5rQ3ZBrCXzUEUIOTqEnCVu9hEVkaEp9lhsXRRI
tGG99aIbPRof21WsxsgUQTOrBa/wPUXPSNK/bHQidE1wuNCwxVSWbrVr1+Kc9wBBOOPCrXCqRC6+
CjVEpwQxmijgTGtrbbp9sVFfsntOiiwTkP61ihQi1BI984XG7tZQofHt7AFQrCP4i0ZfVVRRRIx2
RYV6Si4+0ifXB/B6lLF4Lcw808h8ikYBV+pV6h9EhaMm4AvczUG+wATqWzVbIqjnJwWaMDrEBYAm
DikFVpfnA/AIqNrNzC+9xNPhkRwu98RY7Q+GuPY3939Wsj/GsIUFq/Laxze2SMzYnc7RsCHCeFRv
qSohvN61Js63CyMm7kLOJs6KqsfDr3AZG/+VoRXMJ4/QfPE3+RuZNurYdGGo9PsW+M8eBD2YkIE2
fuWPdDQy8HTgjmQRCZw4VnAVO8CF/BP4sltothDpwLS5clJwADbx7LpfQ6Gib0wTRu/cUBYoqPep
kTy+D8F65UZIJRxiDlv0Mg0qavs+fPsTYRouan8t8uC9yiB22Eobx5u4UVyN9LtgAhVuI7zj+owz
XHETOjfO6LYlLg+ynS/gJ+sIODyS5Q31nwa3fSA4Tw13fsEj2cv0RLkyW2+n4H38VELgvZI7J/Fm
hCvHUgCIue8eUapRWpbaZ9sxRPW85TURctaye55o1A6YHObDdJmYewGBz2koWlyrq5wmsELxkzkw
Q/T7nTKAHzRN7yTxPRbFWA5PeMsCAmvB033DY3Ac/XhnYxW7Gnbo1ZPArcB5QevJ9dj0eJrCHqjJ
9KU3/740M1oJZjyQNa2wXLZbuumIcEWP9qLqHaYnBBSH+iiAM4izTPi8yQsO1KjM2zKxqtT2aGSu
lz6srfJbgX3mXPXPZF38R0DR5GyzhKQQUJl2cWgB97WD4wBnh6LA2pxxZ+5Sdvqx+Mf6kx3paS7+
KsFn1oA2ax9toz5MmogezxXJySdq0FOVdK1qHBEHzld8AASrSgtyglZxFDRJ3f3DHQePDfi+0XYs
lhg3UAx6XFNgBFbIXqeELeKYQUA29kOanl3rtdm2RvnIkTxBplhGPSg5nwCYHEr7w6khxmi+0FId
14paaBLy4rFY9iEjkNbdfVRSItFBhsv1uCkpk2DANEKteYA2+VrQGNzVotmGJLMD7uW2+6NQFhMM
kjmR7aEJEVqUkVZ41JW6IQmV/RWAqxI0qUfob6l/jFsmANS6EwpRlDW6iqUwAZcHUOEX7bBZPNlW
/YAi2J8x2UXGJ1WeA9cHUdtx5mOFPplca0hwUv+QMSDhk3noWDcpYhV6ZjweCKiX/1nsZDvx3wQT
2lzD3w/iB7vAisQjCla/+m9Xk3TvWGtJAxtz7bd/pTrCpweK4zLia5SDhiWImJVa9/8/Dr2HZSct
fyGl8EDzHWJ77BfumT9KIdION5ZUSuaCiavtujvtOzkDpEkNv7qKFGIukBLCtOtn4XcT8kHsj90m
fu6TeuG3QwDzsvULuE58hB4hj84qgmkxOF17FjxCJ+11lGEUEJOlOLMGNayo8lzyjfO3vb7iFret
H/qHF8rXQE567ohB9FBIriC7sZX5i8ZPQdw9LpqSpuTIl7+LXrJUwrzR9pT00E7KmtuqJqhCZWaA
zhx2v2h/j0H+JNQpxazLszoCYkyd0Hd8jhlOWiYqrTW+WR7o2wtpRTsHaAUA+klGHQloCd/373vq
ctwMlL5zyu1oPOHLb2nFFnPTy4BEwVEmUaWQnpu/ZCYjr4uaRUDVvAneF8QXWexPxOERihjNrOpe
9/L7pzMA02FI28tti7GRVyfh+HCEpVcyx3sqL3gkz4iXoQgyCeCl/rwJG51P8k2iIxtIunju2d4H
1EJm2CpIUuEB41H6o/z9lQs5U2F4rGnom6ySuJZLjkqEk8m3TQEdTx665O7Gj9j4fKEMUn3v6s4P
4U0nV412UDsj9J5PekXOGemE/FMbO8G5St2sUnCVP/TMZ0oa2IUc0Ebmn+Lgwbip0tCK36cIBeXL
onC9Oys2iqBWcgrKDPDvKivEHhwnOxFyVXaJMA7etu6doDTA0KKi3weP/zvmdIUtOfYHm5KF8pMk
PF/kiiYgmG60U3B3l19pz3qvnigMq1hlT3U367pILFtYO+bRTdhBNuhdX9N2N4PedsevPjQOllfu
LvNDkLnufBDZfpMYFwZBT8fBExVaih3AlWf6h28rBSW26bWYhFGg88bewMzB2W1Ovy7DwxsNy7oo
XxL3uDjkAyCk5MytdtZMgXGn3qBzQ3VWNGlpnYokdFKm0S0ULwY6vZ6jSS1IsnMwu0ISCI1zCpj9
skC8U2rSYMrelF0uVA4Znr6gbPlIvavkthMq2iQEbL/2CdxN3ViIZdpYNNTx/glrwpTjin8Al5Ej
Ewq3BlMhocwKnctj0QynDIXlXmGz62Pc8T/Oqib9GKVFSc8/XRMd5HYG8hAejdHa4dQNmXVPSdOU
Sr0pPQEKvO/9oS/GsUE2MkSoALOwVKljJ38aZXvjWOBs4Em6Ts5u/453uR8Fyo8NPeTlQr1rxbpS
UBZgl57Oxf7Srf4ckURmeYCw/hxLxFcLywuF1Rxzaz75XdtJC6dPNEiXz1UgNE8pXy59T4dMj4A0
Yn+Tnj7UUgIuc80jRYg84R5/5Qub9FQiir8znj+xYMjsxAfMblw0foLdR+dRu5bl/vONBGQ/zgxT
2RErjQzKz6mqeIVBCNy4YMfRscLdPGBw72mL4CDHG6AM7DOT9oMwOjGN19yNrozkwdtq++AiUOTE
7JtBS7JQOvr2Fcun9YKVd7xX+biTi6M4/zKr9lAp9eduzIjeni7c2WJ0FonwD3oOZ8QYGYhiXNG7
erkXWFd1gqLulkRuITKWmWRG42CGE/9LuSqvx/lLb3zP3KvfkzZF4Vxr7SPaZaRVblidJVtGL3lL
BUxAW+NVT08VRjbkTLs+KYt84VjFaaW+xTLm2QupofCsYQZTMSDvcEYUKMhql1o8pHcarsroHZiR
nVPJdn/YNysoIA9RJWSekxb3YM+6iUU89WgkAG5vU6d4AuI8urUsTq1wHvTxInY5qI0ye/1CXdol
wo6s6hUVWVc1NQBpW2Vdes1HneU3I8aS8kIC9dpgC6eVU80dRhZ5j0yxlIaSnys9GNysYwy3Yi+/
qLFHE+ZnwwUVnpqzUDe71lzH6xMaL9ZBcxSknqSH79wxe77BzZbUTvV9+JfGbZ7nCMrk0aIW9cjD
0CSFAOXH/wJnUwqz/xlbrc/XQC6TCtd0VS5M/3NhucSsDOtcEYSfDaLdLrZTeoUgQu3+ip0ZXwoL
iRJpGPHdfTnvuh5l4AvINbuYot3uLToFDf1dapu2/M72BctHSca2SlBLyvALjaCshaEdngRNQ9eK
DaKTlxRVHTASwrGjMpHSoGSBrzTStnyTvcRTB/uPD3oCB5TsD3KHwYnWOx3ziw1+F9tcN2gB0tT4
O9Zs/gRs0BXQRJ34A1LMvEgsNiBuYKQ3WSH5KSETwDtu/rCLURRSg1DG+nBxeH80jp7QHkCouVmv
NA+4hRO207w57AEG2NFhOJEwLCLtVzS1LyniAETpNbw9MRVlPXiGHH7sJzrkObR+scKSBacaKeca
1q68j+xrxJyKr8vMc4KQs4C+euZm9aPEKps2uEKgMXsG7n2ME6wxp8PXNCaRJgSBy+BiCTdb6eFa
zx572vqB83BCZDPQ/3OMXbcuZzRcJKV/x9QTbjl/zoLtSreXMXd3cXq+bZnQEP8oN+MTu6ftGTp0
yEzr2v3/muVTsoWW+7Ma8Ch+mK+bhDqAivLzReUP5Se/CAz1PBWDUUQrBQaEn6/8iXzL5fIvmCDJ
uoBkrObB7EJz2uIjzTTygM3JBOFAmYGBqwd1nxFrYPRiSIUzBz2GVZymfPTgRTBghBp7msPGuKqb
uOURPakwBFujju6MoxAaaqIcYop0Ya5l/pZFC4Nrx0UD+8TPYeydVnXUm7QA53OzODRN+FSBiuJE
uHtho0gipx57ShxhizGPeJPA49CywLNumRNH0CBHVCH32/2q6Z4D3uSm7HLfU4Ha6OokHoqZjPU1
BXSS4AuJNH2jqufN5Goz17d5sjDOI6GrAX53lHgtpkyl0KzRKv/NvYY1jCti6DLlIdsgHB3Wxe31
5rXFNnXNDROSPLa14TwTOHex5R84qzQeZaU1Hhj0BlQPFZYLz0zirCrPeKum0yXZGmqQrjCUpd4m
RsoNkYJfsRLH8n7ueXNppSdcmhl1GNIDAi2mMwD4hYWLandjKntpq7uydvfQt+vKZFXh5b3hA9H0
qvXLiRr2yF1ltMg0JlU6/dtTu1OLi9tVW3CFupNkiFcTKI/yWUIowbTXqKFRpUeGV4aWrnthqHuB
ifVKlIk7P5v62j09vHC3r6IRzFBkJG5pFf1NSUikI5E+XxX8VLi87jJElsV4vD+383DkoLbT/UAc
pAi0EJHOqQQdLDgnYx9LD8AAQ8okJEqSxZHCES94XLngshi6Ocfo+KnP3HdTe2x2gYt+u3DDwzD2
fL4OblcA+PtHQHnBdzZw9L/nklCKq4oPed543ff8VsuW2ORqLJNxiXZ8Q44dsR+xFaG3ZR1iP+0H
lUhsBdOoqzj8xe0jiAoWa44NqycVYwlgMhitlyI0ODijTHm56OgNhrPxLnjSGAOR7TyYCfiM9HTv
+5OqjEZIWecjfRB0PJsd1QDmnbns+yDCqh1CCf0Hs3jQNeBJpq4FiIDwQ6lbBU/KjwjOWSm+hUOK
t5B/znjBFp4eyzCV02qm/k9bPepXk9uXj9k49mC/gmpy88TRiL5WQIyoEjD5pkQyxdXyhSplrfjL
xaNMAeMD3lZvQNw1A4Jj4knsX9H3tCQy8dy913ceHx6h2mXLU4fIoZDlZ/eIYY0z0dKHhX3kp6km
FBe0leoE544oxtIe9KoLQgG8RZo76Q1bRs+gV+xFN0M6cq1WUoBF9i4lFRJPXJQVze4YikuNefM5
rG7YbORWvCCeCmWsIGiEcjVrl2uowwu/Zj6T1+GIfYQN6JNLMm6xKh9JRjcC9SOL6gV01ZZ2YzL9
r12Nm1tGh6k2l+JJZVx0r1cUG+hIwXi/2V8RWA/Ld4CQtqycQ0ja9icFemzIeUMMXmnlIlRPpQ8T
IytP9y5nNaarmD9otX6iSnzpt0p7CsNj1V8UFm67FHqja/4qqA2VYTfw7e05jPz5Or9ypip4E0ad
0rjhlH1p8xfFOiR+yJgfRwB42Uv4U8JIye1ehdSG3tzfuOXnQfVP78au5py5a3vHtXR07poMKYT8
wM0jYda33NEZJJrueAViljoy3Y84kDwsFR8dCGfbT0qabpCXHG9XaXyBx13Jhsg3kzN9qsqwdSZy
FHwKVUY8Y4/NCFuHnrQF4mpnk3E3Zi/YkN8stVV3gJHFg0Srdv3kzIUPL2CJJBwU0nBBdFWURBVx
jvocu3pryqXu0Y8joz+gExFq+3ihoQy4pF1TgHye01N2q4NYS+/nF0pgXshswzGZgE+4tIO1sRdF
i4gfUnf5xZkmvfiCHzVT7FluYCZLtAeUESrngmazMVUsBPkq+pqE0cVyfm3qc/zHhlskqvnMpn2I
U6tfupnzD4JfKfKUzK5v7O0Em8inW2U7JjOexWO6kMFRiefZ1DFA8/xIF38B6EkrLbRz6tR6qN8J
nVPwpWI853e4xEgobiPgNCcP3y9S+fqRvYi+McTGUjVijlcc9jIjlCeBf4fMJqMCJpL2uElJRvGn
qjy0QFU3tbj4/1kGSLVFD6SRI6G7TGgdirBufcoa/cxrnswt/9x8WPluovbWBy7LDfJUJ1CK4KkN
XIvybnb1FdqTnWnTA4bGHuR2HXIocjQp8Ldoy0Xoz2UzEU4reaaz9h8X81a6JlKaE+E0rjLfAM0V
xzBduEwGk0ktkzyL14fN5JgZ7AhowzwOHIwl+ZzqET52NelE+6UmhEb1zEU5U+7Py26LKz+M6djK
MtXEd7w3GrJD9YATKMspRAAkYG79oynFTqtzGNzEK4EoXpHo3V/tb0Bmi5tUfWE541/d9mr6RTZ3
YocNeJaqkHJWb43D02PQwPlBWU3JTdZ7JFB1YptZPbXA1b4ZjzKlLGo9QARCv0yyRlSe65Q6V+jG
vPSoQoUxBneamkFPt3O1y9fjXMFpRfGpOjKkzETqYouBf3OysXauhroWKWyiFChvqT9+dxoBBFa6
+g9dny9F7QG+w9ICuLGmNWM3SKE9HZ5LNallMGrgDs487IjY8WBjXDipKnLMthQpuC+e7MoiJf60
JGIdKtaM9pCH+Ho9pCxE88/LonNSrpPag6VMsthlkrALCpRerww6h9tlky+4+pb0IQC6vd05tHvJ
MkG+YVUMj0fjqyCK1zmvmzemJwzo4ADfnB+BUMwdcwFM+T+b3uX8VPQKZ/xAZyISp0nK7AcPSKdb
6KikjfiGt22aWIWxZWQ+Fp9Mo4TaP6Ih5wEpqXv8rSIohaKHlYWjF/eQSCV69cXlNWumPFkQ71fQ
d+xP2qd5NJZszCEkTPA5O2pwRSWnBuJmTxiABb1XBU8ytd6XWht6DdHAhU96hBKHhHnft9AJXO2A
Nl0WepN5/T4zHuH2WGJ8c23GW+7iOUmH4O10Xxsue/7IMJSYcrIoCpP2zmU/2hYYRsItwBe1IJ70
G0tCTnYeHg/WouVBrMO8ofqnbQz3mSoCOjLLjFx1YeZPudHW194GWC10slX8Y4cElK0aaEjZKNRM
Ll7Ikqoe3VX5Osv8K7HCzabWdbb9zh6d+SAGMEis4HH4eQnkbZnLN/7Ia10fTYmrCC/R4ous6+AY
ptn1WUVIcYrC+5rBBvhCWi986xa96hv9DWIamxEdJ/NZ0v8hMomCxc6yJ/hK/3p796c4F9dEYIki
KA7UQzEvrQ2jymC9vvn/xbVSGVuTNgu4uU97/O8s1EsvnW2RVz3VXVE7KU7IXfe8fnC4BEjAkK1Y
8Elp8tRasfB5KwBjI34MZEb4RH5HSFWlYORY98xiuO372/wfn/58x6wv8wHB+vFd6k+qthwZqPRb
Ie9OBLH08cY4M01lr8TyM5x8eMUEK1bIwKRuYF8QSG90eOHgF2htelZcHMtHicvwnicP/fupC0l6
Nh4FVZQ3U8AeChS/L/+4EpDbMJ96q8xEuAVwAfsAIuzWI64oT0rEKXfZ4xgPVNl+wg/pIW6OqpU8
GGh2lhGMRkvXWlvchQZ+l4v0d1e1h+8sfrgyubdHZXRlJPKiigaBd5ufImPBdvKL//yIYa7Lnt83
NlaqhKZgFxE63PhthoWsmJrpt7E/59b9pzDOiaua2aSj1mW2NkXlYZ0TntNoS5/2dyjDBdXGVhdC
NXeZ/bJkBD3tO7WUUWKJf5qMvedxBNg/pE2y6K3HKMKy7X+gI8VRlXgedyk0Kewe0htMjQ0y+uSz
J2ZVG4QlIjhHbxoD5TjC7ZA7X9TFp60KyJonsk/sRFYzYBY0Ytwa2IqOUjIni1m0X6Z2somdY4XC
Ev5GmoWW7Zb+rnkQ9WIOOXq8qQqBfbp69jjbl+1p+74izuOHyUequg6iDDqR3HAjdzg7/IyyfkhO
jaGwp5SJ2da7svfcCxEl/CzIY8f5+WV4v6r4QYUuKQFQqEKo+PSgerFwI8+ktGfPWiB15hHIy2+j
zIgqqTIpE8u9xPCbUJhx97lE6A+56X0ydghRR3ZYWvSeMfp84lmvSl4weYcA+IjIhsPGDdQ6J/kp
P7IX4ebJGcJyZ6piUSh9CaXwoBi+Lis7/s5h0ubl3P+8mUjgc1gAPfEZkaT98rbfTM2u+kl3uekc
gtfN6pW3QQNIwo4IJ731qdrQumTIrE190nWs/+wESqhW05S4BGNCdrrt7Iw28LetpZtpQZQYGrqW
Dwnd1z+Ki3NDh2K1b11EuiGrsPdKGVphD0AAs1RBk773+L1KKCa/kQaTmT6IoVOQygg2DP8iY+Lx
Ot47tb2k3rFeVPqa7RePqo9SVNSs1xUTiG3ODJ6wN5VQi7Zm8ev9nxU6JBCcAZ+mlQkoKK88/MiR
uZpIQvUzpacqBx6aR7uJsb0o9DTmdZZ0vZD+bE51CJjDW/veWSn0iaN1c2+07iyCPIb6vjk9PIbc
NEbFdPCGf6sJSh9ikMvOROSF3Vg36JfYEqgNGc/0Fb9D1fMNsjN6Q1wnsu+LbO0kxstsvi8RhQ3Y
wB1BQRW58fVa9UKG1gtaqFFctjPKZ+mh+0yNyB+2fktDvXRhmCTTpFPc5RWhHIbVFcbwBq83EOkQ
HrD+p6Z1Id/4XSVwfM1yynN18uvJj6ga79Fh1EJ1j9z/HngQGoA7c/MzEAFSUE4fVopk91qttuQJ
PGxonaRLTakduGeRgFoD/2tzh3b5PIIfv9Cs29LA6UcNZ8OwYXCyIIbJwNPrgpYezkFDGxO4y6C6
jDemMh9v3eGuq/2fq/3YrodQXANeW7zjEm1722ES0QFjTViE0+XOm5kqzj42HaRvSGdfgrtIRotv
M3xWcPN1FNDpJLiCynyA9KUk85ItHE8GqRRHGoCM0iQUrFMQlECuQg/18aAphtz8WLPmUo8r1eaW
310r6ihDlcrmWmLxGQPzVCvg+R+H0boOF4CUAOD1teNwrOiAysg/QytERprJ9S5fuG9KjMr/+10C
POhfPNGPvi/mcX9WfP7akl+6nCPxkWJirCWU9Av21q2o2tO9l1pWRgFB2tJRAi0e5xf780YU+GOy
PH+pFvUgSoHkOt5YqLyl404OknclufbhrgSdGnn7PuDVbjAWb2e9CE0Za5sGXfyV02EbXtQXd/0w
r3KYYkp6YWsYNFB4j86/tmVtZkhmtCzBPOddxDLDl808EzaDkQsSOcUn8Ikx2srEZ/1WtWNGHsfu
WYZW/JJjJya1ndo8tf2cPz+/CCfRsrCHUaLZorp/eW1JXvYTiBH6eLuOEEubDg9R5sLLyh/rv39M
IjLHVf3NkE0pNZe5a/wtK7lUa+LWtgONW/p41wZHBHyjkc21j43wlWuwhVLXjVH4nljxcIgOKtDG
lWCsJR4Ap87FEwqngtZ7ybcIU3sL2cnXY+VXPKpLZjqumZGFw9+kalgF7shqRUCJ64wxuGQRmAPr
hqy5BIy3K6HYVOb1Mcd4r2+5PQaD7h62RT/GYUqPiOvdB7VovMcGrCvY7ILr1coX7SDF2tf9rgm8
YidF7Y/8bt6yRwcvPVkbXFpJlNJfKaD8XFgq+y0GQKZf67g6lTN6YtMiotAgKmKFxJLNRvAPD9EF
924t7c4fTkodCbCn/2W1/jH9F7Q7r1wqI6yAG94hHPHlWyDbUQZa45XGWirjCTM/6CXUz37QzUOh
Q+P6PExUMf6qG9Hi3N7dXuHW7XEZuXc5haq/9xcjhfy861FFHSKaQ/OPFtBTWyGLfsqUkU/nQp4p
Ty15KO1/OMK5UGv3mKXhdgd9ZxYsT+LdVpzG8Q1Bgd10c9u88GNQoTKH9FGw2OnwQbHUxVB5PpQM
s0g17DvY4ek58Nq42rdV+vzBAs1/upLKR66+r3L6FwDgq/xGBObxmANSKOSyFkRW9M/PeS6HUvES
EzV0W0kw/GU/wGF1ZKG+ISWFgA/UjTBx0pwQ6emzdny+csCs7rFfvPRN9vUDvCsx41fOpiFGpe3N
7fgQrb0bBVl9RzqdVCSZT7VxTG8kMDmTBITH3e0pcpV6pGqlb3xx70+6im7Vhxr8ng8wFz7fCvrA
qOZmY5uByhLXH5AANyS4h0U1nFX/C+P05W1tV6QX1VgqxaML1T6aS2PdC/qY5ImAO02TVlbhRisU
UNSiBVak5HCBgAMZMyHpp18CYnxRqN17rz78ZgohAuJeza5xX/RGRZhojA3Xor626pEDdLXI3Nvz
U0JWhCjlOP2J2pGQCoPHMrDn3grDAc4S4ZXVWXUwRckJ+PqFbARBU+whI6R+8DnokB8mMhWJWWVK
RAd/LyrLO9yENaqfTJ80EqVTVmeXEgL1vanPh8kwVvAmQpNyIdmYhVwIUc++tufmF6Rwh2NNYfCp
rAnmVEUnosgunpYFWhFI0xUnGxLcmGotyIK892BwfI0PgPv7tamZlompZ0d62k4L0B2GBI2W2D/0
vWrmmkhrxi/WoJVCLEDAGkX7e5Zw6j5kFA3hvWBmUq/5mfNT9BEQB+wnKwXixtO4C4MVy2BLh7CQ
/4I9+zZmY+s44H9/h5PFIF4c9v99mQzkEraH2NmzboPVkVhhFE7eigFPXaDI7FDP89EUGZwnitqt
bUM8IBXgbH3bxygBG1+UaZO5okULf4drTQEbPb12pHN1MKL3uRXG9Ak/FhJAZz09l7htp/Ypi5bA
5d5BVFdrUM32wK8Ee+VL0P65+xVcrAttfzrCK7AI9OUuGpY/+KaLfFAibGblwAVpLXLPAiG/RuJI
o2fGx9x8NnA2uH+JmcKVE8YOeHA0Xm516R3FaMyFbzUVDUxEXDxTzvudPOApx14LA9fT3FHgpBYV
XMqlbDijyw4BcwxB7ZzhHooScHOVpG/5Fj2KR/pe/J4d9avWy3Nn5T18Xh4G8tLsVUcy4R4NKvSm
FMuv4l2lra+7fuaR8s/PrvPxcgwr2AUjZinc0plYgNwv0xqURqyYlhF4OXN7k+QNOuBFqn0WV4hc
xIaZfBF9DcdorJKBuERof18c9UcXSowAtNR15ln5vzrwUFLoQzzIR2wV0LelTu4sn3g18SGkzoNv
rnU3CM3zMhgPwAzzqum1+ilwgcs37DgeJytsGHi+ejWUJiSInQ4qXPArePSUC5zwcG7u2j5rkr4X
6387t0QUC+sifmuGlDcgKN2gRo+prVbOJQGiUwBy6FSXhj8Ojvts/vADfhOUKVIVldT2cSCIvq8o
eLDgWe5ZgI81TAVqbtr3GdpVmDuImITv/6ipChbVg101mnQiXMgCcbmPCiY449JGRDWyiMJddIjX
/3iOKA9DrhFJI/QkrkvHmqHUWIOU6rL3JNm5O5CZEAot7CjJbbIdokjI1II8P5IWuI7DTdTptTE5
mTi5iAa88zpYSm4BhiFGdhUrVEXQ3tArxdsX1K3XputNv+4hAdnPwnMx6CmSGGpSw7OeMUG9DoLd
6NybyII6rOPpyAsUvFI9Jjz595beBZ/VwGQjswTqND2ujenkQCnwGly86YQe6FR7jkV1lxdqBipM
32gfxH5PY7QTx5f+mdc/w/dPia9XoYji+IN6B9P9LHNScOrmjTDG5ODjkD1KpbI6YYGZXDM8gSNa
c2jdSFmPsXsa7Ke+gOuiqbUMubdkzIpF1/+XsVr92VZROkgxaOL2gnHS97AqKdoY0WxdplOwcJH5
0u11RqZ12t/blEWIdz2F5+pz+wl9w7PquVrfTuVMVQaijsUS0v6cz1BelvFUzOsCd1kWC9AeoFzV
+WL3PyXvNZns8W5m/Jm7a4AWtXENWNNGxJoFU+US+Guipne3KAfdIJApkzM/G1YK/FNZt5C/4aKJ
V3OASjU0Mr0L0j66UKBMga3GxAQ55ZaeEDKW6Yxlaaw1uDrIV6JJ4PIbkUiSOX4yuWDDXVHRQPBU
S9aoa7m8gxsDEq8UBtCLceIVinFi3XljvGdTQ6rUe2Pirxcl6s0WE+fT8FMsi94PHouNrkBHR7MS
SPt81+vAA7JlbQg4kVbTk4gMaChW5Xdch8h8M1h75tb7xNP5R8FBFGt9ce+5dYUWSFF6eICK3Km5
D9b/5/spk/r86nCBxh8lz16QRML0E8inK0nrEkXJPr5bq/suF1lF5t33eG25AUe59QtKpmmdTx/H
7BnnZg7G/T6BioO+9vAfxZfgUgrViEJCBaSD5XhV1lUEGz7n7pe96Oq3D4RKu0H86MaX2HPmZmu3
vP1V6L9C+W+41rwJDSxUJmV1+YR8uxF7mwADGdA7aNsDCMYWyMBvJxWi1d9G1se3cKxDCDZtcRSj
ymqvgHZ4WlNwgFISniezdnmeLyD+jZWROiUkV+PzVo+SCLsQbhJeEgNcgeJH7arypqi8cyi7JDeb
iyclt1Pesar4HN+mvRBP3GJEoA197mvPXVpk6kuBVfG/fjKHkoamyvJrj+7u9+eNrJK2/em/dVru
lqdvCBuyyhiJ+gcTKkckakS6r69xOr1BKHwRVL7xOCs4HHC/qVochuQGRg4nDZ40eIREfN2imeI+
KQWs4DbV75NxKZttQ9UkCwUZ163DoI8q3KWVanJiRbrjIKcwEknMj0XekHsr6OF+x1mH8WuXfW1q
H9cdvcTmat40wSYLpq/wxP1pySEzfUVcowR42ucPWfFGp4Bnq3I6mSCrAlGo36PW5iM7tVUzg9j4
q/FDQJARxnhFlidni3ybC3cr6wDiuHsfruX3I6KpbVWjohhc+KykAT1fX6NTqIkAkT1d3OJQXrJd
bO9xVzO5c/5tfz6lS8aQH0e+QO6kPZU4FHWWuKAoFOl7lVyTvpDUrepsjc8JaTCCvYzGa5erGEbp
7fcL9qzNQqFk/np85DFncF1mQi6EojzsQc1qCSVhwrM+JK/Xgr0TTTD9ooh/Qk/fYTAIu1KHvclm
AFPpCe15dc2r9MeOVG6cDRFbuSbHqoRQ5Nt7QbuCZuy6jIijXt1wGyFaRKQEzZYeNVv1klcb7nUU
JBhJI0Aa2x2YG5jOIMcqM/kwTUeaad936pxcfIGZ1ZcduRAXuuhNgFR/QGBKP3v4lT2ENlru+EGw
8C9WHUbIdGTz2FD6qXsXBf+dCprsMvlVMTNNULjV2Zc++JP1UfC8LnPmxQFRuZs4bwZK0UStiOg+
T9EJmfrl/CT5gwMO2jYzO9ZfjcaCApCQmfgGvARVyK8s/aJ8LQHXEh0l/Roki0UfcjxGtVTkKkpn
6fs/YnPut77jSz4ZB4EiSukzz0qGeHGvuvRlHX/+WZ+IGMhfftmWH6q00iasSNsbtgisXTGqWc3t
C3a6Vbcc+zsLsbGogqUWk+z41greR1FapSRG7a4fdxYLZlhknQHGuR2bY6wZP/lPAy8vFQwAlM7i
7AY2YlO6T9xQxk2WWCRPy3WnWLthbKCKvavSc8l+R/sEiu4M5ttL7whkjQLT0rhcH/KF1R5i04ab
NBWyt0W9Vup4ypkbqGRBz1cWs4uZJvhCyrwGo7F5T0CwRK32Htcm9yH8TLCPJg4t8CMu/FoffQE5
TDIlRYT7wTxWq17ukCC9kvoPhwv+aw9InYgAvlXIusqSjtjNyFqIblmE8V680+qvbxwBPcYixL+k
V7Ui+0EJiF5LCnhJ+IfbQlZNsPW2WaUxfi2fYNKYUx1OkoXwfR4gcYgpRK2ir1obSYUxtlaIMRtG
IhZm0B1AbVmeQTn+RihwkuMjiTdY2ZQZ5cbzjqhRVXG3LkLQC1j841o883eQS8jZm6wGWPTPpDN+
xgwj1tXwjvr19Ee/NFKAkjqDS+yWmC9Po8TByCfEPzUkR6dCYWvJ7d9CrCHcPF5i8Doqxwi6HLu2
Owzt1ris5JyqgldbyWuYbH9i6UE7bEZNIe/J6vU6pjXRAygZE8d0LH5uACvhwBwc2yk+sWZxj5Hg
DvZ3KuibKgSHyZNHsQl+7YefYBCa2CHm7obHxY3TyxpBW+/+aAcgdnaqwoDODRAhwxN+6y2HNsS/
e6QSRzFwpa62DHzngqIm3SEzDyQHcBdDFsXSiPuaALxS6kexM04r0EIBrdEvpV5DfA+ynZs/A23D
o7Xk78Nq7H0viaxV1nkjZVzfzEr2XSCJAS1ILrxMJYMxbRCEkt6YT6UQlcOPFRkcJzVyXI4qlHLy
D1yf0sHzbCcD88GuZMdfPVuM0s3eJGeG2ZKyJGq6bQDSaYmN5a50c3nm1o3wtxMnuLaoBqrdUvP4
oIhtXowPZhFrNfJSUf33HrdyWcd0nv//eTotckT9tFIJBLP3TxaWu+1ijpSrQhyplOn6GeF9AGR/
7Bi/7i4j/iVzmDPtbMnyltbtwn//GvOWVjvE3QFybeeZftDdHoJbwsCpwN2f6ePF1Fhf46UJoCRZ
BOxI82C9d/v8Ix9w27V1L/hlToYwrmTmUB9WSoSXUAbPw/G++Szn9lZCBx0sZEyhJDWBiaYY4k8p
LvZ9+mr2LASUjv3/0r83G1dFSmCwKiDJEo4JPPCmLw+yd00+LKDVH1liIQaWgpQhtdlzmmgZXXAa
JxffUpdtKCNix+m1Bqqa4Pshc86YFG9IZYxgF+E8rtdEclMOOArObYjcABRNXlgdhJ/hBVJDI82z
3cF5qKd9YpWzwtlDLYw2vN085BZrZj/AWnJ6FybjHAGX686jYZ6QPSGZmU9KkQ8Kh4LVa26SIfQE
dDzbfNb87YTMjlfnt6aTqYGYgwDJ6kHbPVrMhgofcuVHC16YcSxOfaqNbg8AFqpq7iBKrncOtc0s
qhLzG/YEJHYSQlaMH6lCdKF1YS13DKAp0GUda5NbSMRSusukq99srBj1PZBZmVxVgXFU44Ig4CzW
gcE9dtsyWnipRMmFCQY51BzFG7XlZhDAeEYqvgz4wsDMvbqvXcQaF1xQgk9qgZ19McTkpAkdZGvd
dwfenp7k+sZaRny589rKMrOzkpiOB9g0PTHMf0aXp19hYSGVJur/61rDiNZcPnqj/CX5jOfUzwUJ
NUFi4kJLBmAdD+vg6DJPHgtnOZ6RqMSigvepkw28ZDHy6Xmck4XVrR5sfr5mf4AqMIJKjtjvxIru
HC4SpeXOG0atXIOiGwUbTJqm9TnnV7tAU9uTyacywnqz7LrjMbm2ntVIZ2Yymi7beaKccTGMJPFS
OCkdILrIQIeTy60Sal80P5eutd6ESx5zaHUJCzkzRwgcoO5eEDFHH8jzpiDhSxs4rNWS+xZYGRQu
w+NpRgDagQvvC4Dws336bwHpwWO9THbC9x3hdyuDuOZ1yxmi4a/b3nZ4lQ45twEeMVuDZJG6p63N
iRYCQk3w6RBDCoYhw92lozffGuYRaywk0ypJydZiy8IS0MmuW32sc/A4gHxn2NM8t7D+6lhO1ifj
Fv+gwnmdYqAmFeFipxy+lmsqop45mWU2vi2WjyDzj1jK3dTgRktT2nSD36zi4yru72GE1BbIv1FS
+SJkg9yqDcrUMbdevXEmFbX0EJ/rLclPLVLARrrjc2cut8EITse/0Hu1gNB0lUOGaxSPBnuYUAFH
tZNCOHV3PvgvDUg4bW1exFAcXySXIgcA9AxItRGEyjjiAYbXZ/6LV09cUBb3xOWAEftvcurwPppo
4x4Yhgz+LSwgyZioX4UyxVPgVwqZjKQEPmTIhQ3tmmB2AbTiaRiZJDqBh/XApRv37OSeLpJOKpDE
uwkr5oiByeJHedOOcpIG/k9WES2EuLRGW3gD7RqwSmpGbRLB5KDoQRjtlepgAI57xKHVa4pCJfL7
JfhDGVqSzkBswoMSIuqwZMfsNYTDM7uiwqY6dfOZVoWdWj4rKKKigJdfJ/KFgqSHoR3rMR6p00pA
3F5gRZ3qN6aVxrFglUJnHS/qhZGySwYTc7CC54nRCsiPxI/y0+dt5md4RKkNEy00d1fjunCIONLj
ZdbFk4aapO2obZMAVSKoJV3f6Zt5gJdwg10Daq7lLlCqyhiLmW444OY5AjU+1s+Ax4kB9TRhEk9T
NBEa0aMzV+FrzdHqRhfaqKTekpWoYfuV6XGHsGvKHPJg6UvqKcqtXk44CVhQkBN2/kowP+OyMjU1
co+YwY4Xzs842l/mTf3eeZlb8CKRvvGVzxriK0dhPIy5GfEfERdEQghTn+XcZpstNM76wI6vgXYB
QIGstjHIfaTSTS4C+uHNQBNsLaE0+tW1kOYPTg1cmji0zWDULiVo+lSJbBtAFDoB98vd/W50DCjH
RNcHOqYZYob7F6xRk6kWLQybZ8bPWdgSL4SfFSuVN1vfIpUR7PvB0ZNMMDCV0E+jiq+jGKnjGDtO
fVMHYZZKX2NiX9QZuZrT4i/C+gtgxNYZq5Fp7kp5RH97/lvyTp/X3USUX7XfhxRVaB/r0ks5icz2
cHB4xjlYUbY8IbVuvMk/7TRlPNDGgCom6a1WjHqQSaIJSfqFspzoMDnj3LtTtfAH0gGny3foRW40
XC/IsswDAxwPG4uZW7i6MyHITWuIsqLxwAnEMezti22QP78BbJmGZ8ZstmOGFUVlLp5J4qInElHV
FNLk3/z/D7zNoPKOgSTWN7rMjpZT833SUGDxpnYw8CaiSpealFb2KAfUZSwy/DA6/eb+DnQCVPS1
VMTh/mXS8uOniz16/slknYx0jGvyS+kIUuVGVw7zbgg9sxzceGN9mV6q/8Uiwy+EzPE1kGafp4Hj
5zOMMuB4xkAmXGn8jQfPPE3+Cjgans4oLZPtdf3iqpPVcegZUi658Kzy/d1wuZRiK1TAEDQu/zyS
0x5RB84tbQJ9HmXjOmO/jGlu9wko6iiroi0XVJueZNKBa+r+hlkNJRGbTcT4iLQlFkPFZBexjHii
8xhWi8KFel9mxD6svCGEqCzkg/Gj9SCHen0RGDhfiLA2KWMqPl/A9yUGih/TFwX3MJtR1mKc3WSM
btEKEeO14oiMuubkYanE8y2GZYHJjmF5eKDBKZQMx+NEQRVC+Mm4PRbzDFr6bySjwHTLP5V+jcas
ZkxZ20FlrLnsFPSaQlpdlRdHAOgr0YZWhrULzRg2xemrHVySTjbbqEqnfHWMvblAlf1GIvMlBNTv
VUVycgI2wyc01CEJkNYSgXKTWSEuJgYQ424uVD3IeoSKqDifj7hh8g+FO+c9cZb6f2ohN0JL2c4y
o3QSNKAahBaBqX30OKL+Bl5Jpt+jkaNQ1dPPzwifhHjFwbhnBN0Fhs8mbN2S54uxYauO72ezbj6+
BA3iKqH5O6Pk6X7lRJC4mGeolMQJi77nTjdhP4cUlkFvzltOiqXwsB/2EnjQGVjg1kIkPNb+ogg2
/ZJwmqcRrTy0bEO+lL3xAfL9DQUfnfAfuUtEV1NN42sDsShLJE6CXTZ7E5Z8CRI+PeYEsJyVPrWf
ywGnZkz8ybsypVTegVWTzod1Ejdn/OPZxckRpjTZwVknBSupsmmMITqyjfPAQzxNZfTrYkmfA2KQ
q6c6HuvwMX+vdFyjkftC1VoZ1Sezyeif9lwXuEsACfAI1VcUlJJUv7f7wpvTjzPkaM2XwZdIgRdw
iYQpLw1CWE0qa8gSJlQtO4g5jugAIK6TgvEmwAxxOs5vkleLS2AbedKbX+gGoP38nKjAsqkUijY/
9Ds/z4xM1gAlUZwvsGKhqo0LRc1b8GRY0eS4BdyOLrdMRPZZbJulEsD2B4/9FcBQ5sdDr0W7jFZB
U7pOYKSHlr54+EPWZd7ug7FRdsfh6ym075RtPHHlY9zh6cHBX1OMU6TfzwENNAPcPH2Z7d9DYtYK
Pv3kp0xXj2WyxwZy95NYzhpmILgT/S7viR1v2A6QwBAhBkQFqUwCcsw/84+IFrxzm21agO+jVTMT
pZyVeTlaGqsxRlhq6y0RYr84kOePSZEO9iGBRTaUJgr6XwCQEpwBsLF4IkyT3yqosZRoU2Dk07Gn
FTXdZHi9jYu0zNYQNE9I4dXqyBQJONxr/PriO4lsEInt5DjETDWUCdwP6D5Y1N0y7CgvyAnXR31o
pdygX4h0UQNmNMBMxg+IZqJIU4BaGrctpHnajhgnFd1FiAkulO0oDTsyeQA9vF+DF/XfOiNyUQPE
qg3KhhmW/M6dTjZo4Np+/u9wfFG0Ls6iWMcoYYPytHPPKGRh09nNZMJu4lbZL/fVhrx2dERsiKeO
R716fcqRtTHSQ0QNptv5NpvTYPK2zFQnOzv9DCF+CoqQramQYHVPTCIwaf5k/TGwnLPO5//TseYZ
zthCMllDsNUpZBFX+VWOIkfvby4IGUvqR0Ln5swB64yNuL2aavmbHF1qJc3p+CwNz6a7T4wH5T67
uEAXmmBQVqkCTaINwz2NJ2y/KzZ4IC9Nh/RXjH/UGYijJUSD57AM4FqVxmi3NqgLDPs8UN5Zj3rV
V5/uS2TmqvSOf01OrHac9+/JTO/X1oOO+cBXMVEinPIIGaeTPyAufR0K7qhxNnm5KMSy7N+Z3+Ry
TfAlHYExmK1wPdL4NF+vGqV2HHX6nyJ1YHMBE/DlPtw4RCE1zbSNciTUWMZFg3yT7uelapIsK5iK
lZaG6fQ5QLN5gppsFYP9HRz4S7gRFvcX9rMk+2qA9VyKdVTNCsjp3cRhCVlaGS/O7c6/mWalHFD2
0Bw+bwAX0yxrMyEy2U2BVsLSw0tU6PXdLVNpLLSZVESyr2DfeWuwRX3QScH07CBxJSsi1LVA8o+c
nNiPC0WzzMcxuejBbAPjDqsMVuG4yJVF8eo6BHkMso+OroxsOFkk1uAORvnGjKhVirZjhdgW8Baw
4UhsM4qgFrd/SxnicepCKdcvQ3pqYgdPl2/b5c3EzUJN7ODZW/NiHjywjE8hkF/ZFDIXX1S4fAjB
M4wJKh69G3V/63slGEyZX3RmmHnJG4KB+444AYZJPvkP/BHBt40pG7sY3dq+Zru3SjOFXocCj/GX
Q7Sxi2TzFR6xT6Q67LgkmhYZypnEhofy0P0Ekan0h6y7fV2VxJYKBByNUkESxfHfOc9WLY9bzaXN
R2YKAKm7dP9ECtFyy9mJ8JrhjtxlfmoYlldenM29i2BUpz6EL3tMztJV+AeiFjyntyvGMqkjURXS
ckG+NLGGyaqNS0Su934K3u2yGhnsomScCwpj74rgdUo/aAqLUrgBMP440v1ewmnX3YOQWia6gIhs
lh3lMmJhInCv7hKQzNk8p+XxSM4T7lygBwdXvyJsyyHKgK+/WQj6SVREZbIxtciWzcNlU2LPatIQ
aNoBoXf82xDZL4IWf5VGSeMTWk2jqrz4/JCdshEF9LO85crEjgPLovt8X9RNCJU26jBJoRyU082G
M+IEqIRJjQkLKMIN/16O6SASUKduASEgf9p8MvxYI9vBolNiiAqD1b5AtTOWBKK6Fw2JORlDVEPj
lDvWHvulSGcDkXbQS5IJ0wF/fpVNVZsD+HNbO0x2k50nIDBGJOWSv61+GpFyPalVP71Wp4FdBAzS
rG6LD/FDImLQbAYMrLBTwjkGQ18T5XdxX3wCOvIISOtY4WOyIq3pGd6Q0hgdoDNap3Wy3k8AlEJb
6v6RCgJ0K11PGlq7nwFP/TlhiKhKgi4RHPELE/mZlWnTjmS3B8GYMADvFR9pcP+2SfgQmNnoU9pa
0WE0FR/s8pD1vLm7kB45x1V1hf/kKE2UY9XWKlCJelF1BpG6h8WRflaLDeI+UIBd4ueBBW1+N3as
zMKnss4YErz80fY1BV4MDRisCslDKAq57qK/uRTkp6Em1Qt//Q/DlWrZiTI62mO58bYVBQxWGGRO
ahNf0sdKH8ZF5qWH51Kp87IY5EkviiCtSsyvsHATSLpqmvMt/hZvFFYurvqyu8m9QzcMXQDLpZX/
DkofR8A7tEztKHxwxuGc6iJsOU9bo45XB9z+rSDesiwjUJfoZYKyBcakYBWXLrCL9F0W3xfV1/KP
XcyU7oFUuYc58DTpv5GB59p8MyH9asDrbij2MXyHDka7ToIpRGNMoFTiAn2h+Y/JgaRfQIurK0Mw
S5JTXdNyOLqjHmWh042OIXOt3ur5gjgxBTmh9MQe8vsrrJOJkRjx5vjzDmZKZbHnEcqwF9TxzOP4
kJ/iLVYiJDPQPgb6h7yIVwOd+fZ95OxoQ3aQoGp804AN0uOYR7iLt+XJjWBsLEQQyMwPIZmCX/yv
KrVoObBVfRfs9qkuCi2xFXlY6Tdo3QIDHjqzFcTepSPbtKyHQ1QhpEjWO96ao61XSsOqB4vWGTG7
0/8NHxOZu6Nm1lqtgfHNQSqBLNkhe+h96224tAIUrCII8tWRoDgurwSlobwrvAwBCMvxIToJ/8ou
Ud66k90D3Y88Iv/ISDOKQN1XIgS+hJHXPSc36jB2gAO2ZTQGUOyGDbiMz13qIlrQz/xmLGElF6OI
bn0m0gr433aY/3f9ixZStCjQ5+REiRBIVM1FzesbfgGJnyB64bmOniD7X5wTBMzx+sugF9srOxMF
u7SMJt6HGkroAHBoCfSPx290F3bUmNbIHpoKBZY2QiaRLDGTTqEqV0YgikCNrzRJ64IlHfZMRTm/
EewIJrU+7ctw52KUqyYvRl/eCz0KCp9pQ80coUw+K8RUP7CcqJPNvo80lIRskWU8bwMxarM+FHtA
DoqfSLrwdKvAgCDs+3AWDG5Rs/mizQH9ETx4gEiNO0Tef+9YBwskuKXLAgZAPWmbn2Ueh0DwtKIG
zntypJYqWOzs3MW9QdctUaLrfEAFtRn21f37gmhs14kmh1bFQfjG3RgRP359h/n7E1phKOzqWrAc
1WZGeLW5ArukeqB2pQufiG7QP3hKUctCWWD6XtZX/HTZsX95wDD1SQejVTc4HFm5LxqbtoQfMBIc
EM6bTXfLLlTSb3+KFJ0zKblaOyuNs5zBRiixmv/dr2Ym1FEkeX4OM2H1h7SrL2HjZnatoDkbWpFf
v9sdbhDoQH1KcR58+lb6EMq35Us6yK8/1FzSymFhT+zZbEeCum1ZXYMH6pVvMGdc32Ocy1rE0jkX
svrEkQ3lCbRBZS0X1SMOf++J0BYKkCTUqw+Qe7zSLbPN+vYdoW8uNWQFrUzowk3LIhZ5YkLm8fQ1
a+LI8zWKp1+QXr0utS9k9zD+TcCNI4BHWYfHT/jd9rkrsMAEuloKfGZSoBVaVhS0rZP98tDhuuhi
HBSzQgKzPCvTSpGJQOGhMBveAOCKnHAXzO5NaRzzG13LmIBm/KY6cKkOo8UCAaK1lv6H/AH2nGh0
IAKzlNPHTmvwN6Tavdx+LvkmTJ8nJp9I6h90odEPD77mEcXEVVHx965iLT5PjG6/k2PfDmIlVGLw
P9g9WST6DftQi+a17g5uRBtgoAex7Ux8+1uwBtZ4XQZFL2L6hle0pXEFNszh/5TU6/vL4yfKSyZ5
DUg4o5X1LCidYib8zEuIve9rtGLI8YvyyMhOK06D084iUPN1vYXUwm9N9ORLlgPPNoQ07L0yStIq
gOgiscKUtWL8PmiAxGM7OWH5WZ3G3KhAwjOTbPF4MA5m/OsRRPsNMatazveb/pyEUfPcyiv/0P+r
wip/uOGopgCLOQYAmDJ7i57O+0UqtZmc9sFq07Ha6eCbggeqXx6RtngRLENA34WcL7WvJnFD99wb
zfrL0OktSoXwSzHvjEIqZkjFhYX+ETvoByFjJWtIKLFk6jCtWDGVzSlUGw/uWZztxRGvdt4cXk4N
pzNdshYvaRLfB8bfYW4yyzc7Zf+D79bV9kL/okHjxgG0WlLK78oN4hJH5tmB2bDftY7vDggYBISA
agV9D5Ytg+wCaROtKbLibAMgcbOZFaE1M0ln1i/PHRedI6553YKK56tq6MNjgtfOCzR/pEe/zU0S
+PUG1YY6xpDlbcCqXJODiJiNV60RTsdfarHoYhPllE3ZTJZyadgfT1ACjDbftt7EvQ/F9ImvdRbz
93Fg5RpQsr8XtgDCf+yq9omotJopcboGn099KcIN9uH2YywWSijRChlyHwOW+X633mAlsciOa1cO
IFR+qnTd+vNK2gErDTKexXkyV0giI8P9u73b3W404Vu+C9qycBxIYHOSExJBqcDEKnkZL4+5kJHp
RNXNYhJDo6SjAPyW5TsxjQKEZhizsvUhMgvS124Q/gs+QtvXpxnt4t59S74iCBdZK7Bs/MmH85bt
cwXSQxw1HIs9mX2eOuFqnCBrwBsfs57tAjhKNjVnMQ/Yrb4CengZz44vogVgXGEYrU0v/ojUOkKl
ZpXapSMvw9fhQdPjUvUiRXvNmBSivYojI52K0ClvaVlMJyaFTuNuyjbb9kNxLUagBrksmawgbV3n
p7xd9gSJX8IWDLCJoCjXbq4Wc4wTMB8joYa9CXJmTInFCb06DxZh/0UQ8oBlSb2Y3kY+jgkTUH5t
pYKsnxTP2XnTvq0dQr3dF0iwIS2DsX5C3+GA+kFbbyWRQkn6BDG8+MSMNhMKhkfF68sP4UMI9i+n
Z1y1P7pFF5mXYmlxcrMEr/mPmNZDBBC6MKoTUPtLYvCN/EPIN+wtahl8Srzt61xUb3X7ZA0+W5Zv
1PVxV9E0y9Z1iVngsHQkw9dUuKlO3mpQcMyvjrDlHNldNyZgge+NbhHdW1fHTw2PMERQQ0VT/3XP
HcfSGH1CCYnYO0XhZab/3i+SAfNWzE561pvWTUnCm9sr4/ioZT4d1tj5zdU+f8jKvk9R6Pcnn9QD
UlmxCP8M96w/avyisYVDaStHfB+ea9H276+zmM6tt4r6HxxLBhed6oYVFYp9pRZo+SVRlJGEZrc6
O9QPni46o/CDH7AJW+Ioi3edvxY5QNqr4aMsdfD32qwwq2NbypTVwdnTwuDhBq13tKZKJS1j9JYo
2zcofq/72sENWdHiSWxqLsmvlu+5sV4xjB81G3hReLcPZ5t2aoPTrfV/bPA2efAB9kY/WLhyh//V
qLz9k7cC/NKyP037EXxakMu/eAW6G+dI80lZP5bgJnfby4M733dxRUvcCSWYsh9e9u4WKzrUBakf
VznV+snYw2KPykr5BqGOiKuTU+176Y3I4HyBnw7nAXyK7Cu4f369gGCfFzf/3Uk6tl+NxqgPeXR8
eUhLbp3F+fWfA+42I14ozACe8bcKLV2FYFRmFgpFLL9L4Vglbp/KyKN5hmHS9kZ0r+mq6hFd577i
BwLDKcV6HpJNn0y3dg31ncj6HaVBFfkbovUhwCIWtbBgiUtNfo2wrLyc8Lk3gmxWbJmNQi5JIdew
8Z3TQqhfwyHfAe3cRtbsuvbS6gGFrPzarPRy1N84JJmxPHc2thSlrNnbS1GdQMv260V8BORBGZni
hGXEMXzA3Y2J/97weqEjbppm9IgsEgMavU8+9tFvCx5uGucdz0VXxWHmxQsaPjIR7U/0EtN+vNpJ
Bx0UWPRCdnQNMrs9lQEdTUpDySNabQqWXws9UqGe6FDLrtD6flTjPdP0PjKUsIrt/B17qsmWhvJO
9rYg25K+femAtj4cdHnDpYArMH3uvT+IF+TPfqzYDSf5Fz2D1lA8OZCRWxZ0osMjwu4OH3Q4wecx
/RKHcMvrd9zj0fj/LDrVCOeevRWdckshH75D1pH1TP7G+gr7xcC/62hTQET0KjdB1YDkJ7rbcDEh
vZ8qd4hmIl/CarFLny+Wamjntb3lYkrLuLoHk38bp1xH3yd45tcJGZsnf3VkFL3kSDsrfClOUirH
OMWjV2j20oRyR/5pfsmlg54ATK2i1jXHoRV/48Kl9vR8uy9AkRwFYnAcfJx2iW80+yBVs0z7KX12
NTcLr2TbiJZsSdqIa5DCVM+aAELkBRDTEeZGUP9RNQKfY2Ad4S4U4O05ZykDFhukcFXSAMK4EpSR
kYPcymgXRD3ACVssU7PAdaQz5POcWBsnL4f7Ja5pqgmeFN2o9D5lLTKGiajAV4QEwuuzjT96XxKd
v45qY4VFezmqIe9uQf5IrWgKUFoQjHuGqHhkQ9timNfx0B0sNcIoW/A5GNSua0J+plvi/K0/uikb
pdV7YgHTfnd4h0JR6EDexkN9nazw45Q8YaGgJp8xWY2XuPlZGvko2JVIu1rsfml95cecXqCNiHSN
tAVo7Fknij61Jtqr5r9ccipy+LpTu4XPPwakaNILXu39q1mwdDRMZiYnSL+1SRsdtElXf4JoGfJP
8+XToPNXJ4M8EV8otucEkaG2sr5uF1SJLtaFuMxFnr1Itwh0bqzN7fW2ZhaTJki3Uzdb9B+P/fn3
1iyIHRuz47yFRc+zS5oZMm1QzQOBSRVouZJq2k5EIPv5dCfpCPcnj2IAGJaVi7xyQm+7ptZb9GVj
dh8SPw1m9sAsDRAVaaBKqt/mQR7IFwMabbSUz7J13dmDVeVa+1gQYXtgRTLCI8ubKHQL47BWXZqg
8nXh3eODqpaTS7hQD7eNNUioS3G4HwxZ1Lagyexb8c91KpkicjETYKBwBL7Ekj9NyKYgp2bfPhWl
Wscva20SPl1KIhh7MkF9y3OdtQ6tbNgzmGI0fgNedp+k29u/1C7OrcG1eK/gbwApra2K+Vub/qj1
rfNNa4Iik8YwfCGR024tuO6IXvGytkHlpGr10xdq6MKw950pY//dSphD0jUfJHacmmxSQai0XSMx
Du6gCygAoJE3yNdNwlKFFy6qDS2ngZPiLQYtApmZzvX/U8Gn60w4yLrcs6ncM37Z7NXhriBd4j72
xnUcw3o3uloitDldB6AW8gkYd9o9v9H4+ZwDBy3L1IdgDw4uCHa53qYeAQZ6ye/53pcIJl57mLkA
pI4vaMDUIJEjpf2Sg8EUN3cMNEQe8C+WGmYI2dYdWYSlvuF1kd1nvH5qSv3iywYDFwE8IL/9M2SF
5+n/ZNcofh4PdNB/EjGDxbGVJmfhCNnbnxIxQ4dN19Izsi3NJ9rfckivR/9rCObTHxVgea7fRHhR
DZso1AICiTVDyo1bL8udBAoyZq+tSJKwrdcWv2xnlEGYyFctcII6KcRK6V5jRXLcTIFKhrB7pbgb
6mmIQzNFCKM+AaY6uPzxBXnqw/tnr5TXJVfaNHpmeaZac8YBf+fnjTL12BwyHk/FhmYREC5TEeIj
VG4BvPt+BsjRPRCo+w9nDY4H/wM+KlMsWH6tWF8rD7xlUZkP3qPQ4KeUcDlGDCDh1KmrDgHmfMrj
I6bxh8bJjQBQME6BONUU13tdQfQfjVtXdUHsKsaHz2VjTyymO+2tSTB+nDhw0tx7J+5zQzvhSS2c
v2RQ132VX83RGl9uDbJt4AkXid39PrSt9Jz7sROoXQYjmxwRLt50igCTA35ZyZAQg7YVCplyvLOF
BXkHDZJoMHFQ0GTgUmfaKT2khlMVOMLGY/fc9rBN3Jzo2DB+Ri5UQz6aWoYMyXelXxUttxmKXmVV
8b6TU6yDRVvgqoyhGVN8XtiRvY3mP9wHWFfu7MyPh2Ej8IppfrcSLqb80w9e+4B3tWSKj0hX+u1u
BRtsgyH6iOr1cz397wuexBRXX7TV89Jc7jggPQMwncXti0WQjcUz4rMgjDmAuIcEckzFT2TT/qlt
5k656ZcPh+VQjVHwdcj1ASQTrE+ShtTCOp/k0TwbjylQ/Zp1+BO4YPATCqmcfYqAO/q9ffbzs0oj
y6gfjMILkWDgshxMIFQ8X4mUdA8+nKldIFlZ/gDGJn3kUHIhKLCrtm9pe6Mec46IKT8NUcHuEl7b
thIJ3eDw2r6lM6MM1hurQrrL+00lW5IdJ1B2OQH4mlO1c7WYW4Jzin3t96HFSJYfd5m2QZa3XzQh
k3qEP/LrDhZ4JLTaJ4ZR5pap3wh3gxUdKGp2by4xrZNGVT7PG0hd7E5HNdvHq89jpEn9WUjHwXSu
iYX8TmC5ntuizHzkKfmzVOVGKXzIpUZa0XtIBLHWNq6xpsrfJTVGZuqxxXDWiAuyVoM1OOUdVLkP
U+SRidMez2RMZRtY5Yp75w2muHXBpE8PSRnv8wosCsbtJoQvSb0Bi9P1SUFwV3ZeON64IKZmNa4X
gEE5WwFFaZWG2X8jBfJYNWZqDtFDe54QS3Gdz8crs+PcNnGTk+4OxfGktIMmSlXPlLGczIoKjkTs
qYBUgIxbI2YLcEdYT7l0HdElaqSVBPhs1NLOEMcY7j4p3r2Uz15LNb/dg1dzLkEj++Lxihhx7bKb
XpjhANeTmesWV3UyhM9FyoM6aDP8ascBQJfhLL8N066ttuQSKKeo6pqraFhYmzBpJV0N+Shef2j7
hLuhIKC6kg6w1a7C4Tpy3f1NASE45T2wP+TULMyrLAn9CYShzVTVd3l8eoQd1NC+2iiSKXzG3FEa
SKn3Mcvg4XS3j1Pe2V2a/5GvEU1yE6prkEqWEMyDh4gWsntqCbtCarT07ZcGFUpuYYjbX2A7mZU2
ILRY84z5HTIsDOY9WhIzMsz4LO5dtVcqJEaFSjckcRGGc4EoAEPzni3Oz5TSiedb9GKcm1CvTMmG
c4Ha4kmZacP4RUsq0/+5Dszxosmn2PTeQka3ZAydKKsVHTZmhuBUFGk8T4Gf+wUcO7i1xo52IL3S
RJeXfITLyhjcBz9rz1iRaL81EpgEyufXE8Re4XS4aYSL4h/QlI6R0pwa3tVGtVPseimv55OlbiJI
obRqlxlkSJz2BzmjbFRAwiK8QxMDf5RNeSE77EIjecYgPI40sqhnExajxDTkjy0Vq0sZGleseCRz
tLMCBFodDv/BsbD9bSlxWbnG1ED7RgBPXDJKtiYi+jq/UIEdDEIYbRg2qtz6eEJncGhLuWAodhof
yYpza2pbddDHLfnUwsGSyTnMVzcDuRyFib9p5hGXLBNRVVWyxmzo8MliAbaHE36FZtca7nWZtISk
NiAP5lTnbV+vMe59lUBa7SZDBPK7P7SmFLU5It3eePq4xJ7qUl5zJuuVa3zB2pluOLDhXXEzQxr1
1ExfdchTwE6mvVRebA7FndQ4FuIV81E4gM5Iqga09QfIPyl6fK0HWLSRfwGZDmBtGPmyZela1BHj
82c2j+Sv1G5LOr+35IhuikD6p/vpRKalRNdpkNKuKYpKpP4p2cPDztsQtYtC1ZgQte8ENo7lgWKl
Sg5flf/ymEzQNfk5J+ond3qs4KfFM+/wKjD0Iu2+dyPDwUZbSK1ZKA1oP3dH9PVCP0DyMliWuUh0
/nyUZDFaY6tPT0+jScT74dI4T5p7iPggqW6v6tWtKLzVtjnZ89KgWLZQgBUtIeXqs2qUZs0aGXbO
4GNdNW4D/veGgKFB+jN9m7UG91A48PET/7r2QokA7xcWV56T344LUx9YS/pJKY96aU+0QV+Qr+0G
YjRYzc2v9e8MaRxTBjrcXhWCDJuoDTJ4aMdfqHUkKCtFTwgjKzSKxehaFSN3Z4TM0QAFZ9/kbuVq
ot3qJRTJUkn2ElwzjdV5gLUnZl30NEOjb9/BiHL4JyCZZXktJi36X318RbL9KLxzSpVXye/qtlIz
9T9NANRSUZNT2Jgbhhfojr2Kb42HPMnokc2yKNpa9zMqIhSyjX735zykPydqL6+Xx5pNWnYVhUaD
cT5ww+JP3iMqtkpowr8/sKP7OljT82CcMLgZ2xy+8Oc62qy8uJ/6jF5/DBYP9X2srx2d7LpLrQOG
kYghVo3oxBhtzs2lV6y/Wnnv/0DGDyI3mVISF4vMQkd8KPCVMcEU/+U47LZbB5Obc8cVTEPGY3P3
eBiARnPLRwEe9BaE7dJpgUbG6+Uk3OzeyCpj3SExSGQoviBHiFQbReIIqrvO6+LB4G8WMvsThm2f
k53uZCSjkH8zBB0ro2wn+fmQdMD+1G3KwSkQmjgSphAXVeaVBdzKXgjeeooN/ZpA8kdOkBSutPIh
tSlIySDu+o/CIbJDJjtBi5JDYCBkC0uZRGaV4aPMCPiUWO4TQVHQ/3a65/F3BQUWmbEQz+KiA0qr
PW28DKM7czCXwK+U/mD0P5kqlhlkVVfVeiGLtrDqGVrYNwbs4QB8YiMKgSQbqgh96n8DCGj0repB
frcyNLkSXw7MfDh9LyLZDRwXarng6ffY17EgJJw+LIYm9YwHZZpkOgwzAw91I/FO/3WXbMnE9nqn
+XkdRa4TsIfWPFFa3gsvs2B3pKqnZ0yn2PA3YnfNqW+AqDPPdOGRPArq5F/Nf8NjyvWBOx0bHeq2
SbzwkRS6ykTk9OrLqPorqi1IWM5EdVBbo3JqEzf1UxNws+Zntwpz1vlvJqPTJzcbX9eUpLfHHZAS
m0dOq7E02MCUy/O6KwB08Bu4acAsV5YaglM3mK0yqabriTEpun9Wjytsg8JKDTBfZZyTvj0nHu8Z
GQocdaW6l2FCJlIxV8V9evFn7pyALgqeZmQhuNZvkQhZLH/4d92L/2ytzZRmKLYKe7teMeUQh30W
NAfLGsybW2rBopyiVUsYBsitlQCs5AOxEiPiLtfyzeHmk7IS3yXSQtUgpjT0Oc6aAo3FFvSuZtKV
R7Om5M+ii3l7+D2FIGuJrwCo1zukiVRD5V7P4wKudGrrVvZht0hupFXRU5m9sY2S50RLGiHhe1ku
s7rP7RKF8ioMlIhC0SopYFSvMf0lBwn0Mj9cRAwrWcSpRTaGMz3pc0AdpOe1G2rh93iFsSqpx6kh
E6gEcFnpfspx/OJxmgGviaZvx7ZePGLw56RoD2sefeIbWAoc0s4tONs1H7XWb6Yyvi5lIUdxeQcS
jc5B7nR6H2EKo9imdcz/b0E8Vxv2lkc2+Z1XiHAfsW6bsHLJFV9tGbKZKja1brA5FbXa0J7qGNIk
35epNdXofGmx58WFMHfGFF0PqwVRAW38oEwoVwBc6UOanS/ojpQzZWfPCJQ6LAIrQMtJkBb6qOni
/M29hYmIOVXwMIZRnMIWZAib0Q2MDdaBOtO9KLN/OF/MCAxNSaGbotj6JwIafP8wd2vk9amkvlp0
VqT/OpiurHqSDw+hwlNA0UVjtg278g2DqmH16pnAjo4Ya0zb3Ed9/h8ncK6zRgSUMTg0nC+FN1N2
LZn4fM9FHvUbGoocy5ZyX4ohpTPjuvKH2qaZhE8edNzz/qf2Ej3H7/hhHAMjoHatWqAnvrvorFyg
2JbDyMNCjj119IUuzqICnXD+zZebLOkzoUeH6YuOfi9uRoRcDm+G2rrRyoBFXafbPLkxI32qYA2G
38d0y/S9HUxoo7kURYNYV7xOW57LdtcYmFg1s2U97tIjz41P/2xgLZqXD/GXU6v1mXFR4jM9o4FN
9V53q0B4wR2EFGb0Sijxta71DdnV/f5RfbFpuUO2O5tOZ95Oq77HWDySIQA94BnrnA9zKHonoYJg
VK/7pY+HWz72pyLoq7SuS+Cpyd2Xwlpb9DEB5OylFK1TJsjXiDvZlzQ3E5ceCKrX6WxZw1L/VQJ3
WJswRabK7AwY5kxOiJmV86JW7aJoRUeYYmRYluPBHAhyGFFwFHDHIUIPV034eX8m6sTXD8sbLRd1
VeneVSIubBuAu5JYknIgmya9JWR1r8704vcFg89ZTc1cUZi8QlcOzzIbNqdfD9Ft1IjQmY9pGD65
LJ29CDu6TFtFuTl46cqydPT4G+Y2mnSx/e03dgSZCuciR+MY5/7EbwvNUtN692uH1VzkLAbUjPvn
5/lAosNg9IfgVmccqAx6GKzUX5RORC4fQoFZrMRaXaZzOTtdTsA3PDOau68ZvHBagCPAUI3ptAJc
hHWyUiyCN6PIezKUG4QWwUotIlgZsTPEujdr11Nxirb87Z07N0JCDVVHu2GYQJ1QzZJk15ZQR34a
gUakPpQCn+kEjJW0SM5Wl9JNQ7h9y+j2tA4xcc8282R0X/1NDlerM9LpWa+E0vs/PxWNH5LV8ERJ
K3LBWOidhcP1EJJyxw9Y0UOJ6YhjEQs5pwelw4SGOR3FrwCUUkHDTtooyOXcBjBf0wOSg0QzWk7k
nqPjht2Fnm84C2NcaXXtXoNQlfhZX+ljCSEaR0kaXTKNSJVjBpGmu6sjkJr6uEBZKEOf/IbQPjZz
q/kFcRD9Pe9nCELT2vSNjsM1chNTV031eP8jyzJVzWryFPbH/xX3nFY2rxYFa1HWRWByl8BjI66P
9LBOK6z+3YeZ6lqHAoTgbaljZbUfND4Yjuechh915iyqLgroUrIwyzwKIj39rG1hsxeTeEJ2yHST
igB1COZ10IjQwtNbInmrxECT98eLd/5hlQD8WhGuZqBXdIm9P77DhHp5tHKFt2JPkL51J0+a4oSt
eoixuo4shwi3tiU25a2a+NHD037GCjUImCVdDfS5RKt5PkTpf1sj+c2s83GdIlDetETe93JvpnZp
vgI6VFIRJd26/YD2ni95340S+jkq6wME5ziZijQsnrFdEeTXh++Skvkm2O9E1Z2KFXS/MXc/lfaH
m3hyz3gEj8zhNtojizYXi7D0+na+LE+UPBapl3GId5pm4TiBbB8Ud470SyySFsjLoqL0l2fbohch
gj+1jUFt5S9ikxIaZ0cQiAPVBFNUomeJc2D0Cg+8ZljFUopyoFpLWBULxRB4TqMaZOoKn48j4pHW
gi/eXTv+oF/eAcYRXTPyD+hUpJyi0PFfwJ3/eAfotgO/lpTwAMQyEAD8MrJIxcfdOVc0xVLiyOKx
dP1jFNAMS9BqKdz2BCIhcMXJrtH2w5naxONVtYpLW9D7DgFLqzYtFEZjK91ZRDG32Y/r7l0KGu7z
ULwYI85oJupiayTAVDlK9VW5fHsglcezbx6MXLpgUyV9N29Ii7viV9Zz65P11oiiY/VA4iLHbJun
oKOA42srsEpGdeD0v0yIDMHBB1Kpofgz2nTsNv5PdtKHhn8ZAnUrQ/H/EgKJj+7uDOJ4DSZscxew
lLlV6Fwycvec86W86tsAhoC6KD0WqikDMDubQGacM+bszHU4Xh34cOunD5Ea7CMlbTPIxlnla+0S
p3Th0KTyi7j3lRPXz7ZEir/lnzF0SkJhb457b6fyIY6Jy15aFIx3UyGOPZwEmSn628W80zHPN9iJ
y+dMSN1pamoyl+mCKsuYK79uk2rvvBUmsoTBDjMGz7yoOfMLomXRizZHQL5PQD/E5yCoZ9pIsre2
JHR5nCkb0hnR3jb0sc8LuIpi7eFs/UYmwhqyWSFpszddM8+ZglnhjFsVGit0DhB99rn8xaIWufTK
UjbY7NLf9+36WnjjaHyzKH2VZUhptz6ePsfnjGkxS14LUwEG36NAP0FSn7rUCULAofTf1O0ng4E9
EV/6rmrTTMkR7vBFzIo0aTSrJeKx6JKCuEWUjLxt6a5RgyW2MEBE4SYCFBXwxS4eQBGJr/r5+Vio
85dPsc7x5IagRAwtbsnS7E7VGVG3u6d/hKZn0GAFkvr97V7mXGsu+C7CAOZKhuQRZENWoKfvu4N9
henA88+mJe2l0Ahv6/4kuET3n1DFr/JbCvlvDLLdsaQHSJaq8VcR/VymF7q2sCWRLnrHLPb4SCpv
U22T4R4yr/6HFpyEHppSt0D70hmbYktBPWtO5wVa077FyCGxiNijBU42omFIk7+eUlXuv/LrZOiU
lgKmqlxsWS4QChe1i+pv0G79Mw7z+eIrEA8iLxdaxuiqatR4Jn9Pl8IMjE+pdVKLacOhurpXmSwd
PY883SAwBwqpHV5DBvmF4eV4cdNxNnqZdZqCDgJOQ74rlzthKPMgfptnuvdCPUF12+YcsuDXkOGt
Tp8TSsGNUstey9Mi533PTJnbOfRUzZExa99luwA6MY4Ljva2lWfwI9PHV+nXwbZNLAgCQnZzFrcl
M/DSqJIeuDonHkMJK7kuVWXTCYJ/T6wFPgTzcs4EfJS+9AIlV0eFdSKlu2Zli5UNXqxzGH7q2OAf
scWe1hozwlnSXBeRYOttSG1FhXbvnDKx12oiH+VN2yeokILhx2m9/zIZoBsXQCUyCSzxyXL/+O3P
B784zb0Ln/TRA3BAYyJYJlgWGzLXhr024BBcMVOgS5eyFnZuhIAOm3VeGoGXGa4fOO/pAR+cPWzV
R5gp9HkVVs+mwEoosoy9ob1cYRxRaYabKxV3dld4GBayAbwwqN6crDLtXeW+3aA8jMOoeOTRzR6M
6ezWfA9iLk/FZftnR57TlCNswur+WMgT83zEhsSCyMQPgn84W6OJX0xRlbQmDoHSAyuHwwQptrPB
vQ5rRIev2Tz4xp6FycV1LMJNOGGBp2RCHJfnA41iovwWTo7DUHijtCQdPk8IUeRskKRht4u8PFY1
RAtNVEM/6JxJK85V8mnl8TtJmKd8+sS+CP9SuQvpDTDTIe6LNZ2r7NTUuXQXAdNR2m/Ecznj+B4E
kmyq/OTe0ILMVqLGgOdYsXZ7pybhsGzFKaqneY2mwvFpZE6UnF9fuaxwKodHHWnb8VhdVkTs8Ql8
NX9a11sVykfE+KwtypVXhAhXRSwvdll9mgxIxZDeM1AM/97EHjQSCf/sbPVJR0QmrgA3wl62a9KI
erZnJh4iqN0XFSoyoQ5Ip2rYvV2/LG8ZtGqAadRVCgRlaIsGECZuisXPF4yky91tBZoN2wsn1/4C
KhEcq+VPKDIE9qgkegdSxg4lT4JrOWtUPr0NSLWm9KXu+hhv8jDBYLgJm+M9k+tyX/P/8DEEbrzZ
2XGy3Y4wNHeI/ZNeh+Mf7VTuJY6OykVyotqR5QAY5CXCptTnfrLc0SY4kg307qiEtz2Sqq1HJdIn
Dws4WbFPxr89gp0etsoLqRWD+5NipY77l2aa4t0EXGjfVvuX84BRxEci7FsjmTaNawfyk5R0MaeW
GE71xvRzApaO6lRjgtqNM1JT9jJI7Chbg5ACCOT0FJtiAhakxwukJ8Gq3zRyIUeQzK4QyucfVKHu
33JIQjzR6rFGh8oGDPS31c7Qf4a1sFWngvcDtaVLKClf4ZE/X6+BkT10Dvs4GWFcOatKdQJWvXja
CU/RQJq9abC8ovIpLF+Q08J21tRxWmaFhxzkboVSiJVq+s0u5nAujFwCKXakUet6ENXgL72EuCjd
j6LYtvpB8o/fER/doI7h0D/HzkBH8kpOwy3r/hQcm8CFSskJ2astpA2TRWc0WsRpeH5nZj6fTtfv
yJ7BDX/iP68dRYct6kheukAcx98OZ4yTKbPYq2Sj3+T8HI7COajktWvxL8+X8rrfRQmquDAaotnm
BpD+IxZ3tCyLll8i1LPWp3FonuiiZucS8D2lK6oBaIN86P9aIbRqADRF0JPIpFkKwVW4OXavtaQ1
djGqMVey0svRnxVg/RYGV54sY9HjKXf+3C66zeQKLogpUwgoZNxPJkJFxjZzpDhnTOlq7eC2h8UZ
Zn8h/J0h7IGjYOF5uo4SqG3L4p2UOuSP9KX+snngrzLE/eAmWv2ULLqZDC++3QkVZ23cHXlce4h0
y7hOD1fcAbET3hdLu9zjK9iDa28VgOCadznkbdxVoYtk8xRg6AxT0kVy2xILej5xPBRKSSOw2Kzs
2La+25WZfp549ZBwrX0P8ktFNnlAs0vfIEXDA2G0RFZtvqlr9s7vImnsD4cijFsVxDY5uTiCqsRU
C5ZpnWeQoZxhXGYuyDFNisB/dN4zSLjV81th9LykMsx91AjGOMuGxziPnjSbhmNKHnZM7KxNI4sS
Qf8QxaPr5A4tFnoz3AqnhCDfddmlYpoWz0oTdn4zg8ghUO8R/l8GaQ4xqGFfDsrWHrXSashdcpSj
k84AcgF2wj14hyHyDeixmF6dMjB/3CupPTADlcnPSBPsM/zC08qLzwzPHNQqcJyRzsUvLCUtSlIW
wFc15NZMG+zxmdKpLOzN6P6UoGVyFAxWeesFJiU4aC4KT2gj00g+0y+9uGFv+BSgyoX1x+Irezg3
OR+W1RKHZP86upfZnZ9bhMoKQirSj5tFVIPKt4wW2JPRf2nhpz8ZFAj4oN6Zjw9tb3cwuKR1kO8J
MxcWbREbB8upXkndOhgi7bh9i7d7q1o3M1Q524q6+jvHW5oFmbF6dTCIXij1hr7Pco67oooW+Mte
9poA19mKA77vaXNNJA9IzbtGem++gMu4WeEoWlXNitwr79T5WAiu4grOH1BkKPM9zPoszz6/RfTe
5OmcAoLINg3HCKXietLOHlO8gQYAso+vY0eDFr//vLodlEB8O45ACQxr4xWt+RdER/lZO3DKYBht
yW21PZOyOcJnM2jS3F01/rwP1RkyMpmmT/D3fEFlAmJb6LQOKNlbed6tkD5Q5kL9qdCPx+VXrAas
7xWwQ+KK20jw8HfpaXz1Lvc6GGikvkGXG54hWZfBnSS7uQbXx/fwzvxts1my26TgS385V8p8IMW6
/+TofbV1qlt8N+sbJS+MBYZskn8mdFzOyKWjvscUVIyQ+V9NqzYVL7gmgrRFLQzWfw/13GA+fvAD
UMgzG8il94X1KjGkmQ3Ahx2wQUFxUOEPMHK/ghQ88o9WbU2U88LxhW2WjdTNdvCHL0Yqx/BcQvhX
b+JA9/RmYysNUmkbQTASBFknFNXGhLXJCQLRPbA5+b1eoZ9ivxkVHSEW9jSc0m5bTljnfNy2Bvdt
kq85U5ugqTnx3qRM9fjZt6F6QfVA7Vq8BztKuVpVSzB2fGw8mH20XwTuk8OzqyjvEiTLl/zPaP+2
T8aDghi0gmOpCVR8vkE5F0/GVkiHTQXHc9C0DFkPnWdlRJIC6A9LD0xo6KVETzgGDKoXhaYVdHX0
45nBx/FgN9nmlndA3ITXCWNTISy48WXBQ20jAXWMldLPzp58U0RH6QpJUXTMAFuc+oRDB47Y8tz9
s+a1Cls0H/5Q4oooyvcxkL/3KaFIEOgF+YNOKdxcG8YZeL7Nc1pEf/yXW0xwDb+1YN67KgcQ6An+
1utTY2eY5JkfpJNAWpRcpyrt6Jox9S9wV+um8C0FjpuYPyGak9obvVWDQVgXRrpqfe3pRo0whSPg
r8ReaDQf0nqEmjLaWUk0XjjfeLdgjEJ0adltPz2vmGuaptrQdVpggDdhafPhQDG/1yPx3X9hhqjY
l31duiq7o1LUZlawXG0psrEeVtZeBYyTq6NOc1SO1v7cufxOjuzAR6TuswhWg0CVinCPdsHiMdBO
eAjvvcnldGQaMQ4qGBKyhBaT/Ol3io9zdlYYV5yHhDoEG6fKvwXkn8ny3tNQDYra6krYrURO0b7E
TQwKiicZKJUcfMq6tubf7Tyk7eoSowglFFYOm5xYRMsdb9As+h28++ptB3ifVuS7l57oaKKMs4Hh
4BI/uTdwiuXHSs4+Bdig3LLzPLSqHguGCrOiLLdm89AXOOVkqudf+JsdnL1AAG0Sydce0FHWIn3V
cBkOA7qbq3Z2ZM49erj1vmbdB3xGHvK5OWOYHmBICujgnGPxJE2ocbLTHWiyYK0JyRXWsGbdLf3o
3lDV6wgmWYljixUdRWdQ1NtkHmOUICN2ToAsWhe4gzfLK3Vj9oPxG2mqLAaz4H4ffqPFeqSiFWK0
2Dm13SFPpwYPLhHVsBNf6ptFSWMBae+JpnNZel7hegBy0DWIHCtb4KDYIaVJa0Yue7YshurRXAIe
LSOu81K2HEjimhAVO5LbXMUFJ++u9GdOqw5hFjkNxvXpnKN+vg4HUw22WijlNREjj4Y8+wY6mUHY
+6Kf/9qWe08q2mQMwnM+3oJFKQ3iCsyszE71talqclQXWBBD/xfT855eGeU4psWuzZgL1Am8WqVO
gOZtW8ygnaPEkihUanpkzwoo6rwDfs92i9YWg0kDCRRaYqKn5B6fcPL65dnZh601H5GvpFD9U9fQ
g0vT3Fua8vuW8NU4ONIplsuc1F6NdCJLMH+0glDjtA9Z1r3l4Jry8LGw5g0iM3MdcgSvpw5Dehpl
E0qtayPmF2dLlO962LqGGZoyGAwnJ49wwvDNlKgdOpsfGu9kp7y9Aw7mhzaMyK6uesfTEkCAsELe
BVymyymeaMepb7PTWbW7FR1L7QyTzxwSpn2FqnuZ9KjlFuWDVDDCRf7kvAOrVALs15cBUSoY/psf
Jh4Wcjer91ZDl7xxDaiOMayRD0Z5KNGVxDOW6zKg848I+3dZIO39LkeS94y4ZrVSN+VduVTUttJA
nIwL4eQ2W08jsN59DgtNMxKMMltKwq6t0N/2RkFrylULsE14mfg4ufOedE+1QPJnhqNnOgnbXl57
X1PFYONZI+1Xw59gJd7Hqt7ETH1pxe9gTUmwP85LEVaRYf8XU8nc8xUOWeoTxZjEcjMgZa+H53AK
X0Nso4yh7HjhM3L+E1O7rdKFQxot8F36M+Xg3XBt3v63p73N4h9xsrJS883jggrlJ9N3CJwHjTDH
+xaeh6MAHl+6dltmDvJ2o4OYZMjNs1cERbT3h6OZOoqyzo1r0XxCRvW3b1zoCp+NGJOs3cp3Sie5
vX31fPeg8bnbHRW/ogci1hB0uDy2ctu691q4T5HFnCm2sE7Ly6NDFzZg9tJ7y6Huy7bV2Xx0IWWU
c+Axog5GCI/Q/puOamUiTRj5aNuRdhuoICALjk4vkgdq+Jh4CtSEGbE5Ui0KAYoIbrXlKWG11TCK
S97CnrZjiBrUF5geQCbz74J3GVDT1eq6m+K6pSM2EEE+IwdKdUjeouB9c32RTyN5+OhVNZQ7LtQs
YzKbkW1gjJNobJvvUtoXb3cVwZEsWzTqoQEHmpBKQnqNOirifbCO+j9xWHZ5Fc7f0hLeB/nZgx4T
VZ51yDEZxwVtZrJPRY801Jl5iwAj7cBmO5Qot/bQLpTt8pf16liyZg1WCdQVMVUEHC0D8dI50Q9N
CyeZqvgSxVS456yeCNBXUjqtwsGplD+5LpmwOIrzGeN4D3XQup3vD/8TAVNkJD6f2ofz86g4bcjo
x2iJgrQY8iVDYvcLqwF7W0HVWqRVeifWA3ErB9Rzhrd4EkPAhrSmxqhEQ/+gPNNs8Gy2kbyPIeN9
HqK57pYKXh9sSFAvD4dXvWwD+rc1OHMJL/Xvw9FQcWET28l/wnKZj/2Yk+IcpqhT87rV8BY2nQLX
7lBNCNIgL6aIpA1tUZphqWSuHrV9oGyXuzLAiLvLNu41Hp41gV/nOBrg5BW7u25U3tH2lBX7b4WF
AtjKyZKmMpENyRSo+1oYRSZ4UWlPUHYzrilOrpodQE5shNSkSwlNDlSyJwl2awnWeAtLOUK8HtkL
zZqkT0LFOhqN4TKkmpEeYElCOCGqTHQykj+YK2X4ppZcYEwgHiYqpFAoCnxECh8WQLW+fVdqRq7N
BlioqI7JzZS0tG68cze1njsaTLQNnzq+Hs79u7CQFFGak1bbDbTj2Ul07sfmlCJJGa9dgcyVhXoh
MNl86nWdbSWWd32AmBrILR+rRZ+lWv1PGurypZeWOYPaQrxbI1i3NtYhdWw4yUF1+laffhjcEIGr
6cAG4FGrszaojXL8KG2YAyHsnKfUqBwaVm7GtVsD7gYsd427DK/1X/tnxbDTT9Mink9TyvcQhTsX
Q74ueFK5Ugzhs7JaehQeNffPndnxNr7BI5Tsul4eX5bD+vnUbG9LRiHlvfcaATuZmX/b5jhG+74i
68OFAuVVy92nGV02fxcewF/RKhrsJvhco5QAcBEnfKQVhTdhJrLdolwQiSfSCV5Gmu6V9mtddnnP
hM5iqj2OI55ZRzYAJI4/EGy2ZGRE+VNpkGAaY4TuUTFulxP+bip3hEq5Zjg0+Is+u+NZYTNGDCB6
yVj/piuj9xI3O8WCvu76gK2BRvLh2eXhKm4am6Bx/tTe8gJT+8TcAG9hTse8EAF2jSExdPXDI6EB
LttUb1J8eIF8D7KfZtMlcZIbYxCNGQUqkvxUukOxuLxaOCq0BKvph6TMMO4tDZ8WmGNAStVecTvL
/ypS5o2o9D7HYJK0JaRfsbYuko3IKO/AOzgHuYmcuQAF4qbXMc7+6qRJAq4SHU2Mj+wSmp9W3BHT
KN6wyGKhJ2URDrWksUY6PFqqeiQqu5PJGknS2ch0WpeV0F43QvTPucWW7nsJJnVtZ9HUyOSSeIrz
MbVJ+4Gsw+EAaR7L5XJqhQSOZjKffZkByeGbcmlsEzYWmMPcApwKVHbZJ6vNuLwILZ4Ao0IqOYkV
iRDLiMCgeTv+qN+Ab9LmU75ihQSxA4IpxVpcspsm/f1oPw33ME2kDBJdfIwK4hsKFmgNFU4y5HLj
Ne5uhVRig3dSjPKZ0xOjT2gC3Z5VeC9fPglVf1WW0QBl4yu34ic4K4fz7UKzBwA0iO+qvqOGS1fA
kinXnSMMsNZMXvaZl15db68K4ZSm+ucsbXYlk217e0t6RTcvSH9oGlcnL9dp+n7juWkiALOk1S9t
xj42gVAxUj8gY4QJxhkkusxOme5JyCObr/NK3ds4M6RQWKyoGynABMHZZCfFOKCoGuvtFngtqZNH
MKq0siT0DKxB+7xkdX1j9ScCDzn/yaciZfW6b1sIJiKgCB2fuR/qn+CBbHAJ2ETGCAX6W6Ou/732
AW8sdrpwPaOFp8QESmYqrKN8Z78L5647epRdKWU5uPElS9eL7w4tn6peuXJpY1o8Ho0/IzzMWOv4
wr4d9NYinxi4cWPGIXAc1xIaqPffPUCy/PlDaKVf21X5yZqjK45vbp51NuXyP5il64zo36lk441g
KAXNp3rmSbLG3M7Ajr7i6V2STJRfCdI7iIp1DFP43Er/+aBppSiMyNsPktTshNb5sKAsSigbMp1Y
PtI3i8i/8INXH00G70GN9G8ch28HVT37qeqMLD6jXRV5SnoZsUx8xV7Jni67e0WmIlj2+6YqEQSO
yKx6cy3DjJP6hKzQTblaq7seV8fpz5oNO59oH9zQUnt+v6NCFUXZ8oQyWLbXyF3jpi92+1XLd8hC
nifL2V25nMp/uvuknw9GxbIFdfoSzFg/KN7sdgtDJ1GqBHRKUuvQFkIcEwHB64fO3GxC0RAnrlk+
dqRUHYIyHmQ9CLtDFKLCLLipoU/GlvC3x411ShyewvkD0c7h9Q/ItQtNWt/bAhiZv8bqIRbAgyCM
//+B4iIw3OGNMNgxwMZZypd7Js0VgjmFPLhvpnecFjEwMLdKZFgeT6FBTaq7XLsHfLWbps6gXTQd
n7A+mBEfi+oUxIcgm3quB491h3yR3A0OicbyPmAr9CMrBhB4W66wUXyVHT2edf3jtukuVKspTa8o
S1P1naAKlECR24EXwoqoPpLP1ldEeqy0V855t/si6bkYG8Mkoy8H6Mza7Ooj1u4no5emnv6D9r8e
HxmqvA62HFPeQ1uGXC+pmbimuMxHf+muwGONoiDI8WshCLQzCnL28tRFwBnbOfTwRxK2SHoGWIoB
DbEBlG8GvKGNkHzdsMVrMfopwYOWs9Us552LwuZ4hYhD0GyEE0e2rl4AxB5eC2r5PSPrPtDh8Os8
xmEPlyjNACcU6UTCnohnvi8tSZNkA5k/mNIsc/ONB56t9ou6qvCMS6Scx91mLaLMWpg2TR3gpEUU
jGfNXrmjdpvvY9ICNkQBqRqRMsoiPwCO2ssiPdbsppK815tSAulmRGCX222o7EauSFiWnU83/H0E
O+hZdEYy8WXf4NMKpOVs7p0wvfY2ZqVoHcqXzF0EPnisssnM5WlnB3MqsmB5EjCro6t6GudJmpbz
bcdDtppGnfGMGp7S2WcduJyNUpJ5CstBUJG/ZTs+6vAYItoHIA9iepQDk9qUBvLLUXE6GOk4EQaJ
0a6PV1Pfds4xgqR1ckQvWosFqx1OFcu8EUXqmukdKm6W/yJKlfXIadtTy84x8AtXEmcXlamtJsBY
UISPGUsqNDEjtcjxwN7OP236VDP5sT/C+uk6z9mKvIZuCUpH8zjQ7nQrul8004uJLJTpIWs3qI+L
06jWABXl5Yc04LeKi1uH8H/vFUnQXHISptapMYxMKM6IwZ2zMKVt5BlC8EDBXxG6q8CcKwymGOln
JVTyK8y37vRckMA8s5fW2irYuW4nJXErwGH2NrnSep5cdTqe26W7KAr+4EmXK+nKtdHiUs8UbBAg
f72aqIJFwa3aH0lJbMHNSGZch9onZb2bBjCuzbM11l0WAF3NqipDOd04HPRWj7U8jxoidOmipp60
mTiYUhanUJUNI8JW4PWleQvRNWMErxyoZCoUaGFECbdPY+Ip2K9+rG9VZs9h8q4iraW4OmNsH1AX
Pnno/DOAAT/ja4S3S4k33rqqTcf1naCr4Cim+epelHJv5ssHW9odLs0IIAJ9bYPRFf8yeGdMrPHO
nTOhw1he5whuc8pnpF/KdsRc/sFjadsTx0nWygvB6zvS7C9RO+jxiIq+2jJc7ISxrT0OWFWAMiFu
7BxaBAVnpzkFqN9ALu0rgNF/6AepsP4xwoBQ29euUWuX3ZL6UsTKiGulKDaRZnNkaO1SWyjugPlI
T6sGD6Q5IbivI2szfNGuchqJErAPwPkqN2GLEPyewFzvhaYgKNHB0KwdgKMmcK5eFcU/91mD5bG/
Q5Ewp1EcNIlAqvjhYTYeq4kK1pY+5frCoWepsRiZ69uaWqijhHnqHOtR4KEiOmarFt1LFZ58Wemb
198UTesvALgNe55FjGGbrdbO9vHZzOGDw2CP7vVRSiLkaDDivG8HFi6k30EAVb0J3CZGdfzrgeKL
MMOZSHDuDMzvY1BABIYdE8Xb1/RDw9UxspbdJzgDvv54mTVXmNQkAv28/H01Hzbg6snQT1oOlXFe
VIul+u0T26ehA69jaq9bBJd+psoKF2Byvp7c3BOAeJIohG+YoWKgOFVlkZsOym9h19crhOTXifYp
yS1iaVW59TH5j38SDsMOMAq9LRHxKjuVaBSscnkZfk/TJ1PdJFwp3JCGHMXWKXrzLUDtB/TOWI1F
KxSfQDkbe71jCCfk05hONyk4+w4Sq8agyKrbUmTzyEyoIQbaaguvDGajEJ5xpsdBVdKtGepyrOeO
6EbthtHkZtx4OL1vg1619ugQXdzkAMApDE8YM52mnI/LgczqLq6Z3TBPCuCidR6yyjtxPq0CIFvL
TFFb5sCiCkmUj/VANf9KOoG8wFrAx5Uy8DoiU70uAVRlm0Yv2jEWG5mZs3YrLBS0UpTC7Pj43awb
MXVXcNnBwmFX4Zr151UizkJb/7toquIaw+rxcM3UjpYjjiVsvxi0B1qjCK3X3KSl4BhSwa3qy/Jp
zwtsAQe/FFUEmaIMooW9YBFHoLQaQEd4g6yfLzcc4gp2T9URzwlOzmPH/k2uVjkuep0CjfwkRd1b
3NIC83f70f0H0YCV3pcCmSdfYHdlBCzYndYg6bXvJk33qUMB5owWfYAUhhy2zFmSQ09ceW6xkuyD
ZmYz4HuQwAq07EQO6/qYX4GsQBsvYJmoO7CDlr1RfIQBEOO04JE9H8m0y9VX2p7I3a/yLsk+PY6O
kbG1HPCaxo3Ej5K+slaKMomN2n39CDIbl8CygemEZk3R0m5kLIU4K5Ah7mW6j/+K+DEeqSAZ9Tny
eAWRwGGTnCqh+WGMnbUI3T1YCcmk36/o7dMUK2YAsjQl1ooIR++dWX4QF+BCKbahdFKw4tLWSSLH
RqsXW/uw5lU7t9JlJ8gw8+/vHUVy5nzp49ZVeWpEykrDZQjYBXs5zh68WUZoZYoI8McQJNbsYRCs
Vcl1/dgoYY+Yza7y6JD+ULYTZQOMndQC9IK+lBjtbjXPi/daQRD98ZUGv/4ES1zrGasyrIQ9kwII
hvpVlpf8rp1/2N+01jXciXygaBB94PgoYZO5ku5XEN0piroWdtl0rnh6+0JyANAuwj8rwV5MSj5C
Y1bHRNM/KlKJXJJThFNGMXCgt9B1054qn2M1CXeVzW8KByWcDkc6knM3JUAQ+BfUIaQhqMVwwbbX
C4djC9Nhnk5BGKTgBB9zBSjexrXwkoBlrgT/EyBJQh1yI5dN29QQCa0JKBGfxurjSFjUyhUiBmOX
dHW38NZD9rO6vEI9Dw69HCRlwOOGfv8CaCSscBd5gXnIkFZEjk9YdfGk+IaWrghQU880vGWRRl1E
UngzZv1+Q7YZPwhXba/8SsKKWtXzGWW/8BXX2v6qLVk6fW5K+bMSYqvZf6bn0/XKwGCKVkyG7L3O
hzfeKWm6NqyBG1H2Edf6xbjtto/O0MSEjPwHm7iFtQMnDj7g6x8sVJPWixq27jBwmsLr/SzRZMrM
Q9lZ9ZO8jxNasf+W/eW7n6y7jNXBOz5c3WJ0/9tMjWLDKA68OsfHJbnGjJRUBVI2CGcTZavZV1uu
B7IBjWN0NJznvfmeNdMZIQAaiNYGpBGX9K41658X2vk5sYDj6okSdduzBJxCgcknUlxnhkysnngU
JxmvD/mNXrcsDuEbNN6Apb+KeKpTSP2NyiD3ovxWRrW0HdPC5rqY1rEcEdDxVHFcaCLNh9xjnkjn
7IKYMmDClzv//vbqHEopKBsp5G5847IQhE7oDg+fppfAcRntwnt8iqDlObiagfBA5+a8l6aDQTZc
saj+8tED0KOch9wp9KZY3+s/gOW+S+s6w1tFqU8nDpgNEte/4kK+KEtr4mljpCnUFIu+/AkGpmcm
29y44nmIXOaYY+1ItQJbMSIwEjXRu/yJeD/LazmUNpPVyjKdpLawWIqVPYlpAATO1t4JzDL3g4kg
uxbvoK2ZzAIH0aTAZbjmQTFCITStkk70LmWMxB8hLu7k4rRgULKKyot9jp9V8FwX8kNzv9+/bKF2
pdme90/0SHpUTnKUXIMjPkZs1mpfq0mBQ6YwtWE3NN9zFHc+M6v2R+SJ54GadYHCnwSWPP+shv/n
G9QAzLFQRt1GVMixWeytm65+JFWs4+MIYTMdJgETR52uPdvzF+Pz7P5j70+6uZs1mtz1ITPXCAJM
gABoXKUsWCRvhL1zIKdRzzVJXIna/fI95NpyFXrO7aaE5+hqGh+vN5z9+JZmaWvsmRpUbaefK6Ps
6LwatlUMe7T4/kdiwOllLQws10S21GxBh8ht46wi4VhzEq3wZuDzenGNKKNXUDqal0PjNrjG7cVi
jlWRZKtdED1vykUN2usPrwRqGnw6n7pERRC7rfB+qVrDnhe2utOtdCkfk/5pewPUpgXzmx6ARCSp
LwE+0A7csCwZzH1rIFfJyKKvvHbJNGn5//6HHpXzvc9h/LIskNB63mYxJnfxUxiK56+9C7E+x+ds
dFUFdru4O4Ctor5SGdFRICmvPWnw+nhQGkzKMEBEnXDyQAahvclJAIocORHozlLKiRthMyCZf7do
lwHwl3SdqwQAAUWxuU6rxKQfDzaCbtXA1wuIiNcUUSG1uq5JzCij7bBrvoeTUdmoaYANsUZppxbq
YgeodV3o3BcQbvJyFG7vHdLWKqIxh3RQ+eN0QC/h6nFk3QNPBbzJ2Um71w7uehZpKvqGUKeoohB8
a0erVKEOdGg30Bglr9BVgte3mx4D7oU4w3VXbadXc6/pLx2eSxampWtbN+DyJKtesv7ECQV5IL9z
tUvI98EzggzZBBv0nqHYyKeGDwcWoRbEbo3xZKFYu3/6Tv1IIAXfMenXDG1w2bTPj7cmGctVunly
Ac1j8ygOPxeE7Ed+FXfXkSZm7QuoiBH8lQk5RIyWO5D8i4D+ZIjQccwyI64OtHIdtfw/Z0Rumywv
5kNz5+UW2oQx82YOYpUmCIwhHKHFle42iVGrkIXGzt6EbPSejH7orB3twmJDPCIab2Q2MWDN/rUt
mXe1ssB0kyzP6v0LM80q/j8Q4C9iVBqAl82QZTHWA0lLfm6PDBkNfevsuSwMxJIsRO6kVV+w/jsh
eRlpjH1rDf7dGgTEkhpoZQ5ME65Tcja2oEH3UMV7LG/71a1pz+m31kS5Uf9J0Qq82f/lb7cUCWSZ
JKermHs0GJtBTiSd/Lj+Z+DVLwiyaVjUZtWfviQLZHZsaqJytDpfrmoMWhc+6P91o4KW+ka3PQEr
Bb0yyJsdKKUIl8sc4l1opq9zYQd+GHymimbW4zDWJh5fUlbrz/0OEnfmOPKb9bbAftKYk2H7jUfE
/PMmGCmz/bnOTiJ50R0mjWDutEMw9NjjYKNNa4+bSX4FY+ot4jszpwmjv1nypUcpQJ7G1hqc58bR
z24I7/HnHMoUEE3SNaQ5p8GTbrLsIFPxyr15ECvy42/8eaEMci2RFLfgH6ktafCGnzYX4M9PjRVP
U9jj4dBWc7d22IxTJqlKLbv/bqUW6qlGpzrHDKQRu8MMgGFVrO/mELNpe2D9q0G1MdbEfqJQIeGN
xllyprExZ4ow69EC7YhZ16HpHx2gcJLn+PvWb7o6bH6SjXC5eGuL2cra21pzZse/bvF7h6/vzr4s
JH8cURJx7H8xq6cwULZZEv+7ovZXDbB7aDqWFPwWgSf7WQtHzna68VgOb40b4YO/GkpT5bfjW3/C
Cw0J0DJ9UbejxNB3R0gIx+PXQwVxkpeqfTjgTaXIMzSCpYUnomYcbJpIzFoTrbTCO6jmIwtoqFdx
bwZ3akYeaeZk7voVm1x/CS5XpVz3ZYADxWveLtugR04c/wGLnr1kalLD08pdxBeG3EV7iNxsnPo9
GajMu1/DPhUQrJOFFk6fsWi6HzZz/RIarLJg24rxAW5M071enNfey5yPe+2tSroi9caUi0lHX2eb
Y4/bEZEluIPUk9jDLW3Fto/nMvfN87JUO6Vh9Nyd+R/9pFloLZCC7BiFcWLYOOVF4M2pAD/lnj35
qrLkUd75NRbinKCGuAyOuUvBeopbc5BxVU+bFEvhOI23E9gIMUdEQ4e3saWrBvbr4Fb18q2jCyPi
0j83ln8EjexXKEIyReG7z1LOAyLQ0oGS3SZYvFx3UvsyxGQ/qje+sM8uVJ7kpe05yMamD0IOxnjq
ikoS1UWnTY2Z7H2d5Dekg5DOb1FJGPU5SJGMONUPQ1q5e8Hr1QjSvPZHi12WEJwfMtkdM7G9OBEO
ZQMCf/oAHMNLYKiIx6M7CiwNhATOU2j9zfBZsFWFbJUFp0yzC8DSv0JLM5jRyQYIcc1SgfOv2qfa
NrHmlvG6nj9zkfdAW6Sb5qr8XoE4Gnp/y3xi6fZl8V1waTrA4+gqpoTrdrfD9M6O/aFf6aYtMQlW
oPeQfgv9r6c6FIxkstMMh/PdxXftND/kjdXngZeLse8AcKyykZA7w2E6uQD5Za5H7AYcrQhG0loO
uAgk1EDcfJxALZMIHEEDFe8uplrS1so/bgA/2qmMNp6dWfj8TCme6yg9wc5+a5WZ8mv4WKYEXYZ/
NBF87PbfqWFKp8T9PC7gSyjorZxnrkZL6cSnXdKT0f1jeNJu6p4ufW+LJ4TzrWRs6N7TNEfFUy89
iRNu2nzMXtZz3JLVIBwExwqk1KLi/EIdgksYlhVGcw5+2746FWlva9FVZS6y/jvKv8ljDqwD39Du
xMwW1luI2AWxmZsOz4FDaPBEOXssdXlidsE4heWPeReHr0tZ0Ps3w7DvOnILwyOLscOzl2v4/G8h
8BDht0rpaPp1Cl3WJbnm7il7m3h9n8N/67lpRYCFe45tw5VeJwvsWF901fsouIdPc6k63pjEwcXY
ZsiVcUtALCQ4gVJdPR4KoLGHeYS9splJKPKEX3DPM1dtNU4GfQfzZdW+2h7ZI3/gyDbx0Y0UnKA+
MQ5yX8XWntXUScFbk803tj+Z36bA9tHlRcsWt29UiKtrNSlqFkcl8E8Z9WalrIZ+U50/O2Udfzze
KnTduEordcQmh0J61Kx0yjeCSJvD1HIVpgifdmucvho5IsM/u3/j8qaVpfK0pDdwvDu3oKWo5R3u
uv14kvJj9R2hjxGkDqlFW6FR3TzAZDMYRPj+iHSHVJh13XvWCYEdcHIOL6mOhrFx1WxV4gSJJYfG
GH+PQjIQxuj8RPZ1uZ394C8Zhgaf337sizPhcvIAT8W1GXBa0z41E9n5yLzNtyHMAz3d/8RhNyMR
Qpt4H+MC5PPGDmKiW8oCNzR6A2dLvbS59vjPbWg2nKULjhVDL4jWPKBSaHTSOrAj3H7IGpbM2bYV
2UkYnicCacOeMNZ5HbbY7kLjrldbOBX6SrKMs8vvqWQYj1JMq790H8L7EoL8wWmW2DK8iUn7WUfm
v/lpHu3Q/SM5Dp9xnoZF4KOT/sOTIvVxNAtwLWfMJBap5TmOon+lT9jX6RKhVVVtUPs8Svj+LKsf
xkDjzO8mdMQzEOlDs/SRtLeY/2RFOtDrV1s899mlC/+0bDB82pGUB04TfZlNOeDW6wuIkJEMfX/2
zZozyIKrxRa9aGzk5SPAhQT7tUByt1ugrhIha7vyIZlqCbNZf9y9fyOo8t3De9+l+yCcIMEJ0di0
bp9fZ+IIv3OtUaxWMWqngi56JbiVM4f7GEDaT+AwfBYr7YL1Iydp67J9sZWF+o3mcn9B2G1zOy/1
Gs8LsrN2DKY8fWYRvj9ChdQaFXG7usYw6Z0hdlIWI+Fy817QxdN6Y2TdSWbPP/tiwkbRCK/cs4AQ
ATcspiTMy31Ysdr3ijGTmdHa9dWLLd9C1L6PpGgf+R1HCn5kDbwTi26tHt10c9z5kvcUrWhfzK7+
q8qKd0Cx1zP6hSA2iQXp+7bb7EfJyPJqgr0bfPYSaaSUrU6mj81wKOHAbo6p/r5+C8wTpzGEz3GJ
s7M1fHDd6w5yLRCAV+M2RwaufagGTQYLYFAVQUzQbp98PouPe+cC9d7sdMDymBV6ao6k0rQz0PaM
IHgTZvo/8EV+e8ZeVhBRy1TWn9ab+vQQpdHYyb3MwG7xmmYz6NDoNfwIwF6tZD0UB+41p8C4iVd9
2YtVK3/2/fX4yCfcFyfo9zA6AMAGDFIaK8LyZ8HzCnfRw6hMIz44qO0arA21azeEiJj01L7dgpqu
XqYxu9BMYrL1wduaC3ZWpCkozIwb+eIjWm4f5JWAhJMzSqy7BN47aCLPs8o1ebfW0pOZeuA7Gycp
a3H4jVKWR0lc8l30aohXwy/qWlnvsMI8Yfcgz2SIixc4rpIOWXV1VFgiVHbxR6uFwHocFrBmaBFO
HXipgB24l1vfhxMHThWz77qVWtotgDy1iO84VfDHJoFm/fVPKAOw4FSlEbEPpcpvjdVGAEhRpidn
rk2jMpm+/IRCCdHG0SqcCzwieZFQpHKNESnO/m6RBJf2ifECzsuBzEUf3wZYZ/t00aOYfUZxkEuM
uCt2gATSSz3818GQKKtsfuaurD5UMYAOZ67EuC70pzIY71MTuAins4YScdtIXRK5xHQHSJS82GSE
74h5ZNbhGsG587CPaxjNqCVhmi2oNNVF/OcESyFldfttKMhjgQ0iWHSep1hglX7smlPUB4Fci5Hh
BI0jN8vOh2sooV56NTfkGW62NWNFf9JPwQ6QG+eym9cFjjWNeZqaKYeXtCh3SnLYnIHlXMM9EtcQ
E3WpYZkR92NJLCAUlEcgU+dq9jGhuJFKzsj2bCjY/4gDau4nOYFUDFwVmwQFR5YuotYkeXRC9ueQ
UfgXGK1qn0NnLZ0AyhRzVqu8DBBGFypviiYCvr3bRhvp3f+isLO7I+e8+B79iTi+Y5Jsv0e8ed0W
gUayr646u8GZC9j/DPxewTSHR76QZCHuNdABZoI3AcyvppHF6cM7Bs+hPh+FZPfG2PCeuVJgF7Do
0h9KahtdGA+JLPLKsa3tPW/MXcALPxRT4IIftPYcVYlgOT9CqEvrThq5D7qmID0tpd7HT/ZEq8G/
J/COQD0cjgY4zd0MS4wMO6Gr/t3dKfBhWhcUN5k5iH4SkBgZneznZBg8RgsDRTzzU0PTA9qZ9F19
nHK0TknvZ2xdlip2XvcE8jlj0PL8jmkZG1bCgkSfqWmliyNjdLVCzsq/0eIisES9Mb4FkDHEAfQ+
FZjjZx4pLjzT99OQHO4zA59a4ex1XlJ/m3DAoB7wjJHtc6sGIRRbHqIWzXHyNgFJrUTozuFE7uYj
caTDIq+rGx78vTK2a5cUulvb5qoruiew9lm0ef017KytG3Ub/P5idkBI8zZYtQRAWU/sbkdei5mp
6/n1v7ld7iPx46OrmjjlzovhxzNTIi3OLcGFOMb4N0uiWgpZADr5hjQX7hRP1y8oJ1gAp/3eLtNM
9M7J4bXFFo/38d7Z4NDGFVeN6Lczyxq0G9ebLJixiufrISUL+dm3lML24HrvXUOBK2xWDp1klhQt
eIiz4KD3ywtS8MN1SEiZo1B5outYsh0UW2yh13LXz19dKyeJ+79RnbOQltK1P2C5L6YbYhixY4Xx
gVrzwajoJXrpBHXzF9KLG82PPt3P/OYQxQ8E+kobDlXp4bcUkjtxhzCf979mh8L9LLL1G4lBsYDb
66ymLbSr6mCmotFGYYtOcSSPCtGqvI23iOCrUWJCIZ1QIzT58zbpqbAP5kJjgqGuiUSt+sErfTax
x2z7eIgjbRDC6t8kYiVsY16YHeCQ+APEYYpwcdBESWgI2cOeeaCyfdhikeX/Ybd8hZh/JBZeG4as
pfQkj7T4FDPmQI9Ho3R/A9ueoQ61f/0dpqkQvzMsb07aNFg4qIy5zacUWZ49YFUW0kg3cOFGWrXU
Oa8Gj3Xvy4IElpCU2KVmWRU5V+ple9KeWRIyllcdfsrzpmMkfJLPomzlxpoalCsOGFCvPj32ZrtH
mOOTQsYIsHavSz60tYEeslEhKHuQ5qWgiBCd4Voyu9D+IeQ1NMWMkIrAZ9LDS3J2lwzZWGYtTzcn
zTX4rb2P/+dTVaauQa/Z/zrVLZFRR9Tkp01dmjkpJUJCeKtshrVtStUiaVfZKVhcQjSsz42hSOLy
/+HIiFEaDYUqDOc91arWsJNLnB8ghlhXhscNevcajThGCX1CkzFTdHfvirHOSi6JKcZ/suhbA9Dt
GydUcKAspXDfRM+AmSh9nuB/vpaKVWh5MrFe6f+7F32GBzPUXPkYdGRe+KGHepqKVg5UYpuRjc8g
gNAcwlZbf7K6jdODDJFDJ4u7QjI21tyUYKVBqDb/uUjClC3QgCzDS+R9TwOh53sDTjbdiuSkDMMu
qA6AJy9EXNkiRZrr4oOhV17g4I4eHAagaikFCVwAqg40a7x52LDAkS+BhDfCHDuluRcMwnSzaoCI
EOGE4WgIiCdpyf1LkqrNUvW4EWFrOt04Ykd812XWq0dC/Vfahu7N8ZLw6zTb5YrmX4ST7z2WpMaW
XGxllEwQfSeovkXiuf4nTr7i1LAhRe2IFR8ozeF7dwtq2odPgHMDokw8+VbYe2fYzEe/CEXk8hM6
xJ2pL5JEHrlfjU6mgoLnu3tOoyl4NS9/+/PINpgdemwRr0thw8aBv6Xa5ZUp2y6VtJHkMmy8SJjc
EefI7LIExUHXvxs+7wAqZSE6+SLZNfOOngmEuqA16VvgQahzvARmIOvE1JEaNeRoMzXltp2yK0SG
YoIQk3qZRUD+run1W/NSMuF9HHne0cWVSbe4LItHt+AYG/MUWpA3qCnXUEeGZ1z1WsveoiyYIhGN
hX3m8sLyAOJyxkgOgfRhcNxl54xYc3dMSfiKQ4kxhNLPPyfN5Pp69Y8Bus5TaJ6MiAzMi1P2N5BY
JatpnaYkkTgZjIi9uz1vYYIwiuTcvaR1x6QSWB2cDxtnznPKf1+vDSuVhYT9ZMyU9M6ylFqwgPLC
WJ2Floq70Fg9f/E0QSoDlM4TG6Qji9zUgaC+J/ty7EhuSFH5ne8SaHrhgXsVNN6rSgtAhZpLz/ay
pH1l7mfJET/OlxAK7uXt41kPNOpBK9F4POmaVEy05eyyyvfVWzckG7l2FLjejzGYOcGVlg3CtOCN
fwSohFljPloepXz4cA/No2AoIOh6GtET0MCCF11etrZbhW1Z0v8Eb5yssBQ4JnZ6xrZ3KQCc4I2v
MKLJNSWVTGieIGEUTuVcoFBMVndZgJU1UOSfcbJw36brsGxs/gdXRpIULQ9WZ1Na3xZ8WzAs9If+
J/turEodKIsBYI/8oGFAbjdvgTI/zfcB7+OrR7MfLkK9LNzsxod8xHz1sq1cqO5AzK6TLsDO1jSQ
dXUUA8HS7kFB+Q53bjHis7NCDS30TsZsBfQ9+WghqkynGDmVHp/AvSQdIeNtiPCwpPwSiPOWvJ5S
bK9qTG0INtnH/aLUw++3m6ZAKFUuFwNbw7hePkjaNQYg7uQ3padxJwAQUsU/HDVdFJlg/R5SmgaX
isjP9CYIBuOgMN00o4etuOHo3+Um9Mdd3L2Wz8qso5qoCGA0zDbNDh6mrfGE8eSOh4J9ggxqiY5z
Z5or/GkgsKHZWNMAiEn/TiM6M+92Q/zqVMBe7IsrfyZGOhrnukKsoe1wmlHjcbBksnNYAmqseqrf
dTruAmKnJCwM66hwoHfd72uXQIuVjPa+ELq0oX3GMfPTI2eiEFXUXJs3rLqc5VUzbth7HyE2uQz0
kVNZfIVsrA8egaFjiWbIGOzLeDYH9i0Mk/aSHLgFp6Uo2S+CSPCALGjkqA/enzOqRRAwLZZqj3eq
Nd62MJ4A2NWXekC25SLIbifAptSEg8spwpYy7M7Z/eKQziLsElZ7aP3nJeNrnIH1Potfo9gpIBAW
p3A+HMMXI2Y0/DsJMAM/8PS6TjMTYaDBKaHnMtAvZHI6HTkqTB+RwUnEhzxbPqUh/rNxqRI9ZhfR
YyjKUt34MTq56W7x0mAmwnhyXn1ub2ODVwz2/Cx1Mn8MVGDe9IxSJkWrBcL292ii4lLuL0s7+ecf
531snRdFtJ82K/C4Lk7atykaw3Sud3Sr9wihi5TdQm1thgppWUiFI3AirESb21ilLx4Gh1HEq9S4
RTZn6eM5tBqy43cbeYA2FuqkMG0SwDis3pz2mjmIORrPk6Cf2us4Iyrr/D7ORYFeB6ewVfsyAlv1
0m3YbUj+O/FjhJTpJ4GsghpJTjridL0qQ4TStNLmgVNqTthyGTaaAB2pbm3kSAJYoMjlUQpuEIw7
2rBGTWfZaivPo8jWb34IrHYJwPT6LDu+6j+GpIbsqnXK46344I0p35Bcgpe6z4auiUlO4WuVuhOO
ADEofrrluXwh3l4drSCHGvXx3ocDftFXIJ5Y2UpZc6F4KIlipRsmI2clPo20d+n8axS7L0/Rz4Sw
WnAR+PtAFVkANWRFjC3RDFM3HQgdmE6U5xu7AFxEtKthxgWXlS4eV9X8w5IYqDaLgJHmw/5xR5Wi
vfAvnoog1CRChnvj/a/ejHjpw5PTB9a8qgyqLYXzxgdyY+JlYqQ4Pw5ITNJGmBYnt50vMorfLVuw
5SWftDlWF9l6D03wsU1+WqnUZqxq06Z8r4inW4yUbXivxiWHOGXtzkL9ngj9Kt082kYDfjK4wUHI
L3P3JaTvE56/H6GaI6fvZEWCuPmBDinirJ8RktP/pwqmuuzwiCvz9haFm1TEiPef359QxnDonFed
5dLdjeQKbTKmSjjnVapnmqV1K7oILYP5Sx4KvS05rOyKPmaBNkuL06qI1f0QI9GXswuUZ+bU+dCP
ukZnQUc/LC3B5pbNUuJ3T3CQxSbDxhYMM2rSWUabtC2/1lTg1vuowCJzYere5gpU3rBZUAkKjvRx
RKK40D9uDM7AAQBgZ6iD5X2hJ9KM7ntUFdLP82gAUJhjJ4azgRFVsQ2q/yonqKa/mQHBdK9kdICP
tAArlmNdUeAMZyAp3Q5hmi+dzRlgHZnNLqrBZ5wulW9OIdGQu+dYXJZg1CTiAgrLGxAG/TNk8NeZ
kwuXO82CkCx1ViXkFYB2hlrkUPcg9myfHNpsvJ7U6OAyE82AqpEi2eYd/7AlVJwfYW1VJanJVNxo
CUxTXCbxR/edR9DVVU42Wks3ZhwxzHJvUmH32yyqKXSGf79CJzMVPhJueDv+btl5yfX/XaII8TdI
AKDqLo8GcF9qbCV5P7KPBfPATTzAh7fU3qtAh7GGv0PKGKtN69VFNlViL8z3xv1+Kqhefi2jnFcI
WGcDldTS1hzQ7v697ncADJzHsGgqYR/7xfWlxEALkSzsS1a7ej1DAJpMNw1RtoR/uC5PMYw3C/wO
1pdmTaMANWrezfbl/syVOv9kgNmx6WNUmxue5PZ8/ncADAbZ5zom2/OFnSz8LrQeHygJq4BvxOaa
cIQCLjKn52RuP1WTE8TUN8d14IK8jz/TwrkLoxy1WaKe4yanE6WQOD7aOxDwi8DAoDDZnB6RSO0w
StOxG9kWxdeahAwGh+xi09fUkCjIRSQNkb0njIG6Ep5lBWtbpttANcxOihWJoj0AXptfFY/DyAD6
4/nlmWIThM9HybS7oFg1vxWbSoWTkivAC939HQoVm504b3x/kb/s/Ceq2TgdenuA9zK3fFTHw3Bi
Gj0EUS8PsktPLmpke3rdWJjJPPl9e5WtFmI/XCk4NnGSCcZhJ+4JPENg0IoSVYDVORDwU/Al5KBP
+tV/uJ2SM6wmibb+m40WLN0r5xy0z+TCIG3Mm3GEJh2fPv+s23C6AbPe/gAcytGlqzq3Jlmbtj18
d6FyBX7vLQThJYd5jgVn1pNXMpwhzka2ZFNz0Dm0zCAptZNPH7P/6JCQCEO/MlJFdjL6I8Uf9r9T
CTrebCtIQ9ppViixIXrO/iM599jA6Bx+I/eIHSJqcsm3FVsBCu1/akEE5qgPc1dyRMpPKhEMbj2t
S2kJQPEfWqqCdDCCCwtsQhM6EazyHcw8AZ1IFaSNZ5ySTf4Q3EfKite/sJ8+Tvgfm7T9LBFZ01va
bc8RtwCRDZNR5cS/X0fGACFz6dBGqCGa+SDRA7i8fYIOa9ldyn/ZAr9XcAmykkg+HgnPqaqIpo5B
mb/efWlXr/xGJ4OEdvxyY2qbVnZVs/IC0FCUFXA218qQa4NXpVPKFvZ7t10avs1TLpJsZKv49nVm
fPBfWT8M+/2y0bKFl+JXZdYL9pZgncKAcPR9/UU20HsCQNaxvsfoAVGXyUNNtYx+8898nwMemtnd
wUwjKL/a6FmflL2WOGiEaKhD1C5QCAwevNpEu4SMkWdtcNhuhPPVmTH5sAXw+qoUogBcdDhalEJH
5fWuy16NQWgHQQb4u3bZ7L/JpniIr+khTRvzmswGIMfze9pbsMq/Iv/WZa1XgLEfBAKyGh/Zf44A
56W7F0td/4Xo4Pw49q2ifk/ev4Xa+X/Pnp/li5VWpOdKwiy6c/9tUbCjRcU6pmlHeJCfgR3coyp/
Cj7FP6bmSCCOA3utUZbyZBWTzPwbQ3Ycd4+lL2w8uh7OxZCfa49a0YUnR9Pg9uyqvixfcF0W+XVL
/9c2XSmWhxTeZeQ+EatIcM0ssjXapgHN8DJjMOU5apm7opB5QXrZsYvLhlS9wnUBjIwbsrRhNh2x
vZIOe0vClglkIkh90pVKM8HMheLaQX31UIo0qAJO2+iEQ6KzdFjJ5rx/O3IqADTUjVZP1FIbnGUZ
u9MhrUGdidcFfqiWqvNId7g8LBvi432v81MjRx3GYLQzlaxnZe7xhM7Zi4TWIaMAEqyhwN8Gg5fs
uLNLe2IgdoWPUrX8pVOWsT5WwwyqGX2MuGT6BCXhBV9TsbDj4o3SU8L0FOUeN8/x9fqQS036+8X+
mYL2eADjn68MdLQTTN2D4ssWrEI6hLzKbP6QAMHmKYVfiVwKuXuNh0OdkaHtBk88M5RQgXXI2b1V
O+mxc4G4BnUENN0npHxEKTUNqFwWvGnISyERzaLqVoAz1moPc0NW71AUtRikSlwutwq+YBuvtMkk
ryxRW96vYj3jKdhkKYw98+eBUcUSV+V2M8pqqk8POwO/V4nuEfKDaIi+ADQmoBau60uTg8lcoGRo
lU4hdf/IVGSV7v8/re4ai2QSNopAZ3KZ1uyHzmjw4VvCHiYP7+7sB+8O6M50CR0x5/9x7Ext/HUo
9B8hXWH3hDP5Y6Srg+DnxjlDPV0yyaaD52PRyD2rofordNW8icZ+RSJ6lXZUgkcXvZ3e3ryRT3Sd
dgFHB8DoltDoxQ/eR+v8dE9qOt2sX+E4LxMgDnj3r7xgoPBQp63Z+DTLcpFf2gYgYsaFbhE8BPoh
5Ibr7LUdzs6SehAyQtLRagwJBZC24O8mS3dVqJe4uHQ9U1O9juZpwh0A3cgWcP76J3V2JigxDDdu
ocwCnbymhbUjj4OLLFXgzHuD10eAUZe8Ga9ttduH416ab67+sn5KZK5jZ4N9nyeLo3WFGlx+mrsH
ExSb3KR2cS8QhUof8Wto7XXg1eKFZhXx3oGApkpZhY9PyuEcRZ4BZUq/I8maeLm0IvcaNIkJG/Mi
gwi68ZHBmrMno0apCiBg1fLIXdHrsxpySumtQnF0hAUr3snQ0tvFo1K3GYxz1Qx6y2UbuepZ9nbR
vPX2QjR+moArN7SwZMV5YSPIW1QtAdSelHQ2Zvi4gdCVHB+w7UKCxjAhUf7W601xrctPOdiH5RC0
zM3Ad8CFlkUIWpTMXV/0+5LxCYJziVrfTVc+FOAmfh6ssaRINCoTGG1E/bXKRyCfk8NBA1o8fiOy
9MfbkhVpaHuIczUpHBl9++f85971LMCZRzg5TWHC9u9Zgod6W36s6EoIUnpCT6YL1rA5Ye4Ah7lj
jjzNLSHCoUbbLFAIWTDXCdOwUm2ZbnToHZRdQSqb+m5htCN8yDriqCP4e0UXQgBmiA/I9l8YHyTD
HN/Y1RCjDj0X1wz/hV4Ni3ARvQ9d2zSYe2CsTJVh8esHjs4AWwc1ihDxNCqZl810Vv2eyTTJ/f1p
PATOXPH3m7zxOIDfl958yfVJ1wDATQpFbKY1j4ckIQWkOz2C1AY95L854nh2PsSAtDjMsPfVBQ4B
pdwKk2IwXXuK5HcIpuO1LtnyH88OgJ6rLORTRAi9I3eT29RV+HklzEDf+1N1B4XuLFub4tSVYGiv
PoSDhN0jrQAP+OHcAEqg+02Y6eoM+XqKBRIX7LUvG6tNqb+6bghPMpP5CLGARZTBBzkJl72U89M/
u6li08gSXMWEFDSfnQtotWvqE07mWP3pik1rDJG/8IOJpoPLtRQpTXhJCdBVGFnS4YrmkSXln/Zl
TSd8kixemjL2RfmWdF7hE1GVBMWu8eEJGDtxZGJqfBtcoWijm6RAOeH08basliNB5DACW4w7Zbst
+cs916U2ndM6IyAdX3jr0fT0FASkmaDA+S85eeilMFmSFWMng5O7n9R5CMN6FkE3cKbWTOe4khro
L+B2UagltQv8AGkdQ4LCChXwoyUVC1hRVil3yK8nWj16+TTDrhjinPw50Z3o5AcWlewOARjVyqs5
tuqnaOLNLpAQbwdogy9NrvMVO7pll8t+/v0RR8bIPlaH4E1zKS+mrKZBLqEhYBAfC2QXXqj4Z1fp
K7cjGA2hs+RgS8RtpLbymeyG4MjlKO3glYqup3Y2u2qBZalQDAYG6KsBMnRPIkSduGf29wVbe4+8
BoILlR9R2ufWkO0vrfhW1JX2pZkqqa580OjnG3+AmlwiL274cOLj8BmgXkJtgHDKDpqMZuCf7p3q
24F5b17lxQAnSf13iBz5btwqDDo13HKqbGklgPnGAyMjPeWGHOFGUu2vRM100KgdtzRPlRTBqZVn
t4VKdimbWzIjQWL552H1XYdou6TN9i5L17NzhSgW7m3gVqjkxcft6L2Cj9BtcEwBYH3GxWXCyzta
UOVLN2IdcfyaINvdygMDCZEdjC+NlZ4HwF9s4uNn5HzFyqH9f3tfjh2l/98XjwITjy2VfsKEfMM1
FzHXmq0PxqVJzomfwKQ5H4tBFwNfwpHCRoKz0O5+2nQc9ogu1DhipNHDJwD2f/6oQ5J0Ai7pYbBu
RAMj1+Pm4h90YLyBOLHbZeGnc7J8nOQAJ3juKiKJy2OzbpE+4ULvaJBWVvBhCsrPxD5eeDjrAFsh
yxFRBZVPC/j9tsrHfUSwVbqFsaPN3Ag3rzbz8j6E1nOD5yleT5dzSbyePLE+La8qXZO/WIJuR7g4
3Dl2VoVocfhj8r/0pq8ql3rCdYmDSNLf/uC8udAGhIemdTHr0aIDkZHTX9i4zQBEyV0bXy55o4QH
VYoI5iIaFnkaQ+v1QBWFh2hPr/kUYKvG1+i0AVGt0K5knw08gmMA11HShKl0FfWct5lNMMV+cAGG
BgtWY5Tgi5598X7NfErhp+uglRnXcowkdw+uyOvOz6ufbp7JqT7XHSBY5w5bRnMK0HOKt21xwMac
tLJEUJqknM8aq7K9J9ifrRaYNwlzCh+rUY3BD0moa+2q4xylR6OBMIJ1bwsM2srsz8uW1tuzy/Lb
aCTs0iPp351I9HGpccUDQxDQahm/oPXzZlQNinFsmYAhS0R4tOd5xPFONPFA/iaGruCprf/mEBR+
mxLUndGkeGE9fARWmXNiv83K3DNdaGMifEICgN2+v0iJTsvBZ6c9vMo+Q0qddaO+GqZJrmaSUQZP
40BJBEJxVoL8e42aZR8oAmyTlp0IysMAKoX41lDV0frJcBa71yezQg==
`protect end_protected
