-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HGkHn3mSMtKb3pyLwkFKZYGPhAb7M1cD4rMN6zwsIrEsrgi9ZUmG3F4tTuEwtjXxPh4nRYovUar4
676X6BoUlUNmnoz2f/rp8g/CSsQVYax+teqI5/uHtwlLydl45Id9Ktznp++jc+W7mMWbqZ/wkCdN
1TpkABp9nMC/Dsyf4/kiQ5rnEL1RmqjxpJFjhiNxtGS+Nc93nopfEILdW9ANGKKgTQUGXfcn/E8n
1SdmRg/ZdxYfOA0U7vJSha+Eze+td5BRYhS9Vb/d2cr34mlgM1Jr/zvHWDDP98TgY5AtHJ6/2lGc
z1kduTqAMkX6ybML7RQxWDch0H6tib5KH9oAVQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
XmA6Lnd2UK6Jrnp3qJ4mbPMkQEPwecEQAzsjF0pwkBRB6HjexyWGok8Wv4Gl1fV51355zKtJsHY/
XM8Dam5dLdTA5tJnwB0V/M++ekILvCjJh5hlJWvp/oniwaEXu6sOLXiJCxqErMU61dDFrYrBB8ww
xGOV+vW3XUz5X1N9AtaTvDSwcpO9LfaGw9dP3kIONDNJyvhS8BTxkhswKOT6HGmoWDNKVucsmG20
b8P0vV2rrE5Pi4cWW8IhkgRKN+XtV8u0v59WeRfzRPJW7wT3J5cbO2zJwqBBtNDKAmmjg6hNiPg1
kzQMv/WLGwiCT43FBIodNhS+mM7ptrqL780fmB5o9RTSR/UPWzDSwJeUDgfvI1zGX8HzcAI2PmPH
ipvgyBnELGHIj+jpeb7jq1N17IvqI5gLM/7BK7O8N6sxPTSl0Ko4TR9swsp2QJFmALbRcZwhd9Cq
OHc31Nc5zJt79287Mi153EUlylohLi1SfXTPZksHaCSyW8NHVij2teVhV9plpB7XvTVKa+/TfvkC
QKvTWvHZ9zgkoDD7xIHM8aCm/5IVrbpyEdlIVdnenyFZ4voRLGyMf+svI4inUjtr4NDCgO/jWs5t
yw9Np2/SsQQmBL+kBkNnrHMBwSRr1iLg4caOB+6nQq+OpBaPkj0KUkxH55d5os0aHr9w+qZJwqhR
F3HvuS909sIZlxTpevMaF8AlZxWSw1enfbpCVtsGdLjEa1hLuFCMKT8VAb8Xwb4OffdDtIIBHkce
CumFij/zP7T8pbnfgxR+crPP3Rnvj2X3aOBaMNK1IrcZhCJ02K62CNeKLblmtQPFSdSWc+HGR6Zp
MXXDaV7Xa2fVPpt0yrTzC4KjP9Xr3AqtaNTHobObh/j1D47vXJArnX9L7MFeYA+sdaKSFfhxBm2j
AH7p7NDxDK3yoyJcw1YPSgW26CuqaKD7/EmfsYRbwSaMh/ay6v8JPqPAqlQb/0ZvGg6K+ZE9CJui
UfYC0YTnx8oz5RaVu+5UqQ0JlWDfESZfPutEAWdgfEcyUn4yir8Pm9xrh315tH/NZj5fFBnzt6Fj
4mFe+7JuBEABeDqEPT8tEGtg4t4jUDLuz4xEUie1766PtGhrgtHNHFa4K4RYt4cqMcutz4VVyksM
VBcqjAYQUwZgR5w8araKVmxtZISPreFdvgtq99VmfrEp4IK6V8Q7vm+36Wa5If3uOe2cg8ihgfuO
aoqPix00CtZmfHlqu1I9Sd9KVEpFHxpQfiQN4BqbAckXJ7qKQR/ea+C8cuuZW96c4C0s0bk0+UWw
dBJOFtl+NJYIWu11GuIU54hRf6U8nlmVEPvrzaUnCSV6M+ILEnIUx1MO/oQ5D3NBG1qZ5eNVWJhy
cr11VlX4lYvGQSxjmF8YHT7Frz8L0DEJ1u8ClCYj3/5zFC4o3w1n93lacr1YpuiZBgoBPeX98gyc
8+ZIx+CPl3YOJfuStxTPptd+HO83xiKbY7QPo+E1NZEHypfGBWF/iImQ/1BiUvAFDpvANlP3SKz5
9bgPXK5ROoBBxmyHU0iw6X531cNdTxaJ/AG2FRxFQJHZSm5wcTg9OywIwSSKhxw99qqN3RyPXU1E
B0/GxQqkf3jAHbWV0lN31PNqRMFFZnQVNH3e0sHCD/ehcHUiT+CYp8luNLzMmxwbh+zqWd9fxGgf
JHwDrpMReafGjdgWhqMCeD7jMnm/dozspPESd1gTc1cVHFPU6ZeV1kzITkZ5W+5P5nFuODz0T89p
aYv8D8t9cregSazhQwyJxKEyOjLhH+cxNJ0h2vlOhuZscqI9h+RDQF5rJty04J3nrPtsUISxvFhk
oMuoRBtmUjcJ/cDgG0eAH/FUSy/qDx7b9vmgCiT2q+D3l9mZ0NmVus2HBN8YIXbi3mQCUBNQTAaD
zZJ+eBjrqMPDh3mudx8hHzt2Eh7B31uX9dLXi+xILtRz0ACu0YbuyEU46fQiFp07iFn3uCh9LkJY
JaMvURQq+QmRim9oqSr6YvKrl82ZGmwSD5uBeNQQvfOlRuQzHsnQGDjsgCr3LkOmhwo3pwZT9Z2/
qXkxoo2BGacwTNiWW1VyVVuummQF6tGTtBJU/7xt3qDYK+qDSb/fTY7SZCtEsRAKGnFzfQwHg2FY
5FVCIS5Xi9rtljV/rPkPsTL/6Syfdez8RunJo6QkXrVspjGZhkvX48H8QkrOYL4ZIfBjLF/8RIBm
eWxEVkmlS08bPFZjZBFgetDiSV6mIxtXy0PY/H0C+XN/BlnSaWMhYDopQ7kWovgpLZXTonmOlm88
9e7KSglrHGodpShk3drk/yuAW8Zb/WYrOdUvWNOA4R3a1CP32ZR+DM8eLpLK2wFpnspiHzWEO+of
JtUUY0JviXY0OPqjcuAB2Su5JmNM5cEZiANWuLMYPEWf2B+ovrvuRx2ujGDK/ycqN8jIP0fKFpkP
Th85YjZOUJmBMJWAfwYh/03EK3fXVRmmKd/OEgVoVdHt61I7dlSzEklv1MFyLdYPqsLMXkSFxbfV
HgHg4g7y4+7TqXL126P47a9imUCw5+TgHoMI6KhCCbye+KLj/2FARxrTCgLNbW60TWtHmpESM10z
iAgkeXporeSPQE9UOK3Mz7samA3yjm75SrJoxkZVkp51qlH4EDyLhWEx2IjFF1xs3nrialQxthJQ
WF1OX1XCmdfDDGzAo2WVWPeMyg8U5ZUsKzAV3cXWUCwZr36jnNLq+ndkpXFXp3TMEFMX5LG13HVQ
rB7TKR4knkUSLl32K4ATgxt6nzkeEPq8gU/8lw69NUYfvcmj9EuWWzvrb0R+hxAaELgAVNg4O+Q4
e7MPhaxgf8FxzDVn40EFH7fJIpS79xLYuHPhXDI6gUYAaXbR2q23W4LzHpzRjCtcCBcplZBU+pBD
TFqDxptUVHBw4iH6uPLg4r280ewZsmILI0Up2h1mOZX5Wd9aKcigLNe2MkRIjUFF3C44DMwx9T/S
dXJXhm9OR2tAGFFSKppbIXc6z26lWILIeYANfJZ9BFGe7MQIpQYGNaVWbLlTEWiNu/g4ree0kHsj
tjD3KSk5kuB3JkpUoogzcO6TenAycLcSfHk+H3VottHha/+NnTELHGi8mS92O8Ok/95EBDkGlnhV
7RTase4kjmARv5X446NL26x/uLjaI/Y3I47Cqq85sNslZoji6hINfkgoSlYDCLdn2v5eDQEcbbmK
hJWfhHT11gBFNt/S3p3r/SVlGWR9tTp+58wL9Xsm7+AIQP04RduEnLqx5lzAhqfq1wTT9eM4in9E
ZPjTvfZow8YwzOcjDZCWEOlH32d/8jBJ7cfP2cgG0MlCvpLNwGvH9nD4JaKx4bXYZTmaHS4tBmH2
ryBg2sb22ex4qk6L5uCOWmKs1YykEM6IT6FWGJxKi4ViER8c4TDjM6rjN5c6j0L66xhl+EJLZIla
TSJSif8rwP6GMj2cSGD2Gsej1Hb0JLSJC7JUNMjhp1J8s8O3tj7ZWzz4WlByq3agQYnTegjocL2H
daovlDfyYgz6s7wVBxiPt8UBfWQaznOw5OsW74l9R1rhxr56dqb5C4RD4aJ70ELktErzt0joYtFQ
t2I/zbcAjxQWEnR7I2T7DQVn2estwnbCl4MKkNJQIKO3ba0Mq23hXl7YrU/fMkOVHJlbxxTAbO/Q
suJk4I7WYaYtXi1mR5FdASxi/QVtNe/OXDaZrdN2rzxYpSSdMLGaFYAaORHttDnIduqdDxehEUs3
M3ewUeAWKbYiuIZkSuiwCm1fV4z3PBv+Q/tmlw9j7DGC+17ewmCJUDKid5axZCRKrF7TkpW3bMW/
8VGW7GVLUXRoq3xHge4LD7keRyqG/lxGPwuKNAESIjMPWxmGb9bxG7NMipsZgwbGcDZJDR6rjEnG
ZI3q73tVV7I8SrEHCk4Z4jR8pHRzxstFamcVSh6mLuXFHec1ABnoL5fwFlRNcxgims+znlgn3iOV
2dbDsQgZDS/hTLNvDwanrEjWutAlgU2WHwNgYK5QqG24831VUjppUGsVoPhqsAnDbNeku5TTFjbW
8cO2g8w0x/oDI56eSKLEpmvmNIiQyZ8GSBYINI/6CCUeqFeMx9aMmV8GRk+x1e6n8xdyj5EIoYkQ
SoPcZN+2roKR1Alv8VDllfOZDricMbZugjOku5d7EXZCQ8SoQmyHj5aYarWGJrWTeV/CDA4OxL+s
cx9G1eHxvl742Nrn+GAX7qGltb8qNoH6nb7fKSlP7R2TEVyHxW0tjVRk/CMQ4JqSkRviwjdaQ8fH
lnH9VLQjT1Ta2aU/okGmSIJGOBhIQVt0q7ht8IRwO6fGW6Ucm9Zzt4XCePFR3wPOiGj9gR481yUB
EuG+ZZrE3q2j6w2JsaBbY8LTkrQP/J2dsmYJQnxaQLSLq7v04ZOHqCcBVfFF0ukvgQMcvqt8B8zk
uUmWWNsKcRGN/aDsvxXzQqRzTV1JfHlsLyL5fBLeyY0ygJNgPU122kCzTABvaeMmHa1GcZdAq2+y
Ox6rIZXA/F2a4VgjPbhXIUR8ZoVQeI0AMiOtxLE4E45XbTSy9jkpMV88UgfUj6gY2/MkmOOQe8dD
RlSfc2kv13pDYzBpPNuIIS1SSGBrILhZ/7IaA38nDKzyQrsufW+KPl+doW0w1Kejaq7mbwcd/Cy8
7JkGVRQpzQSj7+KM/8r6sedlSY9j0+8Cz86l07+RRRYlkxcD7wXyq3U7ebUGL/vuC0b9sLXwv3/0
3RMtPNAvC4m/2kKUlczT8XSZSnEiEgA0CsSYDW2xo1o4SG1BXBP7CsR9W6yG3Qnszr34GpcCtEeC
ShKPk6GyeQ41SAHyffFWm/hAW5x3OOmC4cU1iCZIgmt/asNQ0fzagKHYEA1iL/+VKfSdPu2/7fCP
Y4XbZhSN+OfLUmIS1Qni1pPFosCcO2sWTSH44x5MkujZ3HUJROMVbXtU/lf4C5GAL0SCYl6Pq1AS
3Nk1A08dM8oZ5Mt3L8gJNx3OQiww735rk9uiHqBtvIL7jxty+xQMz5WyBfvJyKI/JDKD54UilFXv
JpAubV/vl+NTzzAilzHyfrV32qiMOfDIuy0UEeDBIrpfWfOFoVPRr8YanKgEdG9nRJX+EEReow0S
Ofjte8nmA4wP2TlIj6IIisVt6cBUIJSgotXJ/xEfgnHg/qxmKhwhIn9lJr8m5HT2C6gO4pSJ/5JM
fG1WBQBZ3CfAx9dtcGlP57VApgVee6rvGVUaar5YNNaA8YtxPxArLOzTcH8FeMgeq4lMIsQNYH6y
hkA+azpFjRVIBCFyNrBkUC7rujq99O72hr30xaWqxyp6Wl+3fe3LYDv0PPhefXYDVwc646Pxmo3+
req56tAxw1RbkRA8pS7DmR3n0tpXls4NCwYn7nxuFUcKEZUIm5jSGf5asRmE0EUjw3V5k6cCbsSu
6fPd9aR8AHtScK+MBsff4GuIgblM6jquQLKJV1zVUgJOfxt/fIrVqOPG4aRSGv/Nm8WU8wVHFyoD
Z3THQywl//DW77ltrYx5db1ungZAkVC4cn9vM3P6dGrMLEIC8tYkUJ985xI+P6b6xP9Ft7a0Kz3C
EsV5+kuFdIRqBhLefQapS+WN/LopDTCYndO3bx3DrXGn8ehwWy2Ota0M0smg6W911tT0pk5Yh7aS
8eo7R5rnNaasS0nR5azJbB5J8orsbonzMoWnnV0MP4WxyRSGQwuZj5CKZQhcgyPz+sDwbaa8XPs4
ahn0KnKlbv6XwBJ16n2UN8jOO9f2d6uJciuroijkUYvLMMTtMNGNRt08u5SsOsieRpiOtf6P3z/h
aURcJJ/tmZ4Jmq+axjBPINKMDKYh4k5HPg/kCd+a2B1cozK+o5SQGC47JNTqKZ4O2bhqilZ+bnBQ
j4ceHoIlCjtr32VI/kmIU/pnC5S7MbS25M8LOahusXMO46w/2OkPAD21arPfMLAwnvDXcAW05q6S
aIGtQRUEvK+AcSZXSvQasv4XuRxAy96WDYotCBjdPYKHc4pkgj6K0QumjyNKmGA0GGE764kCPO4d
YFB5D2tNUjKssmyH7nlOX+1XLvxvha0dE5j/4oO3k6UY3yzbBwIAG9nO4uyEmWmV5FcQ9nq01LXP
y3A25numgNoMEhl7ZuyKfibZQ4J7isz5eiQfMcqZgePmnfdcItW/eb9gffLIyW6ik/87H/RHWAmT
LllScqhCabHHbnhXMA7cXK8SuNL11AfmlIFUwbpxRT9Kgr6D+ghsckpkoMBsX5GdHb5tDcTskWG3
TCFGmnWHmX4Nyc1SK7IKAITMG3ovS1+1rKNla3oEN7WuFqAmdpNGId7he/rK5slEEk6mvcEyU907
JFff1qdVWscUu6kP+5tFBnPRZLBiR2JNK2a4Xym/6Y/6SWduLzx7u2clKHDbMoQ4O82Su6XGk+KV
PMKPGCME78Sr2nPVInRKPWpaIeaWBDqUP4xPUKSdoyZZZm0Ua/yAGHjzdBMG14w4QQnlYQfd3Qk0
mJECYRNqnFDKT8kDvFLI83tR9vNRNHpjboLbrKNVmeVtb1OHaaKc06Cpj5ov5GyFzBxb6dH3nP5y
zGVO2sNeE18fm3y0rSlv2/AeBWNsemKJQq6xcebx3cHPpgye9rXm87JuqTR/vEdFTbG4OdQP1wvy
u9ZGIcL97GCr4KagoJM89KgFRgQGNRDpyrFiu/gLsD3H9AhtB3MZpdJ0J7IP9k3T5Sr3C3WxdaKi
EK+P/PFIckVttvvUaIw36QZpANoG+fwfwdHhaJSUGj+fW5Nr9Xqf0tXUmX1cv3r9juIYBuXiPskF
tZSFswof+eeGhLgJ7Y7Q6HYxcAzZ41U4RJU8pvgvR4INGmA2SJrGMev14dlQgC8wReywLI66nNE1
wvrkT4F9p7a6VGk+E0J+1x4SmKqwgQX59E+dA1ISugfuGfIHKSXYfTCZVJSleGO4qyeIUiUe3WRJ
CkQTQ6U28LIAEfkH+zAV1uxpRLJ78+/bw6RgwTIaFvbKRZH3AXtogRJie/106PxVaUx1XpJv4P90
AvH3np9PDHDW2+q0e8zlJu0l/NCwEBUJv0r10cU69aRlaWIBdhvr6grPFfh3k3y1OkGTvCHePNyD
QO44eb7FElTsno6FcWUcs09UYlKsDYyfh4q+jdgEzbC48D/26BuFVrwoIyhiJ1HpMEFMrXEDMk0D
SXmjRe7FFXluCRtIyzN5d5mU4kCBTODmtuEts5yEntVkDqM8JgrCw2/u0Rw5/ctSt8FohKbp7yEu
xxc2OsPuGB3itWn7sySjnnd3e4n9NHV8u3k24u092kUBVqC8/WFlipyoZQ3inqSLcjk3jQiYe6oE
ZFusEEG0rYX72TSRmqQWJ8HOFVbjDXrkUjaZM4hbCJ34bz8Sn5U+is2KOXDQxl/4DwQTJzPpS/wK
Ze0KF9ijlbK1CSnCPaiMnaKgjU9mUZUFEZEjk5MKMqZHZ33DxDznSr/Kl7aVqt0jWFHzKxwS614H
10k8jZkHqERUDJyXPTmlBoHUIvJahHDOtLzC1qZxNz6SoOrDisCv/vesj4CJSHHMEepUVItTqdTM
tpXxtOeaUjyBJeHUYpV3STz+vQi/M33t0A4EqTznEA4xETXvf0NgYDqFJaY7t6wQvL/4tkY3WPx2
rGQmW3duCBGzEBezWb78t1cXC7Uz4krPGnMs/AFXG7Q1kycdOhcNoyeE7/ITajtCL/TaVBsXaewt
iBLVIBAUM1Iuu7ApviHdu9+fktvdHFRR6td3z/M0TFXcc9xX2my0Py6ZUdd5xX8sJmCmUHFI2eax
GruJr3LuXySwvVsnmt56Cddkd9jBQUCudlXTxXKWGgMwLbk2zb2qhopiOKLbEZ3o+3CjgFYFNGnI
pL8FnYAMJIiTtJsG26SLG5SHRiX9ptozHb1JhODhIFikOMVuJdKPwlNjoUVwM8SfQ5ovedo5v/Ie
da9dU/2UQ3f9g24p55YnTL93GR+7Z5wYLsHrodc1tGyjAeWx1n33OwqtcCw+EA12Eqobw3bnzWRz
1Calyv7Brh7cJql2OTJPgzz81M6GxWKqT+miw8cAuQ6gYEV6Q++N8FuTEXx+U6g+HvOT8NUWW3TD
2AR0eW0MuluSSCApCHzAAqdKZkBMWneIdiuw511u/dXr1jYKM/+OtGFG5kwpfwBiU+sG6k5D9bFy
y+0py7EAxOYQI5jARZYejjOy0AJdxeLzy1aq4eZcA1yGh6/30Y29Qs8de9Hu3PXlU9qtgz/BAmqS
7Yxr9KSjNt5yD+M2PtkYu287FYjs9F1EYZd99u/n928m+nmzYqOjQnvsr0i8dW+gx0xl2JCcRy3Z
3l1sjsTPcwY7Fs2ZYlDlkqIT6nUn0D2rlYyKiv+v6F8qZRsLF7jaZ3ITIJQbt9FV5jsiYC8/c4pd
PW0+uC+6pX0Wuz9X2d/V6Us4NmVSvY87QlzELLfgtnCBXVphE9PeFHQf2TZH1STtU2Ns4bxJZwSV
KDhrsum+eIVlUvjjhzHbKXIMgVncHjk/4g/jvZrMQmEQmSaZ1NiuxtUBPhcDhX6vllFZ2nrm2p1b
1TKtYnri/g/33LrCYn2S8pzDZCIJ3drNyAYl9pY0MdWzn4IE3lJA+8VtI7bj6UkPSiYh5VIG7/qU
b/LCc065D7sxTBHy6WA4qagZdRwBkYnpbdSY9F+UeuQBkZCNO0kbaGAIhFrmEt//3s+aPBF80O6O
SmByGWVb88Df97PKn57KjEg8gAXaZMRIxt42Fy1bKECJvQ4Jgp8WIxvlm+87FmuWWh8ASqzydb0Q
bnOrpbvVrgFLMZ+A2i8ABHmhQTOFJcKBOenV4PuBfo0IC6B4jviNh5YKhk2lfdKo7eKPJ5W14Ukl
m3FgNULfFIie6I16hobGBWv1O++aF2CCrCdJ/Y2bmbPkSaHauGPHMVmsYCixcnTLs/JYEahIsdBp
pFnYfV98umuQx7f+ItlvsN93s/krwPC8PhxQBX1UWp1oWIJ9irSvgicyNTxRvLAkyQP1XLbiUPhm
b/iXXrv13ZrnxtXVlHMG7sU6HURUwbuYfwS3T84TWRp5oRkPdX8EfTn0Fxbvp7zjS7s3sKZLDAfc
5vLXKAtYdmv4XGP9ijx7geLkUujnDpS0a7VPXTTAmvANOPK6toEM5fGny2G4Idx9B5jRkCMQbqfz
al7V6NtIbVyt5slyVXWS/A/6lj86cXRNfOEl66XhuoEK/KGJoXfK4IOET1OSgUjMAVx9T117TFDZ
3A/XN+tkvtVLzLZEdrc7/WDmN2gGt5c6D9c6lusaWBlViropvIR4oRQvE1kvOGNPezzc/NMUi0FF
D/Hny6/ikY/Mcni3LaOQ0t8PBJWa5rgJLfCIInrkzzkIVQQIx/LY7rcabFPjGljjD8RV6uZwfORF
O+XGn74fH/IHL0ZXErjS9vBWfDrvl+/q0E+0MRXm08fJAM1qYU4/Ifl0rcSCoqf/aDQFwwQDSlJU
SA7WJjCYFtzWHhOjQyyt0KQD7M+CmnOY8G1m4Jnpee7h78LZu9esf++pXNNUEYvv036+H48GEaNh
JelpEwx21RbizIgmjbWVHhcdHs/yd8yNJQ64kG5INkZwMJA8WOOXwc8sFyv5K+cgLoGt0SaCB2Zj
R9euBnfIzVGw8zh5rjEhfsKVUpmzTu9yMOxIvCF1s6RLf9vPgdaUigQJJZvda9ELwi9MLLOKuOHS
biqfxgmOP4JP3NoO4pN4v9qNmhI2zmsq33aJqlaOD7ElPA+wbMiMOXvG4I2uNbXhoJYq6KZyGWYJ
UxCzpp5N/lKYRXd2Xdtotfz6KnZr3ajwZMWAUV0ip+fUoSWx1i8JPdBO5PuVTR4UDeCUzdjV/bFz
d7WD1rWvrRs1VIcl0Zt/bi5pUp9aOkStK0vdwkB9E8zrSmE/v92QXQWvEuA1/CesbXr/ZMQy6xkq
FCTq12o1vWlOsYgzeqUeJlanXKyciL2tfVejFTPEvMXOXXoxdDoRYmPIHl32FNIuGW7BrcfCftzT
f5Y7nKAWzxTC+zkz9G05mWp9uHIKFdNDuVET8oRqA2Ha6tdH70g9Otlz9viRW8viiLfbvGLoU126
yGZqwMy0oeAqoedUYPSntQOGpwYt/Z722Y5OmkwPz3HmSBmIGTHIBu383M2hofv7pMaglZFextMQ
yJa88medXBZz4Z58rhmg+ggzdQDfQ1zZz2wyPkWLV58UalG4lpcDIY85KhRt5Ltya8MwPI5tL27G
S5Osx/zlxe3stJAVivjrcqZOXNCEYKZSCR/b6y4lmS3Tk7UEchztrRLs+HD6zQUaoz+dBOIcAJdl
mk1bA2IQV0vix8BAkRdGxdkemK9gez/h+PaTFUdB2OWrWK5cowzEFmxM6SXOyxTbYUJ1BJISp3dl
9OTwD26vXquhiP7GlnMwAYPdE0rnp7F11JlN0mIRD5+TY5HWKmq/KG6fGwI5cHLWP+6S0IewsQ5K
TtZiCGIjVTQtSEC/RazJgyKqLlIandp8yyqv+byIko4dOFvI8tHgZuNw/KUC0zWXI8lrsTjweOAD
BlfImSsJN+7xXyUraMWsahi8Xwd67WfbnTL5SasDPfqoRUlmgI9nROWnzHc6MFWvBCU7r2GT9h0k
/o7lzBxfv4GyDvnGIgR0Ni9KoAl+5tjsquhl4a+RzISEmHaM5bxxdGPYL+lRbimQDN2ViPkl94kd
4P5mjBzDQVlJNgwAGp+2/ItmC5mziLexvN6lZEjMvRv/LM64DLfEYLDm0DGaY8Mbs5qZ228DLPyz
dZT+7H9wo8VsD9tQzuZN0lXwN/vTtMmxUIRI8xKtgt4QgXZH/aR2/uFdOG+CqrVQQ+VWS94RvOkP
uZUP9V+9BJvzItxxYrNcQTuDF6BeXN8ZZJG2cpiwwczD4LQWluYVcSnnSpXreibGCTRtBB92NwTw
42VCZBiiblcpeJ1SXLEsGbW9cWaRKtENxu36dJvwTGjNwBQUUWTYJ6h6FyYx40x73zHjgYSwUk6C
Fh37nl7C/Ql31ATijimEojJm3K457oFCQ2HkM1mUenKsMjF0xH/GLkkQ+C1fYg7GQCGc52r5Xfr8
0PANjdAgxm6UTl5h2/U6/d33+BqoxFmK2LzyD3egd/sQ81TMlFFiaFebuvICX0enQDehOgaYpz0n
QO1kAqBaJlnBf2CoB+adwBW1mQtf6Zi+XrKrTG9520PA8FhsTtemyNCwhUqBZpgn6vu7yr8PevoX
h/tKowOtmu76BZPb7WZJdg7TmdMtWPnR7sj1S8EjduRJ/PSUHvWm877pT7L+XVZ7WAcs9nZk6As6
9dFRE/vWYOwETvJ1ktG9jFhWCN1zN28QP/dnTJu2sntU239rBX5YDCA9w4GZqF0xcBZhyiq64XK8
qH325c+Fr8RmGB5c1tGpsgwmKdkyjGF4+LMCd+pZ+fKTR4+YvleyO+IyOYGqdc7L5fxMlQ0OKeGG
i9N/DoLFGk+Vp97PhO5Jvwjk1rS7u3sFaES2EHRSiH4PhNCjSDSoBYsr2Cx9I2EgoAnAuH0ZhTxd
BWicFwh3je8tdEH/LwGgSjsbGz9DBOXyX3eOwej/kJjUPGfIm8cdP1/0NbXZaGsUpxJUMdSYGFFj
ELyzZ2AHRvXqEj/V7psD1HrBGf0q/tuKw/kAv+ey7/brtmmvw1BNiQfBCsjKI8+vX/o9tC1tR4Fk
OMiR0IjdQMH2TRIuxCfq7hcY5e7McJFXhgi6XZVOY/v4lDV+WLK5YmhPulTvaAgDUooegZXliZGK
wWb35Unp/EBQPCP027oUlpFYnynCe+8HaHORROaBlqhdEGtX2FwJWo9/ZobXxdAFsIhiqhUWUWI/
j2EYbzKwZUnPd2LbRV9BS1ABZrMegBPVj38bijM6LpsbNjE+qiWcCAlaP32BRLESeYmP7HVcjI1Z
hh+Ewh9kODfkn5HU6o0HZV6AKUfYbUUVntZt7xhbbrLcwpNHAyDCbiW1biAh5z5H4p7ZsLYdAFS4
oPOfgPBxLSy253TYRvNVYUpLZl+V/8PHVxebdEhPqSsM9GYVM4G89LQVUu4eN5ozi9ppzjrFKP21
r/2m8TzzW1Xc2Tq7Mme/QsIH5QNlnH0jq601m2tVHLa6LIukB2e3jcKKnaXoakZrcGZ43aWeDfkr
6pDz6w6rAsBIyCwGbhI00KctbRbqOujHFrI9RNX7u+Aqf0kMxHnt3V6yMdTPHork1kllwJSY1QKL
NaaBOdJmx9/KhzExwcLjIZxDgNcmXF+jOKKvQl8nByf8HYSvEhwxmWuH7e2GWj+1vry8jyiRhtF2
ba1lwkmd/5ZqCKAfPfQymBVcHzYDqEpDAKesObh9yX76or5aKF9BfgMtugiGUvYnC0ToX8yYk5KX
M/K+5GuklpsYGVLpAVuhy5smabq83tAvgYqGjgfgoMUW2i+2Hdxgqe9KummgP1VAqYEqDQa6vpd6
yxKWTDEAAhvpY+bVdMUA9aHuvAu7fUlSeH5FSUzabJ683scrh/uOeo5AHUWAik4eF8M6gOPm4WbZ
c5MgVvl07HYjF69rf5YxJw7cceXy+HVSBOkXJC7ATL0WEpPaXkEBzgQpgefGm22EbIM/JUSy3fpU
FxeekYgBLHW17K+X/H01yBuT2wfMTlvzYETCnrMaheEDMqSvJogwtyMltL8NcCQ9s3w+n9IK/10f
VJCVpIM0K0c+Nz3a+mH554Vx442W2b85puEWp576wlIT5T3XgrKevfv6QYBD2wIR0n4ThZKSgcCV
M3rMXYiYUBGCMd6MuSoO9sGT64ilIzmGzXgevXkioeVdeX5O4NmRhnYkrQJmPYhT0y9VPX4VsgMZ
8wgnQzkzwQ62CvvQlWr3OyEuVGQ/K2H6ljGOEYAF73iYlIYtPISfRGkVR/E4tdhG09gIvicre+mH
MBTkurhIiKSP/qsifEZrD4uNloEWNWUECA70E7uPsQVZZyFkETOBd67xxIVbhsfNDAxTzM9PcJfj
yOW2NnQ3gOMU4PuY6CB7QUxmAYXD+9JbAYCDbGnbuDbkzY79oEKrdmIk4DBrtkdiOyIAoS4tSFoj
At4OcAQFbwGH8qGkNo5eGLTAoCBzaD/1mhN+MXjSwEGUMyjjYQiDACoTnH9wslwtfPJvCVGgyA6o
/AMnaDMlZlwg/eDTEhaTFJaYWuqCz0AZfbdbAsMWDueDkcGGUtoLcVA82BMe07cy1gW6nViPHvjJ
5xPSs3FPh8XYFCYcMvp/XlgoLAXw6oovdBdEXXzCDRFHaUJUCs/jFcdu/A0izQbdvkf09KwvAXiE
XMytwuV1931KPDP/gaOf85Zh1WI/b1P3nBbOoTMdOs+M5TDJ1sDkflGoTlFH4Wz4fHcCy5xRjTcq
1UumZtoKiSnRABAWgUI0aI80Op10gQLI9dlO1mydaxHPSZlKiOzMladDAy2u3zJwpvHLL/xq/Kpy
w3+w7aCqG6s2eWCTidIyBSRsI7zuYzqY6+qrqQf59iCb7J6+vRgCkfoSCZA+XWqNZB5AnDJ3zy/5
yb6cLtDZ/fSv1tjwcCNE8pMpzLrKNujsEL5CeNValXSweAFKlWgQnAy4PnCLfw4jrAXyOxVawgf7
WNf4mmmGKmQ9QfVG+EztYQHXf9t0/mKkerD1HxaDfsdZdOWrLPg7wcQJ51t4Xld95OlfIJwFfnzF
5kVrye/DI5QL7HtfXQ4KIi+sgmXQq1FOwv6YvWvE6ZzwFxg026YV5dus2y3HyF4ywLULLooRqsek
pGPuY69zVlHhx8HQsjWfcUdaXka0uk1SqfnPQHLON9Umo5M6CUKiVLRQ9Fj99zO6wr9lQapLV3CK
KF8EWCctcBsfyeiNVlteihgJshC01pKubT1XSzmwiQASNBmS4DOKyn6mMoWFuk+hqkHlR/5AzQEW
QAlCHG3T1Vs6ynn8zXF6gdfMhMI82n1ZiM3Zf3RjrDGd1MX+pAcVHbK6EQNOJpqle4cVnAxi8WHl
cYKU/Xa5NtHzFn7Z/EmJm/4S7hMbfijXxHOr4NV816O/8p5YV8ULaJmhd6g4VrO+mBgHjh3mD8RO
Njdmmq1Nb1pufJEeXA4zZ+ljJ23kjMZbXeyh54JR+36vckDmkCM12FX6AdIlhpjSH0uoNTPJhO6i
IiNf28fKlbzQWBaL0c3eenUiMCPf7XDsi+BM1yZ3ofGpOGQrxKUJrf5J42tL6bECF/GpUEcjjSqP
EnJhpe1tu5pAjfbx/FB1VLkA3IK++xO8KrODo+DjAsRg9voHAMYGBP7+u4I1y4NMNM9yCfpadUym
+gaPywea+ImmX7bJd2mzHUpZSkLUDAeu59lfU0rU2i9J2lfzt9+bfs4a4k0C8Zpvwdindbk0x/O4
sg2IpD3Kfim3nyxP3gT+7hUE7RrUFoB81R3WDifEpB1vH7JCvUy2dKEE1q48y6cPCzq5yD47kSQE
07DZEGBnm9Aa72tcPfqE+8xhcIcDtG8gTuUchdgX9tsoPeFBpPH1E3uS51LFnDkil0yUnhXR9wwI
Of1Lbmfts1Vq30O55R6M6LnWhC+5HFvsL2GgVlagz+92UiTNGRwxhR/cIM5ApI0OWANGeG8wTGLt
l5HIyQCtKU292keRy0g1TzAPZg6o5745RMaYjrufPM+gKG8NxohU3DVcXOG5F3sIZ9wR37ooZKXH
SOKz/+Uvg1WeoLDfNiv9/wzTTGG5UC/fsye3gjSu2/Vm7+ciK3EVGBih9vleEvm4QrbkyAAZAuS6
IuxztWM01oNYqhoWhPgI2C0urJQUMYtdxSHU6FbTC7L6a1ySEQn8wV+k+s6OuUZ+RiKAd9+R9cbd
wgz0d2TiLqpxwXMRWDO23DkzSWkJV0L+laD9pK5If+P7zhbRl93crKBXzNtmXXwnU7yenVG+gimO
QfHUminWFWVYxiX2AHwVWCZ8XIBJy/qPla8t+23JX/2CdCyHZoySaXKa+zzFX+Kb32UnaltgMiXd
Ay9NVLHHI6xh0VKE5gK3fKqGlkMyzsNQ4Fu5agdRtkXhDfe23NsLO4j87filkb6bj04BcRcOpk/c
RZKz7l1RvwjCvSD0cKmib3JOn9cVCrEP868PHP5GFgPygqVKiW9cUo4rsNi64btBSMT801tyfvCL
xyfW2dbRxrbfzaRBw0oBxlehicoc4jXwdseMeab0GZI0lk3Epcthvfn1qh0uBE1fkN31md7BdV8H
jDkyyVqEr0se+CkvULHX4vZqEh0hbNOU31yp1EoJ/NAEzbxRSU3GwBGURMsSMliynNvrDB5smtqZ
IgbnQeahIo1ItwIVXFJ6KSXpkgV9JwRzkh+E0KTlEE497dO+MRHPGp589FapAYqd3piUXRVaxLcU
nRq+NW2OSJiwtKCMjRQsO43Ofs7uaqXTUkSZZXgRpb+7aAw3yfxJCZU35Q9cfILak/L7T5LGXr3B
nKfra1umb0AeZlSNGtPoD0prKZgmF3P/WjM+84iq63D/EyjAk/Z5a5m90edjCNeaNVJwBthLbq25
HFcy7xj3UZraF2DZO7IKq2AlZ2++mzQ4TlTFgYQiZzjNYhicZjFe8V1bhBYzRH5NfRu8sj0SqTEz
lFQUlA/+qpnsJYQ4OEwS/HnJLRVp8Pc+fH44sChZy8aVT0ygwYkFDiQprTkRzvC/647WCnfGLpRV
XuLKZz1asNtxYdFhEMp5D9vNX5EeewhC+Dqt4KptC4FV5tQMIGsZZivtBOlzNHVcDg/XYQwN4YeI
au3iaoH4d3vTnAryMDLGIboxWCwoCjqBv1DN2xuWMOKB/iuo+xH0IElPDpxuv2yClvlatNdNnhdp
K0eZ3SECk5/+xbn+pkmB/uBy8OpiXMZstz+Fk7Cd9mpgs6Fu/xDWYHeR8DSlyOSqtgKnqJz+gQUW
+rqTJm5kBAiqiFdQT/FbyjOXpnlqnQHDiOrkWb+kDxqkF+Octuz5srP604nOCPQHzLnZJTykuK+D
uNF8O3ybxyYwp3IgbF5QOvqCr63TLQ3Qo63+I0xF7uv7yo3TnCjCvguBLj1wHs7ZMFbP41998AHp
5qHDolmLQ2k8aI63g11EI9pFZQbgsDi1B5vjWZEg7wdgBtpxk/yQNZaitSUk5JcPl3hFvQK0pJtC
s0fNw88WOsAwy/7+Mkk5SqmXF4OEwduxKb9PJUGqjI8PQUFUuofcE5fi73cOLFnYSLXfNsfv/Nhx
BJqpjJhzSJyCzgfCmFcna55/wngoUy7qoRBHidOnFksYFyZXpFuwwwQXEYhE+IcxPdKOOPA24OqM
wYzGZc/soVUEePaf0JqQRB4A4zjov/Ia2Dt7DHMskgkAwbfk8Y3FtsO5MizL0U+8NLa08bZKRQK8
YIqoWjqqixiYxgJ/Y9DLMfuqQ1sOq/QOELEjU7Yhcsa7K+VtDFooR9V+xTqioISgx9VCY925Kt2U
PH00z8FOCN8DY1aCc4WgHMza7xRjjAeF8kNqtx6t3h6qKHPkcZXKZQ657qoB8W1HVz/b6COYm9wo
ULYvNwwpwXUYJjGfXoqIXqVbj23htLY90dbEEhnrc9YDpWVx4ViIriHn5zY5OJdpwo1Xwy3a1e2t
6VjywNSg0OxCQ8vNXqmmebYrs65yCWkxZX3S9h3qtV8FHIQgZq2+Cojw5Uowe5yjgBRDARhVekrE
yK2CmZQ4LKuJEgz8MAOgoDaj+7NldDBKYUZTMHYfSRzlFQbRGjw5ItmlZ5BLBBkjQI2/iSth1AWT
Y7Xp9MYTvrIk9aaCpEfNhkF0YZYYj8dgfUZdjxazNc2QmyaPJ6tslAR3JXMHeWukvhMl/1MAUhpK
aXwUTo84JWZO76aX2b+4s0h9kj/CT0LeK4ukc+UY8dbiWTZlN0K8yvdobhN6CfAyi0Q/GPE40dSz
EjAwBtkhlsocn3A5FckDHbJcXXcTUvpeLg+H9EX76EYEFwKzs0URsZGqfVo+qKi8EnMLSEnxiyBS
+Tu6i0dABjovaZqsnkxk7XmN9BUNY+Nep/0/eylYYYlC0mz6f/fsQMsgQGHeK3/paE1yQFLXd22G
OOKL68ZWybthTalaXOt5jpTUZYATQrb6VwaEmoBJ3o9/R9qBPQ0kjKPSyQEDwkPjCRaBUQVMKMRh
JwbozsbMjWB3RMF1dmd03Tw63NJV9k1+MsloG5OIvIbEQKqogZVKHROFfckLifGQWfZx69lq+mM3
v7tXybe5FMau9gtJOkTg4D28vMZFH8oftwxZRG7IOIGX4BPJe68AKzsWNQ8IU7gGo3xbAKxiGpSx
fZxBbvYJ6GP+iitYWgl0iU55MMRbiR4PSZSCX35LCmWw/V+KnIrUrPv86oTwM4pPOIfTVnPI94MG
1cObJq8tgpQQSa02CW9lxYy6TfDp36mMXNF681ebpK8Xi6vrRVSOzwHn0QhNyEcwHcPZEB4jrP6n
pK0LyHfYUSmpnkWDGc6g9BDCqXbL4RAMtbluMzvI4lOhu9HQTmdIZjRkafeLUmfE+nUKuAH3DAhe
1zLr0RVzoXaja/tYPT/vt72VJl0WpUNhMhZ3zRwjYesQpp6YIDo2hK2iKoR85/pVzlKQL/YiEdqc
2WwThjPsBMIgCHd6RX+8LVN77E6WmI4GI4TtEegEMZbas8gbLCoj2ywkR31EfdU2YeSbrYdYXNK8
/TmKxQVo6jmPYCKmWpNMzhk43y3+Vmg1gGIGdBX+V2JgS+EBKOrRbJGipA31rBkgIoL8jI6k2ATm
BbSs50C5dYMHguWyt7m2MPWaV8d3HlPEDcB+wFLnu8xmxNEVEgTfhjbuRYfM9WUFO4zL23xp/Q2T
cl6h2ZZWJcnggO8WTstSkcQoWJbu3zAda0+u+aKVoU3fK+0061Y0wa4t/SNFfDkVMaBKZSbCqEwF
n9I6GWdo0v8fYVX3HV1Jht7wdeEjMsGyZB8SoF5FsYmbdb6l6eMhxrMqK84isFsjgKbkxR8Y95da
4yVUysOLLK4LSXw8p3nDZqldrGhYZdBwMzVXDt2Y/3Aj/qsZxZUKecsiRMtnjxC5ClAh9djZGWL9
PriRwuM15uyFEZVUdR7sPgezNGh3xanPAbItq8PxeOBYT9tGPwKopMYs6NEd6PwUYjC/yvobLl5g
7cxANnEiBbJjDE8jbBUYs0dYld2V9uFYkjBdxFsSzgGkYfgJLNCGcCMWi01zjNut64rq47nVpIF3
LL0uXyzgdj91gbm4699VLTjbTiM0Hj2oIwpOhXqK3XP9UVeC7lyTOmDazZXmtRv+GWBl5gFj/fk1
IC76Mj80ywqe37GCQ7JzA2qWK71FQSOCJ5u6P2ZUIpziOaepqT+gQpHxBab5raAu9oZPem/VXFgQ
7rqPOkg34KDTSmsZ1JmORpt1Q1dqSCxQzdLyKGXIaZ3+PEAWiL0vQANdTjAs1QWvjrETNrAevs03
od/z9mKWkcK86l3sKpRMl9rFsMy6FP8mXHUtF1OPwEei+0BOp8Qg3+vFVsItP6ORaPEY5JomTpfJ
9c4OseuOjRsRxSHUDikNpQ21YTufchSt1IfvFTJwIuBEA7lIH+2LgqJvUPqY3lNDcty7MROFnxNO
pX9aOfkaoWUNFj20ZH82bBL1Mp5wuh9ZFKc/0jm8Rn3X4Cw8NhRnECIjdYDlunTWOnAsHCkc7pje
p3DZpfw5Fx9SwgHOA0chsKlPeosY+3tLLMHuhAmcBQjcsk9Cq2IYBPEUNoks2cbKYbDLqhnF3LkX
0JxnQU/YzgNwV5MVSZZP+h7NAmsf5/BXPuKdFzK806AQcdBlM8ih71hbGf+Q0AQHgbEKVZjZNBo6
Seb59u1Ijvk3Adl91HB9FK2z6rfHhNToDO/FJ3h7t8D/6RGeQJzuFotmOMcAKOqew8QXwrqW7JWu
58MsymrNvHfQyICcaNm8k02BOO4DZdNeS3+afbKvrhSbQuv1cKo9YBudxJMuINLaDx+8FlKXJMih
uyoEvsRR/26m62zzHwcgkGeob2W3U+83mQ/NanviLd0e5FObO4RogC83widDPb/zuo/9GK4eVKT4
48TYdIlqp4f26HbPM52J/cRLy71jQdjgbyRQ9o55AckJXypE42/RHUh4JbGPYJwKQoUwYdQbdXcH
s+zyahPGwsauKDINWYf0WM+tOdAh2NHL0UU+7nIy4TbDuZD8dtcKTBC0kyi2YotdfaCMKefPPEkH
/bsYN/x5b6uWfNWDa7EF019RRyqcp3gBo9OvPj2rtHB99fyJ5QuQrzRhpgWiHzY6o/SmgeXQmbms
/rAMoYIdSZzojxiPugSnOAV0SC3FBeOlswMEyWMfHgqB+0nf83x6dHYuULP0aZhV1gCFhKj5N1Fx
xTEv9OMSWZQNM0K7DcY+GXxYsrqTMnrZwH1s+DUc5cxhaqFbYVjO/sL1y37d16fQugAg8Ypva7Mn
sEitv4BbzecncorDweaGkvKEfIgwfUU+mzEk0qcq7zR7oqrFA1iQFLjpZcBTjrWc4Q9WGTeABbvm
QL2/EX9eFJTAVGrMESKoEbdLnccmWglIwy4IokLLKBmmm+rz9N11sZDQi8NnyFpDlgNiDjWijVck
ec5nO7K0MdpjHrj7hKhILIlLbPm/2a++Z0eYQeWpM0ca7ihw3LVrKmKrhRI73gml4eqtZxwkWDg/
qNDtKp8upa5qEwEBevtubkBKrGU0Fme0jxX7jfbLeA7kHi4I7hjpFNcXCJzeNm3i3Ee75laUm/JL
57k2A8nsVcRSo3BV5yyG8wRcufvfGXBXrwIxmtGxPZm+LZCOA6/kYOEfFK9GlQG7FGwhTFGNqoPm
zkpqprN+jQNJ6tvjdioAR8Mp44bJcRywVNEDN3kBw4Mit8yCt1fBE33sXv4wlEN5jgOeiRfjwwMe
3gKzLfdPazhjuDrNuMyRPvD/d0/U7M1B3IUK9hNuTgFEbCaSSauY4b9OrAl9IgzcRi6FTkPNOHqX
JTFZgReL9rLPjRatIUg5r76R463xMtNpEUH9sNZ66mNwEmketdRS6BXTb6sXTKFmdRx+LsBfiPPc
a9OXoHIABn2LvR74fNDbELkK0sVnt3DtXK5Z/LF35ZgDFKvbz4ADv1GJIyh7gQVjyOIIQsBdEz4W
5M0+CXtmW6oEQ26+kMTOSzmsIWctC1T1PEku7dHTkVEKpIBUawn+zgObsNg+3IV+rc8m6LL47hN4
weVNa+PuH9h3dwCqptCkmODqudR3DQ6zlOkiOq2NrUWk64RhZ3WB/Sm71j5ZMm+65/DsYrJewCn1
XpioRdET/jlQaUgTUcH94Apl9MGiJcQfOsw4Y3jrLykPpNgRG8ukzeXJ2+VcK1B+/ew+tRdhptqW
WR8mrn1nZj3zdfuB3iTvsANdLazpJa51xbxcalr4gZPGvBR5c5LQfSKAie2LWGeJeUiGb21hlL2u
ZDmsmGONz89Vh8mMWMVWJWpYuGi+CALs3XIajksz9XOGDf5RTvIOLq/Z2ybKfCU5mieELAcl1yo6
jb+nGbJ7Gkzw2pJmcn3Y82Bq21K6S2IoaFXq+Zy65YnOWENf/NOEPAPZSFkZfaaDgU0I+taR5jZv
Y/fG539kZOYv2PpKAbQo9mMTIA1GhY4107Ii7lyN8V9RQFIaJVXDuEUMejB+LhJr3KZ7kNRV/+v6
aZ8UsTmadYZpwmS929hvNAGAPp2hnI0zbujy6wOlYEqXWVDkx16Xk6GWAg9qv6G+Leh9TMyOsmlb
wn+IRKfM3a9aJ73YDDiMIViwnGTZ/NiHml6daVWrSdwYirtw6DvCXBCt8rUIfRKp5f6QF/ZSYn84
0FiMmr1OO3JQA0B4hlE4c0THMF4rkizQbi3Pi5vdn0vlmAr1Kh6rwdjDKcQDhoN6aTxDer8ATY+N
tPeXfvj7O0Tdo5B50jU3BvDz9gS7OSBikg9Ogk7ciQAYyith9UIehjHQfuYqKGJjfA+LclylqNzP
taJyftb3Mytj9xDz6GhcLwrrfeih2IJaF7rRa2Uzx6LtuHtgI7+9mlRwdNNnaUFrUtwbwNJY9O6S
a9fl6c7C/27AbYTlTIIQta4567alqMOpEWocOxK08AkgHuiAVB3xsGLZ3dBBwkRMzHE3DD89aa6t
vamTJtj5BLq4wS49+lVA1nyK7HqQhYdIQPbHuuM2TeyOtkg8Ihw//WfTW9YNdKeBuWfrlW7iUfem
lcTNWmSw1Zy00yQwr5lNjTcKepiiqx9MbCdU6YHKXMjtOiQaNC7CzGOR5hgF2ILNXPwocpvG7JPT
OrH0ZeA7fI2cSX5LlRXpvvaDQ2F4koETyBrGBfNerkRfmJ/M6/8rxZUw13pVzrVrJD+6d1pHTMFw
aJCIcTnwgr5XuQ1z91IKJGDCtjWD5/sUS40mtBvYrskDGqTtKH4O8Yy5MxLF+KLiHqvv8FvIM8xq
E6oISA5/5mXdH7G+IZ+kZlm2+20P298uI8qvc5SSZQA0NMlfCKVQZPIs3k/Lzvbbp+j4UJd+XSmW
pHz2S3B5uvZCY6JsmR1rrp6ROMsTYQ15I1OmlKKiTD9YbItMVbt/NNhmBydet/SswlRLJjgMOXIc
jrv+R+F3dx1dcCHPLRjL6tMUA2yby9B2bp51iWBzk54O9SPbc47JHgeWAnyD51mD4gC18JWaSxTM
jVfUa517BTsJ9LysBmseD0bf9r4HQY3X0Cby8fnCGJuyxjJc87szQNUdLLplFWFepaOm4YSmy2ob
eWukJ/P3Kt6ZXj1572rcIkGMj2m2g/zhMiP8qbXknH39Qs9R+ZaX/uUFI37da+WSY/QjTVF05Foj
hjyF6MMzJLeRvkouzuMHAXw16uNZuoejV1JkkhUzctFu6RWPgTn7wwKFDkQRt0ClIgO1bJVQ7Nw7
rxhKNQLvyRSg98waZe78I6MogIN6NWDdiNtm0jZesiXhwvGeh0Hy6k0YGJ9ZWkXQvjWfbcRuDYiW
iIh2EUqgIeYUC7/ErC0WPh155Pe36jiS0v8RWdMP1DTug0z2TS3IR9ZOYh/I2P06ts0DXM7Wwebe
p5buWHfoE3jUWeZE/ft5SNE6pevEFUicA9MzkJmvw8Vc0bJUnz+megBFawjDNtY/TwdjXIfbhRCd
w/aE+JoTf5c0WbyAi32z64MV2R0jRuzS3xpV45Yb616luhV78PaXui6v+qkN7kvkOhXtalSsYoED
FTbF5EbQTv/td/+J9kziSpgsGsah0KJiCuJItLZym9c+um53xOkvO4mql5hQvOWQV/PZxECpSTG+
XkJ7uv/AqWZgJrOLkuRKvvSdA1XhvXQWIR3NZ/P1lz8XTEbcHzpOWMf34LJVs7vPA7SMlZ2mgoE2
raNfkEjc9u969P5+vGg3MHA4/QfGJMio2xa51ul5csE36OuPG7tASZv+8o0Ajc0AU45ic/uSvtYc
isAwmvzr5o1T+STtnLJf2CQn0noMPPXQXN5vW31fo5aHbygwcSs8/z+AxXGw01vjv/K7tbgoAk8r
YAcJQizdRa+vKqqbvskpTz9CR2SNA5kiZzjZQOeBv2crxf7giAX7noCWQn71yr3BsPkfg1EIO4yF
fKl6hixMtTbc/7APIOQw9l16YJyxnHUrdHUNQFeSy+ofLZ66dPF6yZ/SBzDO48x2qMiJmx0UjZOc
FPkmB13gT2GPYW5VYBF1bHt6raPebKsIJjLsze93+QySuA5QPBPgtk2cbVIk60mrzOd5+dNORQTN
kWxkvivmgc7OYM1phXLbkYaBo9L4IJatu7//bm9Hk7yeQTYNhJDE43l4/i6/y57gXEhfjnDDnxYA
bfsg9OjCyrU4BubQmp5laQxIoHm+l3CgaEv/AONpjXf4EyNGgsceddYNlfXm2DnNrbOdHOvL+qfO
F4S9ggwHcw9N0T7ImOxWOENAOjMDW1PC9b41ukMgTTNJrMEpS+GUFKdiTtmn7UxC7LeQZdhYGM3U
ecQw/w4j29O1zinpZOwuqxkzWPdQecCCp1n9XDn/11JwdMlS/dM23bxYoD1PNKwpNotvPjAEDQNJ
zJAcsVsWJjXIqsUHDBpNxRtxc7PuzCYxcSVxf0JO2p70u3cqmw0wGL2HNYMDVMuFosBWGlOXOl59
NZdrlMK8U0uSS6oBaDqXphkeHNcuPC9L0VUOrzcVf14V2tdAjszrC6IRoPCMWFYSk9YlmTtsiUr2
4RJ16ZMWv6gpYSlxZ6yCfD/lZDUVdyKnOPxc7xPNluwQlyGqFpQSCocjxZqLtFwiPgunJJoeBTUg
jDR1a7YVPhlT6caUAcht3l8W3bKly4gNR456jppECaAuy6W9ZjKZiJnsdjvBf6F8cH/ED/BfsUAx
aXdvo9aHjF4a3ECmhckWJ3ZHY8vyy68CDpuh8l5uNJyaMaHsWU/CchBW4JS+X2lcDCfjP+NEoY+M
p/b2Uh+QJC4FGK/Pr0qb8vXG1IIRiYtvR+1img43KUhopSqC/dxly+mwfitB8BGE/VWqRPVyYcUP
UKX0O6bj+daeTW8/Sf8oUIzlZEcfEM7a2QawovmExAuAS5jFKjxMZQRrJn0kTIc/vKphwg3Lgf7d
unsgY+xPc13c6vH6i44LNxJ81RItePACI+lcIpyoetC0VeclndvXGB+Oy04695FOLIFhu0Y9vayx
IiuYPcOhys4QsvLsQUHNbAny+FXLBnrekzd0/G4RpLxq3C8Mm1CKydQy4dH0z/7djz6lZKtIkeAI
MZc6XERu+eZ2GHvHLVcBiXR5L475cbgOvcqlPhNUnQjU0eusznl+PmAlFfIm/TlRVbWC546vBLxA
UMiOeP+3gmK8rzxfL0JQcegvekS+XuGbr1Mzevrm0kT/3lDqT42bHuuLjR4AH91aurvZeS4Uib8w
9DBGqoStZ8OhbLRG2rZt7G5eKeMbZGW13g7QvfBzpUoIRzVqPXd6USTXPSHRHdTFhTromROfWJeW
3BWRHDw9FePTXMgsuJf2MEjQ+TUN0T7CiUTZNNZvYdbdUWyTgTGMYp8KBuc2NOrJNSvozccZseGP
XAXnBBNti7hOeYZLbRT6a6Xu1d9m9wu/nvd2rhCtdrUh7hikdfdmtCVUC8xV52M5gk0xOcbvRvi/
8O0sbVCRjrC28o2InT0ieChrVmZjYfy2OwZ1+GFl+XwaXvZFEqF3aFbP9zPRCByWw/BFHUVJaboC
gkHWu5yg7E5Vr63r6N4a6Zk7qC9cBPC1pO/lf3q+GGEYkn2P8z/jpKmb84f6617UL3KC+3vL8upv
0LrWRlyoU61sl1AfUIh24KKzKtW80QGu8Nd+kInJ//uto3A34LB+KXx48OlWv8MlYDbe6hBPqPOj
dbw547zVLKp8SoOUrxMLMuWVuqhfVUBg55AUQF32Lm0aNnB3xy+luQ0vV+CC4J3zSvdX71ge2e7l
NoetOq195jvVhZqtZz1mKSRsDuqWgYtji1cLk4wXxLcxeuaNrUqnmEx7TWtGyTiQJitcZRXQzyGI
Pfzxe6hJGGZACDHuc8hAnEtZzNozcFGX6yipzQAM2B15ZYoFuRVQ54/4FXo1K2lJHLHMxmEveL6b
/m504mhxJ0xx4FK+w2WlApfIqeVlt5xJj+vaAAeLeGmvNbe0vEEICpCuJr/yutBpf9w+KdTI8h4A
yipEFONvsr9DxeqJjp1XTA6Xsw8k1lQoTWOrcKXTpXR7ffq8M9T21WKxNR7IhAX0dedyWjPMGSso
28xrpMcvjdj6iyg82PEvgS489Q02S6TKYIHxtbCpb1i6vHNa2F29wOzY1sNfLQLMreRtRWokK9ee
ijDKg4WUSCo9qvimim9FHCvcxy+OifvPwLO0+eqz9A0V54wOSCMmvdc6InhOXd+W3KnegCAJ6SXd
aIvSetgA2PG9aupH56lxWKmiunWMMDlXtyE6MTSA+uv/Neu+1y/GTicTSUbJQYgYD9v3vOCey7RD
EeUij7IHxG8m8VC00ij78AJseoRayQ4PjZf9khQaRMDsKlqDV2l26QA0RbdjG/hqpVeGrd+rUQH4
KL818uqp1Awe0BdaG3nbvt5vxpgF+c723mz8Ek1ffgAGIDFdOdpWnZzk8NNcSEMx/V6WgHih8+I3
MwOt146UE1QWGiP2yyDyN1eyIyhbL8mkNpgcBVuLAKMD27pOV49R1f1OIdnf6afe4yPuEWJobcOT
UYVBaZ04K/Uj+0A7RAVFj1hrbFULHbTIYax7zwqSQ4gXy8Wy+xy8Oo1OO05Ogxf8FPWA7kXr/GVe
yTUowRy1hZbH3zdOZ4pGzVQwiZrP/0ChTxUZfc5JD1zrL3EGDbdXaUAdxj22aEVPYfQp34gG/0uT
3+VcUrHVaH6Jws+8CbOXQW3YQZdgXG/gMuiqWAx8X1LWusz+ZGKQRvW9QFEEg/h6qwEXHp3t00s2
5yU3lYWzJkzaRQ07e7kXuAjEhl/S+JjbmF5+Sb50F/qUpWTgX2ATsL6vT8XEH2qWXsIBLtJlxZRv
LuyyTwfxnmqvR+x4I5rBzrpdFYGrG3NrvaL0oIafbj/mr6uK4UyE6ylHlzZAEnKCYTEFb4X1cdCk
zIu8uRdfp8PPb93eAfBiMsmRKBnVNrZa6buzkT7FFFNjBz2/pdFGejvnkabYMtnYYVg88zrN7gUA
1huu937L4CUA0/pFG4nQFcUTRVoR8YK2gld8bQSzZQ5g0Tc7lkXqVXsvvBCHORgYJAC6tpFu2Ns6
O9kVEzzkiOcSfSsH5GyA5oY+7Hvo2LeWzKjd+aDe5V0WWApsgo+67WErBZ21xLhJYFIOWMP9p1cZ
JWhjaF2EAVjCV/7tAus6knrq3LlczrTn9+4SR2I8lzR501PBAinD74kOw5h0uzBM8grfyqGckkS2
fjVI8NyRuNLZmwNtv6cw153q5TM+dIcp2gfQBH5PFW6ykE1sKluPLlkh95DV0JXsmiNIIcW6X8mQ
vg2tbhzufC/frOJ7UZPDJ9M8sO313PE6RgIh27G5vHEkEXjctGj9S4Yjff6TgD8IkqDAltXUQnjC
P2lmFkXG/ikesKsNLWlYnusoZYJPGlMA/spyb4OakLwQfYf1qacE5+42RP/Dfy+zRdnWd+0r0YgU
zd0GIgRxuNNFcYvHn30Q9DKlcsIKo030lJjiq+Jo0I9FjNLKTPPCI7xR5bdSovEBJZY8nuFBLQIs
wJI7pkQyZtfHQ24JOYsHVT7pyfCzo9U4CvFuivst8/1uX5F2xnAZqs6HPSMF9406tvmipcLrazX/
utnoZXl93phayVAB0aPWGXYLLjSYq4yT/R8lL6lvm8ZJBACnR8U7T3l7sRyD7tVgJZSl3Tkjkb+W
1cP5cXLS1eygM6vuPzFL9O/7bz2qGx4cUMx8FK1eTnyFlsb7TQiQPxGgqDwR89qsbw+426yQ0PlT
jKjpZamebKjb2VeHbpU7QxH+HzzCYjzv5iL9rylcoshUZMvvO5vzzQPJY+PZMudrzv8zgMve40PC
JSxuqfBTnbuyPQi7+ZFG7zmUWsZCfC2Ju+FZ+iQpFfU9KcVixrkbcouMpqcL8kElZUX67tOS4Udc
bgOyKh5Mpa3ukuNTOrf9uPVkET64KlZI1pMpStsqpOE0R5pS0ETvgF1UAdUTHZaakqUL62QfR39q
E0TQfw+xLiQCvlyXLr5Ac3dnaM4CprRBfDnyXlQeUxeF0YGGHjfjrb5YEIowyjcQji4e0u4Fkxcq
kWXd+Tpl5kFxHdZ2mzZvTDBJPbNPeklDEU+pCStwNgwMVoeuYqw8jYu0OEAJGlEL0zafiORJUkKd
BrW/CVt6+Qmv/SFu2QTMcCim6G2LRAd4J0iCuKE8V3E0z4BiuWZVu7k0f/0Alja2AYP+nKzqLmGa
KbdqlSivNzuSE/ZYCi9PksHeouyPYwJ8Dzpaa3o4irIyKO9U2flSYrUXZIeAx4RRVyNTd5Bsfr/y
xj2AhMf5XbnRVr9n2VPNIrP86l1PqKjSijx+A55kEG+If/WLlbCBRaAj0X/T6WjSX4/JAGEyVBbc
g2x9A1rRwvJdKdfhRPRFRfvIy4xDfPVEF5T3VUlBgzrdmakSOwze1bIRv7o7uupSdxSHkPQxeEKy
KgTqKWvx3g1I7ey0Mu2ZgbWX3L6VAygDl9jUyN9B49xT7di755/05ng4NX9QF55PYmd7aJflBUlJ
h62YvBJLIRP1op3lEWVm0WgtXYFqIJ60DNcjQ5A9LfjhFlgPwzwdB5IcsxVcljdpsfBu5FgEJmsr
mJAiy/Y4u4SV9VP2y6J/Rt9d5Yg0FPmzHcdouKAtUV8zp2q1UqdZNU+/IxSDgbcd4XwKHG6Nxhj7
305+gZvtwYawCuxdcsS0Ro+m0W5WosNupZ+kG0lSoakdGMlc3g5lrZApoY/pjrXSTpw9FsK3j6gu
iLDsz8cZ3aapdDuw2X3tGrba4LeO8j/0b+FjdsktdC1oQAe1SeI1Zf3kQ7kTkHz4H0rP3deI5zvM
bTWGcjIhHE3wi+fLQEu+4MIi27hAwuuC0xmzPWST60905dIcBRucwn+KsFha36OwASyTVxEyYNOa
oMV9Nzi6Tsn99eH7LX41M5IfFucy/yMsANl2hV96+U0U/dlywo6Hf0etOGJZigkplICR4879yfcr
doBL8NHxihT2XsD3daMhfrsTinnMDI0Ia+zGJWluTKR2FXPcDEFCh8BYxsQrba6iRQCn6ZVWUqER
d9ValaYERvUW5na0gu+fkrvod9jI9Nu1NZsXq6tcCzKGvkY67m4p69FgIfkMCsnIrpFAUboi7wYk
tQBnbSfOBUhPPVXtzFMcJqbU+R83LRcXhOyyE5AQlyeT5yjhgTWLu7pG1RbSKLf/NlLvTbEqw2/5
lusINtCHiQKpR7eiYGVfOKxDFg4ts7PjiremCmjw+D/6A39JP37lc/DCOS0OQhOIziJ7MG21Bjy3
h6bmx2Cfov6WUuLM26KJWOoYMiKv4SDS3K7ZF0O5lDCrgF/SSBi/rwiVWOXpScfYuhpp2D0hJP+6
rJ6uWSgwC0wAKGuhoK1K8XTCYMJWOnovR4tcSukyla4QZyVnO2Gd47+TGeIy2dPnqMHZGp6DFm/J
XALm9QPIPTJND4jv4cF1A5SUfM2o3Hm6LnfS1KwdzwSLg5t+ZjSea2xXIptSEWY4fQPyRR8nkZ0x
mpptFCgP3d6UJvcNgYBD4HFaGNS4JAwuB2qwTQiDfF8rvwXREQUpVpJJAxaiDVKlqeIcfHTnuetC
Nvc1dkIggyaOul+r5cuz0xkx0SsERM8s/qcapxuq3eWJJ7patUF9amJsMAeNgVD90g+OH6+BBMiS
e4NxZN9+qh0tNlHcYvIAQUX2WY1KsLbKZ6H5gVFEMg7c4smDFKyFLXvaklMFyL4nsEp+EQOJXnaw
nmnYOtBXZlRccmVujqzs7m+xac1TJjCLK+gbc3lC4MJe5lcrF1DywB2LXskDlBfFuJEzq93i8Suf
aHcRfguT8d5p8t9FbJh5y1jb+GL8E7wr31J9NtIGD7BF2SgAkFSc3qRgIzKHyGismFUIPMdzLWxP
n5m6WrBdrfHvf78oYpYOt6AgmJJp0fHTIUakWzbvxPYFz294XcY2sacOfoc6byzYS9EZZJcorSJ7
Dy+8wHPqiFlUAaZEl+0Qd0VMfWgPyAhKE4GzI0KZ/WO49tZe8VFCrQfj0HDvpVCuLyLgrHkQQOIk
0+gaFVC2wE4hgymWeImWJ/pE7fV9aHbvoBTMf6hJ7t39rIBqkiFUyhJCypwLTHpbSb+xXGvfFWUk
fFx4jpmjsYqFDkF/qMc+3KaRY1y48xieBSzuzx4tzKgCFUZJQ6vp6X6ZrRaGDHUC7PZESXj7tTfX
f8u405t5n2y2iJDl8NWGTgjRQmcrjObjZsDOqCvGCSqGjdQ1XgMS2u12DLuU/ok76EM+ybAZ6CF6
CnLsSsH4Sb11Mf2/gezolTUEy1cHGf0GdY0oTDncqYpCMIaV8cuaLv2sIV7dlvjg9tpgSuNSOSjQ
z6kPajz+Zem8oCE/JElBUF1Jfa+NCAi6ZtiyiXeTq/D8nwvcWJxfnjzqMZHC2xCon33TUby01hVe
n/ejij8FxAXdxfTLGpNAUT30wu4TRQPSeX+RcjIBrvyTiplSIv8VyjYTjBKwaH4MAgh3uFBluhaP
XjJJ5tYgEjCKzWth7b9GL54TU1gC8pS+h0SFGv5jPeC3Zc+IC8wO/gIiHabPg+oCKR4exg7uZ98s
cNtsxPyHW1BVRBB/fGYwRsPP+jDxIYCYTKg7IuIJTJi/L0SKJ0c+ViTJtBJsruqsrJ3O6/uTNhPD
k0+jN1dANEqVISX56FTuBSoFgULKhfs5/k34rMdYPF02gXiIbGgNNGPehryRva1eLzK6WBMNPA4B
4aCGhh2zwqVg31N+9QQ8OB4k46P1cSovzMZAQP+Z4WkL97BI4PRRS0PnlyCyk1cZp5+aVLNTaTAH
SNxnjkzQKLIhsZso9eyZjIpmDMpWHaeCwCUTycD9tRJ4Hor3z+kXzPPSeAFlb6jlqoUogQ4YDA0w
JZmY24XCo8fjRQDmcpevyGkyIgsNgYzhHOe2vOojunC+WnimDbgeSSO1fWXDwHnPFFcnYwrgyjph
RXY2uuDJAAnZYf1wXyJC2NmIEqlITHsS7cHsA/arCLDMwcObc8fPedGQRWwNjr5yJOnjOfwUsIxm
niOVXbDBklYfqQ0685VTlxzzZ4dLKF+SL8r+L1NzqPWMlRm9X9eKtKdbQ84GLzJFSI2Z1nPz5j10
4cuKFHKz0QVxFeWnvFuPQe0ugAl/+eGgkuzkbUI0Zu5N1ReHN5dIM1yrrabGz2iM1edXRmUAl1J8
PJGHiTg87zEiAp9uKUI5dFMp1ZThk6LJt3SW8gr9wmhTjc/1vsuoy4zGeUmCGBhiFO7BEDC7CtLC
ABwA7//v7pd4yRws6wbjeKylSAX9PMBfl196QfQPK6dRJmvVyYB0PkxBORU2/FZ8FB6MeoO8snyC
Wg5RtnrOmvmf8dJt9jfQtGsM5MF/dwqFmX+oo0C05hrYMxcPSZBibL5yHvvCcdP2N2leDV2NFsD5
S435hazo5zAQXFcy+Y0H73zbXo6ZtlsjHPMmdJVJqLY4E18r8H4UocnSPKVjDztUYAdnjRUjMX3i
ggPHb3yXDvvN8f9zIr6XWauVqkYXGzRKnjooiu+UUNViYQ2naLAFC5aw8IDwy/SF5JRdMTeE6VoN
MIpVyEGOWya/e+Jrm4D8ofZeLnPiOcDqcwLdf+JUfANdi4KPWIFBs18Fh+/wttRPsBxjt9QjfLTx
ohnT+pAEZgaz5Pe4jU9sFvwT2XdakUJlzQUE+P/3GbiMQdx6x2fazqWrFZMu76hkJcg6zrjqYIou
NUSXT7YlI919ibQscz1JANoo/ZKSgbnXaJ2GmV5/ACFTTUNQjLgASYVJ35cJkZAlZ3wDOHiCY2tj
ZEZ1MQaHdqxn/p5TNi42yodm+KuyUw9GxV8csYv+Eze504XCarXjd/8zdlLWtQVQhr8e1e/cqpqC
YJM4G1huimObphrb8hYdU1am869FZUz5HrzPFpqCZAP/C7EHSonRKytqYPt8R8JuRgKiwvcJQ7hp
CNEBwYzvZ6EJvhrbwxPNftIylNsIuIZ4Ga+k6uhx5WPaBfPs21Io/O88WMUancim0/AmCs+RGmKK
WZwXZwynDMQaRMHqzudX+H8v2DejGw2GUkvfNIO2ykLVHk3dMx0fior5FEnIjLcs7tsjtwwFATp3
RXJs0kCCDlrZE1BeA27GEcb7QbGljq/DjGRmoxwFW5Da1sKB1NgOdStjFyWIgquXIITzyynrsVmV
lUuBbfydCTaalvgpM5P4UAIW8uMTtG5CbxHLAfSdAaH/LzHfEolbeLJ46lPsd432uRqOempsJBYK
umuXsrsbi0glM94Tg3UKJ+est37y8j3fEOLa8m6SmSxOeyPjuW1mx7waYcR9StniS27O1DXgAsjr
c71LOjWsxuRibrFgnnn08BNGHD478MPBOzkXT1/9fJCJibNPjH+oqdN5Uuk3q1afXCqja0FMHW5g
P/nbYSb9DOF9IPVbNU7PQNnTpFSNj20R5i9F2LJ5auUzolds0q7FzKc8I0cvmS5NFP4tVtZHQR5i
P7pa9OpAfyiIAuzXfTVQV2/qyTM1+bz6v0iTgaFsVYyAXiziK/mmFNAi9IdDq/r2h2Xdh6Ku3p/2
Ky0AynmFFC6ZipaxcYzow0+rhMIquCAk2qDeDHB3PcQwKRF9yrPO4ba+n5oaF3rDNY/k5nlYMvsI
1lIxOShcGl/idfepHvRoWjjHR4dDBebQlkJp7vRagAd5w8mH383zk6L1ejEsl2O+lpWndrmnL9MK
ZniXW4Yjc1gP0SWCSg5cH/DHiBF7R68bYVwzbKSa1loV5jlNE+RjZ2Jf709iNaLxWyhk5Van/pZK
JFxe79rKHGiT55yVORrwGVJzrcPm7nhPiD28Sjrq5McgrWUy/IdHGiQ+YHAu8/O5fSRHScF98l8H
DB5zhsfaPAAljpmU0GYQnG6dXWPM7mbzn9X33gMPut5gHTpknmp9MsIFvg09CQmy1n96JcA1Ax4/
eF6rpsPBLbXseqceAvGcU/mHQAswzm1FMvA31inpKLnNUt4XDcrkjtqVkCDHFdqHD+2U8Hzpk0it
mefTt8+qVTzppNmELLyDRvu03HupYl1BidUxhx8rZyhq0uX1tslgLdJ1fl88w9pkAI81wMjboSID
g7Kktm80o+v1Xx8/ZYI9KKWj+E/PtBtPQ1w1AY3ors1ZfUD+JKLDJE3zlFa+/SOVPOSiRD5XFaOp
kKcLgIdb7MhZbS4k8Dlda8qzPnSA6b6GMwuj4tznjSwQqkkk7q4dHsSAX/Numg2scc2sS/dJbh4l
GPRU32GV7S3qKtTZBD8q0meDkVmpMUQeMwqB32gZLuoYfQt0Uo7/2aop3m0RwelFL+rEN5WfmReF
lRT3dJ3vNiw8vWYyJ1VUBTsHJEjagXKsXwAhZw9eELe5Tj/+IC4rZjayvcBH58c+CYvTEeH+pWSB
4InlwTVW5Aq91dViwwQKTuQHrbMsfioVDa75FusquDk/Nr6Fknse3uOCmau5/Pv/l1Re15iH7SFA
nDzuRNrMVqDhHHVbXfLjnzyqDeveaZn0/jWD/ApLpf/ccDuQtyOR6YUug6jt0WxDeuckam7QtMx0
B+Jy6Ek4PXgQkK18IURG+UABqHi97gMqECQdw7mMjxNqbr81/8vMEMfL1C9hIjGNeXg05e66aPg0
NFei4OUEk11+DJV5iuJy8fX/iMtpRAT+E2AQZN4SeTmpJ9lBNaNm2pNRcsp0OpO5gnN0QH9a/sur
AuI5IIHHRdG9nDXB9MikwFVQWa2R1xVHB4HxOO7NfQPR8dWtSCgjKO0JUUmRxk9vnDFx7rALGJOE
TvM0nOx1ouTcip4rkyphIBMNJLoiuIO6Ub5DQVNh5vPFKprY6S55PiuW1IX7VlyqSA28g+3jzdVg
Jl8De+wYiidHoU7e/o1HgDkbyGA+Ha5R+f61tMHsXP94eq6cLLCOC/R+ozl4qAYSG0DC7LnOyUPG
+YRTWKnu/hSNDURTmBEbTKsNNuvPKwpW0ZLGmrOruHazl3HgNoJSgMbw4O6nfKeyua1c6yuaUEzi
OetYZHDrxm4cIehag4TaSDUCtzhAdCMvh8ODGZE+1EAqVeRG5lbfoD2+WIYFRkqsIK35XIxZGpXZ
qM95oqOWxuAIx3RQthWbPDWrYwzt5/oXKLfrQsgMEmze5HGYqMYtYP6Ma8TxW3d5X1xEgZpQ0Zzk
1hfsjNcT0uRj7VhIHPHiUqqhqm99RmmCf+EkqZN6j9ujKyZMrPWNlCxyBP2lVn4Yn01s37HlPWKo
ecVtx0XZIjgv4cE7xvUUErYDYGdVv/5LB6md8tHh/bKZm2P7w6pTIHkV5AQkEeDcgyGf157GfNqp
j4LMY6/SXHb5MGph+vs+92yerRg1xUOsMsA6wvzyVS5C/nTI6k5LLVWC0ITgfadi/WlPzmc15dx2
L1ET4xiKfV1Oc1jRlt5IXhNUWJLYKe6ildY+tDxPrgIbi08cSn9J6dM4CLVN6A1eyqiqiYAe5gdr
r7FWLXL0LQL/UuBVMyQEF2sN4X9FvlYeGIMqx6vs89tXsOpryF/vI9RciElwPMueSi/ot93/4sNK
PeV6gLxiFP9MwvMi37M9JKBoB8duaUqskWBqvLsh7QEwvBPmuXxCxPRFjBcNCtvpZfzD2LBFGnFa
KZfFMCo0Y7noQl391qdb1+U+dBc0gLf3RoLaXsjdQvby5TY2B9GruBRMZIHNMnTLsHf0FJF8opTq
Q7K9QvhZwjKGJzcqwlbyBr3QH87shZZcOeZdRmfDbQtgrtaApbjGUKNvvy6S3+6LhtRnr1j7fUPM
byvOnhY2zxDy4FnE/91ma46r1d0hp67Ofqc2NNfX8J8tZ6OBuA938cuUkGg2eVK4TJy1AVs2ThU8
9xmYR74wtXbePOz6wt/xNWu01GnHXtZzt0b0/lI46Ci3sxLnxGuVOHjp6ZHYantRq0b41MHCZNqW
HBrqa3w/F1lUH/TenoswJR5qnFfoRDVz+Dth0HbonYxq8XHfNP6x/q5PBavhA2dpP5EoU99o5TXK
+48Pg714lVSUqe68LGBxbZaHcvQEnIYdjNzerD9jc8zuEkJ5BoHXYkHnq32bSr/qjoCPxfdon/R2
V0rpN05EfOniT+LinT9+3VG/AqwbCnssz11MX8Zj/Cqe93rp6EvwiwvagQzDUo6nCiuuFwDmWvUl
O9/KjHU9oJ60hY4Cm3N8xiH+ydlpQhud51taN3XOlN3wpo+rHmMCemCzWJy9f6ZJxdtOJXITsjbb
4Tz+xTfmold5YAfLWoi7+/DUmU3TOEMHgbypVMXzQwiMMjhCedjl/RzryfsdHTellt4Xeg7QORPM
gPmnc1mQXLRK9VNMc1QcqwBy4nBIsrq7dhScdr7VnT9s2YFms1xf6QjiZeUqW6nYSnIqC0z/tfHy
NQmXCoP1H9x1+bZBV29dZbladly8HCFgG+zoDPB7y9MTYOOVjogFyzIETW7//vT8ePCvRpZMuIXM
RqaiURXiEgXAuP3XRAyGk3ZpAaCuD8YOwJDg1+/AJsbXVVCETrZqx21soHVeTq1XMTLRfA6BGfSQ
6Ibph5Kaqx2jTQNXt8ff3gd/Lii4BJYLLIVLgZc1rIiR/PaBEbV7yNiEPxl3ZSMjR/i72gYrxaRD
GIDIQOECxCKVgwkupn81LVUfI+e0XyYZvg/6pL7cDOpaj2mpH89kIiDQpoHHQJtZUxhN/SVNBhkc
VcUYmStGmj39DBc8yDhcNZYaYtcGunNsoRYWZJDZgUBr9QNz0vfpVnTqBmoSMgc3c5yY9FhQqErE
+ZYIu2/ipDI07MDXWcsbVO4XqUyJKLxVJGwVbUc+ufHqpIHeKbH6hvF1sLKZr/6LhqC9mTUwuMvJ
pHl8fFyUaV4ykRhJ9cB0AswbUk9zb0KKHoNJclZ7oA/pq3iwOvQ9WaXh4F2SXquaJPN9AqHHoDGt
Wpj9NCJ71YF6sIV00q1PuTlwDy/3ml9YVk9M49hh5G5IroEhOHcWBSDIKtML2rICVTustVNogJsv
V4Jf4eHSCYEnLFFaphgPG9e+ZORnpQvV1xigpopFTO9aOtj5DEbti39/CM+gYHYkeA5plcd+SD9y
Ic5cfZUQAHHWlMk/pLQdiEfrYV0+2+nv5gq45urtZ5z9UogWEGGV+EQdbxGLVtwm5Tp4FIgoWlcH
bU67tO57yGT5eq0neddEM/UmxYru1mUVWlpjqvZU3Rt466kRRcJ/NNwfGBBeww6m93EEDPesEvwx
0iQIRdE2KUOQthiFbFqUW0p+sk/5hUQQobSoS0nAHJozUHMai7pfqNtoN6I5VZIkqSJ40THXGwE0
fE7PlHScySzRfzt8HrwuvTcXukVo6c96PixS6D/nQpTVUIeX7HsWJe7h311v0uLFUh5XENubd/sz
VFG4hZ0lfutou7qdhEQiwVi4rjBIusFrOLrMke+qUBeIfdRhDHVyQ4PFNtya48ylIQfy7VAflgRc
ZeAAkSDYuASZTIoK8XxpDdrVQ/M9FiaTztdXysR92gbDzx/RzG+AKzKhiVowzw8o7Y6W2MSRAMc2
B9DmJK1QKGE2xd/VFU/B2FO4rKug/Jl8t4rgJN699uoHMpIzIRdWK0icQKYQszKLOhlph6ynybey
x4qEbLdoUBy8QAuTeT8+SnVEG4FkdWrebXnWoNTVqfik8RYrqXu/aTYrzBDgFJn8KDd9Hi57Fkb+
0Y/j0VwVeHuzxeeNY8EekCMx+F02/4ksP7iWGh8tMU/MIZ8vr4LzK3sTLE/ZNZ92HnulRWMQgxA6
8wd0NqSHia8ekftnhw2rdGpFaY8gmVZG6dvRGseoIGJ0PVJZ8D+6zg1WiF/N2Sww0KSrEfoFOZmG
Ep/hzqi5X2hbF83fiNWX3MECXCb+U2/UgsQt8AYnF9g/CFzV4bxdK7WX3cufx28k+dIFaCBm+zE2
5tq+7m5iZGXJkqaLO9bAztw1OrfHSoG0CWVNqcHcmNBTfK9ifbsdDFJJ8AEknxq6fF5wfwuCns0A
g/kiDXu6NIZbQetzi9LxYHy7cSoN3WkVxp3fNtUzDigC16wQGASBYQCS2hwNO/Nbj4Q84Tjj+t6p
xRS3sXbhAmnGqNzZW1fXoW/Hz5ZyozXw8FoZ9UvHLZXBa1oHCcoJTgKkRiQt4pzTKPk3qyLlLjXg
k51Lhpg7S9PUOd82rZfjBuOZChb1HI7zYCFI7W14XNyALoth++nayfZrF2dgUlPsaDXZ99AnH7Ub
r0z2SWtk9iHtP0EBswnD0c5gxPyRjDzPs8FiFw4bocaCMrV/bdrAamRgvMu69ZpNJGsr1IWDEbg2
m2mee9LDANX0PA9lyU2fLZrFOTYqsK03jqQu850rlan1xQBLBxDaaMytIG7VwSbuUsfCKRqN8i67
z7yUBBBh2aXdeq5xWCKWOLWaYJswnIEDIwz9nTOJau0Sj4sAvzzell1Um/De1AVyOxkcnQxl/mkm
iNxnNwYyapcaYpHEST1GHccfnfOFw9DF35HxUvJF2Ix4G/PzjH3NyxEBJVeyJJ12R8chkKGX2vwk
ZNUtilpnNilajjtTpfAjbaeDF7H+12O08ktiI4rZWg1iP93PQFEYfK9CYlybaDeMm5D052FXsVhV
3GnkowCJMWU3SIseXzGtvS4q7/k+iCZ2DxOddvg8C+rjscUi1aTrKvVyGBp0XzCfQYTfEyS9p/q6
eMHGDjHMYPB9uYnVS5QUFOktstdYZD1g4NNUfIN8+IliP1F24wn+x8dKdpztYB06X/5WjfNo23xi
8UuFyQD6HoB21AM61IkvzA10f7hxP3UYFrKbKI+iEw6w7PKEEwoubi3BM0+BB2hfghYxm56yKcQ6
ENZvGtxGJ4vZn14ThcZ9ISw4hJ4EA2xSfCejOCi6z/hEHYCS1Kmx3Yqw7S5+GV1CbIyZeaFu387R
jf8Lz8ju0TcL8rN+YXGfTtnqdWR+jJgWhSoDUaUigbxMMZbmS7mgzA2bNpT0eGSggJcSSt5b9MQT
SItHhNd0q8zkC+nsh4hHzImg4jEIPnOehrDH+PqpPIogjty2R8Ze9hbrPptvLa9V0LtV3GHPGL7L
IpX67AGIc8+M4af1zs37y6ZrUUf6zxu5iwgHJ24Ed7zMUUMijZgn6NC8krfuBAT8Uv4muFmFDZYr
5v5BS+S/PJg0Np3HbQdFkdPQGXzfhPoB4fFd1VScRayKBL6e5F+BnfbdTmDtjLXuAoID2i0BcpFM
dCzQbv2FLJ0ztgGYvNzfBwj6sasQjzahBCCmEOAnHRWny2WCbBf1eYFPVOpt9MUV35jJiSUmmlYa
qQao7HrYFq7MhiItfuE6iyJiWWrm4wbiaJumHh4ht1/HcnY3iWp7vRtc9x+bIosRSILJ0rY+EOqE
nRdidkcBQa2X2ejVjb1vtiowSHC2TgnR/bA3F2t1UAZwTwEihk7lErljFvg9KK32EBbKYNZa1+ps
cvL0u9XGYM5SLFEAVNSk+ehDtilJTOkk0aak+kFnjWZQxgBuF9nVxFk/Qr63XecxZp+JIMlfY0jn
AZghoeA4TbgIRMlQdET2oTXTaEDqm0yixdV0/Rv+vA9XmIflkvIhhBfknuL3vjeK67KL7RyI3CAm
qlUJYoUqhyb4mxEcmHnJ3t48pTCqZY6TkNMLzB7UBOMJQ6n1DBVSIFanNQntYX7HCNmXf0QLA0jr
4taH2ASLhNb7NGVR8xNggM06nFys0h3yngyCLQKWsCYQRkukWyYHC+zx5XAMCVG1/e7zvbX1U7MI
pU0pvrqQ8MLBpvyXVFo9Io37JWN/u6Jh6xEqMvDS6Gd212cmpE5nqWWz/GpAGaSZgIodtTbvevxw
aHUpm+xZ9BOsjFHXsNt2Np94ARQgYJNF3G5rRRhlRCZslyEwqOJl77kizaUZ/+S7g7ZIi5XDQFFI
rtzJlVUryppVcBKa0QY7IhakLdSiJyqUsHwp9Pt+q2NQk3tOOg8rFSKj/2pb3CArnsSgNl/acyvG
Ztvq/6J/nNceIl+Z210rfCLUDrPLJDv7DYyiLhyCaorPpbcC9hTexAbpRXznX3WKtTh4p43QruEy
FFdZ8welGvBJIq0v2sxciHaiIEgmpHPocm+Kt9cxjyBXVaQmjRJ8b0mQpsikfegxiuK+vS9nMIUV
Xt6U/qRxi95lLHyfeieTu78gVupyy+lIP9+/BP983bME2IhDWOyr9UN0VsRks0HAnaum1xs6gY+N
SdBs8WzO14VzMtVor2yscGRHDw7Ni8cW01rmzT59ViofMv4ex07tbubS3oV0IQkhEhUDoV/mrTcF
hsZOpMBAVWAIKQIWrbMnboKoSx9Yi4+FIN0h54s9gUwqzcR6J5dgQ46TKfIZLP7w+oOz5i5++Dt6
dNYarH4sS7Uypsn2N5xB+sLiZgUXYb78o+0zZY0Zgc1tZ0pbWNEa+qOihp9ev5+Bf6iB3PjnWwW6
Qdowzrg5sjn8ao5qgKMGZgn6/if9pw2OOcAVs81J9suRpcMaUNpzoLBWb2XEUn57Lju9ZfDrgfMg
HyxAGksVoj5m2u8xp+rHdgnwIGdIlkgRp7FeySpKe02IHeFa2Q6r8FytK9+Gc/aWU0m5Ti97f3d8
5y9cnveXZ35voVyvgtW2nAWAMFAb0j1iQWgMvB3jEgisOCVRHbEWfLF/Q60+zOdIzQuCwAhi2nAd
kM2yqmhF0IvuT3/Bwe0eNT2J2Ngc1eJlaV3o2+Nsa4lqPkoW5jDjmVjw51qtScm2YuWiduMzXZzg
4W95qnfRBIJiWQhkH/aDbDZeFLEdXjm5QkCq2a5gAUX+tnFxQNfcDt+DYpqfelz3Tpqtm/ZCsR+P
U8+5/FG34xQaa/aoD7Ucp51m9M69WS2PYz+0psjv/52GlZhEjQXxox+08nvF2uSSLZNXcELoXMs6
S2UlK3aPvEiwif/2ol0oIEt7I+eTj19dBWGYei7QKg64gkuk+UbaN1EL423GmVUxj7kjU3EC3jCp
F/1iJn/tjsQsdSVDAXvtpH2zRaC93BhlQWm386mjArFpT9WcTC0ujqwX7+IPKiLbRK7JJmlYKdt2
P6H1M3sckZtNfTOwLqTSLyZuTZJCpGtFfJTaX5Tq39SDZmdFlZ92bHnDUbIOKzyDrbZJAl1ILkU3
g72oKOtpr0DCGl3qRI6JrkciinpqT6D3hqUTNiW8LWqIYA4QXJTmPPxK77qE2GA3yDeCJubMiE0a
IrJNBSxWtMlW61Opwi6uBBytwlFLNgMvDL3tOhDDOUWJc+vuQnRFW3BtWXcfbBSTf2kymOh0IWmH
17tF8btdo4lRgN0P9Ku1j7GslxOYTPY0Nfb4iY1XF5k1FwccBhgDwGwQGMQNUr9BAa0KR4W5TH7Q
8Z6JPeYBzQDT48wCj/lp+LtumYBVEn4wzn03BQjivO1ykrxdNYzmgDDApS0h3i3eOgGmTtp90oK3
1+UQd5b0THFxlGqqAlh2R3nV6vtat/i24IL7g6cgayAyWroQeS1wTV3YmLjtfcI2vP4FDCIYQNAw
DVPhJXL1va/SBBlWByASLIWkDfPEyc7eyXgl4FD7xblxsYXise0lPElyVkGqNthsUTncycCH7vOX
L/YGzjrz4GVqmPSThHQVAvUBCyP8yTPv/RCmH7NKTV9aQdsNN6DHTH4QxJydM2BUCgHCKwuqaeUt
YezUFVPrZQ4x5Gp+UjRe+vMIFhfc/1clpESR4i2Nl2KAUJfRgXwoMfoceeQvZjq1OuS3JXak+rmv
MntybIievx/408zr61jLCVgTRjUftvdrtBsugI6iKo2HA8i5MFtCaQriRNSLGjZASlzmHWwpSJps
kiYhSqzzvpEeGlNT6ZzZ6mYLUJ68NKkQF7tB4Mrdn/uK9rCQQG9aFtXWmwsOQPkH3t2brlOZ1Njx
/LVE/AegF+XQreEvYAP7z8zBil6ehDbWdyQKjdR3hwmvIBk8Ir6EE73ynfEnzSSUC+353JfKSykJ
7EylCnt27hZwbDAtwL2n4QtCGqfLlDBdLl74M1IG+FdgFWNvsELtKGfO1b0KQUYAiPvC8644padW
WPpgXPpf4Ojk3ETOWs/IGLlLNW2uVbCYUIxm5Qm2lT4RpeLtOXz6Gj6I/2XMg7GUy94fiqmqHL8J
hDJBtar1kemb6XsSwKyk+VRxdadNvhQ1bN2TxikvS645EviaIea0Gf4s/PotpxbgphqDEVbAdigS
VMPYi0PBme2YXcEKHtttLrDwnlpahDBVOl2t/rVNdoeWfjgwlXSQ6mnCTb+LKu3ngifrG8omSpls
Uj1X8gmaOFRkRMQ2zVjG9N0ncqWVwcuMI2FJIRyPX1k9ar7KSNRmkp6rM/oTrGgZvmqIj86t/JJr
I7nY8scIYTqgOQ600Qbj9me716ZZ4H4r2SuqTtW0ddP7ycx1zk3zhHYNKgmhGoIQOLkSTGptBsoH
11ZC8QMOx0sb/EBbZEv6pecxX0iFlh9YAV4KsPnaW+qoUmWWx3KmWs25igknw1knxHq6T+udX5qc
0wHOV9qYdQkSRAhoGqdmcS5Ux47zHkXdHrJmYo9C1RRhapa2DKpqW/xexci9xgsq67NtUWEjjivB
bTVdh08rjetG5ns+Njrp+w+VeWD2vTP7j1K8g5DXNAPmHnl7/RepdL+e4zbChYooEzoN+oui0hup
QPrEsk9jzyUyp19plc6ZPLVwRZTHVftcJIDo/Kp75blip8XVe4iH1vh7+g+DCgJY2J8i97+txkWY
rK8Te/c1LCJaLhFAeKpQcLysXTGKRjtEAowAIKqemMU1H3b2FjjY1kQYGcv47TbbZvGXDooQ3Hfd
5d9IHMQ+9LHqrhuG32I9uIN8Tn4//lqJJh6kcg2QCAOudQcZ1hli9KsDDcD22KTwyCq3t8QSRPrq
WXgcSSAG5ww7tXLxMyGbV7Y+t4xkyHgX7qpVNLTNTcr80q4QelzVWJ1TesVrPeoF6ftwB5TCyfyw
Z/cVCnjFA1lfj4/IZR9MKY+apZcUvenwR8F1/qR9hcjxWxjejbkAXIPAlR10ToyFG7HlyhadJDwj
FmME2GxjsS/GlJN4UONUA0OHPgfT++qNENdGq/Er5Xoj/DpIUu9kw7VDNzUeQVNSLtIKawsTGO9/
cymX9+RmwBZyyNB2OjxFy7YxmHggb4W6Z7W2wxe41sBBbriyd1sTWNuzp9RjnYlTYw5RfpBrfjrL
lG7JQiCP30aPatWZ9jOQdaFDQMohFIh0keLwtWPeRNut8KVTk0N1VNMdS1MvnxaUuu9j4BtFThWN
S8jQvjnJtVAdV7/rHDWVK/aHHcRn6/KBnVpcp+mF4sZc/LzDRb7JyQoEhTWFdWButqAc95i9Qpyh
U/+VjWWvXaWCHjE58GOYJPWG0doqIu7B9ARjMtNnq0PKYLx4DAKq80X4tKYPobyazfKJ9PnkPRMz
s5HqwUH4Ltr6Wif5L4JgWj0Q3/T/+zFYsYVKL4K6Eb30FaIjN6nUmj2G0OnomPloUrwuLog+Rr3f
HbA3/hJwYlrLosnLUZliMDKJPt7IgjTLrbq70XHP9lttCPzcliSqfEFWgF5l7V6hqvMlY+AOLivB
JSVau0fbfDfuY3RlshjZyzgQMTFMKJjK74XlWiCzvF7MUqXdSvPk5ayTd+d8lm1H/MmS0ZyQzZ6H
ficAmaW9O2dPaAQ/ezAOqOM2/dXsfhWANVSNFCx40p/bFmvGCMUPNTXfU38G7NXffXUOMROK4Ls/
0eMnGpqL73xlU/0PxIn2p4L+tUIRgmg3DjKkxumkaHukEUiYtxwZpjYxZGr/m15Gjx9Zqg20hBID
MtxMhMn5BhRijCccsBWPmrX2ni/DTBIMn4OtoeAG0n2xf7GwO3uh15AWvrczhS9Sw/l3sqirl3k/
y9jzn7f1SEK6Jj1w/FKWdCdmZMABvWDiUwfR2Alok4+AYNc31qyHNFnfN59SHiOJCE8iZ4kI5UGR
xN7RoUMsht5bmOtr04U6w/IyFPPiNgIq6BK4LiV0dKYemFNuS0dGUPSSh08tUQ1TYsIN4tgdZLA2
aZkSWiWf9G/Mkdwto/25cfyan/Im7rFmBYmrBExlCXqJKrugP/MItqX7kH8kkcX6p2NmNoSlu030
HhjZPNmRLlZkmAhi028rVhIo1DT4+KgBVdStmNvL/A8Bd9rNJHWlV8BUW1RbvPKB5IJl2FDkWt+9
ztW2KEyjc3dn3oXOOKfOeMgSCDFxW+KQDamlcv7z7t/oCc18A1jBA5RTuq9mtwRsIM/q8c+3LDIc
d800H5ySZFgnNuwOiYP2C87JlYE57deTRniEgcTuuPxuotKrUjk8HuwW87e2h57H5/kSqi+ZYy/w
BWG9AMd20DtWRUUIvymv4i/cMct1IrpLCM5bl0mjl/EZ/6DML8Wyl+ZqV2jgGPxzDXDRywmbUrko
LMMNI7pjm2FmCy3GD6MLIye8B+3h7gVDzbKcYxMkufHOZJUJzwwro2BRVUTdUsCwk3NqI9QY38cX
lYpNvcrp+vpulTrr7Zmi/rkVGFjQrQ+/RHWcBtPbUE1+7yjNMlnStW9BHWmjOxnMEI16hGYnbe52
j1O6xfp1+BCNVjFNVmX1N/2Eu2cS0fvntGAXi4QBbxOtMhpNSzcF6aPxTGexU3UZIY6SFB9M2rdi
YHD3jKcsMCExvPvmrVsQsEnZtSE/CjgcwyfdGQM16NSPhuyox1vQ3DYqv0dpP5d+pDplW0qyofNr
ECk8tqLDOPJSghCBlSZvD1sjofTHBGQfFpktPFZtzDGBxmW7HVl5rwOCJEA2awlpus3rHmu3ATlG
wHmRpgCpdAAIdACgaWGyIKRdjUrYy+/V5ryeXWUBo4J7KnQIX30s8LZpmlxkwyUWfbuVxUiiC7Us
5PH4b46s88i02jrmnhVQnOSZKbvN0ls3JUjCHckiTLzyCFLf8srFAzAzD30zlJKZzAhEkR4fWF++
8DEYKWmH3T8aSghgovNb0HBFHWrNaVO4VW7iUgjBBUnHBoi1cVEkI/lCF7LKhg8EOIfjKQB9+gL0
Z8Q3RuKHTTn3ZiRC+IGkSZn7n7uyIjyLQZ9pgwpJVv7rW9NUaZmi6WtCbrvi/hSmBYRd/S63AfHH
5t+m9qKXcXtKkURSjj3t8gL9QBZBbeuR9HyOGUbcys5k4378gSa9mHMpYOvpksvbTqClnFnl/kVI
eRnFYyDEWvFI0ZkxFk7un2L+MX6ZgE7BiO/lJF4CIT/SNFG0u/X/150v1ess/lUKic7w+5ruU6H4
FpTdCZBc02ye95HegDDQpfJZOBoRRi9cdwqGgy9e51y8jBab6LHqAPgNMrU9Xu9S1MmxyqB9Uz2U
pQniKovK2brsT3DAq5Coj2UBWWh5KDuZsLu1q12r51VRzQMuQzzqPrMz1iqNVYhh7kBHiu+1UYoS
HTPbksbL8bRo0KUhJliSrgc84jJn7ZBhpKH3IHSrEuh7gssQbPapPAVMQ0WmyE/F7L5fru2WyFX/
BShaAsQzYQkTgZPcb1dZdL+Fs7MxjkYoA2WaEXhuOJZ8qqs/A0UqEpZx+4ASr4CP7x9bIOfrUs+P
mFxcvfz3BU3SujnHaD8x9/uB/90MxoBDuZ8SXEekLfLjbX93xsRu0WRhVxrIam1TfIkBN0ievCTT
jKoENdzJEiqLfvgAvKB8bPuGa6WDN8NMbZdWSfNnTLDjmceJ57BXYXAI7bTyfNekMv5cyo4Nd5Vq
uypyF7eSvue4LxsaSEyQ/fajfKNovtFYoFowoEDSV7OAfDGLFKTe8+ryEHXKkjqXyRHOPwMh1MQL
EWbwggynA9+2mBjHa9ZgB9Q8uKejNFD2xhkwwFZUJam4h1FVZmKNxN5oLs/o2gMFbdOb4ZHPsHaS
4lCQheeYf8o6WyrEXsBU11O31RZ2h+Ge1/h2Le7d/6KZynSsiSx81QGxDUc2bh/vCtaqCtmPNw8L
67zFYuMmat9sPxfd43YqISqOtbK3nlS+UmY9cz+ymFHo7xo9yYuj6nz3K58BknAUu/qNp+yPJ3oJ
Oxx6w2sVEVnrdB9Uv64QSti9SeiDp2tqWlie7FuRs8K2yMvOSqLla5FfuMvmLZB7kq0+pbWF3PRJ
wWt7eEOjWp/xigf5v8boWTho7cRYWPjfDXWHxdf0Jd7lJwpX58/QFi9+1eXwY1QqD2lMhM+0srwQ
r6Eweh8dmfaJLzll/+m2r45eIu7G49NLa0PTWW25XXZ0l3PD82d2hyOqhLrRl44n+LmVDkXKf9qq
ARKjGijmnQm7p8iJjfJ1E5YwRPHepcGTNL4coMrBhobYOy3Kwu26DpZDay6bjMbbPOquo9NqBws8
fDL3wJ8P5KlmPkQEeGr1o6v88vFdoEZtxZ/hnL//GVzpT7toERX2vBDVbF3n9emMWBQJh4Zt2EJp
l/dsLoiCr4WVVQ/7rq7kuA6CR0l0wgzUjF7H2SeShIdbpfI+miEoLUCjWHYSAKaESZlPu3T3aVD3
br1cApIn9IAeu9EEFQo8rJemAnJdzYca5WymZta1JjDwMu7aVa2g4vujiie/cigy2XYc3quyCXSO
f8MV5qDHnEmKJ24sdy5hIzEDv5JEgBrO7TLbYoZGWTQZpp5PFfVub9LeW2bUJyD+pdUwZbRdx5JU
SUQbNmRqVBeND6ZnS8qmTYP7NmOrYMak55AJtIZTBd25OSAQZEnQvzIeHz7RkoWqu8PCrWVMxLZV
V114wYypAgeT0AHAXc5dPLsx8x/83sUMZRhDJOZDEZiG4FlnCuLkyw9HyOI4ah1lgiwD10aaleQo
EqeQ+vTRXXnktCFYftbLHFUR+FqfK6V025I4dUEIQAHSY/Nvf4F+gSywzNNbQ5Tvu+1V8dwQ9T5/
e4B0YXXrveR0qYO3Wz/i98/nX7PY84Z5XRix/kuY+ySdiDccmiJN7mHHJeQ/eQNGEfnEA76ec8gE
7M9BpmAKAV/VNA/n2P8IYHuun7FVJacc1yl0h/PknRlyzuVYywQA3sb4pD0gF+cBaTvcY18jobfg
TzOgH3Thtth0aaP5CXsX1NBqOMKqPxkujSO5tkp4Y6daEnGtL59Uc5mbyrxIagnu/MW8WWb/K6TO
Kc/4kOCEI2YcGpaf41Ru7LuJSSfF0/FKM7ECbpI3aBaachDN0ys9XPAFydCaPRVzPel+2k7pRHc4
GS7gDiHba7OcnaJZ6eaUPykbHwIwxyopKo9y7nCADszve4qBgTRAovoLX/gzwyqUNNzDzFw18HLj
CaTUy4B+KPFUyP6OWe59rCdu0TwZJByK0GSTy6LJyKhCaqkdoDhVkrbWraFhKNTNcm33YFUBc8kA
qgXsdyjddOxpIcUipJOCyzXz/Kba4tgGQ56rNedfgZDIx2A/V1LiSF2srV+l1FDpciUrW2qlCAFc
mNaKmlS2hXcLPP3Ki+m/LSijAo9nqUEFfmsj3APhJI/0nWQ39slsKI+sQQzWsPY87d37dSZkWV+G
JMotLapcgW8veF8oTcdQ86UfLq9V3IT0EMOTjVTK3MQJAQQy2fVK14qHD5FGHCviY/gBtDmS4wWP
5r2NL4zwxPEcOjdZzk3oN+MOBCdxh8jo9CP4H2wjzHnXkWLLUG+1cuZP+Xdsqcv9MqoPox1qwer7
2wHt5SNk1miqegsdArAMFHatkvBp5exF/9vEdoE6prkj3fI05q+kNEK5reAiYWxcxDigWY3miilm
o9yZaJdAF0p2uU2AKMYRPOPvEN80EHBIMB6AX6PaLhH98xYWd7+YhjZhZuiYXTHhRnTihACLMSYF
DEki8WOed4AemhrKOxXo0PCw1YJ+DjOtwGuq/N7GbW9u5OGGZ4U0dgc7VcN5kGOxiNjSYgRgJMif
TN0PjU5n0i1tTI0P5rYTsrVX8CrX363MiLIDyMh000WGRkr1xRjK2A6V8EZGXl9L78NE3q+7U8rU
uKv32S//HTvddiw6zFCYslg/VGeS4gp618rZRturbuclbHSyrPj454xisMbV2JpMf6O85mlWFY27
SpGPawXCXpbagpjDPJ1xpxTzfgdiMRDKxFTVukb3bACkFrT7hL4f+0ic0q4dRaAxWKZIJpT1KTTc
//VHJNLCwCYVx4HoUZsQaYyGo0xd/xFag5CrD1OD8eBSKGY+UxuwXfhb/nxVv8aOSrzAtnLL9ose
D6SVHwaeSaVif2eYKXHblv0ppa5n4avOpLQPxRODRQhEwl1urTxoSA0ebzbUxrfhgSfflAaFG2G4
H4AaOTL5Tm+E2p4BWTGu6gSi9oU1xqey+gRWkfbG17LzDy2kfRRYewQ+Bi9VCAz0PkEC4VJB8+r1
fBnxM4YEZ8llcRzqoEHMQXkpiF0wguaN480QgaRDgrsuezoJadcmfQmjz8wmjFczI7tXhGtHaZMR
F9s9CyxonQR3/8FyaHkwAtEppT3bWiNMu5vHRZLNSEdq8tf9F/RbsONbq54Q1r4ElnVkpl4hMVla
1ASIEGyAVyfbruuy9Gb3k4ZSxaf2xdA5CabKRT5fGYD6Y6GOLIgsNgHajLsU5vIOqxDUIPg67OF9
T7gxClf1/R6oEysqEYuoYyOlZ4xZmhX8khYN72nXGdOw4vZ6qCgIyuQN9CmXBWrlFKNirurozDRE
jCzydwDKLRXecqQCIT1kF2VTtfAV1NA2O40yl9255N8OPEwCoFFy7/IZM6nTnrVPsJGhaBAxZ3oY
WPO0jtJU/6MPBtQ1brOkFn8ZgI2dIhcb9Uj1r7q2spiRCR6icJDQSVs8dJzR6QL2UcZh7GWE8Tsm
mtQi0oaaWnjBk8OITwvHuiLE5s6Z7PhX+y9jWDr0lHueT9UjqicR0VLIlFilcG6uSoiVI5osjo0O
APkLNaFyskF/s5yWtxLqWEUfpPhnjC3dGK1T8+hgLoJmOyUylKu79MznfT3ZzoxE+jn3JnYRWLEw
SFlmysR4BRO7eJkG+ic1AykKLDFN8vEA1Bozby74yoJFRdMV7TC1aU31gv3Gn04Zw7diY0C+VQ80
u2IKBW/91ZvPIw4xkg9Q5vNoO3uIInqsh/mQbialLteOmo87ZK67sEeVN8BXuSP24rORNbLLZO/T
ElS6jNCSosKSxFq6fm+p1wha53oQSLtoXp5X9UGtoDHxkUF9M3dWYxL0CrKmrPjgx8U0omJLak9m
QlE6Ge5asX+Sy4UHZUjsmsUkQIDbFu5h3VKHs+2IlpIVX3wyRLLBOdzJsnTCcMBJDiM6KdP33hZz
LH60vB7ocBZJIOXYI3iqvE1YtCDsoI2vJqQhp7iu/Bp5LT+88RHlUYdfYwfARKi/aS8mPZMbPKGZ
V9pPjsP5IHGuJSTHOhRfo0pZSf8cc6TqJRsD9+Bas568LUqXAuCqmDtNqZEx3jYzGIQZ8gq4FdKJ
MnwHqvNSnfbXzHYYwAC+cmlvDeaZZQi9nY4tZ2EOEdi+ei1ocQSq9UHj/43qb+rCIQCaAuX5Xm66
XUvB1i/BCfzmOzSOS9QhFULKiuq6YpjEgc9K1RGz1DzntP4lxYwvbdQc1in2zfaKiUwZO/WAztux
EAAQUpUrspDikDUWzIzP94pClbR9Hjb1soxgOh4dlRx9oC69l8abcNiKL8b02ywzEovLKwQZq+ob
jpZBxu2W28pGiQrHJ865MAWlekW0bErNkIENmPuwiv2ol9ZjFGRmo+4J+y9Q0ybe4as2GzLozlVP
3RSK437GDAB4wJ3OqK3GOcU2RV2pvacsLaoLBQwsXVpFbq9xfa8SZ0zMhgiMWOtsvS71Hq5YhsoT
iIrFixp45VJik71LZg+nYm9zvConhFgo1aseySKM99rPF9oVsl7jzu47q3Hd9Q8TTHfcaz2kWmRB
rzwxfGcKyXq602civMqLHQzFiuQq1S2gFDrkHBpxW97fSKbw1CjWQ0HcjDn5BEetE50DY6YYoF0S
0R+7Jfi0qV2jis+ujolSl0itgC7hcCyfWDb64aM5DaTL2JDFl/TgpmHoaM+LwluKw3+I5FggsJkA
jJJ9FQIqMxjnvvVcTebm0ukLweqJkei8vzn+NGmGAfEjVm0wYy6gfSdRuyGZa4DinbJ1FjE6BAyo
yi9CwW1v9bgA0oHq2ehQlZGoxF3/fMNduLOPTCqigf12K+jbPzWCke+J8fkUB4Vlo1ge216Ebdnr
59PDoZVsgDet5CE6Fm7MPhAIs15+r+FNBNcVSfl/9zQJAFwvIrOKLHjRzYHX1I+bYiJxIHGHi2bQ
BYzZmJOVxoPhCN/Q4DP2JgJASfO9C5CNRyyizRyc8zfdRfXZMi3LfoAxAvTbc4nZ6zY12nqpG7oa
TX2+l14s3VYyHRcq7edomzcrM2beGvnw8UP+uCZRYy0nylugn1rfV3IfSXkeHgLbRgd8GjW1jrOV
IS4HrQ29l806wvBri8TsJKsZUbZ8T+roBMv0w/iURysqOpC+jvMhSxG5X4U0XGXZNv2WUJTCMDCo
ARFd7a9X2pTz41pMvETgGGWAdHMmvHoE6XcyJQ3AxqIKGW9QQScAXIIPwCnICIW1xxe7kezYrwYE
UjTfmytEYAhWyVkF2+QeWnIXYnGvRHPLo5pFsZDzBPl/lOLmJwOuyQzYwS3Ln/cc6lfAmWVA0gPz
Y7Kzce/4oqSQDGcbX0mrxe+nc0YQNLhRP709d4Z6MH43xEoMUE4guaXWdstIAJPqG74PdbQzTNd0
2T+gtdxqFv6IROX1EPZtP5BFDDT3jbvgP19jbfq5ZzUDDfhAf2pLBMtZcogef7vftGNIIiBuAIwe
cmV8/tZE9qs5XGvZrxZlypoWAUxG5dI4yibjqYmSKeZCObJC4QxNZMrZFt5rUTqE1g9j+gHsZJsk
1QTAdmw8WnFcnWEl9nWBZglPDyJGLJI1S1kbF1XB4PL42xmRT6o+J8FlxvgY66FY7PQ6RwMimrV1
KMSHEdUBDG6UEGRnDKzXU6agDgBTtOOCwUNqFlup+Asl40IKsfAu4RStUYymuJt/RH9mZXH/E98m
486iElW47TZd11zUpisbDgcf9Ziw9k2S5aRnd2y9NhiTDn574sujkxMqpzDtkXBI1iHLK2PLKm0R
opDqOtcZix+ktj5C2S2nGo8fel7BZIyFVPs1k8ERjMoOpj+GdSCXf7XzO+QM109SLF4tWXKqxgDm
ZqkCCbolhahV0mfYJR/cw5rKUe5DkH5jXSnhEzVwtgBjM6F53SRnbyPpTQo2bUsunAiN+PQS6+Vg
Vhb0C6MYuq/ScBRMb6SuxmwNgvEZcKCdrVmyundP2YXX0n46Ul3Oa2NDli0wDy+D+mrJprAjbeDZ
rjPHzaeUcdq+Me5SZnei0ToE8cb1lQBeft0sYhhQjcFybeRh0ZAFEug0p3fXhqPuBSFwt/WhOkz1
9SMAu1bquITns49pndcNfWMo7BVyXsW1w8ZOt80C6VUj+SjAsNZ1ZqRdzZhL6Zt0bYcH4Fekb3Tl
ZcDMF68hnN3B6P/M90dj1Rr4vvqnJT5q9F9ViL2onNZtOvd2HqrUfz+mZYawLS1JnuDP00WTO1fS
YAW0fYLkajouQCpJKMFXOUFhtFVWiuG71zcYljhzjCIBY/0tpfjEAlI7lZPH176lipv3JoDyycRn
KVoW4Vha2HxXF3UZvCbmdmxVh+YGijPBNMr5opmgSG/XmOnrpSXK8CnDDOsEv4D/XgxJCNmlShYE
K81GB/xOTb9siCK3W6OPNZi81u6JRe6U4QR1x/MBRGL3RMY9nnCpun9TYVsAY/gXNeOgoKJFSrwH
EPYckiqS+RzWZELy5AI0wph3xoNjpzargM/WYXzsjEEWr4R9WioNYFQDfYYTgdfvGlThtyU+EYGs
cocqb5/5B+vVgKc4/ZN71hO5BebNohnqU1r0Yi4eiM3LQxxRNNgTo48J4esk64Z5ksy+PTTw+GYQ
6chQ8c1T4hDCuMik+9ae5h7Gmjw11LYEJhbTKu4ChweJucpRlaO94XgqfZzZCh/HEfvJ0GzTc20R
tMEHq+6hx+cNNuOgim7diO9h6iOF7G6bEOguqWoRfobpEOj/cdAc6RVsm2/kxNUMJyaHe6zTJ7jZ
DzF+nOzbBAYT0CTkcmX/ef0wqstGCHBv2rIKAfBe8J1J3FIeeDlDKIdlVyBYJJO1uIUVypDZkqIC
JPJGLnOk3cuLGPwgPkH/QW/JzxLTF9xCMDq9iqevvMAz+MxQUAO8emseqWqDgAyH251sTW8z9a6+
EaY8ugWG39roaCnpELVqwny/hthWU6DQK42AAtOafILNuYAfiZbNDxGzQbrmc2h1KQvLQnVfi92R
Z6kVGWwXdXgqrMhSO3QdLpC2q8lUa1JvSMn4M1Qs7np0y9VnyoNCkMWNCcy8kscYKJFd2hnlNDqr
uUv5WwhsDzrVwR+1p+T606fOw/68E0IVtQOS2UJ8N20wEBwh6D6tbmMJgXr11qL6pjST4Af4CEcY
RUQd/pO3XVk5zwpiAnSOgqKss9a+nULt9oXkEjn9+XRKBTL1X5ujgytwZOQIIHiCCS34/e3OuA6i
7JJy5JZJ8RdthcOUoZjCNApIEFHQzFFucVSbJgRpPhkj6meuOX8PgXXug4pY37C0AH1VTxSsHWBB
mfBpUXs/hsuTMS7ihi+uAaODplje7pN9yIT0dOVkwha3G760Sv7PQo2wdJd4Mme71L4MJJhSpVyC
TR0UUCwOTAXo28JRADVrEnZNmllgDIDjxvsaEolVtfJoMrgzniCxja9B9tiN6UIKvIfkFx4miqcT
W88kP3qPuUsOO4hyS5Yxc/H6Xyrc6k3w+QKTGxYwFndCAIYfmsznjbTMdIw4tSs7y0dEl6VZhHEv
sa3zUwzGNBXdcsw5EHRbZf6ciCYIAuXEbCZsV563cWsWx0r9SLatDOgXvbW+nhfUWINIWmEPxRYH
ilNoeE0aB9YKYwRNmLSGJf8O0E+L8Bms4dKfZUlqnOakmXEoOVlAxIwKz+3UQtyRdaVj42uBzhh6
4LhYbtmu/Sraq9Oy1hKzwowf7AEbQ9McfKY83/stTeOwq8hvNEsLh2Y4UG6zJ4tN06bpDlTklMlr
ZqKsKTMGNKaz+HM5toRptWpgnXJ5vNLGIIkxBZyA4/67pyg94FE5qlO2+J1e9tji0xKwmRzTSauk
7qKl2ejyYqOl/3IcPTKUysv8CCShfvrjRPVjCBYCJaqWXvymZ2OCihuI1K5ObkI4acJbZRqo7gqR
tJOM9lYOiEoJ07qOFvVnVLLFvzxo8m7O2SnK5Q2gET6aV66n2NOfu22cPQ4CHs7+dkPruYPsUKLF
2pusDxGxEAgOydMlCAUfY6J1M3afbIyEqJAzPDaqDukzTtMxTYjRq+Q/rnOypp5MKD3GUBnaySyB
Ogb84oeZyH+c8gWAHPXlVZuDhV43ob1wWRBkAh3/zNWmTVQ0czYg0MbE+qhNINAbCkEDSp5Xo58E
PuulVmXkGPhC3Kwbf8mRNaYz9sQ5uXqWOBwvrp7nfK4x5oL8OJpk8qdZd4vZ7ltvo9kN3etiB9DJ
QVtn6nplQJ7kjHFLSR4uMfrRW6PsmgWUiy3P/YeHbEil3X56rqNW/EuTol/zySZOWfCKclQL5yg+
kI4AEz9/F8oS/UX2vYCG2pcW/L7BSS+HYIecrkhUuuVjqlS4CAuQHT6kcFJ/q8JSrd0nzHSH+XyB
HWhNlnSw2Winac0YlL8PTHPraZ+otYnWPTq4jF+UDpXZV79u2FTxxR/wTOQvcCYYBdiQZvE3bONg
ujr6uuyxwdpeyIwnRc7MI/PfFJyg5fX+Rhw5UjNOUKFCYsf28injromytgNH75mr88gCM7UzTnOo
k2uCBlKC63czf/UEIPy7G/OKhsHTBEBXeBosk3qU7RBpBS257g93NQq2yykrBDgg9THcy5chiZpi
QrqzWPh08ta91FgtNYMoxi0xlKgv+H+v1JVKUYWe4EfudBA+NHsL4y3irg9jfmm1vBxbO+Yk6OWg
ijilpaf1sGYYAlCXi+nQ/zhsvMZA646Ipmq8gJJSGsTDbmGCAGTuDuM5mUZX0na2fbGzLakCpf7W
Vq+Vg1/1ECZUg9gap06ANSZigVTlCfMpECC3XF6ivzBEMLifsE6tdpaG5ERXCJ/TMJge0fqb0c0E
VmeqdH1H+c3ij1BVMpbRiXchL5wxfLaN561M8w+YJDt+y2i/XP6lh8JkDTnfo1RPfo6jXYxttUKr
behplDl4nRADrFrBHQFlGQvaVL7rzY4JDN+FAx23ES9veLEtfVuWUJXqizaU6VY3J1y8OVvLSCWG
vIm4f6mgd+iLIMWsgdD5E1iN92WXJMwvAt98moPyxuyOBKcR6AY1Z6BPHXQ8T+enwXWl6bWx/6xq
4rEJIArahMm0hnj62UFIilM2arffIZmwKwNvLeDHcvACohO8SyLDHx7Yki7oc3tqz4k6rJaObHg+
dj7u3mLlR2BZFjsCUy9PLrGQHGpkRnCklpn+GMXtMgDNIlG3tuPMTSfBXVz6/d5Bhiv576nK1U9u
bz9Ri/B6Z+EDV3Vyt/0+6GBgVfVDHlPXj8VwOL/g4+BltxSMxaCvxaMyrniC1Fh5R7+Di93me3m9
zMZ9JStxqM6NY5rCmJBTfHdDjK7RM0PreI0QRm1pRyKBG9TCDqVMs0eIuV4E34cQXJTcr/3u8uL3
IWXaCpyffIxPg72dg71YnLiCMXpGOoFxoc/W4rOHhIejhU9Jq7cs8nI8/WWuUWMBd2lgtH/3MaWE
HWeHPcv3x4O6MS7X7ou7m9r9bLi/mAorEZyyEMwMdMejKqu9BjBZt9vsC3rhDc2shxaMZg8MHUMg
CpDa/1h06HjtQY5ZZbieLCbZma+8ZT9uUycbkBw4SGNCkj27qFrMecwaDrm/yLv1UUvvZrLDQ+EM
RT+r7XHqM+eTJo1+nAOKBN8rJ9+Vu/YmmpRLQWvvsbjDDTg+h1y/JXHSMvmqVuQsW6sgjQERozlM
epHczuxzw53xPoVPYYPGxlAJ0ekH7CIkaQo409zRuKhnOHsOke5eAb5k4lhVb3bGPtBWk1P4pgdw
iQFhl7B0WUApCu6n6vJ33WNYqXbmm8QzJpyTDEcZYK6EE7szKCX+RwLOk2X8i8gdDKlW3hILRyNE
qluI741/CjcsBCOcux5wxF02qYcK2dw9COUvCbDPJYIHAFjA3lxUOvrB6+tkb0J5g4vd8HAWYRS6
nUNMhsX+yr3nTGoMBkvueRR7Sbd2H8nsNMRJxFfVDlYvHC0IS4osMGI8oI6pkV+ps6yUxOsfhl5L
1K0Qp/PE/ZsZZ6aNjaJcRQVGU3qzqhu53Sov0bQXE5DHoQafUgREuky0ymP6XjJC9ZRrTmLUeyKS
c/UQHRAf9WPYjsYjw36XRgLXABdL13CODwmo6mY94VvttM1zgTvlFx6z8goEqAjiu0kQK8YbKgNj
8kVABwJu3PqbQGPA4CP17jKax5msa0pZ+6p3OXVgUNyHcTMQVn+B18L6Qq3jtOxhgyHTKoAaxt8B
eP+Y+rYxvNaEACF5qi6JvvRSdQ3YdYlA8FBYraoFlBvjsQLqEbGXSi4NWIu2bUsrvGJYhLNA5MdI
gMvv2exSEOyEUqgUsM7dWamXVXN5boV6ywvM9TjyNEXJI/XC0Q3zHkp7UeJOqidblM1W1d1Tk8Mb
/mcYfkq+EzK+Xw6jRjHNDjcL0J7EAnxicoQkaZ9LaLzKfZ9Q/ww+089mqa6FjlQ1OL1QDmONxKCS
LfG2JMDX6VwKl4+jh0SckUHODOGjGUlgxrEqVUHLvWfXLky8UtkTEk25XyUGX7mCk/S07DMdopra
mmZMxTc6AbXQA6VohiZixweni7ptZYrTyiRHtft5hMTir8i97FPl/uBaV68P2Hq0jEpJFJrjZMO2
Y6nsubq1ibR672CYm+19Vo+StwvDPOHBhgjeJFF7RMIv6UgDfxX3rWs6OG+HiJyhuQlIluMiMnJx
ZNQ+i7ODe1l7Uaye96DP0WwzubQ2fPnDkBdRrPvw1DJ73QSEtcpaHrJGdBUzfg5MoknMC7fRYqiB
437T3UQ7cwU2mMSAfdvSxqvPBOT+T3pBVB61E6hINUtE8TZarw0nwbilc+zr8Q3h1wE1EJtNIPvN
HCzofR+9HyFnYFa5oyikwXEEBTNb8fYaMav1+t+UyaNOagbsdyFO0AMdzX1+OwlXTXqqLGVsbFRl
OMAaIpxPsffl7S4L+NGfL0hPeSMTipf+G+ZNHvYs+ywU3KDqRLBkVsB2PGMrQQ1+lmv3Ge609U5T
3/nb9s2xJ9RGlOwsUUyg5REDVil8y7uYhog5esAqjn7bzDW98zXekjPrqBjb9BLUtNKPms5TYXKZ
tNhq9AUUMTjleLJicrLRvSN0mdDZl4f7VrWFkeyk1rSZztt/EQvC9TAuTq2g4wX2vqStBuNqFdvS
NZf5gH4PkkGRotFatrn3uCv4xkXwCzht+cQsZCBAMoyfSilwQ0HUmApaiWh0u2VAPHk6FFsw1HsJ
/T6uQSIRhryz/RjfNGxhNdzOW4CZ9ttTdd6y1BFCIzbq6MXmkF3cFAIevoldEgdDb7/HacYQQQeJ
/Asg6rHDfqsq1gsiaLHb10UB/ecUHYmdejec7pclh42ZowmnfYlHYZ1XS2QmjMZ+wWJCZzN5Z64R
WZO1pmnMy0xRgjxW/tKaCsORVtsAp5K32peKZEgfPaKFVtFNTZhMtYy6cq6+OVQQ5V9f0BfTk4vf
yX3MHJCruYaBjMQ8xbuLlXOiS+7qOFhrLrNJByZK/gdVlPm7ccTBnP14+Ccx55M+7cSEWYj7xIG0
wHvWpKvGxgAHYtWzzVi4L0n6R55LE6KF+5O4rG6Gs9fy+Ojl+gnxfO0hE38SmaOvl/xO8Lf9rkoG
miJpzt1SkYwQEnWBHU8ZmQQCPc+5cWXVSTzTmNwHAVAb0V3+YLiPlNS7zj61nm2hKmyTpsjU4uXp
oqJGybhuG1UT13bdIkBCyBhDHU6cFlWbIk1sktSHXQJVZvtIKs0uaCJjLZWYr5yar32NFUXvOPY0
fWflcrL6MnRoU6w3lfIQUmj+1UQJDgLfULoWhJrL8+2EMsiz+9+BNybolear36KmHMTYrINeXWJi
+iCn88uR72jdCixZj9xQFZYQvzZj7RWPaSiL3afcTAVagL0vU5wysBD4zD4HudWzwChRgvzHA172
yGFu1ILSj0kZhx5ztuQWahT3slCyGSnH+zI0fFfaAJ69E8WL7bYuwfdgU3Ijmb3O1MDPSfg0dYWF
myJXWTq4bd4gIarHRibwhQSA6Bvn3yRRuV98mMfqu2ooMGlmjvaW0s1kMVhfxamHebsSiomWoNM2
XUUPG9W7vJf07QYjAxkhJXSGsThwkuEA/2xr6jDtRc9SAhybK74Ocq2iJsxrkb+1mLMQ2K0ISe58
syPJFR2XISurD15z8bDy82Q1xJBuIjASpT9RknYr4hb2/0zCpkPejRQhmD44JgOQtdnZjC90cQKC
Kcxu7qqaqs+xOLighRYoH0Q8kNbTYF8ppibwg+7KYE8amHUur6IRzLNEljubgDyPvKclD7MBAoAl
AGBjBaR/VD6ldlslbP63YSPGWlTH3ESDcbL0scYqMuSfElKrD0Oxc81/ZZordoYomXveiRslo87A
inpkdjbOPlWJre65bxMBU0Y5G/Kzjhe4ycMSLyBgiXhvuaCBNPsvOt3A+DnG2CnzZl6sgAfGzGw9
+11u4Nd1NkLPKs6qz8UpSQFCnNwTJ4gs0KGQJIfzYFzagcQ9eKJdgonIy9o4A4snKpczl1pgoGMG
90cvqk1nVQr2pNNOo2iMMD1wwTJOPZ1Sp6iIk/Xn8FU/7QES22DT2rd7MszJiHcZMo7Vi9ErnWma
QVDSHIexEnHz690vHjLmt0C7+5ba2lQPVuHgHPFZrQ/89BXxl3Tbp4h2HNPc3ElcnceuyOlOm3sW
AC+gCjr4ZBUOxNn0WRuHzat3dBBuT+8YWvyBYQLaiVvW4uhjJIuF2oaMutdJsw3Npk406wlMgZIU
03dQdxhccPr/ycGsz+eo1LdhI8202DttD1tpOfEUhPxM/PVU6d6rHpUIVXmcSVIsl2Xe+n6eRU3w
aNXgxCbPoIwXqjtAfqU7fBid0inENCzcgJZnrDIcvsoDHsfBoJBnKJ22S49eQu9hYCLo3dNWRT/E
VPr9EfycJZdBFTbDQcjasCDeGb1cUs2aUVc/j0KoP32k3tA+yEG4MxjC6UJrcJe8j73jHig3saFS
7e6MW9odWRzeWEc6gkToVbAASvgKj/+lp6FK6V9zUU5VVTM4b9HAytzPx3q78BC81bZ+96TlYXzM
Z8Ay9uCWuw5my4+4WJlMOSJNl/e+u2fedoC08eFB1qIzPLUiBEib0CzT/LHnTVuFIgKPNy4emV7G
FUJgr6wdFunho2Kzjmd8gW7TTfbPPeFqrz8oZgXqIICtGZpEkw0/T5VuKzhh4rbTpMmu8Jyxdmdl
dcoqWgUWlM9aOKes+EBs5lSZhVLtv59mTmcueScPth4yCciREl3R0U3w4AZ8QGVUvZ1RJhY8+3xE
nVuMPCl3CvOanuQGYyUyk1MpCWPaYgBeb8upcLdrkZlZ4JT03AfY83VN3YmSHm8jgTRiao7i23KL
nTl0dxeTWsOb3ZMoo7nyfj37v72dycJGj1UgKAJsKrb4OW6cgYn0Cb/Aq9y6cdQHUQMQi2NTMTyz
mJ+hBX8ngZOSHH2EL0yti7KCJIJ4hgX8aWwHYiZJc/JpecFgkX++ZpTk4kEkQnpHYurgIPnff5vl
6oKreO9SIkSvQn4PlkSDIAGxAzSj26zFJq6qBlXD9gZVvRIThCf+YUSrKuEjyyt71n+myAc42PQr
knZjMWKyIzEYO4nuToflWaL/6I3uYZtV1KOQazrtAJ+sH5gySYNas2Prs0L5z2DO0Y4VPiZaFH0m
d7PQNao2evoB9ieEBD9teUWjFupLZRC+LClfCZoqJ3q2dVRdxdxxh9OgVszOmA6L0U3PSU0bZQUj
HojMS1Uv35duOQd1IBRt7Jcem0g+Q8FWVsJKag+z8GAVfvnIJLb7eHa6vHPQDspex4dnVm38TOSm
QqwztFgpKruf7FOEUxgWXI/SkLl4Dyqy0Jvn29wlJfKrNMUIp7DQbYj35Gkkh4m6jlKkmy4Mz6wY
yWS1nAr+UFWg3hXrz/TBiV2Tsk6cVkDC7sx4mh/lbq3KiqlPoNj2kSavwcTRT4/5A4hZ5oy4otaz
+46ENNjbFoEsqhJf8ssVHCD+LJyDWBkLds/e2wp6GHe2uHmGi87PVdJm/plhRt4gDT5sfzyDSyaS
o4uZCTz2yCNynpZ51M7OOxdcBD1eHQv+EuU6uOtAFGSSDcLGN7G8lFUhRB/CQJ0SrJh0aiWzPmE2
e5WTc7dHSz5Z1LyLy7NMON0nxBPzRRyG0dGawTJpR5heP+hnIifWtzqQ+yAIF1xDsK4kbOfNLtG0
T/xt/nOOXZFv7XecluXnV/j3sGU3UWy9rVah7nHILImBwZxAOMaBUbIO/vKWC7yavPsMYdbDFDEe
E4DTMS2PCHYDg0VU6oMaNyICn+s/oaxtYGl2GAVXhiD8DSlgfoncP6UqVq+AkjRNQdP6CgAr/7Jx
YandCACQLaYDrVWyf92s9COprzFQRoQGKAwfp5uE3eQg5QZhgcENfCqeIQsVkAnI0uJzkmJvtw5H
armELiAJqt4jdD14PicQPRcQzpODoxvYXcHy6N+uApvX4PPFrXzdvnJDFVTbLIfbP5FEixHKTieu
tIXBZhnICOYyOTgXG0V296UulCBazOLW5DexV2JIPio7TVzAyuYJXvR0UGKOfaHaFhwvl41nkNrK
vrVsaSxurHmIGSWqn/juNuQ3vB5KCaA16iTtN9HzMWgKrAHhOol5FY67ctPuFnJByEeLkv6pTbRL
w8CK0sm7IUFxUDoKIANRNg7V8O6A7zUL+aF0hlLVmmOBAty2lUz3MTXMcV0BPRUqQ2AT9qGovk4T
5x3kCbG5F4VAwfI4H2xKAWsLjCHesCXjIdTbH64qyaZW/Ard3ecVnSVnAQNYUw5jyqQGDqg4O6qF
gzTWT3UyROHuH48I1cbPhB9fgt7BuoWoCnSqTYN55ySyRmPMM7hdx+nxmGjX/4jjvTM1G4AN9x8k
5VrGS/bnV2Aj5kB1OxC6OHUx/24Om+W6IYynPeikuIGz38UOsUk59+UDDyiUE6DMnidwJTSJt7Sy
gsdTv+e7/wO4pqscU9XEobt7mroTvTNSbWBsZBvUQlm1NqcCQdUTqRxmOM332wN21qw/LZ8j+Hhx
+yJkMJe6Wq1tzbKEDPQ3t/PCUH454ki11FnyIZTwj+Dl6YfNMElmMqnF3VFMcWdSsTk7u68tCaHp
EYGgq9uvaNYRcv7E8ZCdMgn7C4ir5xeiJaAJnM81q/zM9B8NLXUqBnbJH7sCDCrblmjJL9jwbPCp
pdiyTLIChcPXLL2DL3q1ego6DPbbCYNLSTFla/wyl02rKQJHkpmaZzFtsjjrc6cW2FJse7PC2n0p
/67QDkQZpvMgvtJLIj9nl1FaXoi3wrG8N5iJRa+1J0g5KACkkvj6/Q4IRxwr7Jnt1RAtndzLqbqM
17Z4/JL2+WOtR6KBA+jLJm2xRLQ72xdIXOOowDo9F6IzK8MXymJVLl/ru0FwvRQ6YK6WWVJQn61i
t0CLIVgS2bO3pPlhgBhAnlNTiYm3rjS+CigoMXKtKG59Y5Bk9KkS+23MWrZZrbwGF/7jRbdzOJtK
WCIHi9rRlMbgSuuwzAMdCWzfqWhkTWnWNoj5cKAKQM8ZTh+xRWYY+c5V7wPGXlDs3rt1MqNLt5F6
NKXRGld58muxOzzPBKEaKOkkzPjFAPR7Sdt9jF9dMLlVDiuU+zWvHRuPpyiehqdwbpjyBAca8euS
6O+BtyPAc8DxkxVBfGJBU0W96cKyAo8vVRl7PtUwLqlCVHGKyMqzCUZi5FLPcU5Ql6J1MAyfmPkL
kqYJUZzjQy1HfMEdo6Bra8/jiFnmcapN5v/NexGrjCmOqRtKSs5X5JIiL7hdKv4kd3hAKkYlzopt
Ep2cOicAVKRUFyq17WW2dAlQz2rdVFZJGp3w7TyTol/JXao1aepy5+UONeY8yg3GRggvK0hMGtOO
x8aQ4oj+e2Vh6bBZtKg8C8YjJG4zu9uy5fIsXWhHd4ZVH5Wr/wjEuKXmZ/v70+CODZS9onesi7Fg
uNL+czi5xw1xrcejaSPuejYBbUDn4HAPpG4Mrp/CVNeEZV61JQ/cn9yQCFRP7KlfkENLzTtDgKrQ
/BedTNspGcdaSEYGTKWnoPXfk7eDSr5keDHvdbkSo/9Da2NEth9jMENIGFO5cqV4GeadI/1r20sc
ZEmxdGscRlb8EwXvJKCf6wm2fCE6O5OTWomuCfPNwJOKDHP6xLuDHBdxZQvzAuzX/60uFwg5LXud
Gm7wKoRWRmYisci0aLZJX02OdToKqaJbHQ1eA2sqeFtM4HyUoyiIa32ic+iq338YIV4JfU+PmIP6
mqfUpfzO/FXBdG6PwOSs1XCgT+RB/xrdBc10JgL8ss4pxrq9VwzF3PDEa5cDDATLBjtsKJk1Wk8c
KMHGsF33j/KhsJ67tEddmp9loipRyyeCYE7enDm1CMTtqjysEfKxKJ22SuP0JAxdTaXNtEfTS3LY
cNykBtwv1OY5BQBaKyCKe4aLHB86Q+d8/c0ACFdhLNJT3cI44s1lHeLVwY/xoaekzFNndtckK1Bs
eKoX1P8Uj5Cmd0l0mGbgQJaxpCZdZ4zGyqqUsOinKKQvXhuBdtnGOcHRAXnbKRL0FyIhO1Opks43
pjCLvFbiiZwNcE7+UHutJk4L2KAEugpePfSmz+ry5CeIU2tsfzUqKVvmCFcE9d14rgVRS/SE1lID
EzyfoRsusOa36+UYAfnkyLY0DuL8E6dVL3l7FfZCL5lwoKF9f2UslUrCwg9CVpq7lyXifVy4UOGY
WQ4fTcuqh+mIlcSBoPer5XsBYZEqMkBW5tILDa8sKMi44h7FAMZ3QaM8NIWiJS4kYCtXtbnNp4m0
dLea4wAUGB9v1Yro8XuqkpWYUk9gNsbJJXG+ebqcWzisxEoGM7B7zz03BqASodkrMyfMzzfc5QQY
HCfhijorgflafNFpe/BuPCvsfEbidA850gOUDjd7yWmNQqCeZOFF/mHULTuN4cWfzQuDGn56vMdY
KZh/cGYk5QltwjhvaZUk+k1oZM2fdoQnwoDvyfyVqBu+6UW3NQAcuwU8z5j4jfgmk7DuS0Ru82PG
77EVYgtGs6taPzqwRmONdziN+98y0l7t4T2QXgj8bIqxWIgThLfvFTqOmFsBRIr58B/b45yCbcAw
S6QMMIs6gz5LzFe+mOFbJB4ZxF+RioRRHRYvWJ7UzgCRuUxG7dwdVwSuWjwzF8HGA7FE2YmdzWu+
XewveVOwwrVwPZwGUJgxJ+fO3E9pPCTn0/ui1nIUDG+Ph1p1YPorydyUonQwsujyC3Kphx5lVtFq
VBvQIYY/EGIkpd0xfiK3ynJbztmOLOM+ridgVIwRhLLh83YPpY2v+zZUKzs6WdNdf24+uGG1l79J
emEDo/EXtAnRnWJu2xMxa4ivUHflz9EDrF0pXWMleYvF+0VhMNOmDMi8nynE++OE+y1USXtTfeUF
LocrS1fGKlBBeVacOnl+RFKxIHOdymZZJIKu3DBc982wFUvExjy9GuhmLC7eA+Dcao0fwgaan7x+
Z9t66LsZow2arIU03/YedmexH+i/G9YhbsVh9opVPacFMqlhCgBGT4DFN11Hes4mXZaDSH4hkZA5
u6VEJ1aqnc43SltXaOObz+OZGkuA4maWqBiB46sykhAC
`protect end_protected
