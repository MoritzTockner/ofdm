-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rlEPrP6ZJZL1XDqFveKCzVKXGZduM+DzYOV3gRqYrfSCnbkMYNYB/CTyKI/mQdNoK8BiKonNwdPm
P/rMXR82tgYmLUhJA8drOq8YqQGjbpsQ8ErDIRTnFCzDbCe8eAekv4bjLXJwhqJAvl+GPugcLxlX
82IsIdOK/2XGKOlO5AG06PbHlrA6ehmFL2lHx3oEjZdpGLrGStK2d8fDiQqFL90A8/IqCyYtUwIu
Bj2rSAM3hLXscsviROB3WimN8e6vtvtCNvtq7mciz/whC3Hyp5GGwKH9nhNKDFcJSbpMWBLBY0pL
tux98eX7fDAorvQTf+FOYcj5o/U0fHgwcO8sRA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
S02bhgwKY759ocXGlCdbMTojm12UwMXTqcWb7/DTaFl5BTlrc79nEk3FL9VPuXaQ1KpEY0P9o9fs
cQyk3Ot4JjE8iNEVXEgUlLNtJWRQEPo5cJ7dcbnRT8MK94+oj5M59C1icJZP7MpBoBjXc0rvUprn
1Qyw2gE9EkivCtQrE7DBHh8iZ/HH6q5WPfFBcYKLawIAO78WkfVaQfJc1m7Jfo7cKlrIR7KKppCH
vNZ9lIswKY6AOpWC0jZ1APZPwSSM/E/Y+n91Lc5fdH4W82gb8khhp9BganDzoBzc2niSQf1/Yrbc
ZoMvgHyDG6jq/0hkTpM0P/Y2zKacoBg3zl6mTXg6cv4I8QQr04Tx9/xa5M/dBZnGitBFRLyuk92k
K9sDrB9Izg3HZq264Xsz0Ux9oMlMhE3UVwOsWsncGsSPZp5xF4KrbuxxjOjAB+/xrElNtmT9YEyh
yafpBdrsZlWvvRrPtMoUBkNZQE4F1h01z4tTSeRcIr9f+2IMBzc0ZZvIhmvfeNt33DhS+Zaz8yUA
Hg1jHc2WNzBGTsuvSn3m+TmrLNuUxh65qKvxAsGFK9yczHZ45ijDNf+Q/TN16rDmHWLXvY7Tnx8M
Cs7W1kFw6Pt8TpF7713MRVFvFpA92J1EIJCUgIN4JxZXLJv4veu98hPED7y68KjtaKE6+SctaRxe
68RYxHp4uXRjBXpS+tPi95F3/xkyqZ383yZes/jMJVsgNWoIjlAr+QF6Tt0AuprjzD9vORPZqEYd
LzbPcTVmOnvLxuxTaAjRGzO334gYu0laH8f1pjjiZWXolHMo4Xn/aoEj/JAP5YjrToUCFtw+ReY4
VYRU4IW8AstccSp+zykHbsxurLL0liCzYS8mt0R5g8YYeQNQUV5k/GC797FvEHe9zFk31uyczdyx
hVsHKqPkTmpGyjToBaUjWsAEfNFfBvvmB10qw5eSMvQw0K2tLPhtq9glcWRLeoAfHkzdts57OEbZ
HScugeUNijvQ3e3pVmkiDSZcyfYsyd/7Z9qvzNKjk7twMLoSTrFqZ0MzkvQ1vIu8oidFp6AOBVg5
iY94IcgbWr7M8E3CRc5lqrlQueVDsfxJHVDgyeJ/W7i5369feNUoYO9dSS3yYqMjNupGe2ElBDuT
eDLNylCPTpE4Y6HiKxaCpGI2IhUPGVVaNpzMXYcHXR2+/eAL82Jfmk67x6GXH9bATc9RWlgvfCG/
3HGbLiNaDaXi3q8DqXLFGydrZjtfLfjedqzlSLUax28XvKq9fZsb4PUNtAdpPrQDNwFhuBaye7WT
RZO7h3Xe1vh7oDwSL/sahNFKyP6IB5RsBAWBZaeanoHUNUcqxSPsazXkF8VivAN8a238yjPUXIt4
ltztZ8Kqv2Nb3IUdHhopF3M/2NN4l+nf1XKfUXV2waHiLqBZi2jVUXmkU744z/JV6pSghRispS8C
sOvDlzp/p1MI3apzmMVEgg5QJcblF9vSB3vnh5QWy5MdJiNvCIskMscG3TRWU0X7jHEmwT2YyLKH
hmA/mTqxpjOaQPaFL7i1POFPB6I/in4VA6GBPqifeCF7sXxMPUqzwDRekHasPh/wnCHNRpsnIe7R
t0VjAOrHn+DlxyWB1NY/eJ5d4L0HyrUAgeA1nQvqHA1KRrkGhYtr0pv+6LbzDdhmqUktOoKInh6Q
8NmvXYoe3gROXdVFkZN7Ob+oAMF0eqAj6EAvLEsW0olk/MrI2M1xNyrGVXusgkcu6nHNBz5/3Cvp
pvBInjlCdGS6YStxHMnhSP90a2iP6lVwt6Bl1v8l8IitH1v7fdP9yUp/Q1QRRB1ZelaU0kUEiF69
yfvjVk4NN4ojZ7aDR+FyFgZJIKDBSxuCteQ7P8yhYaWfAS3LY2MR4yMBqd53WEFq5u4eDWzev/b0
YGBl5tTZ+K21u0JmsvMkpV4PPJoV06aewWM3N4iCX9ZGCUOdeSExKPo010ii25sJUIItWts/65eu
9bB9+sjrmTlGQzS3jOXkIHhdyK5dVqgYZ0PctCGcsKvs4cKrq+jPU1yCkCHizaL68aSY4nKDuOF5
Xwnj5YrE2lNqnADp4yR1ptvztqs1NL3ULhT6Y1A9FixFCTCtcyFa52O1Ulu9Dfq4W5dSvmh2blEM
DBMWTxyWaSz86ak2+/fLfRkw4R6BMwya4VitFJN9F4AqIowysUOuT7pZyalcK3tYrvGOmeUp8frg
1vspQuwRLYrZXgHuA1/+3juOILKynP26UHNYjMxfCYA4AGA9kJI23n0WG9TCp+9URpyLLKkiz+Ng
pJQFGJ8LyyvxUggdInX8F+tA+sFrbI1N3LXAN13d388/R+AFXi9TgiGGztSUwCG1ARZf6JWMs3Im
6QMIyBQYB0dwXTTs18wwXRN82C0ClyhCjgbPU0vQTi2YU0YoaN1fAvRw5hxcQEqGcbSrVl+arYlW
ZrP0neBW6k03saKFIpVcZOFza8m5k3d04vDyZiBHoylj+1FyxJRzjtm9otVaZWI6OcMKBc/ACflg
xuezusnTV2QwgDYlcg08r1IIJYkT32ln3khxFvMbN9scj0hZcfZ1VUp8ySxgyqv9/GSXrzBMYNNe
W9WCH+uyAZ0rQdFQ6345ETclqf13EgpoHf/98C8RB4xN1b2sND6zFVyMad5VCsB8FvQlraGrhhOF
bHrRd44kfhyKtlJiZdvlyGeAqFx2S/66Xvq9q0CPR86K7qSfxALNOosKq0TPMyIqEz4LzVLIJHvm
Uj0M7oIC3poq+EyvB6IERZmH4eJz6r5fjl2kpN675N4gzG6ofbE3dzefv58o6CWixhyU9HCXyVif
T8Ynu10nOgsOQiU4DRcxfLo7Yh7mn9jxJlwLHF0KMPJ6781qCO4J1pZc7KQCDujcrbIYiXM3eb0G
pM68/Di+emNqtcbQCMtoWfBvbrvBgLGQUQxYSplBOW6M1hRZofdl9e6EF35EnQMwKM4QpkMgVx6d
ekNnskJylGIuNLXSgeOIfoM4bjq5ylpSbyXR60AhQpQJtlCTVU/zwuRVMiunpJB5hr6pBCh4fqMo
z3rBuEu2X+f+Fzu33/2edatopkEzCY687tKt6eRuFqv1JsFBhhhxxd/iXv1t/T+ka/jTnNdpAGPu
BY49Uk9l6mhCE7MubggbPht+fgC5Ts/PGMTOvIwzuM3dPxZ5olhAnUEWCWQglygh3PK5L3UCO5rf
c1LJwukd+x8hNtzRgY4eBhvzRVygorWHFagbEcXKbuyRR/mJHIrdhNRZT/R6snPBSURl61cA2L1+
vTt36CV8fDqHVTjjAF3nmJNxoczTxRgV54CUpLPQiFliqA18brhw0d4sPVixKK76suzT0OWzskHE
ITogqeEvdA5LyKgx7yBcjzB0SX/KQWuQjQ7dPqViWMkQfKhlZJFWOLKD+8KhVQ4VRAojczkKmNc+
B0jloLSpvtwQYB5DasnMU/LzCvQEArPhFGxBv2r7uoIjmfLkEwMXhzJByAETQ12arXZmGh2goVUP
VZTn4T33hMZNC4R1IYIebtyiU2kJVg+MM51jpEeD/MbYoE/Cvu7sJWap0nJvzdyB2JIZUI9GuiCK
5rVXWjzBKIaGnVYjYfc4KLnUYd+yUxvxJ6vdAF4fQUNG7kjTnHaI++ilImi4IZhmY32DEtFiqZSS
su8G1dZq1Qo7Y0c2FSwPI5VjRNvkpbTgTU4+3rn/2H86QohQov6ygrr99Zpyke83N+4OvIdjsFQW
pNtLTnEUjCbf772CAJ9kvDJ+Za4zvw/m+4+LVwe6zlf/0Q3vP6KP/MhmqJutlFuxnUcHJt6Qs0gK
xFFdElcnZu2wFouSy6QbcY950WJOLB4yXSk4ZLzu1NEaln9QdobLOTysw9+hhAwCSyn/97eA1nDh
zMA1/p3DHvO23QFzwCrSjcVugpY6tgrcHjJDvzj1VadvlPXVQgwlu8KjTTFSbkU4bTTbbTxk/zYr
MMNcoKIpAIaZsjZKPLNapk+cTkJlL3LmIWCr05eMKiiwtof6SmGoiM07GWdIqHju9Eb6KPo2z2xe
GAjuBThaw7eveuryw0ECs6b8XPa67tHflQy5Mz4Vv3aspRvSief/EFgLNhfmkC2mZzyT7MrHtUfD
gw1pNtQBoKoXcBUcSEuBrpksbRNBSwLt1vCiFeFL9IjLFK4FwzfynWshVJ6LOWKcFkzbzTZS9Sa4
Jz0SARAT7kxk+441j2WDVdJe3ud6tNflNfeZsALcvQbtFdOLtfdxAXdSzEVPGxzhicH5/rJJU7vU
iW76MA5WDc78ynAEUHvYCPrrc6xbUJ35ET21/uSL0S3Fzj8SHnwOQWpxM2E92NiDiTjMzAsFPcIP
oOrlAM1nrG0o3Duk+Nxlxc/W+iOtU1WCwfPwf7VSV0HLz6n+pqcC3ilHeITNZeDk05+xvINu3wrE
MsLof0XAxs+iZVGNOUxemZK+Z5GvowLvcqitaA28CnR0Un1epoRLIIu+FX7AoorSO+gNbq9SdS2v
L96ZCkUQI3k2QRHMTDngKc0U+STMobGdqTduf5EviB9p+0mvsdmEMMynHIxB3VTy3eOQM9vTOnJM
bNFM0Do2Nu/nNAckFAmVl1FXvk0BxL8FAZ1XX84Nt5ovF4O1JTvVVN5072b9WeSqFePaSHVAYgi0
CGhlYvZEWfcb7uUybStReR1mv5X5nHnIYOIKf4VuZIXzzVfrm9qLbdYXBhBopq8q7q73eBfZEkvc
54/jJ81pRAdGffTRWWGio8SVN3zfk9eSAaQOpfr93X28DhrPCHRA8mNN1+/vcejjPQwKNQ9OkR9+
I7PlVKYt+7JYX73Yh/WU72/i66krFsMGWaxHuEGCGysTtuVjsm6v0Snbsd35ONHkrxmpFU0/7MEH
ifhy3pmAQRLihO38a9O5eXSTkFqB2jkGcEtRoks6L38LUuXOgvpmMBcJDm/748XkDSFJVCHDM33b
WrK+mlnPEdY7+bwaENMnj5zqIBgCL+f7O8ORFCygwLlkxWRZUm9rszMGV5Uwd339Yd5GpPBkAql/
Ze1ZzD12kgAzR422qbWfkgpuSNIAqiFMZI4M1wmuEHO/JJ/Pb5mYgyMGmoB56oJpjFiQ8+bb4nRy
zvQ6CtveA3MKsobZ8A9wNXizgUA0THZF/JGgDoIA5fXF0VKE+CdQPbGgHR16aQ6LUgaKx49GI30H
VAj4AgIAGejJ2urhQC8polPpebOZqz/ohzD3H5OsHXVAQ461zcsK8fI59u4JNtVH2SyHWXjVUKY7
wCKHvmeztGWg5T1CO2njVUIj9Ob8QSH58yoKkDKr0Mx2iA8pLdkzouic0gbYUlotgP6FZTvnTjle
woC/GrJc2IZXpHRTtZIKiY/Yg61JT4S7/K6FJBKDP3SizxjVwi7Cayj5CoBxQ6WuyTMWIw9XQ+o3
LQyMl1uub3e/yUDwRE2OHGDAUy7jmwNWfvvULXlNrHY0YjHKh+8aAzTD/oMtZbILAvhhaPM+Kc5L
a8rPseecVlmnbJCjosl1iBPrUOPCZJGNZzQjJTbccBrOaNoFhITIuUCBcToD0/ABVMeSqi89OHsQ
3lrczrzHz9ppvQNPKB8k9WV8bnPbzcJUhzH8LFV1aOdBYERQGittQjepxz4WnjUY9jlXAvA+Z3Ds
24LGn9Pmz6gaRbVe4FgpN51LieJjmtp9Pd+CnP6yHjpPLXLMDPBehhaHi+BjYk2dcnaFKLnQofct
JcIEtextvLX3vKKmKnpXCYTbfXh6eJ2wmGWubMP9bA+9l7r/VCEuf1rDewsd1Q/JxPJ2Qea44pwx
q4MIdBmAJhPKUD7YMRI3ncWM0B+rSwA8qAHXMdcNO0Wk/2CsFku+69jy0llqu/SpycxPu+N+gvqt
KdrgmZvk+vVpElPCuy1wt3DaFIIvRf8f9RwSpFcdlXFeeOBIjkGXD+PWUJ7oVpla9Hj8asKAuqQ8
3HLmIxhxNBpVV32M41uJOa3SWpUcC30pbrHYUUhC+oMt45/bFvou5uHOs6KJ3acdscDK9JNL7qYK
dx8Tm32xzGKSjhaFVsHlCI/HDgNH4uAXaxcvWQyivw3yI7DCNjd25me9+iiKLKppRISOQHhqM/c9
mpJHxwxpcDXB2+G87M0TOWTFg0fyDRpUoHSSD7+8QGL1q/+i27Ip8v62K6ZdyP89FPqRsPlneGT+
eol8jZazCL40F2bh15XsaPqw2vbseDpTeVjbU1JN933gfzN+B9uNbMI6xd4Z6sBuwxoFK4jRnQpu
Qyuoee2ywNviVXpsQSDhpcPB1NIALvEbnWl0KvJ814LTUuwu9YYDuYTioCxkGSrV/EOSdDbRprA6
2vyiuxrUomvfrFIeZyyZneTyVS+83BjDpFerXHLpG2uKBHXy4LUJ3OKFdMNC2gKwNhiBLNIWKLFm
7Q4yF+uijd7avl6SYk0iIrfPKpOjm5AMy0ZIK8nDUMxGD4u9Ll1q8EcdttjhqMrIAG9i8EeWtuxq
reuLl/X68zFr68mcbDWpJafUPBprGw8juVhCZ6njLmhnQCG2L2Bq+UwmmDMwv0zBkUflS9xhpAzG
o67ITnxaVb6UQv8sBvQjgb2n0tnzCt/gWWQF5jjDFEShw7orHrQB33oZ4YgsUXK+/xVoGK2TlXmB
qBC/0IwOi2C01m/J2/p3Z3kLs9rcF5VXcM13xIWJ7llByw63d0+G9iKNBz7iPQ43iDLm/0qCnx53
xDNrAVmi6czTY3JUf3MwqMeCB8H66Q4QqmwR0Z+vPnoaiur5tatHl4ZxrmGW3FY6SaxbiyVhLJst
MljvjTCHeykiuo6ZdLh4sOMpE+sEYal/zEozK46ganKJKVxMO4yTrMAdVpEJW9AJFkkc6RSUkXKS
h2UeQWuPMnRlj8ZcLlgvzaeVOe/RJSAqov9pkcCJNi3LDqxzS8mkhh3aKRyKxvHiU3Z62pDztM3e
gOpka2bteHui+NeYlDHNZuEV6EU/4xFLZ6PYcYUB4hkGw7UY9/GbSXztYje8+NP9MNh2wjgL/AlF
trIzYCdODRiuzXkl66RQQLz0i0gd+I7PjaR3yn6MQ6zShxkDLcSx+k/dnhISLhrDM3m5ZftFqIkm
wgQKhMI/Du5eAe+L6K5mqA+qvHpYT9rvkNwFBx2JN9QunlHs7AJsdGZ9rcDQJFKNbBjP30mUN/uq
D0+QrwF2fb2o8TmLcpeZJC29QTgr6SdS2eqh+hRctsyf/mP5Tqcg7tS2cIUSvjetukfB8BgoOUQ0
oXfNZ323RfeXRinUQ5HwzuFiLiKnhq71W7zgtkxTpooBL+w3SiMV9tqUx04ccraB7RYBzPWNVSfZ
uxwjCjrP3e47M9BGQaZJm+kIt1BsCVqnc4v4brcQ6gwzlzqXle0hmkNQbfpMXash/HqBdF7j32KD
XPPQ/n8dHb9d6GG1Dbz4mY/X1jXpZ7/A4wYfGbvxcLIA7s6OKoL9hBRfSUybwGwG1cvaIxGViUMg
G5u0KT/Ug4qGm84JrsENva8xJvE/FK89HqcYHCwJOtF4AEgRqRdR8USheS7rZ3sayj+Us6DbCUyd
2XsN+ZisWffYJk+yPDy87nL7FNRMQ1CaZAQ3eTjAt3kVy2RnyYzy1yLojtew1CBlogM/EEDC1r4g
VzabMQK0k7tONHTj0IqKQwyLHYZfj+6kU1VoTMtCXk5+uHDCyHTE7S6A5BVFZRSbKgosJe4p1sPU
kmFY37sn6HkMEy2+ehHKruVZmsNODncp3KF8lK0wRM+wn0SZxd25l41sHK2c+NBkp57I1t/c8uFq
l6Cjr9JYGB4dpeLAoIk9Kpmqxt2Y3IkG0AkFUeSrO/4sPF5Bq7V16iL2aVs/oDDRGEhpwxLLySYF
VVUZve8LyCRm4MEcjNkxfX1T36RspnzpaR1LNmC6zwl87Be3j5Lsskt/vvD4vXvrf3+F+kkTGOn6
HNoMDw74md5jfFVskNzZkdC2iermT7vUW5ovJ+81imyLUW1e1gXBFtuYpdQhFzVyGs7ApB9vC5JT
p+IjhimRna9KCq1eX0KlA0L0V5VEOj33slZ3FDyiAycI7e2OQhm5DLp9LQtrNViXY0qw5apf5WXl
jwSgCt25YqQZfMaCUgXRTVzrI8BWBOU/WVy33sqPQgGHEanHLHjcYIYUXZUQjRHafKcQOPMCHPwC
8qUD+ATB7ok3pvb9MGuMY/EpjUteQVE0ogPxxqgWA2haJNKbI3C04m8E/5Db07CoMyNGbUluRuTa
qL+Sh5ocF1zQIb0GGueht6DAOqjiSn4ClZ7kvHzym6Ag/gFaqFJ6sfXVhGwOpcTr2OoQetI5j/yr
HhcGS5kDO9p8s5SrrnynU1KDmTwC2blK+jCtLOKoF6XpNJ4DhZM1Y7bczREZX4JaA6TFfK4A2gDe
OEDi5p+He1T88b0NDyYXgmiMLy5T+gUNxFAcptQZaaawPSlXVgEPDLSQQgGeYlC4Lp8clnuI82oM
dzFI3c13Xj3pPAq9H5YojnvlKL89I1bgQPXyaSW+gJfGTqjRga/nvxVJgOQDnD3t+hum/stliuPO
dRnevxuRoR5tTp97llsZ7g33d6fnXmNdd06s0UnGMgTNk6aJC1MnAjWsPtm9Ygl09ZhMTcF4Url7
eF82qmombQtzpVIStPzRBu/te85BzTh5bAlZCt8e9ZKTr29+WTsQt/Uq7TkhrVxAMSr/0U75wG5w
le4mvhjpmnzkmy8/mjezaLsmj3vzTdYW5PjLF+ilJ0W93UmtL/TgvMrkOjUyBQbjVfuGSte+tqa9
V6kDki46NHP8rGVfW7HJAyKLMHdn6ZywSjeVfyPkmEelxswZQRP5sHGDR0WUwQHmWaThlm6zulAy
0pdLFaSB7WIgPGY84LTBgUMkszFZbJYsagvI9FWa0Ices3wN0q7Jr7lpSxBG+3LW+cqXvlbEnpOc
kwv+uYT0QYVpMSAaUZAnZ62A/0lkAAaY2lsYPjJOfYe7cONu47noeH97FHoQOapsqk1Jr+TKgqV8
ykK+T95IX56AZ6DVqfsJ51ytl6OffUjvUSNkX93d5YDgzmPsUUCUZvE8YSwEThdutxQkCh5s+uLe
hayfTkOGwfvndRjPTKCrE8+AFavWLwnlX4RKIFFDS8wTZ566KnLevdhUzvkALQAELTM/qObFKt8l
JlTwyYB/unaBK+ZNhivmRB4P/UBjM56Ka5vOTc0C3neRIASUdIjNF9K/rgSDwhx5ufDzOVylbAKD
BohMZWdpRQF0piGvcc3sPRS9FZgXROxT+PNXDhv80NBrE0EWhcLoSmEQI9vJw3DUNYJqmAqGyqEx
nPj/y8hrNAk+gsG1mx8SE3dNbbLIIFjFWphp+e2FKe3F0ZmPRGbt9F+zBAAK7z2WTGd0/Nv0t2H+
BTl5rG3YzbPAaffUn06kv1t/sNV6zoM+iVwdP9899qPkSeZpPHuuqxfaPjgqcboNCNeqYoxwAJ0u
mPI4AG6AGoAHEjXUbv+U9o2qvoDKG7b9ZVmKGnZsfTmdlpANgePjZxsfxzL/gedUgj4W3c0s3GZB
wpyrzVPyg/DD72ZVrdH/M2HMVi6onbkyeTsCo5l8aiaeKJgQCU+/KKeDEbo/kkCmwDP0OIKYmtlh
gRCPHdQwqELIHQOlA7mIxUgwfDyGyNXdoZs9cp41x5o5Qiju4BxvA19C5TynFmM3ivHgoTy5M2xy
ATv83RrYCXW1IxIFcfzQZrJ0MFF0lmQS8Rr+D3KPyWOZApgbU0rq411Ju17NfDkKuGRpeKS4fBJb
sykr79xpFbqQreDAuI886FEmOp+/Ua7GYBV8yH80VRWm6de3HkpkQi7WqQVxORzhhztlZUD2cHl6
FWWMYMaxSwuDDMJ5B+wU6jglpCvpTs+xtsBu+5OqI8dpfIYNRqSXFSuP2ANMXQ1q/y/ZJZrVKXih
UkXo1zCZDiTNzO7nbc8PpY9rQqPYARjCdSP58RNLNuuEHa/noeHXWKvqfFU55qX2rs1ry7Awpin8
nLu5Md/deVnTOkjUEyYfgsi513HJbi0ayGsDllnRxqfPTQG+TE2bd+An/X3mk2BrtP0UfIRR7bj4
NurluesuiBR7kHosvVAN/9O8N68fRWoI9B+2JnLCpxx4YGkrVEj+r8UApfYZIXbxrIYdih+IUue4
9oHIf0rfNdBMG1+XnUhKNQRZg2jTbsnzVbPVQnOL0bWsd+pg/fkp2hYIKSxCBmpNq9VQp5tupPEX
+mXAQtJDPmtfQJIVbtnTL/SpgN8NknLCYjSWU/qCKuStzAqkcVW1kANbdQh9JLpj9Kwsc1Q7eQpn
JOHVSxAtEP+W/zmGfjoI8/5aF5n4YrtkUPJ14YLJqm5clUCDV0pX7KQP9Cm8EUilCMfV2KAoX45T
Nip+XJ/XU6hfluphgAK2KilENCAc0b3dtmndCsoRgf/7th7p7Tb1U/JWD8Eg3dczcrP/RntVATPz
d59AvWDOv6tJ6OuK9Vkhl8vKCtP3kaUHUkzJ90xrgZddEh1Lg2KXId7d+i/tzhKsBEfREXFGGsa2
D38LPkbWYA4KOcAb56ugiDpvoIyP20NVMMsE4IzSBPxdDe8k9JiaaN0qYdwzhXHt/Fn1qyW8xiRS
58QMjWxPJPPcKWqlamjFOJnYNEgnmKcPMfeBeskQHH37LeSEel+B31JQh4Ev1pYi4GNVI8ncsyo9
OehBGVaRYAMlD3dzbiQMbDSCXajUJdpy8sDDyv5Nk9Bdpe/mts/s19wZ5dlOYzWbbEIl9wS80A4A
y+33x34BezvT2xN/mkiiJ5pUZYfDqXfgzmHM+9/adTnCFovz48BnC8pQkW3yiOKwkbClzLHu7xgq
QJ1PuDngx1UsOYwxwrObF26oW9vTiaNHrxx89PufpQ2Vfb9J2zbH+aUIbuk0QC+gRI2GRuGsbBHn
B15WPR6GoIefQB+l+J8wbBvpjiq068oxscgEChv5cAXCOkLRhbev7ywdq6jGi3EABs3H8q1bjLR2
pBSfpn9Ny63RTDMQ9+pZsa9Gm0uyCa/os3B4BxkI8R3T2YqAOxQ84tBJLza04qzfeiSvmxsAfifk
IiEd7K+fEKH4xKlH19m+7QBeBPBn4355HtwpjkZ4GTgf1t8tc2JyDClJMGO299r9FqpFDXkyt5C0
lel7CVzKAymjTmBk5/AFZQdTWFkmL1pkMnq9Y0IRT7ibiNe0GULywDLaJPHn5Mujwr2Oe9uVx6yw
N6xyo55GlpCX4OKAdJeefwuQz2+LxCkXT3IBCxXexbqRoqzQMF1/kaP6T5JIDg312ESMf69ayWmD
two6nJkJQWOg1sVRTVD2brybKgSSgd85wiUPyxBgxkGkYDUYsq1JEYHlk4txWHOrNoHg/9yFvbCi
9Be4187RPOMdLHoVsi4zgoFSF53tFkd+yZfn0khroD56xG6r8jnml3OyoWcudu/bN4umP6v7qW6Q
Ai8jKfr/0qo+7WVFaeymki1mdSfOT+pXHo8cgy6w0VoF2d3x6fZVbMsoRvtZVBK34f5NJd9DTqZU
py10bO0GuMvqlI7xzJcrxyhUSvhJPuklNa1b5lpy6TgNMl9w9MLZbR2WdODm9MtzTKYNJvpVJteC
rn/G342gJDEpUFE3+F6OzcLv3gsrrBSMna4SYJTxKncX0hQXpebgbcHxmxJzi8YIVRJb0rZpybac
X6lIts3W0/VPaGxzqSalXcqBX7Z9wKUUB4hDDUDhR5y2y/9z8y0TwSOwhj/ijJsKCBJamTcb74SG
t9fOBaPrGld0Y2P+pL0Iyn773/Dq+2seJhz5mGTLgeMj6Tz8ZMJBI812woiQ2zm33Z4wgIF0aCok
tvBmitmXIQkPQX2s1g==
`protect end_protected
