-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pmk85KjoNDZrY8J7lRWeuSJcDJQ0iGnpHZKG9dkUKHYp+xxBuldH6wgt/ndU3x9EevGH20aKB8hZ
UT0S7UzMx89miJVYl9kxh/qk2Zc20K+NnOp4+0j98Pj98kxC6sn5Jqwv5ts90Qi9hb7s+hP+Wwdm
291WBoP+ifLhZNuz5E6vt35maZs5vs33zWxgoMt3iOoJfVWxZiaVYoCW12NA8hyqnyTT2WfMulU3
9/YD5yVFOzYRqEWHhlmWaY2YshTwngSjJFDzMz+Uk6a1GQh7ud3Ja8itqg3n4SysOQHulpOy1sOS
EONhnfyYKaNgRbdrCT6kbAJopRmojDJt5jCFfA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
Tc0HENCb8Sy7bP9TJgzfyLCSmnnTmNUJvP4HLNxwNun50787uZEV2Wim3XcZJG1ifhDiczGfYduV
oeCth/2FalyoWbIOlt2uth2iGTCnKqnJgR8LD1v/FpcN56JCq7I3M7rEFKLsQhey6J/chz9THnwB
H7hv4Bf/PfyBeuWWG0l5UnMmGBIuDj57w27LH0oBzuw7gkiieXLM9eDZZ3tsXTGpt0wK5murac84
4Mp/XLMqBprbcY/Pz+vqE3wEZQCb1Mhw/bMY6UNAMR5jfAwF2VRkQ20jz6ixkC5d6jJ/yYIoFSly
oPDXM39R58HeopmeXuNPXXYGasVm9Esyu/Q9qVw+haaEMEJXb5rIXuP0w+//aFloSAjmbx0qPNVG
gZkKHvcolyPwDY7/lD1FN8EJuP91alsGCs5GNVTUkn1qeI2LI77DllPfVyjDx183psSRWPY/DP5w
6EPgGmGiZrRMhX50YpM1osA2M8kt4JCpTVKF1V9cqe59Udy5P32+GDGytwRg0GmikRWWsWPMH7xO
kg1QxtzlIVqATg9FHY9H51U/yDYenLKZD4ONaKFFcd+Mv8TvCPdNk3mcjNBaAWj/Zs3tCS8zKK18
uucPDbAmRutWNVbe3XVqSyXVx4+jD9yERKPLUMrqZg87/rfehs3CLODFMD/e7IaC3nf8HDIxA7sR
AIAByja7rcZpWqLE+eHrfN7PhIa/oUh5sK/y/8gvQdAEbJ9TfyX/Jy4ahtKjVB+6InJaUI2BPWBo
dKQnz5aL/qvjVLPcl5RaPTOA1pYwoBodpU0VE5kmMYprteDqCpktWpwwr4s1LMUUbk37942jSSLR
5acev9sVYbfLxNIvx54I6hUeHA0gMJE6MSg1KqqCZ63bs0R1KVogLswH0wZFXzLEFowi3h7l/LRE
+QEyKGAiXaAAcCz/AQKvlqpyxAjhcu4RMbdb7Fsg3Grbxe3cp0oBbMwhvKZ/X6D5PdLdxSw5kWIL
4AAZ36QSHwXgc3xEGiyYswCSBFXmtmoCLKMHa4IUjZWfuqqhJREmQKl1KkXpzGH+0wgU7Q9UZfwk
xkthz5NZKz5npQWBwAbQZRahX+ZfzWQ+vvFuVy3dMxKs6HrOZxpFXK+FD4o5Vo4Y4iaav9KU+mcR
icwZVcHBcRIDHGh1E9YK8mdX73tFqLoKvOIXqyDIPLySqhPa+YBKRtkQuL3VLi8NprNgQ1ujJ8yl
HC5VBrDrAE16oerudK0P6+mWuoLngeVCEQqh4fTXh3V8xGZXNWIpLpvkPIndCuVmy63W/JanuJcK
3NXrMPNU6L952fIW3DjnLi+4iWogl+g5OEguk1YenqqbYPd3h6hqx0axQ0rpBhpGGrTFA4g4k20z
bZIqCafrXc+swZ4uB+a016MRLxhvzy+KhCMG3W3ce1bGftUkWY5pSwqEg2Er9UTjV6Mgb5unShag
UqcJ6uelRGklIO+f8wsPSyNXNK5pVESfw6wZFYnNi1QVK6zw5nkIL9zFzVl1rVHOihBYjKRImpmn
MjbGj7hKy8KqfzzWmIFzTm5gD767wEOlIhbkGEZCB6EqvicCmjf+ZnAC8EYvBOPnKRwsI0a8PdPp
PNX73/NugNifC4lVF5cTIWst1yvNTOZWFGiFgOSXyu40NA3x4CXdqElO9J8pV8T/Udk+FPOmiXT2
8Zzk1gYebXA+SSHtVvZQTDfUxBEibWuYAS4mIpVxzPvFBqfeQpxXvoEK2q62XBqZKNzUJ9vE6nLV
fmJ/vY7cYJgRskboi4FRwaoe5SK7Ue9N1NdDROonVNxlJwv26cNroE6+xaAJuf4kaz/VdCI6DrFd
Kwd7BIgk4P5HeCYda2lLpeP8clX2P4Eo0VwK3yANqWMOjIsOdP7AL4qKMCRvsTl9sZW/OqeTiJmh
FhwEBdflxgjtaQ0B19R3rCnpMLfLGmr6AN6jd55fXJPUVqQldVU7ZnuT+hyVXh7wH45h2gkQUoi/
iGr5NKjoi8DqvLd8Dik4H15nVkKXCFNiQCIDgah3FYcC46BTrNrU7WhjttpgCYvNHB5Mqs2USN+/
3TAuOAH+xMMFwzr/dwDcS/EeIbjnKZKhl5DdJ7O8+un9jOzveaRDnolLf5hJXkba9sLwTfgetbAy
WjDxJmN6YX+GVDuOTMQHpGtInXJIa7ICD3Ay6zGW3Zo7SelxL6/LSrih2L1GYa09o6BPe1gFXU6e
5cJTniAfhtVFVbfBnFMvN5aoiCqghz4s2PGy4aKXMF8LkfdeKMvsnbYHTFgbuqmUoesVseiJr4dk
bIx8KNlwJtGHIBWYvqKOyr+ozhEww06UMo64HKD3dl1LECkyrhaxrO+8XfQaJQTb3qAfgDgcchnz
ELaz+zD4uTtkpcd1M9d1ZaCFnSk9CFk8lSr/jtS3JmNQsZMuOw2k9SIG6a7XH9C8NOp5PanO7S/q
WOmlWG8xBvcUVDEeJ/RbjVWaUAS2P7SFpBIm6uyRaWwqjJwLwg3XG4mxDA9SSZkvrZU/0ZMyJSs+
3o1ZX6c36R0WiqnpWBWNSkwWR/MvtNg1EpWkFPU2bZ/HLq7N5BaUGZFhX6KgCANhIkeiiqp8IKuk
g93RyLkq9/35LYfJi/hBsRBggwjFeUHO6jg9hgdvA6HbyHnqI0bnPGape3yVwDrk/IE9KZO48zp2
ftXJ3z3PI6YSDo1JE7CjVk78zt6WgfAJVf77d7hG7qYSHl49NjAuk2wBMWHcGrunUGq1B5wwFIn3
uqNf1Py+dkq2VtCgVYS+FUqZZYrW+p1zyiYT1YZsf1feBAgA7PHkhI/M+YBNruovMgv0fo2g6XKf
+t1EtRCdB5YuckJC5iAk80Hv3VcT6kWBpK0xXA5vJ27Yq3palle0xzcZxGanZ+BiHZ6tVSnI8wc0
DJ9XaNzp+uzhiu8VkkkRWH7V8Rjz0tdW7d17qTPQjt6lOagC92vin3jaLtxD1en7Os4AVck0aNrV
5GgjvibDStJb3qBhfIBHENcH7btcPFPigyPvY5czgXyE5kd1KCDh7bnsGIBP4PYVkspJGfS52Azj
jaXUsHE49/TLd7lKoLT7en1HE2m0WMMVpX0WatC3alruQpKnNRq1nswtnAXKb5hLEbyykewtRF3j
igDg+0FlylV+DFtvcRSDHcsms+dOtUc/Nv/8xw34zffw4m7Ntzi5osZweVIp32pwgesyJHDZ7jnm
DYVFvhGuXjiPXJSMMV4amIBGHW19IHcJp1v6VDMCLzpvGx1tfyrBXEwLXhSr4XL116OsupuBTnTb
wlJqwCr1WKQCuDx+TPPJMZL7+Weh4IB4fovrAMeU2O/2KKSXRXfrc0xJCtLXJJB5SKuJ6vJ5MtND
j8/0hUNNNXzEnggw5JAsktwctja5EPmnmXz95dxt2ApJww21DeDPE67kVdIp9LGtLN7mQaS66e98
FuQSyqtljOnf+m7vOKEFIkk1E9md6RTJD3Q08uEuaI87HqfiUy+Mkk4io6NLPsnXlSC/+GRY+ADW
DATm20qMnEWLfC4KbYLRmWg4oDurTS4VhrZJqAakb+YxtUB31PhBN9KcYgPpYGAoboN7WUIilOz0
NdWjN/qn7K60eDGy6Rv+/14NOidH6tUd/n4QZ38msvglxXUbwKAzvI3F523hsN49rsBkzY1ViJL5
H07RxlnvZGJUdcnSkyQvb5qdjI8A+jfLbF4WyYo11GUm19HToZtaJgdNvn62V68FKiC7vePHimDF
jygpS31/vzipDKOHimSLnqFSpbNFRHLOoOUbiKk4m0LEi9QSh9rWyfuTAz5qwjJ9JFmPHUqTwWDX
uKXATBjmgq8GsfcMc+f7W8jdcniSx5dKl44NUumic3I8RSG60DqvF72uxgPZs+zYN/uMd8C73A5C
HD0z5N2ImHf4QbOgT9h33/xE7vfcU3lW4AQmWNmlRHB7onwdSp1NlAQL8QdpU70aaOfmeRp4AFcf
sfgejoVL1MWR2/7pPc/TK/gkl4VdbfD2DOgX0FrQ0rSTAOoDypgcvHOFu+9VO/WSbXi81r1gawDp
3VIOEhTXa4FzFA82jaGjwMQeJbdJdmPWeXfgYgGsZ3M4tPD+asstHPgR2Sy3DELWbJhj1vcGXfYv
3BswysBVXn3BbxEnsPQhvhrLJDojwNzhVhHDZtuglti3WCG4+I5s8Gphjx6s6DgwJyIIQsR/zChT
zuyoo7jkRjCfY7s20Yk7AlXfq68PdZIgSqVSMw6qRFSyjn8xvWqKVhYkiwdtQGH94QJX+BYrcmYI
Z/noj+RF+cZ8GRhTeBUftpxWrEbD5+jnYQ6MdhvqdWcWbJutbd1G141rP4Mj2zQYfadYu3ivB3oy
hHiuO2HwZWOGtzXRatDpneK1F9Qvw6f+NYmadAELsOCh+wxyV7fito0RrfeXy6shWVtpyjZIkjFs
shU3BOTyensmclud/uR5pZpsFYRA6a9oQBWXfZB9orS2aoe+j4FlfAe9HLZ4pYrzVEvNIDRDmxhO
BnUpPd3aqB36sjdprWtmFrTCOGwNYndk4VUMTFi97Xq0H5W26Xz3dgzsm11LOrRQ5WaT+bTcbma5
dbRMQhtDlYHBBQyK42rpjV5JmAFLW7Zdn43c9saXgVesRMY3pYthNKehtgLGVLdRzFaAcJcbscrW
eE+TIFpB8HZElGH8jacnmIQHIfq+c5I1hrvBVOvbHd6CjkDQKQDCPUgmKXQaVA0e+kng1tLW/JJb
ko6bNbZfj32WF9TLC9UGmbHMLQhPUAipHIHnfI7Izd6R1Y55aY4o0IVgqHfUd3rKX0LcJbuypLbr
1Vn01oDJigIkCOUK5Hnc9Pw8bdT3lmZuRKRJ5fzYmRuFjCdTQeZEfKQ+m1ciqJwYpAnAONFHd0Zq
RRh5Z4fW77brY9K+eHQ/WMsqR0GD5rU/fnMHLlyQ+prM3Or4ZLgB3rip69Q8/tt4LQ+iB5Oz5pK1
dIinz7kTdOflcvNZgkmZ+m6TxN/kXMHm2YsE9y5iWJijHCCK6rqcnb6lLv7Cr0OrR+Pl19dF8nEf
qHSF4yx6gSkF1f/hNXw4fzK/fsBDz6h6DlSoC6FH0mVpPXwoxcsAVTB1/tv1HGmOm5AnORR3lX90
TVk+OANriseuozYW15yNnQvuFFbUG9WKsU9/+Lc6u+55WvtxP8BPKXhBMcSWWJR+pJWdwKNLyU6P
jJNaVStBE4lUFmHZCJJOwWs7YV0tPM0Ybu2TjO3JjalBxqBf9ppvUrZJvgQSdT2xUWLnkDP0ByaY
miaA6mKlkdSx202lVkzODnW4uQlxO5NVJPiid9noYq/6FjtAjNq3twEo5yuNKorkdWwu4uXdbswq
rBUGjW76ym7lJSmFRKTttbCUhQNdHmm7NYYXetyddCcchUu7zFe3iOGFIAg1CgvgjWL/4IaTamgm
J0ep1IN62/b8JkI6IThYDZN0lapa2/kkexMgpWrWjehBvImVqpDEJrtpS1uEngv2T+ZbJHR+GJsv
R4qIUfqr8A8jTbjhIhndXDSEi20TDRoNn/z/TGjD3BctRr384nobptPPzmgugXbcWAvDIf/D7N+l
ajuWEF2APuk07SqjSGGBYjg6xHL9Nvl4Iq0qFDyGhCozIN/7VI35tztSnaoKsWSi1/Lk5IKr/PeW
071fuk7PB7jrx1hpPSyjKaZm/liV4g+4V3Ab6yNcXAb1GSM0nR+6yiAr8SsaDURuh/0pw22aP56U
NBOI6pYyZQevWjsSWaroy7XKcS3zQyZ8g4YdBfha1m6aFGL7p2UaDxEDXb0YGgGgynzT0ZkL7hSP
XDVUZtiirfN4ppvt+Q/5Pric9ytDj6HHJU3Zn110E15QoAeu5TRz1Z8WzqyEbpHu/sc2GQptQ9tb
kUUN7p48AdpXqse4MOnqSM9eWaN3imTHB+c9IijYb++MiFrcFfw7Gfi/RSg2MAIbC6s0vvxd8m8w
K+SenbqPIkik78HJaI/gcpIJWN9k8zKr0xbptrmxuPUBuC4vq0MdhIiUG21xZuFMlllI4U8L81Xy
+og5XP/X0mTuyoPThS/yT1lYMTsdII1EYQbY4PngnWLPduG7cesqCgbqhjQ9o58qFPw4P295H4nl
SoC5kwxHwRhnLIGcXObiEjJAm71Bsqmd9IMckLcKHv1q82Izf/RW2azPJyv+532HUlDBVeoMQtJo
qzp0Yivie8X2K0kXDpjQSvEjV4Nanqb1iD10B3UmTDS/FPY5Yw3OjlrxsjaggY5Uv0AgfcZo/M63
zGFiNdnvv9hV75I+4N1sRTzJAD1Df9qG2Hb5L5ohARwDgmbNnPqfJkNeaOuVl8r/cOmATqGShu82
4eo+wWX1FzRgKyppurBo8PrUDAaTithZk55zC6VDscRAPkdoXbMZ4HXx8USzDL23gwjPKnPwpipK
KTIvRwx3CtgbXapjnHV+z/ILNXtp+pfrzHMvQxULIt09fpEzcyTCVP/8rAM9pLBYk8ukxQieMdvD
RXVXF+4Mz+8pO2VnwmHFWj17QK8G2KXY1EuE6bEO9sDKhEN6x9tOjO4LMNR35y41kyuX+WnqYi5t
gZPKloek/huiShaJP8RHx5WKUYnWSDMS94VKaxGX9HRn/urtS77ntqQI1NFS7zz0wmFX7xB+3rkT
tua6NYDKnq6kGfORw7pwyo/D/3aO40ucaq9E8+MVGzHpDHsfhzgQmRxeOK7NMS0qYAONnWqstYZ7
Q8uX8oYgVpg2LboPp1YTMEhrqGZpl93R3Jjg1L9V59N1rkSwxeMrXfJTJiikZSmrHtbaonWgkvPU
brLyFsVZ1pMX0ylw6C7ZiqttY6lhGBVHjez3hewqKXj2XpLN9XgyxQgxtUnSeQgg3SGYEh1U3ugM
B1S9SAmZwyb29sAKf8aSZcHZqARSAyFfzQ4chspRw9476dGycUAyRX9khm90oFiyiOlxmRojVURK
PMDeD5QRmfPPyPN2c73556qVBDP+o9HeIsLPGZogJaZGajRpecPkABpoPXrhHp2k5eEDRnHgRdfR
efTeZ+wod147j8cyuszZZXoXlKT3OAMqWnvgsDnSFy8EDbiDJ5y5XVEF7MXNhjfXlIyGhYZo13Ec
x9chqRcdLC5U/bKz3QfKVW0nn9vVNFZGn92vCf56TpI07bU3L/QJGr4jvBP+XzjMRbWd1YpHsemU
Fg2/PNgnTm7gC4G7G/j+b6Q7E01weZcy1zebJhmm8djtpGvObdIfgSNBvwNiA7puX1f/engnvBnk
ue/Bw7gAKBg11GIbDqofQylT1cia16MlpBbhZis8joYPPOmcfdqHQKNrGqzfHig+8YP/vKCxs+mb
N74fAos69eRqy1WBSABzf0FaOHp0tlhKFugTdN/aomTBH/NudZfO9riLxFrgSk37cqjksmNzEDoM
ibk9V4dM47CKEbkXa71e3hTuaPyDLr6GXlIc2l+U80yABDqbhJVPHA80evtnKAzVKMr0aH3FbQXT
plDvH3nXvkPz5QLpuQw0kAxKO/KGdM5VYKp2J1/ksdVU5cgsZSeaeblMufkH5oJINAvP/rWBuwPR
mvHnt70wHI0GPaNibfVTwevYozJcF+qksese8Xn2sxBTM2ug+s0fPwH4g4YJUU+wEfg5PZ07A0lD
L4EPYdkACrATv0IabyfApacuO3mnqvvL4j0ql+ePnOGRbJE6x26VOXiokMUBIDtOCVTfFTdP4g1L
2972XRE7xcakiO11zXwHAOpu3YMhS/Ve6Kxv7PC11oPjU7XPrzFDIHTLHUIJwfGxzRhMUEUDhaV/
yFpLMkTLnHJxjYUdFPzABui+Ved1A13LNCgrLEk9SJXlPVxnKcUSAHOEQGORZ0OaWVJAAWjY06+0
v40ey8lvhVF4foaZRewVhRu4+p/Tb4jmmdSc4Uc9NBr5tiL6gHRDK5BGhq7gI55n+2xK7HQiqW9f
gBzSPzlWQcVahCpHb6R/0CcGkeYcy8UhqAJSUIZ0AlDaxYigFG+pArMBQMjlCqxYdi2r5Gy/6Trd
6yMnH4rQ7MfiwXvIYqKt4NHVnLbk4MhgDNnr/PE+WJTpIhwmDdLVuO6HGgNcJGUxCdhq2oi8iWTh
Bp5v7RjISMh39eKsRn/R3RWXjgNdNOAB2Hr3j/+MEaktYUnED14QSQ7kL9NA0NmA+J/SX8q/uyR7
neF7aQmdrmYQZQnD/+untwLAlzg21HxIA6pt0hYXhc9v/jYXr7eOl3ntOQU8EpJuRRibBz93PC5v
9Txe60QT76aUKfvRXxWc034SJiAe/IiakzvTmbAXLvlOF+QvszxMbk/9woshdqSDMOQRM/pe+/mU
oMkoDYCqq1CbNYockZiEn77QEqxo55/icthXu4CoccXNTDKJdFq8o5CCJN7t3iFIUezcQkK6rz5y
v7Cnq2Euoak8uQoDrLKvdPLzMyLy/UizDUVGXC9UI0V3fKEE+PYcMaswkKy4YuOTxmjzTJHjQN5v
m4lRU3RP6zdFjmbVNepJl/KH84LOSVWInGUhjAywpwSnYwdDMwbaVFnm0c+WoNIpsdwptXm60U+0
OfWMqdzl2DpM+/qjKqwaXpjrXKAKQqO2vx/YMsqvRZ4Tg9pURdO0qVBffcRok0zqQqTy8M4631p+
h+xgCrVss6hyvLvUv9gpNcaComY1OA4eql/eo6TAsYq+4H6ialb2l3uHh8YDcwisCt0aeIzcwuXT
XB1h1068PU5ABwYby+VXNUrbvYnlILlELssbLt2x7P/K9+TmTAb4fWjbh78BSoo/qMze/oCNDL4u
t+o0MM6IuwAXwpemSPxdOJQNVjG2os/eqy7R1fY9Zes63AwZmBfqPmsQXYfU3xmM9PtytghFdcgo
tey/6FBsi75q2CLUamKsflnhN4rbFQl767k9Mo3ulrqRopGdoeL1xKBSLkrqWM5ukLlfCsLRe0IM
PAa08BfNPXt9sW394tDA9dLOAfAo4kC+c19cQKQJjNMkv3251dti0U4F60eFs/WvKb7nY9kUGtmX
kUYznTjXzgwR4XZGDUKf5t6Vs1XuARsDpZ2tzY5gZ7L11KBDCOtOXLzQ7QRqvl6StICDsJ9EmBEu
objoNTWOyN3SAH7w0KmcXueUodESYBgRZXkE/LxwXu9JaqK3TReZv/2kjRcR5fpP3fREk/HlwMsq
e7ASEUH7IArDHVgk0mPSrxCNulmsZupI2NJK/U5w0ePhRc56expiLHJzQsusGSDRZOuUyVDxomMc
lPNWxxxHzHlEwft3eG6mcmFGNij4wqpW1L1Y9aPuBimUAyApml66B3S7/drzu6OYeLJVwUEHKQjX
ixlEpTBhlq4FyveuKgj2MAym6PzKxXk07BZXJNiNMLhbwwZqkiInSgDYaoV+CUbXAieSZOYwVZWK
klEzEcfs28P9k1+p8jsB2XBJGOyFGQEUcwgsoOh32Agqp6XfbB5YBze8JOy27jg+ge49y9k4EEov
euokAAdCZnLCFAaipdAZaLKgi2fpmXr2Kh99bIqGx2Y1KcFs/680nZTBTY48IG9YCSOBmUt/8xXm
LtSUJZQMpjLpdPwbKLYXPAlBcCk75+OZF06bE3j0mWf8UB6A00o8lLsoycCOOqVBU2YRu8WIvA+f
eVnBiPuo/hog16EIP8DDDHtUvcCMIqmTLwedoLMpRYcvGnbyuaL/WxvPm25j0W0XbkEKIt5N5O4b
+Wo1HlWSG6hrEOwBacBlTw6zoT+Ije4qUtNIkYSH60UzbwL3EUP7PwHgmvP0GqIkIVKjofDLiKSp
Z+fEczwQuQY9mJG6AEq2PmdwswMBnn5wLlzKLts6YZfRZOlX0sIZKWUAxXKPQ+Eqo5Q/gymItDRq
hvmb6fX6DYHhEhb6du/MTUM8YGC3BDGHm5Ok3RorHz6wJhnuxMsrPLNdjFiTcS75Ig7CecHpLwqY
rAWvkY6BXvs8theE9rJK+zzSM8lXSJAe+Lo/GIjNNLrw2KyJ5hnrkrM1fitD4M66vUBToTgKxw4C
50wZ//+EUIDHaLZba5sArO/jwK+zsKZyHVpU31MyFuqfc8u80uyu/N3lQV/Yf6WE6Jtn+qoaffOE
2XpOHomw/s5fNiM5wsRRSaW1197xhqxnLZN3Dhql3U8wpCuQsTQkfdwQ/Yv0aIKVWXbr/Ksbu2xh
UZMWwtl4DWR+JnZ3/RpNjzm6mNPRpR8BYfFq45G5RQvDHrg82gwUVgmVuwwapVlKxQKajEfWPNtE
Imr0XN/ivEaWo6Jrdf6bdbW+YAT7TaTQjGX6uuq9mDKcxxRmxb41/x/71z6/bA7G+iGlE5Hktqz1
zNFsD5cHywOI/F6/gIM+G4ePgf4R4XEMxyKUFuPmZKmWFGeWV0yNZQ5VXcP85MJGvrijJtLTuub4
x+/z9In72W9lYJiFnJYrp/2+UihHzbp6WGPZNtjkqlXKl96lfLjnR3KqlQKUOANIbYoX6YsL/Nwx
GvfKA0FohnWRFQslCZcRgife+8MyoaT69OZzsQvB+PUIVsaB4wwzI75Ma67LzdV9FrW8oIv8fUrp
VYIDkco438xjwFZTzJi+69QeY+I5B7SVVWI9z0eDIal7fFra1c22RkEDm6k2hi1Q0eEosXDNEgTh
nvrclT8KRqta2tvIOaF7lHSmcx3NM1EAQlBFG+uypYFuTCGumTH6e4N+mlm4i/PvGDPHSeLAYsoP
3x8f8s4TUuEa2xQX+IiLa9MjOgX0v23/77SzFuSmDZ0S0NljBghKmg2FD1r7uJMtaLH6mFlbtS7p
A8dA+y80DOpQWSm6qHjgS22R+//LgvnYdZFVJzMq96sXmdMWfnHfHd6R+1XA3GdcrXHmSE3c3C7s
w6h/Zmk3buRKZ9jKrllV2Yzzw9LujNIWvVQKp1mjjOZSb7oD67iJTktaw82aOJd+P45wvw7H670h
z4uNIgOadvriS2niB+J+APJ9wT9DZLsyRYN1LMhju1AssRJYmG6p7FFCYXuhuiqQV9RX4RXMzaLN
RmAtThHDeFGDJdI1D2LEBj34jZ4AolRmHmB7s4Pxzwq+obJhNClX4S9m7z+zVP+5sA+o2MDPnSKt
HEICbqPBhoG+c1Ot23ufs32UHoDa+XnYt5Uu/titgDXFzlTpRyDE5G6rpANrIeTdGCd65X+ydzVv
cJoNgF1TYoWHJEvCvHByxc1cgelMaHtKs0itaGhti0cmI2KtiLUHbPhlTzhGkmPUaFl0xjGtstPd
vNsXcUOicy0F/Co/peTnSwwsbNJuvfqWvLmfOiTQ6qAIokmn6zMabBrn+/07BZZAziUdbruWU0S8
QloUdYjOcU932/01M3MtzcLZg1tT4NGAxEicjDGhKAHqCjIA8DZcMhyU87ghiQUn7dXvgFLQPalN
+QYbsbS5ls9TXCMV0NRlAk06lmR5Aad/GlTdbwC2vkyCnS2pEAGQoyp/VWfBgxd5RcEiTP/KRGWP
h0nSFzH2OluxCEUSlBGy4M2whqz/hQUY6cYvma1t4q35rDEBRPZFar+b4n0zyWkL2GgoLmEyDVE1
1XlBLFmv5hHPVLPvmyhlwu1qBl61/kL+mjO+Y1mb7mxjZb9wJIwrCRFiXoUL7Slqx27GxXH/qUHq
Xrz44D2R3qTj6ifeUk4fFd14yVBe52QAUiUX5Fg6WWXHJAkwIyhUb2pxAd808gxddByTEoXyvc3a
VL81aCfKTbq84Sp0b7iHaPCQ+bjoPzYAQzrM+aWpJijo2FRBLebQIVFy8tmESZyjFvpgtu0kUKS3
vk7KsJggv4lscZJdxDFHN0VJq9oTVszeqo22HHDqR4h+UB5jCqCmwaNa1qrlseg7vl5g9GJZa6Or
A/th4r2/99DWmB8e9QbkJpwzcTPO0z0CxgYBId6LULGyuvy+9txHV7V7d+/o37IReAfpnorZKF3s
JYyBO2AyBiKEXgKfEY+wem6DITJepQv2nVuqPGDukSVNq95XemJU2SCq/cKLVrmHnRiAIZxNCwTJ
JcFDX2hV6U9jzQfg/CO14kypLSEb4M623IoE7Q81MICVQzDivbYryEcVTItw0xM7tJgcqNSsCxzp
1lTM5PDdSwqjr2qD0zGT3wsTX+DLXj6o5QBGZpY+Y8lN/u8m4xl1Db5mk8SlZiaOuTxMIl/R20PE
cTOv5cuNH9yS4n37t3rDbw/rAEgqkpQRcWoU6YP1a3gItjIhCB1Upfii+qgXB/BpG2q1cj26zWQe
Pda8tW+DiWMpTZzj5L349rFC9m754fS0twikT9IuleIT7adjm3gcqwsc47vSlns8Yustd+2uwe76
kHku6KOSVQVo4UI03LCK7Vmv+Q4XZdgnkbw+p8Y6LXdxT1YenxNUavgKHYQ+AhiIBRTixm0zovut
6X2OKtSb07kclmeLdvjoxZ+SJituQs1XX8D1aRcZClu350wpHhuJbWmPYkDPzi/PjdR2FHxgwEgy
zp3cChjuIDc8WW0NLX5MDm+uqsfXEI65Wd6L6gFqg+AnA4xqfQmkglaSsTpVzm9ha7AGklsgARPU
YL7/FkIjeW9RcjvwYACR6ViIVcN0L2W4z3KXTbgqzuKtlaKQZxNmGjMviK+lsSE2ACkZqNGUWk9M
XTWlnVIF1BdNwuOVVcO0a2oXdJsIdcK+VZBT755HchctdyC7zgm/l+NZ7uCTAQhV+FSNbMbpYelg
ZLkuFU9U2rSMzjjaKlt68M/SNIH2bg/gQiWSB8SQ7u4biaRbbmW8JNmZC37uPcudh4esapjcoY++
aMlfHdOG2FONm5UW30hF47+CZPZPBUPkH53l8lrbYe11PK9WwZ95XJkNi7RkUZSsqIFpjfK94tXW
uSns2NlUcw6k06RnCsMiZjXUrw4OFg6Hfwhh8e12vcx33FBqATMMSJeophYI3doBVtAUS0jf6lbS
e8TpyQ9K89A1ZWuyJ1QiZ3nzBBN03x8aY+osPBXRTnZUtIGKUlTPTTCwSdQXqyP2mgSB30kWPbDi
k9a7tj0rfleFWKoJ/2aujm8S60VIxq06j4ooxTVQERnlS4ty12kcGDSJSV5lmGUx6SpDSEzHnHVR
3Dv6Nv1QEW9czQLm/VagPvtK8IJgCyC7B6ZT1AeEgi2cIpJKfX+8IcWT5vrJEf20gEQHDJR1Ubuu
6u0NMSKmEV0t+Iyb5TkzrdHFdt0zmzEG4zwqpJbCOaJJWFIY+HEfDRtXlso+kpVnMkGuXZ4Eg5IQ
qLAUDeJr+y1F6S1XXAcItsDzzX63FjdiMeHGirUYLp3IsnpzkW9+6gCuleh2FQC2hvz62Al7vGH+
pV1lzWf4UbLdb8CerDYm8MPdaS0M2HQxbQiK2MB+RJekTrokucX9CejYeXri6NFnzxUlbr1HbYCU
Yn1MLM4VXqdz8oNpMQ52UwTn3ivv4aZzRYlJ6V+8ytsolErBJvPnAkZxlfCA5LHGfxS+4wHBGqSD
rgbw3EfgdYHbdgdEht6FMbO4HCC+c4ICyOOtvrDTSm20TxTLDrDcVStFHYQVgDtC233TImsDfEE0
uc9WBDmt2RVxtK8Qctb1wUrE/bFXKQmyAcdmK+k+KL+ENcM977RAX5VByvp3+0mJ4P4lKKcIBYAM
uwLGfKODhn1Vz3r85pBHA2k6cwsQCnocieIaf4zSaZJ0ksPxZLxmhOb+0ENIcg2wTQ1wyonB89d/
haIvWB//hzvzEdD59FKHMhb8aTN+vqenW4qrqewfbqrdFio1NAZ+O0n8xOE9ZRk5W97zxxalifje
4PJqnmKG7oVPpGS9eYTm7ONWJPwxL9QWSTISQAOWvxmKagblbIqSU7eL042Di8IotZwfpEMHIK82
usrT/sSTd5LwooZJoVz2CGzLR8CVSTXZONCrnP8CQsOG+6TeIN70sY4Zu0vrjZfCI20Qx4CkPIHE
o04mdc+QPvLXWKVC5t0B4rL3rNYNgIrwY6wVx7e9fdhFzYHRpNVvcTlEEFaeZbDoQg+EAHsdWP89
QYTdr3e78KyZFD4a/+6oWwDpxwsVbk/Nwa4dr/jesaS8yI+EEE/Re4pgkCVw3KXYt2ly2YFXtZJ8
NmGZjCk1UCeSqgx8BBQ9i0VRPxc/63Pau3fS9pdCt74sa5hcfE/k0rK3TVmGmiNwUgbkUrgfN9QU
MlD0kx393az3FVScETjWSPGOcmkAns1yfDHirnMTYV0sUBotSj9UH1PhmjGp3LeGWEo3IOekZ2oz
jRmkC+0ia4DMPXW55yK7g/ixx9AbHGb0P1XGU/Fg5fYa1/lorpka/smGJLK7C9vVgEPB5cKvuVGD
j+mntSGhS7DQ1bNpP9RqHBaZuMZk3yeVvG3OxwGDzoqncJ71AfQcRe49fui533reezfBh9QjDCio
BLpXOKKaXNL/nMYwg5/DB6gLVllvGUvDHjwmikYuULIyh/zvotN+gjpzo3VD9sRwmDEy2bDlhplN
j5dumbqjXIbRIkjDwyedcbXP1e/yCduHABmwtLKkRMVzeBxqYoOvHUEVS/1aocbPZmJ1KRI2vTO6
XV5iLGuJeLL0QROrpkNmWc6uy0swW06erAmYXw5Fq9MIHTEegMMo2bL+xvcWoZXFfCv+x1mhEs38
X2FrzfL6U9aTx1LaBgN9WQlWncf3cj0PzyhwFHjCNPuEQHwKMv8kRyLRh9p0j+7JMTBMEakK8i1x
uCJpxt34JQYOYERGxIiuVTb8wGuLyi3b9BeFVXydwZJqJxfRlbIs4vyuR7LlLBzVRMuuLavRuXnT
r602ECazno7OSxWUDz1MKP79Qk+6JAsQf8kGTOtYeXtxMZnQ1FSa8r4wr6weRABAwEiYtID2cC82
Kvzt/GbmvDxj94bzAp3deSJ2+OarT8vBpaAeYhJcVypN7RjstWRTkVh041+Pa+RvdiQxZvrgbSfO
p9ZLk2f9FedjDjJKMLi3CHhETmgErPbcY81lqxQb/1xhv3zYtACCDQR2P5WZEoplVG4kFL39F+tV
7/RnylQFuonda//Nzml/WDPCKn4gRuWOiWNqTCFV3MX7hschIQGMWoObriKvdfQqv4iBzjBSQNXq
NaGYmQjc6kwKtwEn/ucH2gN4iXOsVBP/MyOZl+CB2xya7q73O7wQgInggw16pZgoPqYX2r7FcapN
NeD2BUoejE3Rn/iqTdKTQMNxZzC5lWGU03J/+6m76z1rfbVA3yYCWB+Zenb58gvox54JWUgL1Hwo
KZqiDPhqpOLyIRGIW0vPTjp94+WbUbZobzBzSUb4Q1+gBNjJkDjWRBcobN2H8kNYpGlDO0bLmIab
a7msjapKINHvDePLb0Dyo0YpYw2ngTa4JtiwG9+9QW+fezDUyCQ1e+eck2pB58+8s32FVgIZCKwG
DvG1FQ5RQBR1Xk3lx3CDMixIlWZAN3Qjb88drPvKC0wkzqWN9vULWHYQXnlCWrrdjq9FPGuNLTcs
gg4GXrWKvTsxC9Qk9km4g/e2J6v1thMMkp/nG9yX6HB8SAo0UCcJUAIGHffGZ4qkvMFS03ETHEtc
oleg9A6T4J834am3FUPLLFoTHhv+b54etpMPpgEGdCtlToiloIc9ANuElvnRr4FQUQfWn8JIxn54
AF6pIVaA2um6fsUw7ee0euQkFDpvVljIbH//OQS7jScmZwZ3bs1Pv8pqGNhrP8cBQV3C9WQjDqLl
CUruDXj8qykqAu/oi0UnYJZ/fBx5D4SVbJKAidojJQhqB4VaKh7VTJfToafpsZdxNZjSKLrW/2Id
aYQShev4pw/VW7oK7TnkxccJwNP5OE7/3mxJrQP5uBHou1ARP/r8mN8ZPxR+ri6/rhUeo2fALXAe
zN6OuD6DRtoqsEHMO/8S4mBwXGW6T5wnwpEs5/eYDcCHQpavcu/4tp3dLI3vQD1a7k5l34zsrpvJ
4X2C1QvT7J1w8Uug8JpBY9wUPQI3/eUofE8nEll2jQHU1cNJwNDxBxXDLAQ9FRkH57I00ohcIVOi
/0k0H6Hen74+p7mW67a9nUC4rbgAdI8rP/nU2WYYyPrftgl6btDI0Jowfm5kENwgQX3KtoyxBiPV
vpgMajOmohiEkr8Kg7a24mrkhTE0XganmHv4bffLy/nhT8dj/xkq5u6FrbF9rAHNWSnjSiR7TGXn
Ko6QD+gF47Au9WECXjseSDuKtT01eIcbaHQcJraq06q6en5dNBWeFsu12Io85pxNgX05HxMiz7kI
T8VqKcGwSjxgJaxbIwlvZRdq8KCM77zNKlqiCOoQQNaMtR3jy+gwIOmCoZkkFpX4XP7ODEcjM2yw
pohVCNi+5K3nKz9461qUf+no558HxeOyw+CGfNHNuGcYRL3cLDB5CAMjU1MzFpTfzW7oVsfCfS64
iA87QycrgqbQLHzIQ3RcvnmxgbIXg2YmSwNON1QxjseHXePM/ghaWHnK2K8h4wZnsCL1Yu8K1ljw
8DWlgL8TaXvABOkH0g/6WR21c/GH7Jd0NkjkkFEnjiCSUQNfzG2X0aftZ4ncukfpqAexWXTN78Yc
ivjSK80sJ/llXzynqt/7IUEdHBog6cIfcETal52YPyKTEe/UCTr+YN1tZDNQk9aVYbWRMwNFCC6D
emzAzQQfDKBewUjgy14jTNOYvh7mYq/SxapqDeP1G3V4Xcuh8HxTY3yzfauNJOxVz6knW+4SHJGJ
YOg/0BKos01ns1gcrgfrZ4McIqFBQgbmhq5MoADRXndEZLPJKqXwAStRAITTgmeuiAg/yT1LrGV5
AcwM/WoO/9xPYKEr2MvbyqAJnASRmd9OZ5QORPue/PSXXZxGF/oEYlNvPD+9Ez+oRWg0O3G7EMIM
Wng02XcQgsNAfmDQGQIDcSX0HcsNbax16cZT+It5yUGx9pHESmlDvgd/jjrPO1VsvhTxKpy+Z9qL
oRDr+fBaSaD2LjpMjOMGSjOimO40vjPClRhLIlurexgSdNL0zLHcC3NRUp5tJHIdZzCxnHYmmqw3
+yJ4skEeB1+Sq4oruhLPaa+Z3Rq4M+b8jnSveIroBLtqEO16nVN8rcm/PcxpZoLzu41xjb1GIlwR
kW68BuEQ4BFPvW1yM37xXVhur1iYRQ8o3F++revPx4FR+vp+AjRn6pOL5IHdlwcSVjM3wl50uaVv
+QPS3OLasG8FR7xKpxVQLU8SY3Mw/R5t+LumyoGYGarXgTnseeDcASZeGxS1DQRUpoiskTLg9X1T
mBuVpLFFWSVWAiHK90SnxHMtvRAGoLam4P/cCAqM9KXneQqQ16GAOKvMLVsnhLpZ9f7cn3dgv+lA
srYuRs+Hp8mXkvEr384TLHEY8JOF5OxEz5ANY2uUuSxKguAitIM4DrklqLWHTgoyu+NjcgXNT9o7
1BJP+74js2baHiK4RbA1obKaph3jmKMW35mCkEc6moBS58MRvHbSWsYj+JoQF3kiC8h7Ellsoidk
EJT4swraonQNi6W7VvSdL7K5e8VKJWoaxAH79S8wrtTKGyQ2uvIpHuWHbZXgSMR9g2oEQqPE8Fei
GajxeK13MSIohK+0zMch8UKqJ2YMvSNnPYf7wLvTk8aVXTyLaiyNyrmyAO6ACODFP5HGcoCmg+LK
fy9ZycXEywnwFM60CG07znERq5H+p5nFGBl38D+qDnPF6obt/UxaEutIGvE1dgCJI6DWUSr7J74W
FePBfMFEhobipPOfccGvISow+QfF2l9MOh/NPmx7m26RYqqRDGUqvcRBEAitdHDAaNGV/qmVljsG
hxJowPo01Y1MGqGlys/+Cefb4Z3m0DrvAOfBs9nCh0J39cGM2HQKhad1oBS568M8nheZIZ3iMrtY
RnXueFRHeF69UbGBCPX5f4cBGknopMIeDB/j/9KLHZgI67OBNPwD7A8X3gNve/ylZ+a5EUpxLX7V
KRQI2fp3p8QXV8DD3AcxWj4nStbJe81WEWGMaXM1XqKZXlpZSD8unlDNiRziG9mDYMN+PA7+tCGJ
X8rcuWza31xLsZL4hT4UOoj8q/C/JSAlbr2r+7NrtJE7Rg/FBvDQRz8rCx11uAz2sIh9V9m8kzHe
KvCHi1SB3gHIuAhJax8iokVNgVjdRpLrKJ1RimwqysYaw5wA2m/wCYQLZwwFRJZZp0YsHeAoJGrh
CPtrRb8H5Gqe+EzWQybWehchXCt5gh9YKNKl/DqnUXVb6SxmeeutlPtC7d2o+rSQghkKgYyFU1lW
9XUisO+2rOp0eo6VWAVzYMtNmoSHYGe06vmc+4VMZkHPD3fPx+/6I9DoPVvMc9KiydkInhLMJpSW
3d9mb/tyV9Mx1mesrzASgp6fFFryk6Mu62yKZJ+3/9RfviYuxhQJmIx/twyHgbYzi6U5OQmonZx9
NgV56hvsCr9KExOywNhntR6gosI/S9ZapkdfibvlDwtl7zN8oGfyWAqEE9gehUJZwQ6gjuXWLQ16
4KAnXxQ2E4YrQsgEjbbJHNLHVqpffKq3VTQi592XyiLC5h8XaxulwZCqH1JFinRELiuNkwELufcT
DvJCvS1H4aZ1hyV3UskQJuKqgt/oIC0+U3cua8fOQaVtE6riBDXglBO96xw0TCVrS0jHUM4XhO4w
hRs4pNkmBfda9RTrJzm13YoORQKtiZx7Q32pHFhAE7HmBjvDP8edDqo+KhoPhRBTBSjak955yFBH
yZteLZD9t51HNDWWn25mtWzWDyb45AZ1JIv7+pTC7PvQ3YEAhrTa1FRFGrvLa/dF7Cabj/wq2zOH
N2ezWZ/1MXd53q/P4a8KAWg6r9G7val/McJdN3LxCutfmYJImZ5MKdn+IHJSeWHNNGb0iJlNye34
b1UhNju6QfEL+2oLBYAbwoZ9PYjGY93CmIl9HlW8nWsVHNIwAHt/Alum9AD3IiqV7UkvDWh8f/KF
Dwh+qah6uBa7I/+gH9RVX886vd3RlWcspx7tM7+dSzcuhggMEbGNQi6ZHNBIbgXrFtx+pAhofXI+
QsAh5tO4HHkJk92so199big2i5RBxBQa40Nj3kysTVxnXaq2gi8RLpKSRJQIknfKXhDRj07kRe0X
OX1auweJZGDWoPUHflmEmdUZUNUd4+xwvi+QgoKncZJw2Pvz+nbD1Tu1hs0RtRkot1so5xsYgb8b
adBAZtSZmNUI93CFs9yqGzq5lvKJ1ZpNzJbGks7wEDlB71cPCIXuw44zMyOzMsnK50NPXJ9AI6Nh
2rUr1e94GeOv1CH3GUZ7Zp8rYQXD1HU9SAOZXIsimIYUI4uOYimXATFSyx1CWoFZldnvSDWnjSyf
jvJ1+x6NbuYW6qEVSrIHi72p411ibiZgxCrCoGK/SPEfIRuMYw4KuehCIBFzqFRCphb/kXnaUcg9
dDtDTeE3yVJHcR+pGk1NCbP6FUQ8DsCUD3pNRC4SVEi+cURuPMOAgns2SOROKYfGFeUrd3Tx/zMS
X1FxIarJgMk3rahZWHYKvj0RhkEW0vEcMB45rh9fTzypmh/tv6tFo74e9dHz3ZQTIIqUAh4LxKCJ
U0a3kn0SGnJKnzEyAEctjMoJGAUhH78K8KWAQc+grmffl3itdOeWf1TN1JeeGh67GsKDkY9l9vC5
FbJMg5auGvFH0ZOQCYWINBjau6SxNLdceRZPInLs9IlUfzFxAnSKEAI/z38BZTe1GRXCSnZy/Tuv
14sVsmnbPK2HffADCVfV+4AQXlg6xyqp4RGuiTfJaAJIhKjhF2Hfnjly0AvlUlBGm2HrrJKIKJUD
8e9MHi4TzUzmJbEpAQV+zHkBXFe3Ex7X1bC7ObNTvJOywoay5FysdncLXKOL3BqYu6WqDVHczASh
4A2EMKZhuKQ0EJNUIu7vZWaab1WwpcPX1ycjEd7VAzd0qq1oEK4QU3qIL9b3hZH3nheL1Pt3iJ3y
lTvO/hDBopvrfni0V8J2cAmjfcDKIZl3TlvpfcAhPwwiO3HudBTjmND22CfhbkVXFFzn3g2FcxGz
lvtFJ14LxMGt4VgAeUtcHNg3hHH+3CfgvJ99s6Qcl9AupSzqfOO8jLQxeAW37A6peyJ5HlQw3/ZL
V7mRXqI4llUvnxUo1MuVPGkZfqt+ep8UrsqBdy7sGwR5+sawcSTsa5plX4yU43WOAkTcoyH3jSmm
wCZPTuQJiiVEHuJCaXj0GSK/TwI1EsuIALL2hKc2xYC90zNrklCFanDNas0BVoNl41KsQT/ue90P
IJ/cUkkxnSp7EX7pjZIg9nVHMaz/1hA5ousOzxsVFnLiNFYdYL33y7GjtwQDBQJNKKv7TdSjG1oT
JjNXHjwLssgJ4WZ+bbTvCgi8blEGT37arDtfdyHi9hPSLZblTy8iUhcTyFIcyRLRkPTv54hK30eC
O2Y2Bo8TATrM93+mCQ6724LYSLzU1f+cIDMYnW/LUPo0orRKShczG/tpx4ArJje8ypW9UsfHLPpc
lRIYwYBhP4AifVbgAth8s+3V+2MM+SvJNfwvblrwGI/Vd/r/4IABEb8PnyykgSzE8o/aTM4LvM2s
5RAMgk5CGbKqs1LRXUQz1UZef5FEufSE0q40hvqBvghRpRbB4MFvXL29gv0ofxO9HgptSGYtdyuM
Q64+Uo34TCp9o4vMZp0LBnXTT354tSIriIenC7nP7qdPsUv4FJazPeu7pL8PdsWL9nPvuc0M83N2
Smn6/mM2GgsYfcaZesK0j1FTuOPIykfL3UFvdUhbW/n9jk6DPp35Ju7s5WYvbfkGXxPC9Wn73ZKl
3TZ8vyhRruoGjGRmTudGnlKSR0RRwGCVYzQ3aqETxxCkbxG5uRu6xhKjLrjYblp0qcihs3UUOKba
MnWNMyLUbSFOYt5QW5blsz3VVV5TpDLoaHq9rmMBtS1OnuTWaTMa0BxH0QwfImGfa6RwIbY4hTXN
83CpuOGb9M9zN2IM+cxD1b1KvB1XNX7/4rN0Y6uetm0oNNiE8JkjoImab5sakvog9lNrtaw0m95k
YCH60lL4nw3ZP65atT9J9/tRV6/3vPRm3D2AxaIv+BDt2Yb+epL1PoEf+cXqY8cV+r39CXvcJMEP
4vXInMBjsdmh/ZOCquRo9wf92PtLMQFoZwo7ZGjoMxn2td1uNcJvUK88xB+Y/JCv8QMeXZFwWgV7
zbg2GStNFVKb5tUJhlcBjYB8aI3xFh+/iRtLQFj+MpZ0bce1fyj8M0C5SNmW8dWJsYnoA6YESX4G
DQOF5UP35ZTIexPvlHZt/kwQB4wD9ZY2l2omPJPn66pFqEGGj1R38m+xJs8E17aIMzXofu6hGxWr
07jO4JyqZKsbLwX69QPV6av2FwqQJzvjdxIRDonYJqCK8Z63uGtvv5WqP4I1t8QKfXxazGU+VzQv
adtBFDlwkxkZL5eR5+Bkhdi5UTQvZmWg16EqZdqEXmejUUTBoufYpW5eQFf/nqxNN7/MZnWI5cpE
Xybjf6Zag3lRkYaw3PPnPr6lTBwWFq1TMJSHq8H8FIHa3iMKHCSgRVXRjiE1v7CM0z/By5komDHB
sY2OWO7k3M2UhnlzkZayJzw49nOzvkA3LjSvLKchFwQeNQEtrcsiByX/Qrp8xF07ZiyO7bAYzl7E
kSEclQ5af7LMcvFNKRohtrewHvQeCZjQIXBC68DbwnVXVYQO0ZWny53rvX71VpsztcgQKxqTlT+d
IqoqFifY/EGD1Y7Soy+abtYgztE4mPFOS5AvvFj1elODBPV8jKUzJ6eHCPp4e8tap1TF0AXTwNzG
Wr74kXSinl6qtORMnycxAh/07/Y6jrVm1A7Ii37rCgA3ka3OGFF9eLQQQDHmBGF7pPGhG/HLBdTo
zA4LnKWCX57CsjV6sjfoUjjP55l5gxXC09wvAtl4m5qifRyQNpPCPBVT7D3hEEfh4Qyi9oQQxOHB
8Sxspxzdjj1oXW2QD9mgBAQq+Wb9iU9xejgoVNFAhbt7ZOVhBeKnlyNNmXrzB31AeMV4s1uZov0f
S5tyb6ui7teODRGugPVjIcjuIJ1I1atKYeSeXmCOQuuPMdWYhEKqcX+2xW4M+A29z0C3kcSErjYW
LQ4fbIbfrrJPVk1Uy2UO1EvuM58FyhiGMrxsqrRf8Nk06IaJ6/CA8Iiwfw7kBGsg9ZxYbL2S3imJ
O0hQaNfubn+TlVqv3BQoXMoH/Kbzn0Z5/co18b/hgXjzt8dHP2qw2MNNA/eLvYM7WCsRyscmL504
jwduoO+O3sUkTuuCIxtw+QTFYf5jBnjpJrOiaQSegHgvNCU8RFiz34Ca6Bt8+cnSBvrmkxbGBJtA
MiEZXLHt2jvcBU7ErZO+1MoA/aUWklbkaUc1ZIA72Y/mfxrl90NVYItFdjYTNV8dnW8X91xRPttH
JrHuV8wJcTimrSNoSOsHGdHEvV7reChJ6SC7PMQswUeVxMnJm+MIVfdynwJ3bjhpYTB5pKciGaQb
2jIQah5hXt/0cybj3FEfJqKEv2Vy6D1xpoIRRVY+Tjv1FSQILpuP0RFTjSe7wz1qKccGWhsBuepo
994rhaHIVUNo3+kUUUmVgreukWCAL+0537j3VHeQMY/Qe1v5xO6uPxBq8PtQQsEk09HOW3+rIEu6
G6aegb4RXSG8YzCk605e7JNF59+Ev+BJk8hO84LkF+FuHWXAcoPQ29BXlV8b5a5qlTZ73RI84Ex1
/8KdgSNFnimh3FU4caMFvBuNYTuIrDrzO/NyL1LB9v7FdkSUnBsCQgA3BiSVXT4Hrwk4oHr7uvT3
bjTSHtUCfObsXOpdgzEU/z7vQFue0AlP8zLn517LRJKGAz5UneKWW3WQwTCcC8VPUOFP3pF9J92/
qWqi4Xei1ulPAcOdo3mjy4cGoBEEfyLKK5N4q/K2PZadqucZYQ32GMHjUgNy5Il8ts/IUWj4zCmv
M9exeI0D3Ja4NcCUXgK9+pokUd5rFAZ0ohGyjnflFva9rpo/tc+Or5vM6Rzek/vXy2dzVs/mvg3D
lSXgxDDG6g0po7qcuVH3bFmzQbHxVCPQ0Fi82ceVayU3IzsU4Aegj8KxOTby9uhx5pk0gpMBfCyq
vGLTKUQUhvnRCtAXR5cWBviTIxL7aKNcyho6eDHXQKli/2ani/WyoQtArM5yyQLvCTqzKyo1AAa0
blY9j1n4m2jOcutZLkY2k8pB6C/bhvOqWKFClUBZHq+F/2x5TDufONGhRzBtRs5KR7H7707i/cuY
EUM78myRaRS/sH+AOzqRPOdQ3S3AHxrCyboBynKVho38nCA9ALECydYgo8h+imAVo4xMBfsZU6zy
R7Lx9Y1H8bDEfyLbEtuDk2J8FltnxvTP7+ZjjN2bIc6VGSpsv4y+xSt4JCCyBmUaicEDSBanpsNX
0mcdkSp1nqrqoiDSLlZrJAYAjkxCUpNoNztWqeEALr+aFDXvjlpDTQATCC+8PEFQfSTW376ZhV3X
/NYKO2gnReoTA5WR14e73juJ4zUbDm4lFfiUvN4zEJFeX7lLYj5kabprCuwxZlaczRvMxbuAO2HH
VEbNcEBwZNnOuX6ft2ijyTABQB7UQfz6PxrQWUc/lCe5fJ25Nmq9lIGW1z3wKQ8Mlj2Sb8Btyh9c
TUvoGZ42poU+MUNqvg8xECLSGnctQYzANTQXCTZFf7jih+Xv5w+KGz1xNFR5fCRMmPX0EQLtXPV+
pG8o/9172xBH7ZuKc8SIv4kydEKb9QiKXir3DdTqlBcLyKHvStmyilG9/18SjmSzDbgqw+sGCm2i
0zLuFunu/Vd6I1Gq9bxQBpKK06bfLMAnVhPjzrOo6VLYTHaI0SayEvrKZvGyfdA+ST1tuELrFC53
mwI00ICYYmRApUFkJn6hEwiDUl8JhWpqA0USKxGHLRKxIz5bisCqfrrhsIkNsZRAA6gvCQLNQ5Nj
7vzevQIPa2Rsfd8TsMNWNVfXZBbJ8IApDa5T+IGVAYlridh6vUAu5BukE6ReIq/iuM9j6j2LUjRC
E7td/l3NggtMR3e4Zol5pfeUY1qO/FWfWPtOI5W5SkSIV5K9n0rs6lIbdoyQAksDbbgtc0oFtDB4
OjkAAo8LZd3cqMhIX9WRPpgjQzc69OKiEIXGG8pZHyviHrxJzDbRun2FyacXJkoQuTYNC3A9Ha9I
8Afkw106KGdPouwttJvFuvTaxMtAq+9wLH/ft5PO6bpuMzxqHzeLcYckG2iK/jXRbci22dSvRe32
+2+VCm4HRaLsl69IDw6GOYrWdwnVg9LIW6c6z0xUTjEAD/SLaxOA2IbJaKQxXGtkx7myG9Efi9cC
LGWiaHazTaH+WSih6tHSAV9iO7SGRkJvtQSI5CowBKFP79U9UfaFVlCypHsB8XqS86ZB4d0vN+7t
EoZgbY7VulJ5KlOF1xyJUmfU/h373TZ+9VPQ8yOG4FBE2yXwuUnF5REtmWjtH9NntVHx5eiahv8P
pJnHVWOVagHU/thyYjgdxpU4V5vJT+pHXNKQMMI8TCmxugUsZDa8YhsTDEWfqjGRCy2GSa72ApUS
ujNgyMrGd+ONpO3bgyeGV1ky7b0m49lyXilykVz5Kq7+U3bWqA2FI1uaHIGUFen6EyD3KQRSA8qy
5C87E/BctCaW4JkUB2YE1HSWQKbv+8fjak32o3yxMRornPzZCw+yLgqoGD8RErgMSQ4YrscZP/Aq
cdXpjtarRCEqKG0UZVuEa9Rmvc7YBaDk5hfWBRGbmyGp+RzM2mVwVms6zFVEZnfjKa1PNoMpWZ0i
fEPeWttpneSPQAgUHh5xp/8ir1/tVCRjvbpIJNdW9gj8aI+4JLmDgKFh5oL/xnda3uY+hN3Iomlz
JcdOFpYNbNnGo/YljC2PmBtGp2FvB4wbFO6Et2sVsqF4QrH0qN2uphrwfLRo8yS6vb4IhnlFTG14
1hzBjjHwvSop15377AwrvYTIccglC9WlBLelC+N6fh0lqiXFzF2jYdDZuTSr3otUpFxoJP+t5IZL
P3Ne3VGwPqLZmoNwi6vvaSQuJA0oHisbSfvV2J9yVL8d+B7gNCNpTt/4mDh4iqFmbrfMysE8Gc5q
Levskvax+XvDN83Q5QLVmEFqOBnntQDQI5VNkzO0Nffha5MprPxqNm3GljcGvGL7X+k0cybZVZYE
eqA+FTUFNY39PGcCupYlTSbrDFzcVUnWHxSQr9S8jbrpOvPl8K3rDOXz3GghUOYA8llTdspF4AB/
53i3qp5U1GeRaqfILGvR6rnK/Z2F1v6fdSNyc5Gr+xbTzhxFtt6XkcVChSQQxjN8l8qXrmt7JUtg
aQiNs7j5mtELord5k3imP0PDqJGA21LrvuPNaB7gtgXogl+7dX3brIqpF3nNJ+BbiAmPFbNYNxwN
reuHQgtah6RAImSidKeNcKDNlv+BH47vzWKbg38/PKU8+3ddH6hHmzMX4pTXUJsLcfoejvK0tv+3
DqEe1tLXLfIvWCqJk7JM+nQbmZKnn7r33vdP5SSloh+NRP34CjjsplupFtmejluf8LncZ2j6wHzF
xx4rRjxgsHj6i/4giU5gucGaWWSSrdJJEUvhrdyiF7txXvdbVcHIw3KAV7WqEFwZ3w/rdjdPaNj5
U4Rss1xQ66W+YC0PWFBVtCThbKEu5HLtG0PV4W7j8ffy0YlDkzviKNYyo7P14wf1OBoEfHnnfoAN
23IJ/5tO2ldXJ8MtLONseaeByHqIogxZBhn+wmLhfoSjG//K4tpDM87K4huhbroZUGBDsjvHOKs7
9a9Kv1Rlp/dR4X0Ymqp2XEzxHDYr+dmprHJPuSkYREDMzYl1uTn2pFe4b9vRH6/CRx6m38sRU7rz
Wm4E3gRUMO6HlmrTtR98o8KSOjbfhKcOEo1b/xUi4GQU+njpErPjxKd3X/HlbijgckbkOdWPwPXs
/ctID9BhmbRSr6WsvJDr6ZICQlwWSikaMn6kgnNlyGDedLWl5bZlgKMtPYQMFi0GAKVVx7gRqL+F
UZRK5matCbDf5O/RRwWkKW4qs0s2rq5D1KWf57ttp1OzTemNCvJQ2a0Ag6FzWgAQkGsRHmvGQtsq
gulzz+iP/9JOYPf9xvrqkCzQUI41zfMEf6s0QZTraCBdiyrVgmJfOQhtvGRzmAvr95ye5KZYVEmt
atlkxhudNYw4zjBj5PlnNCm6JUVaTWK7ipIH+bKDp4VxjxFsZXhny79HRrsIuKrHywqKJ1RpqujZ
zdIlTc/Jkl8ZlekUBRQBbT+JEOoG6/pVtJQdX5G7kkOX8YAa38WiqLpikIrdL/w+gv+JOh+XdaU+
a0FQrEimArEcYkMzchWCxQBGXcsnMBLu4RkDQJa6Qr0T/t2Gf20I9R1Amx0nD4P2S9T3G9nOBpt5
TtbViIBpwbgMd3CeR3f7HQKH20ix07YUHPkkvZxM8mOIGHdc0LUjdu8iBRB1KsqQDR2O4A/7exRA
jge2qXYWvPbvN5dh0a2LXBs/Edx4HOwQizlcOkzKwaD3uPR+DokLQ8J8LKpQ72whi9tYJHEuSXR2
IjAX5XXPLdMMD82GpEHHyuM7nXCfJpmPbzxG4kphiPElVZku1wGmV1aURfkCk3/3hH1JinMVWbWM
byYVZ3vkFAAytBPjaBH1PBkA80QoNBhc399gxr7YTstkP5W19TYjR/QeOIST2Q5p3mIJgy7rPUns
WdYFycDYFEl8aMBntr4AHO9gkuTetKLpifxTTCCwzXZeQUT101S10LU78JqUoCNF05kkEBJX8+L6
+Jptkoqz2LClNhAKkEB8u16tWwDnqVGCM1tsNoV1ttRr3sH+SBRLM5VNzyZ0mrD4YwNMDs3gjQD9
iU4fQsHeuqBbqThhjD6byFBgspTR4XBoLsB0DwiKK7k/py7lqscXiz8ncVihkghsN0gnYpa0qZZ4
O3zHgwNSjoow00BVAyjxTONdEGHGbUFRETROMqsJm4T6jAMso0dGqU0ceidjtHiv/1D5gOUKFrw4
vBTI+VZ6Yqy1G+H38UHc2nJN4HEnsK3kxyBUYgCRBifJFnkuarjd5mfBjjMdoPv1sxAQZFe0fe5c
cYCSdfCJ6kcYEXBX9t2nLUy+rL7zONNRIbFoPqdE5Eg+scDwPNPcM4kMDyZK8AOLALkZw9BTJzjc
lY47oODBe60WeRMHX6Ikmw1HNbf8lSR6LbQAU2B4uwswBxNS+3QPyqCr53BwI7cV0C6Nc4G4Urip
MgCGw+O73lWM1vLc318AsMMZjK8lq5flx2VfXoSr04O00aU6dKNtbk54UcbxLb7O/918MP3cMQQt
mN007K8DWiLvz8bd5yhYT+hS+U7XhoDZHiZ9tmnNVznleXSPz/0FJ2Lz//Rto4haTQVoPs4xjC1i
LaOenNjax3Jb2Drn+qjp+Qfd6iMpjpwOXUt5sB3oSDeUjQbtt7MJCo8k0iy8u9A7xEfnh4C6+xwm
vXFF6lI8YN69Sht1B3GpGBJkKYOkA9ZShFhlahled2rtO8k/r/v67r6llGLhOFwQ5e3szibcysfR
tonsWuLcZyXMCH78gbzV0378HR59Qt9y7qSLPNcli2UQNOFoVh3dMDyMWG7ofW1B4l5vvF5G1mKN
I5/INVjXW3ux3AUBFfEuYz1rLaj2rxj3hd0PD5ZAW1MXg0bO0aUMQLEHzE8sP2Uo8DHNMi29AchQ
82FhkC9W/W3vVUOmGZ0xiRItGZ+E017EdffeTAXr2k4z+a9PiIst3d+ijdNrtYl0ghcjr60n61f8
qDQ7Kz6s+dr8w0S34b6hi6BewFuR0lv3ky67p1v66oBkzKUEMRlvbwhDtXM5IcgsJZgmjlTVxRkk
3yZ7jW4satWOnaVVHA1/F00EVtWgA+9ptbyrWawluvTEIE4jlC8zyX6pgd4HJ8FgFHHbR8Z4/pz7
RTHRxZyf9NVVFjyAufs/1zTdyzyHBcdsJ8Vj4KCE2y83zNaztu1E5y4DzANDUkm7kyw8Mdr8rSwG
9n4aMa1LcW8Lf/yYusWHGg5AsRzJ34Kl7DniHHdqeL2ZYNlymdoxtpuoQsv7HsSoUn53/fW7tzSC
eX6EhC9BX45z90vwaHNY1nRsfaU3G4HCCWMMzkseJXDEDJMFLUgnXVbo54gFAOdPqv8P688Q6m+r
2A7vEG2sY2uUwct5IRi+9gWQVkg22tOl4hgo6Gp2PZe4+jI0Ksq5wf0gp8vwIKzVNqSJs7XLPzAb
mZkUEW0sU9fK6ekU7bs5ttzFT+7OMK/HppngmPXR1YepJnAzCz4hvC2FL3J7TWOSSYGPRX3b6lhf
T1ErWZp1uFJZgOYEbKQptkTRUZXKN8KvZKHEkOk0aSDOITb7JyaxzFzIw+JWhpUbHSWKnVL9T5xT
bnly7GmuwAJtcc/x+pONpOeYJDNrEBpd509neJqnhvcNvOXKnpW/Z5h9YK4w1I2ffXhMexDO0tC2
NkZS0ioCxd0Ek2z0QQE4FfJCBgMElbywmn/a4zxJ8oELPs7EsqMOteaEzDu1Z5U3l4dLVhN4+wt4
iIkZeeqtqyQ/qm8brTQmHvhUA/QOYSlWFmVs8LUsdcBHXHcSIyOeMXDhVlnk9OZHhRvdFD8ZhLNx
mc7FJzH0uZZrRoGJmZMxXUL5+vmnCgPalgPi3X9QPrE81dNYx1U6o/LpmJEWGgq9/0YjlVz0BZ8v
71ryj/L36N2RyIcpdQMgYaUm+9+1hWbQEk1q2GUXR6QstST6FW79iCEmp1zkMXZxb2QtuLzwfN+f
FZZX4VsvvdHfiuR/yQzp7/faDxSUVwreuYnLzxfNDFW0r03XnjL2hhJCsjAXCN17A9OAqrT2GQPY
ZKYvlcemh1dA1UQJzJayOF5FR/zlhpaJRxO4b93qOWiNyzMCoNoYQ9nE2NQbPUQ15W7kzkbSbYef
rXaG0gyg3/fwaLafGtxfO1sAFlj6gkrNfhn5uYAbmsb2u4YD9xIXVrzIXdVgUVJUwwl9/qtiXk9N
hL2dzFB+z9JIeIveeOwujacA66LT5wpF5vfu36YjrfJtMf9UnHqw1foj4P9aO2ea7OCyfCZBljAD
rDxDeFWIslKAMOJiu3H5DgvP+cJYvvUNF+SdNsb1oSF88cszD9Ma2AcVV6JWkE4Q+rqnTnPu/Ghp
WzhbyqTYHZxJuTY9/kmtcf/dZxXEE2OLRh7v9BWEDCmdHmtur6XVFyewMFRpWCNjklV2ZvHpS/My
7Uaw29Y487G0PiCHUJqP9QntI/4+b8C5EQM033Y7tPr3EQhCrSdldSPOudke19A2Qr5y6eoAGBch
kMceXYsocBpZsYcNkdrSzvZHPd8oFPvS3Ef9CQUt0QP9xNRKuC8VK+pbuukYQc9uM8qgOEP3mcgc
eiIFtTCCAcg6rAaM/6sHbh0yTRL4W6P3DVnXJiLH1NPtDXsmo8SJtai4C0R+kLq8o+vU7V92c9et
a3iQvV7jc7iaIhfNYCkQh75ook5pCxPcbVNZm3t+Rn+VgU9eTuYhpd2FoswZlqPHZV6HXOJ0omi1
9oPdJmCm4XhGwtaSFO+hY89wYFs7Ky+NZ7COGxLpGo+W0E7tFOmEqNLpGz9U8v6AAbEQk/PTFj1d
AE/pT6SMyGXjLS/sVAkjwvwr1OY122yoBV6Xww6WMVSn0zL/VZ2rW5Y0HddrPFs1ez4pgCNY4b1j
XwEdSMYYfK+qsexA4NWicfEYdHv8cXQQ6iGAj9Zi+p9eipnZZedLBUSzhpnWVZLVW+FfyPhegFO4
OwoMelegUPJb76s6S0inzHtg5f2LfsqJ4MkH5uxo9r85ql7Xh0Fq79iPpyhQZ1bXGhEwV4YCRqNy
U3D9W8vqi7ZluxJ0+dAkPHu2mOFQwhXbOPpNXCEBRikMsEw2GrSxSBnWxl7DJNb76tPlUk2k6G45
7/MkLmM+W+3oE7gB/LKdmee2PXmBmo8hesMa2hYsFbXtJJqx7RgCvoENIVQkajS1ORXrFJJoQGYP
673ursg4AG/6jRULbIGuqztBNNvQnqF/Fevqz2GKNDWpJsClAsP7MBIYP7lNpvXpi+32yUeuxAaH
Q4AVdrZk8SZp1zFaZeIMwDgsdmk8lh/yZeGOVriW0/YMBMJ6x+y0GS4+4C7+CY2Tkx7dXUs6Ob8/
SKoFP06p4mSDOh58U1JZUjMRdczGK8tZO+PzoocqfRhbZVjY4Xe9Ed9NSraW34J6vbo92O7Oe2bg
e4CbBQRBd7ZFZ+OSAqABlc2bcHTblT0MqErK2k0K6VMLn6H/EVCepLfXqGWSrr7NRyObkbkGlOSV
XIVJlTpP5jClQOp7H6jB30eqlD/5QXJxgPDQuiLf+1YJD0yk3Z5PA7PWYmnXIURvsx6EUpUf5qcH
CIUMm1NgUgxunrMjmMLavIrEYR06q2LJRa0l2JmGTheWMdTpi+FN2MRtVXkm7HjPvXJdUFflHaV+
k3DfT/z5oaX+prNzruplv+lsF1j0wMvQV62QLk4m0nIoSx7rdxW/OdEjbu61QEVFLYjXaIvmm/Jt
7QxnCrKi5tshqcPIlwmilqmSl5FHLEeIjg52Jkmbhk1ncteS7U1rtDOss+pRbGG3+2Y4oj0D+95V
HE2BY5APiLRJRCrbx9U5cI2seJGHIpYvzS5Wf/R+O265BjBugW8xd3R9Pl34oNM3e/Hp+vIKZdgI
uu04DysuNtNHSqvHsghrxRB1lwSPLr2uJlg2so4OigJ9Vcs47ks8E/1xk1GN+vG7lAILLWCRVxb7
Nk3pfaTJMm2wg4JqCq6aTsxdKpmKVYe+NhrAVdj6pKstCpzXZPs7t7wTxV3Jyp7dnVL171fy8UkS
U15N4vCbnuHPeHY7qIBozEwnz5Fzl41l4OTlW8rGObTMRzp5iRVNdTmfv7dcdPemE5EKtLoM8mu7
8J7/WjsumzQgZ3OE38/1T1sdkNmnTonXUDSpiYth6stYGElutcx16B9lTSKCmpC8WLKhSq778IzN
nALqPGLahAMjUE4SiVxlgbTPU4QVGK65zH+YRoPls1XuGlO5ePNXyRVEJ5Kw46IAlTQy5WOlqbGK
8dAtB4RahYmTQagCVe80HRCieiOtMi+kRxE8fYX9FfLVgLpAfgNSfTYHxLdJ2tglRjMMleYiIVTs
XKahodP3JpQlrXCSH+NXOkl8quTe21Gt5p/kv40IVMbBJJxqbTodReqBU3mH8Wo8X2xoGTZOm1S5
fJkSRrnT51ePF89/P08LF5nsWbwDyQnufv9Mhw7fm8G3wuMlGn95aWmVgDZKADXi6uKbs/4K4xrG
oxqJFE9Ndrenmhopn/eQCyeZpIS6h9r+dJSYj5Jj3q5TWgqG8wePWi1sCZ2NTYDJG7k8q1bF30/l
EPVgAQSZPNQCUYWbiHFlVR63bWBfWC+JeThIj7bCZAFskLdfb2HGrOYYorgabaKvrLToYi4KnqJ1
hH443IEpp2VTyZMeA1mYD5nknLdfEB7Fx2aFacsvPZ0QgGUe78kzTcBjQ7IFicNHyBO1ZC4d7Xub
8b0rW4LqNYBOrXiAHxMdTVdHhTbusQUf84wQIwmZ9bg6ncMNfEOWcwwSnXUt2QV5ElNGGWXjCO5/
xxCfIXQd2Pv0+OvC4jSwgxsXPeoINxPKAsRpPxi6J0t2h30epFVsW22flXuw8l442OyzRUKI9b2q
V5B2U7+EdO/lmuAlM1OHMTOmqHP07OJwemC3ui+zFEaA3DWvUwXxILcAtSGw9SGkmiB8CNg4tvkT
jtimY/zJz5IA4tcIa+eP2UxzZFo+Hq0nMTUhjF/6F1vuxBtBrfDDRfJA/ueeccUsVkh/NbJEsKlF
M2l6HB1IIpL4n/G8JLlS1TcLyACRFPzU1HWTXZU1CcoG0DlC0f7z2S9RhppHwQFCSIj/dfB5qO6z
871b5NzfAsFiBaSG1bdrG7/H7M/E28iVcbn8gjl+yknt+XkSM7XW4pbcNQhynLaBPDL53Boz9wCb
/LgVE1emmy5MSuyQdQO4FjQdN/BqKn/ML2PkYnFaPA2yKyEWWQRS4fr70K31QUwCtMS4USm0OdBL
jLwxKhGi+0d/UKbNjV0vJelLtU/8FziYId45YCHileTlRdnmaDsUKIizyP6oH0ltRDnPNPp/LulV
99lHHWvmbv+WIYLI2njFTV3yLq4L9HKIFZoFZt0rULxHE2lowyKSJ0up+wLsEOtZC97di56a5vcI
tJUNUx90m1dgkiUXGvLlvuZmkcnxgRUVGSC4mdrHIVnBwfanRPrThdxpNxSVAAEQDHbwVFWmiU0/
DDqU+XX2T5qinRLl3rnVEjrW7/GE2r+WMMGRv9KPwMr5/q8VEkWH0pWfVaZxaymVtzs9mhLuCQvW
4V7RMvwpZDsq5HiVaFlMA9+4pK0su/zVSy2qfj+74KAT/ADMrtSoyn3MlgacpmoLtq85s8a4iN54
DQ2W+tlM7TSB/stkzSPsPnexSvCUEOw4QyHm8/kzaO3OdtPsfkMaEsW2LhesKbjppKXHxEUX2sCv
db+K/9xLmkENRuklBC5jGtD1EAoCsCJhRaAflrb/uiiBj7ozWcxiAA0Vs2ZQPdgJa8WwU4GyJ65V
cAxhX6Rtrgdzn2u1vhTtQ6R0a3sR44TVTjhevpZabZJz4YIHVGf1l1D8jplZAq2mQlGGvuodhFM+
QzfxD9EsUO1+ynTuSaTuX5sh/TgLvmBhjaYcNC1eXcsDv72a+6AXwwKnJ03CFEOW0gxZuPU8yhrN
1F4H/JwjD6qEN/EtV7omOgW61Z2gCb2ao0bvx03Bmkgca1mJ/0PwLtqV3eKiTwm0U81qqO0QUeZ+
QlLmc16o8ULL3f9gg5jqqi8lqBHGyxpstiUYE2zCM2iQCmUirW7QPr9O9GngLVDuBQCxgCXtDII6
FxUAtK096ogKfSFvpZW9q5zHl9cD2hNPTvOZjv5kZPw4YM5FG9udKQVzYJhekbQ3RqMN+1AvQV/9
qaE7G0GTwnCUrNs5BJmIi5rMIkiI0gIaF1hiOSJGaXMo8cLPhEkfijcNFzRxgreIn6xTeRL0gSOt
D8PyteNE8ITtLcC3hY2nJYe0jG0LCkCfICg90kKyGX+XREbrhJjP/rmOJZvUPp211u+5mgD+fug3
0lMPZPManQy7QTq9kYYhB6f01oiGWMLgahc0HOCMq61a2KA0FUC1t8br/BEkSXJD9LLWrIAzsRZi
Kd8L3fWyZbON9UrcXkcOUFsy2aUJLaGcmuhAzQxL0U8PgXSAm2e6B3Eml6CF5qu//hdBPs5NF+Vh
e2SRC1t9aCebrBCzmaUxUpGpNa2WzGzjgrkAm4me4Lt/CNEUScN+fEhDCrQHNkv6Hn6IifU2D/my
JdRAiDLqjW5KBcFMyfnEq4a+kbn94yxAVjHxq1POrgL1AI/GlHWTzGHN+U7p2z8d1s377oX7GoM4
URyRMqNJMuSEBj2i/3gHvEPxlElxyQDi1+v2UqaDXtkVhUA+IHRsBOPGrX2xmG6eXEYO4B2lNKz0
y2riWJnmj0fw3SC00dWEP3hgEOaKGeestlH5oXbIN9+pUoAOMYfuNFxAbWXRLgnc3R5GERoIZR+Y
HZEju8xRbdzsXYUWtWK7taTUbFUpUN+6oSbV2yFMY2LYxj5oR0OEmGQv8YiHNGSrKtaOK8yOP6//
JrY0ZdokwGtRN+lGGprgKTx5pGFJoqikyvlA0WgcrKPNvdxQDszZWsTlOCgRPgcCg+dgGRUfRkmz
vqhdwxV9QtjG9on2krSWcoTqpf8z7TjpQGaNynC4R6Quy0supe+vO95POLS1+pMC/+0jAwhEW6m7
gTIcIhi0Pdgegivzi+k47Hv28Q0eDv8NhXLrS+ZFXkGUBsgtqwGAGZjDliGP4wf8/F0zOE1aHV3i
MWkLaS5Wtny3+QPRC+NX0ZsCfCMg61gLvNVP6ZWDHDtsNZI6u00yyQc9mHOnh3A5uyZpm2pTlir5
m+qPtTl6HKncZWwHcuEZjs09jCBgyntO9/iTGQ2ZJMMJf5552W4GctR924VxqJjw0d8xQWO9/snN
4H/fllmaRge4dDmbhaQgbPnUUCNbsNb2wK7ZF73aYo7MVjrXigggbRJHzk1G6AEoCKJMXeWfRDGf
ryU6myc25C27BGpRziYzXglXhC66uw/PVA4sKlKxHJDJIDl898HQhh+Xn6EyVNcWRlbR8xVBaaau
kDGVyxQbXuKoi/fx0gsob1Zj+Uwmf2krmUkFx32MMmIe4s1+Q8lDqgSnjdLdLUXj7V86Iou9q3is
Q0azPb0QJMPlGp7lMooYv2VmFQf13142utMWpjDiDyKI4Qcn7ipZwT3b5GuihtZUFAQryfTvKIZ8
H9QJp2BYL1Cb5KfUvyrpkWYKtVMHnDg6pNFPtBVvdL69+hdPCBWu+uyxVInSBV7etkCGbV/TX+os
EVL5E7/qiCGvHg32H044IU3jiYHZnmwI0p9vJXJD4QTuCophaOVy25HLiYhGuEh6yz3ceONlzQ1A
wjc844AALT/0oXOVGCKzjinhaJ67jcd+qh+8T334udqdJqAm61dFWnHSWEclz9QUF4YqOsNun3eE
uDXqBcYPripiSI2cSnfQdoCaKmNudxZoKEv1L82RpMdt1l1zhIFBmAa/0EinTQVuX9OAZtdNHZt1
BihryLidxIoDY4v085sc2FAx00KK1jN5CVNUBsj69B6FZButa+KHeLcnOjl1+JPAhwaUZaawdQbX
UlfAeg3jAgsoiTkJo/WmD4nptPbI4K4RNvJysIy+nktXorTgo7l2xzG7fAIHK5efSqhknXPYN7no
pr1JlLDTFVDweweaKjrEfOsyRQfyoqzEfoWZkOzQv/GSOhlyxx8KszSxx8lvK6JGZX8k5fKwO2Aw
i0wiFp5ScbcYc2YUlVy7d7CbgEeMrEOZ970GDdBe09LzAtDqq/wzlPRzyCoL2Bt4B3Po/gCfjHnq
MrfH+SvtxOy7elleVIo2ctS+HYGyYSYvmzd29+grRAWgiBXIYD7miiTpSjuh+hcqK7uO+mdTBVIy
JAsrcAzMxaa+AKpRWSCOVxQPPpVowudArTT1nex5df/14WTUMD9iTIZXMRTiOD2YGoAnW+LRQgsl
z6xRiT1IjypUwLKMB3P7Q0lYQ1ECYJXu+xDbLMYKOcRRXvrdgwzZFdKx/ThHvZ1bFwdLiFL7Tpf+
AH74MGESe/YMWbXdYy9FsTZGaeoID8PszwcVHsucfrDAw1AUpG2x+INQ5ZuA4F64vYVMyfmdsshh
KsQGh1p4daL5avf7aJzwu3HSP5W6eR22kO4d6aGzBfhixT515wqC01TxvCIjQCnHoI9hlvN9G8SC
mxhSizqR49vPyMdXSECQ8wi4NrWYyi7E0KPAeUT2BR9hNQzzMuUv4esIDSlp5weKRBwoFLNPF+At
pothT9LOtJ0eQRRx9/wi/Xb3vfoTc73zJhqMfZqczeJEE2XEeKkDbC18C/2DMk/kHoiMGOhW7/0N
KudMz9Cl09nxfs+90A8PGfa2HV/XjSX+F7hyB0SnM9ihqMhb8VA7C0foQM5BZtAsIpeTbvZUHuNW
+exx6IWYFNbOfX+sr29yPPAiMsZJSliei+KCMUB6PC0kLsM5dJ1v0o5R1hCTqWG6gJDFDA8QOOn8
uXELhCgd4Oe7xPTkFlCRoYkShSmDwmu/4ZFvW5CROVRpkTIjN/EFNllv4MVO2vo4T74h53s48esH
EXT/VHL1ytLS70DDSzbk3V+HHN+xY94cqVWQ0FYaZlqKo9VuVRs7BeqqY2SSJixyDPOW4/G2IYBi
LSvtEU5vzYzniVsoV3h0jExAWMbYTeZcnJJyTs7FJeGmsVW5K0pHOuU/aeGWsAZX9QBjzpYnZfu9
BsXq+vt9Tjuclzp9LJgjUeC+Mgdu2llZ0RWewahTOzt1lOb/kfXCZNZigwi9FoAiOgPG+Zz86D6f
xoOJG2eA6FhmHZs3XRpIk5B7vhZpWfi4dqYBehaZK1J15WaCeB3EBDVsMyXPtkdROl2VMiV5bYfn
xqNqB9WqgYkjyJ0dox9vYK44ZvqCpKOIYshj6iDwsPdDg/IUsPvxFgW/GFiYFPocICpgPMk5fh+a
lM2cXR+ksHpytvC6d++SZJdhDl3Ud7fya+EVgXbVPJN5+Cat0/rUSru2nHG3+1OfO5HXbPG8VAyJ
iZ/DWIaLTsCbO6vNasPoskUUX8n0PanTWZynRwcEcfq3UmJXJWI8lG8qBZ4DE3ndKKG9pNotJnoP
7ah7pCylJzM0u+J1gS853e9bkS7f0n36Q7fI/JMpjP2QKln8J6m+1ShuNEkANum/xcyubGWRIU9/
4W0iM7meexZpfVPNExZq81poziNJSrRT6GO5+fVDFsQztyfF//7yrJnmPp0p4tG7rPnEedyHa2Zn
lf7XOIp5cFcFJVkx3SwhIQ6V+udc8WnzFz4ZYP1Fhe5DuGe6HLhnrodJeqXBCPFmjrLJO4WgWNG1
n5cuii52lQUbMvaCmg1Vglw5qhFUJrlP1exJjSzP1M5BqgdfhcvjzRhGO6+LchdSEP3ktMIrLPEa
Yknf4LuM4bIQQ/iAkiSCYu4wbgUCG+1cHRoLj3cAsPxdlfoO5dvYTtyzATF/oQ80FH1V7A09heIY
P2ZeUgpFtSvxQKfqDffxLSv7frm32pEHANYjGznSeJmFDPsRxsQAt2afoE50izWzKxrpmUsJRatO
e4ra/SCiUvIDgMNBxjPddhY3A6CGpyhYu0MAr8jJyxa3ZznW5EPid08BYepxGDTDUK54nD3fHiPv
VWImHXO9znI6SGuuBuhTIiHxzkvUW8tXmP51KQVVFzanQo1Ldba4yhxyRKwcFYVp0Kfca2TlrOZn
VmGIfGo1ZHobF9t/alyVIZ+jzi3vgXuH6RVwh2sFidtdou5xqfEFG8+JWsCELT6tQTo4lY6S9Qkp
K2Yg0l9hANjz0iRTdIAMNi4tDPwnAk+oBpy1M8N8deP/KhzXR+EglF35lLuwjikTyk5+e6xUDU/g
9IOpfhEAhzctea3ovtIadyjez5Rk2cyV6RDWak3iqYj+VMBRuOX7SnMIMfcNJr1Lyg0lw0taqPdV
1FZ8yUuILSra1NlLsWGkYHcJRio7PXfwnuOjYS+iZ1Ra8VM2/L3M7SsGcRqCuH20wP7KB4PRoh3S
UOYu6/ecw8RrcvznDHrNrgVTH5IRtHmML1+vzgaW+3YJz3776FT5VGn4z71yAzNGLYyDTy9o1jDo
qqItgizFZukW7o+/l6uvr5ruAe1VGhQalInQVvKh+0lf/LJMfiSDEJqXNmvpwj+fOBppZ/NpyT69
lSmG+o5uGzRnfgN2fs2zIKPAWd6txfBPJNOh5hqUi6hGtTw/9g2LCyu6x5Mmm8TKNz1Dju81jiIz
Vm9yWNxhllvjb8TNx3DPpC+s+71SSRFYJncailZiIleHB4WMVD9rzKGryLxiN3tdsZYmPUhXFRWe
Ny0ifEGzpxX54ha0CSSIkH3TJzYfhSKsVdMhRAB+eDj7qO7L2FZa+nIJAQ1/s+5rwKSqAdCJcm9K
Jh9oMTdEdZmHHIvmTqxIEXnUQCagZEuzxwKz1Qpb2iJpTWfCqpFAGV6y2O6tqd2sC2le8N9x+a5V
zJGtzuKvKgC6Zp5uOk45LsYtimcwhvEpDGk40Jc7FJ9sIRcX2XwePXf+ISVHICsHlbErYMkenUtG
UGyg734r95SoJmqtmuCYaYPJcUiM1E9tPKOlL6kh6X8vgOGoPjrxS1b1SiPT+1c5ZO6OokGnsVd+
mPNcSa2Z8/nQEov25i5ghuxgR8SNgo/p3TBAXrufQstVgnHWIkL+2b4P+uN3JB4rTRRPJUg962mG
PXBaNaWtmEGQhVhH4vHsdidxR6PijGMYZcBGl80PXGeZSd1IE7q0PxDCjL/AVaRancZt0rSxi9fR
qUWMq0yGeXpX1AQx00+3NJiRVluHmOKBAzm9cfR3eXOyvp0nmEN0f7citGl94AmgazE5SXgG+xDA
eQupzfaPgm3G/8Zq/K6Yv94YNsDIHUnC18gTyqwNVvc4g0KEMsMFQ1uH3gpGUbyPSupeu4lJjlh5
uqYoDRt0A1pyCNUJq00CF2poMSxDeaFwXAWJZfCqmdhHbYFL2wtNRDX/gD522KfHYBvdDMOQN+ij
VgeyL6vCPC0JaPZWRqVRQFgAQdH3rZFEX9ju5JVAO6ugr//fNKwv6/HL4iSEBR5h3hILloXSdLhY
gzHJ97vqk4OISDn6cDeqVAW2RYBRitmMEK/qHR0bM/QLkWZyLJ4VY3eOLG8Ty1dMAs/dv0s4Fybh
nG+DxIMkqsskpJHlbyDI9m1gsBKezJRwlIzCJGgWJff3DunYIha1pSQF/XwPgMwfg9SkqvfK2Y++
YSst38Uq6v6exjkaucH1juQiitA1YZoyqqzeIMJMvwR+wEkOm4t9DTpo+unXPcp38g2qqDi7SFwT
22Fz519O7mu/+/3gZkPAv7VKp0ma/gjR+VNit3VbAvH6MaT4pDcPSeb4xzEgT/xfQEZjofRCzBw5
mvzUWoEj1rKObh8C1bUEh+RV04cFoJ/FradlbVv6QouuA/r21ADE30inXosybwcL57Zq3hWifQyD
cR4xdPLNtWZG+CxE9LboQDR8Sw6cXNFzuXgfEX20d0E5q4QuLZCL8JcauqGOA113aI7fjgKwWaAn
jix0RXSbyJdqTAUBZ1R5EZH88S15WRcDoNJce+QsjTJhEchV8S8+DDY5i8xO6NfzJfB3+CNSbE6t
c6PaTpV3eh4XsHYkyYuWjtBAhFN5376UN08BXjU+jE5i7iB7McVG1+DUU/xEiObz22Khi7uBbcCj
QzA1/YD5OFbCwCxRIIGrA4xhxj8UvU2bnAH9Jdx8K67nPfNvNTVRyVjEkOY1DDDLWKNI5v+ii8CU
5Ru+40Vj00eiOZZyjcqSJvs7AzRXIoWgcu1nr9Qe6T+/6oeVQCTIMOfrw+nIyPfeMVFnJqxYOoKD
C/9xdnvY8hrlaZT/g/HbIxO6hge0+DmLlW0yEafCOulx6WJf3xfGcHKTkLJ30Jk5OPtGKcrugF5w
nak/bOKvhu+/8LUIHwfGd15Uj9KAgoXcbZOsJSEyI505vEmE//GhankIyPLMLShArJTSdHYga9xw
gBksF6zLs353gAE0TWxaIzcVV0ePSqcbOvJiEhBeQoN08fjMB9+W0tJryJz3SXtL2rMH9wGp9/xz
zOk7rUgtxAT/noYl4uaWCVsv6YLIxlUK37jiqMcvUKN6RmcEarwDMXuARkDd7iE/EF/P+upK076H
IoJa2fUMd1Kaa8MXXILjbcVEAvbFt6iLOusOCpGn+32KUUEz9fkhq/SPSWRQseemkKPXctoRpiNk
7OHJPaqNklD5AILHNuS1mJ0RjjarzH9OhDSP14jtwrB4XPcmX20fTOTBNkd/DXCymS372OeDfqB4
UpK63+CUzl9VnQZWYPGS4stgWIq8m2ET6Df+kX4WQya4cYxrWg1DhDSIlA7wXktxsmKY6IBNjkKc
VFFpwSvOK7gSb93locY+VedBRv7ZIribZbuFrBGTpOIvhmnfRCLDA83VCWKOWn7acF00+jwoAuX4
TIbd9kUCIRboDU4Wkbmzhf5Sae3oydCyITl6cpm6afIVTjNDbJyTYeI8HQAOQptabRKUkaW7R0lZ
gc0gCzL9o6o5S7shnRnHqApNSCLvPdKeOQGa7eCeYAEjb0WHLpU3CIoNgAHhAaG9IkVnE/WGuKmn
M9rgmW3GhM+hoOfsucbI9Tm07bDZq2/rabvx3EzyJTp7b6lIxpg2evAfPXRYgZDI52ERE6OuPDjo
QaYinIFjgCDdaUKbJUwTbwDThdGFYNp90Mn6kMIMASBfj5rdpoQ8zwZNghxaSe5vMOT7T4+ovw3E
fn/rWLtaaaI4nD2Rff80e8ijOJbOgjd1hvWtqUJwZLOqPcqtarRKP4FxFafqOJiO24KkQu04L4el
bMkAR2WX/4yxLjMsprkSY5O/sG38v7YGUs9Twy5UkmutJCrS6ub3NhJnfvb9cmy8lkFkIDo2f69q
qfqaCenUaFBKtehSm2vEfiaRQc9L7TkIwxB2m1/hIfABde/NKPOoueIcD19QoUSjYB8DxS/NKmlr
EQzjE4s9D8XXUHg+NQM6vHG8lshhMOogfoahnADKBAuHeQ96zb+jFkQ4wj4vRHHx6JGP+STDiM7X
0vSFTEEARpNLM3n+fpNW+Q2XDX12qUIdILYnKr6OQqrgzCfwOpfMM2UI22Kyz2zyqD2XJ0Y2fgE/
W+bnFppPHhQUbn5G4uDCfGu0mjliLCd28B51SzdfD8v1A+QS8X+6r4pfvd32+JAJoQjWFCBJUiPV
8B3fuRBwUcre7g2OxWyG0W9C3pkko6LuWhupkPtm/exLNtRTAJ8QS0Oh7lnUDMBn03yHi+qlPirv
RvNAi6qIpSfI1Y8NYaQMLS3DdBkK++FoTl1w0ZgN3kUmrIYtVoyLVbCk60rBUl/AF89Nqckyj4Su
QwLnRNVyFdx+X46Kf6cFuD08TDOH/jkMvnTWioz8AZpfhf5wlkZXKp2ohFN74totbLbNf9N7jfC8
dU144/DUkpLSpuW440b7jyJ1HRAZQupuzY7mH7wBQcg8tzdynmVyA+4sEQk8Sdcf1CgKkZvrNlJ5
tyU7Ywsqu85RK2bGb26lDkUUd+RiVIhW1rxAqO6P5Ebd5jeZdj3j0wRSgYD5G/Bgdzo+DgPqTRbU
tnLG+CEnKoezUNP1uFwRJsdY2aJx1srtZrS4hWadWQvTD6NTghAnYVc9uf6eGrgAxV+vyl0dhwjv
nBNFoMz06VazbZWX/pJ+yw1nCEbEbULMO4qUMfH7xOaMO2WF4g45j+RQyDcU1G7CrvbquBydYaUZ
7jmmv0icD+3/mIry0DONjch1pp/khwZ+igJFjLnIvwSI5e0WnGdz3NC/j31Q2TN9L4smMQR91kwU
5WXhA6oC24KViP0dp/r3agR5/XyXQ5yWr8lBNCjhdKso1xYK/gW9e5zbvpC5st600j3aBG/HliQR
Hj/GDLL8rNUlrBhEBpirqn6P5HVaafitSEmxNDSJHJ4ccvL/VQNfhpeaMSjd1zjv1yzFiqagda2n
ksjQKmO76pKgF6jFbE73x4U18fPge4Y1D1TW3c9lvjAOwVFm/jAZlHq32d/mg+eeXPLPri9wdCMi
jjVEYu/KQn4g89cAPPqHb8XQBsoGlajs9eWRi2ZkiUydQeVakRGT0oIH8KJD5Kiy4ViIywx7kc+x
LT1gSxkUvoN15tlS7Tnw/zGjvENUKOkPuE6p9w/JJ91GpvNO0IaJR0aUjWBSYCjRsOrpUe5DZMqn
tOi3Wv5BBkHNxKIUZkwzytcdSHLYt8KP6NmeIZPff7OHcjoP9PzloXRsKwDli7+0J63t48G7Ka3G
fxrRhSlBXuO3vtKRrWmqiSD16IC8tYsyFT2U8qRr9vIriCvHyR/C7XBqnZV9Oy1plK5L0+ZjLxDW
FG05SjUfqV5AljuCzDejixJT0ttWV6y7d+W24DRZlPbprxgrX9xmQDrIqGQW9xNvG9JVjk131pox
CAEAKXcbuTuPKugPu32FqYcabaPQdWzg3N0bIXEFdqkhFb2ugab6XWnrpDi5pVFZqj9PQ8Lrm6L4
b3qOKvSFhOqwaXtNYEFIWFZyaXaNhSxT5xexYnsmyIU7TaO+jJaVY9EiV37KXwALkSmAQt+j70Cl
0mxq/fj80jbvchvy8Pnp2S04Bpa5U6rqfZANpei5ax+fKbBCjtzcbNz17M9eCfw8DG/wEie0DCb+
plQPfzgs7lF6ZcuExhzMTZU3RuPaR6AcKHlVcekdkr9CemEHJ1CJRp2n4SmGShlQYfeSRlQrKhtc
h8Dny/zI39ZU95p0i68PYmNbIp9V/eDYeB18RS/kr8LPwP/N8KbFDAyA5dplpe9a4T9D6ZAMZGO7
OPJElMH+1RxFG2UXjnkYuBG8GgIkCHEHel9LC7fBEDy9cyaNuQUGlXnnFRZtUUMPqYB4o3tIY/j3
qHvnzrLlg22UAby2z+1GNenWFqb3GX98GjOhC35Wn6hY2BE0CFBzMoKS5pmuXkw2hdyhnqobVczB
FTBVqVOX6RF+tSrrI0jZ+eoeLSAnI/p5ZVpiSxma4UcAVKPHiY6XygcuBMPQvPbHEpFLBAcSrc1a
cCSA/wiJTNfQAgLGSDef9sVFbb0RPqI7rUfgkSQZdOTomyhRUkqclHIHNw4bSII//8IieWo/RMh0
63S+PUfkoudwAAXnp63xRM1MOSeCpGb5wt7eBZjFwotaScav8aMzTA+S5jNJjNoabjzdcl7eQOEA
jWKCmz0W2qt9vFk9QCcaUqYtClk2Gob2wHNuX1vou2rBKChU1sVhWMkZuNAYDEQVILrUTwq5hSVV
yaraNH6RZ8DyaLcH+ht278ZvbqbOcKwi/tNZAjqvBFqRzVsN6HKCbP3pcJDPil7Cuwm/SPhEM88L
xtBpk2LhfAoactERwND55E3DXuXZgrx7iDSoc/987+txdD+Cx5EsOi0A8XLuAmX3jcEP6Rhb3j98
SE2fir8nDRTmlY3WXPdFDB2e+4GHpUuoGjRh3DXO5zilriYHy0X/vdf++MUTSVOVYKDZO1tFmcPe
jHx8/zGFaU9sCSCBMx6wkR7suwO3warxnd+O59dD/itFzqCzMLLHUIrvMMyky80swLWdsWo6oFDL
kR71j+Q8pkbOh9qGlE8S7IkeF1+8DcKtXXVIRCBedJDhV5Aezto93TA1Dm19YEcPL1a86FNfvBl4
kEkhA18FXO6YMxjBFbCxBhk/LWdjcHMnMc8GDX0Dhwspwrct/WMqPI7xXZeKtPTduWhmHhc95bmF
t3a5O8I8QEI/ElL+iQfuJ17MEEXhU/S7VF8r7e0Rqqceib69hKHIOgQpN9S5g2UjCifK+1tDoMoO
7m9lu5dPAfNzauyuM6vklrpRkEMnIoA9qfOva9wp8sQ80qjrrIynOs8+6bRL31tIT1IsFewZnqsP
dAXIkA7yYZfCyB2AQwG84UMiNbuKa6q+jEWjYeCfTPe+dg4nqvyUOQZwR3HLCUDd3js1ZYDzR33Q
S0+LOusEFf4zbEEn3n17Wdh+onIXc59Gv+JwmiOq0wd2MJ1Y400OCwL9FHgQga2Rr69hu/awnfUK
mR8pG43qG4n4hc8+Kvn2PGuIab/zOL+fiMjf1kGLk7bRMSaZ+bpdXvwxzIPLaR9NiNxdtL0f4jxN
QteADF6qh+EyI9QVSYLQHsO/7+0IF855P89s3t88hQZJEoNJlGPqC5JXJG0TFGDFE5XauKsO0Rdf
ZIf9McadVFVthyT7pL2iabsA0Pa/WO/Un858tH8G5FFHNJTU2oRMR9aLMa55PFZvxLOfWSbLjvW0
Arj8UcJFzVx3aRNDzNKk9mJUwp49DVBtFt6rVar2W2VFkXCIMwGhlA7CrlNatQsUUoJ7gSbX0c9D
3748dq12dKNKU/SkJu7ybf8xOIYiqs72boifrr1BBm/qhxBUdlHyUKaQiMd0eo7num5IXbHVbHgr
Qepk8GfZBJAXIhvnESslYC4887Nbia9YFGi7H9UFag0ENTwDiW8IUXyP0Hsu93cIA/TALJvCpjOA
1z++M/2WDhJHvelzb1Vy7Pu3g2gB6lqNaJU+jIjaPj+/JT61F1d/jHXJwU8FFCTCHg5Kx+p08vjl
VpJ7h4Jr/JN7DG09xnIPaIGmQjrr66++k3cuP4E+jSKw7t9HEfQmH8dlBSb2Uk0ai+d6PKjiH+nq
lfhDCVTHsGiBDWX637/VCdD1cBWtocHAklLFMl7OiU+Ww96XEQXnKOzmShqoQi+Y++3z90viLPkY
pUqwj6eHLycVwr5NI07mJmRsxZ0GIFyQ1PaGzDN0DTGaXobsvGRPEhfPXVpxawJdqDXjZAJ/5YDA
97cCK/aafhjn0igoOTXZB5nUwqj5p7rbIJDvrKDnVEyVpaYgbwkVUAHPBMLB38+Kdc6riqqEu28U
mQbXZ3oxfAQb3FH1WvV8epRi9acaYHiZ0cB4LnXDJvxxqcaeaOaQSD3iPSrkHFRYQhFkgT00tvwj
0WGHPcBpXQYsuKmFhMD9GwkKJDZYfM9F07dCEdArluf1uI9tfD1lnW4/6ncoYgbGSmqvarFviI6S
wsllnchTT7jKsw3Yri/er/jPNiljF69iHtUu+ymDtg8QJT0dolbweGT79lh1FrD92tYKARkACKa6
Hp9B8iFC315zL9vsJAzCEfwEx693BopYm6m3/gRmS38P6VQB5m6I/ipLJKp4ttMGGyei1qM51eWZ
HtJ36G3DDVmTp8nU1/c44mCnHT+GUMoSGIAFLnlVwW+EGFjdqU6tVjfoTZJcjtJiWNBNZqX4js9z
8ql2WabRhhrfOEdFt8bLuXCSRPR/TSZAIaUQmmWm67GoV8rJvOCRL87kRAXqK5QEyIZ3UvK8LxLv
YdS6WpMeSs/9DCWZ0RekDpuIBG5lHCb3fE0BpcwsN3sknwgJ+Dmbd/bNCxeKPSdbND0KIVH6ZzbA
oCS27xuX0z1yPbErIm/JXY4sdV5HlouEKvAnRfj//QdV3O1dQNelyvhzq9MriOfBwuQRg5DjcYwp
pbsHhwRAiUMJmrkS/JvqsZ5WpdgQq5kSWcFU85lXgh5Y91Rq5RneL9HWE/nMQ83gsp4yilXgp3vq
a0116lihIwxcR4dt1XWimXoVjKM1jlYdzeATzo1DcejL4Fvpxj/SWgWVSfiNgxN3Jqaw/oquXKCp
XImTxVU8xT/uUICvOLWmj9EYwPiEAJxnYfE8kPrf2PJQrZYLzL4a+ljPThyV2fmBl6C/X7Vmnjzj
yMhocloOTOZk/oodEvY2FRnj0+CbKlBSmadhGU3QehU+PqcpWsSE0KLoXMdV0XJr7Bl7A8qTfZ2P
B4orhSybpfScu+HikEiifg4NZppL4uyApST/lZxjby+qm0rem+uBDF449sAaxcRDkGdmiYXxhmW1
nxtbllNeOSjLLZ07zg4JhNmijUiSxfFvCnco4TpOOebMo80Eh3SuA67y77/0FICUgcOvOArxaY1N
D2OJFHbQppBDd6wFbq6NaOI4lVGneK2WD1VDSw2xIkLYJ9pWCbfXImIKPgRsLOk9uJKOIS4sj1AO
JDxB7fkarYbDPyXnYQ4LwHL1ra1xjokDsgkZfhvvy0G37Y2O2Y0QykXJ7eCLwUZ0fsGJOi4/68iz
H5aEYGAOKA/br8CBw2sQr72wNdsWXcSs1XvA3dvR7NADQeHze8BzMSiIy/jKBSlmBZ2upTJvD2y7
Md8siGb9WWJDY9OeaQFUDvc/B+OL1WJsK5arfCuvgi+cEdv5DcwjC5XMgYRA6VCY5ijsNHDCy0sS
BVg8P+RLCHBQBDC28+wcHfDe4nZ1aHz+h8ocMzCl6TXb7vDZwys7WuaSpqt/bc6gz9XwuBDMh0xT
hZqLKCMPDLGPcM9kWMX45ELADwzaDEh0XWi+2HOeICUxOdMf1OlUIBR+pcugEiXprS4aN/JbK0y7
/blXGRS4mpvTTNm1bpSJrt7MaozROutolWPce+V5yX/lr4BOQHCPUlpvW25DmXdfviBoi2dUdRZ6
kS3SqAe/zxK17DnjvOZiWVAh79z2cFvLqLE6te9dkygmgur7qYDST2aB+UQGpUr3rjpiegI1xH5N
W6+4Zc3AujO0uxBt6V4VN3KiEULFsUcfTIz8DEQTMW5SFtc5OR/8tDtIUoFy4nLgPGZNhkfEZkyz
QhqzpiUnIC9EurgoBa/PpUkmSejwIKFF3nrs8QJgsx1CYMPN7BCBQ92iOnVCa/wXQaYowDS4nQe2
b78EyfH9jVrgTYBOVOpa60EIpgbyGh6nQ3VkeHDQbBvQMWSt8yinrHX05aRMxzpWR6h0K+x5haGd
c5yVM75SDW+JoCUDfLww5HW1b5HsAsYc/6mIu6QbY0PyzVt1YMAoo0KAc32pZu0flvoF6k6dnaDt
Y4oWQjI9Drpk7L1xLqd4cFRDi2rfYHovsf3XCk9ljlNxDv3+y8fAiMcgLTfH8Ee5gcysclpVOMSP
vqPQwLLcJlUv7004XqbfgoY0Y7aACUexL9YWML8VuFmKpY0gQn7ILSjM3EPJtka/oWQlFXoNvyJi
QyqLvBwryn4FVkpVT0+SCJ6efyiScQgvXZ9+kq7yE6dgxC8XKCK6IZa5WGZO6F26uJJtiKX00pDc
qvdnw8ittoTcsyuNMgRCnssyrWe15alAvIKATvE7RLW9hN3CE0PIKT7aunycJCUzYokxteDy42xc
1cSOVWznDcX6v7GNeERX22EMTkO33AgE5BRNo9IBm6zIF0fhvm0Co3WVfJcwgOLeoXnijq+4UbN5
VpYWqAvZYpsMRnUlhyS/48HuT+/2rcKrdRrI0vqKgZByWCWSR1lrAD4yFsActHmTbHI6LtKKvx2k
vclc85YCY0VpCwHeH5OgJv4Z5Ni65VcUx/7p4Riq47pA6hpSGH8anfKXkGSK2y885bI3sabEAzi1
2oBuA01SCXNPARwu2+ctc2KMqGk7Z6l+f7y/mqeC+loRyRbSbsI9PoKhe3Mk3/jlNmAv+6A9tD2f
PovhV6a/Hn52fw38jD0AH5VL8CTWVH+3QBonWsMkoeRbGOM4C8lCH7nWUMPmzt1vGzQvMX1HzHp+
aFJyE0nl+aR6JqQkoeBIsTRfbYHfAG9LoitPklKiQMTsez2VVQEwXKJvwc4RE1Lw/arU5qjcxQC2
wLRD8Ht6eyGEZVPxQlA0IpaWSxZlMoZnjYpAG4IbVOA+4eJKJG5gK9Hb0ndMvSFTllKwmvPi3/vO
HYoRk5WkIlWQDprFHxvcArXMy0FpIaVPTfchhLm0rcLM6HGxkJzafMjXxKPDv6/P4/a6OoHHk7bE
yQl1zVZjh4P6xB/uThiHiovtFc86ZXWbxZeYH+IvduUHhx+clfSbDFPRoE4GAHPl0/UoN3GskYEG
G3xmYu9Qt7N8xUf5FtpkJIt9gFGjETi59sSmKaDy2l5oIc+Y5S2sICs21+aD7Nw+jYE2BWKwched
ANV2ajbT4/ClcldZPAmkkpYxgzSKNQQFdAcSyx/LFwBSejYwuhdjt9hgiDiRduLNeL8uCWkE/LsA
jKJyFQqaZlHmhPj6Mjw36hOoh1JcOsNjs1k9lf9mGgjTtE/Ydr16FrKHQj3J7l1zHEp1Mgah0Nst
i2hoHZyQvRlVuuEg3893bOqpVcUq1KaPAZ3GeVZNrXdOlDGZimsyysIderBNDTyqPYLNhmtyqwfB
zBnoXGzf0EQCDZTBxvNJJz3ZUgxDLWEoxCXdCIVxes3OjQRv94rzlOCm/8y2GT7skwEXHeznStv9
wLTVtMefQoD4N3MZMACMvZMeVxlkdV7oAPjleyE+RMgQhtLdm8Qe7pSbh7FVP9ERkMOoHz2gWORM
5kgMmss82dM/dl8Np3b71F8nOuI7uMyBQvLZnQ/dn85EPkT5n3ZjHfyn8HePnMd5O1WAjbfXaK0D
6zu9ZYUAA6yjmFAyfwVcCutsozTTSCsqQtAXv3/T6Q90WaZA2pG8wieH8z8gh8BhONLRBEWnchFx
XTF5ftGJpnrf3A27mQgu1XiUtscpX/5lFVUvKwWuOtgVNIeVI+ZlYM7igiy5WdY4dC8KrovOCO/3
zQClAM2hGunMzNXZcc/3qj86qVwH0BQUYZdQ2AazW+IvXDBAjwzUdlseiWPRiDYBsA7csvYk6mOH
XwI4WwPnkEqkdOteDEQwXg0p5i4j1Aqer+YzEkR6A/inNHL8K6EKFPyY3TWfjZL4/S0yD5/TBGX7
E+GrW5fU08Rrfld8AGG/rKedAyNEbQsJIL6O+zSjIPEzjGIbgD9srDeK+XOGr47oZcev3touGQmj
ySh7l4HTtWFdkssDc1L00sYKnBFmggCYYkkcB9l1PZZ3azMwi/TpPxZHL8s7AFmiPHFa0eto+iAK
vZW+6XNh5cFJUuvv+0cVH170Yp+GXoGZuELnpu8NmXbeA2GDIEGpheu3GcP6MeqZyoEKBisgUkGY
b8TgbmnQJMrNFPpObgS8VQAJzVW1eHvP5DuTwvKVnN3UqiU+VF3Tie4Fge3z8MwXZf2ucWllu4Xy
EYjvK9CKXLLR+ezpakMIvKsJTUKW7NHtWB0RqhfiESvoNAPVgTW/hT1I9bVsbCkChmoIzDWKGpw8
kTJUlOXrR6HRO7lz8nK4n6oTBDditwCtBr3ROoA4HeNr2L2x+AYqe2Gouzk90rMukOndCqb6X29q
K61aXFEcGrbDXFvFGF1JUgzG07vIvtTIlG9iIrwyZBfJPPj0dVyfe/7gr1pKoG00U2kFbBIqD8N7
sNu3pBM/0/EliJb8JDtJVJAluG0jq1mCtUqlX8j2rr3G8kAZgFuQIkb8fZkHTwyjn4JVkRtR9NsS
57nmhikJW6+k7VOR9OtxK4vX0fMKM2uJk36XD7H2mApndWds7jPvXEmmaVBnY2AYTObGr1uKkJn6
vWilhQ/+BvTmSLxSzobmeWXCcunKdRkEaF4J/APYCseg3507H93zFxIGIp7o7A75LgC1+C0A65bZ
OXhAt7++6H01VLqPI5wAlu+mPi/wy+igHByOxmq7LA+bCngDt9GaIHgNJBIUnUXyRdOenO699rQ+
aa6qJav0sABq9IQy6jhdNi/Prk/J1ebv05doGk0jOxnX2wf1/rW2zunmatlmhPbBVi6OTnNEeQTy
Yp5DMZdNjyhWE3eNvfIjxWPsE9mx/9e25S8GXy0+XEhirxWkO2IGFPOIrQHxcVbGaXigThUH82T2
+xEH/HVNIoKa7u8w+o7TnMVJKmEr2YxzjKRgPyz+jUmMAru1b9cfIK2Dd4EK+uT6kkoufyQ9qx5g
XXmvB/tnIp9LZyCzve760DtQtIG2EGFYnkmwxOfhW/wsSab7nA/8mfChlc4E4iX07ll/9GRu8oBV
G9TQRU+/nXfM/+l7LUk15a5O/RBTG1QX+31bOoizUj4nyk1LVqyNY2DAuDHrUn++uxDslu/1EFRB
cthbsL6IQ29q0gmtXRfOWmKQ/Gl+yqEpWmftR+zLtC3M8sjJvKsZEoiz2PgeL7UAEyB0THK0uhLi
EWUH6r8Jsz7VeM5469auWJemSZndbulbseP3YpKaVWwa4eJ4xqW1YjmwqKlE84n25smLFwxs6Qt9
rXZyhUc6fgKMWYgAd0PT2NntJ2Js0+q1vsKR0J4hH6MFVrsivF5u39Exxzktq5NR7BqT08VrWkWt
9uANxaCfK+xrG/es06TWfP7+ymqoPSF1Codd+J9IPG3WsqpTG0S0w3luZGv3EQ9KnxW0ux+xVfWz
YoeBadqa65Eg+bgm5cqTAUOewAlLvzro7f440hC/Enz65O21sUCykOrMymFsYX30v7RVywT8ct2z
oHlxUhnVeD4GHQYmAd99xfVYfqT1hwMGgY78ACeZCPpiah++8t7CaALJNqBtSKAxLcVcJkRO/uYO
HoubTywIWoTPXz3PK6BiSBTbdJF/76Sid4OMvTcYNowaA0gfNx77nRTK5IodbNj4FoFlvyzYPF20
tLjoacEbWnYkCdJO35ShPcshIQo9oCq/NeP4Hg72hffEBtq4nGaoj2TQcLUpmfllYalW6Fd99AeF
xNwITNL3hjBFPHghMDSrwTJfosCxay4NXmE9WN6xwQfAck23louyiFr3QHBe+K9f6KQV8y8q/vuh
Zs1t85fSXe19v0W8UGbxu+IeeHmBIaaWSg7EKjHF2A4rpV0iYHDNbKI6ZtTnZqpAf30oejMwM1HV
4BMJIElx46BinjwJhfACfBFN0MxqzkhfbkZsJd/N39oqAVT/Mh0vmJGbHOfWBQNNj35cpmK0rkWx
NNDA49fDExSZ1AHymTersnpog9M9tSxw8wsJrGJbRx0aRT7aZWU3LxyjhYUI4kySJb6o6eQUA+cC
ASMwrBEnsiqQlxYeACD0O1hr2WBoczzw1sthkMZWvpK/BR4ikqeID5kRmczcSPPdCv33Tr+KECtL
7MONZuhTaAysNU8r6+NbOJ8VnXdc8NWcOWigR3+osqBY8Fh0jZCkqeTDxHzkpbxcs7Sd2xhEMxWs
TO3fLc1eFPKsMlqeYzRdsGyCvebLrnW0hk26/SfvBeHV6cO7iJ4WXAOvjkvxJdpJW8jccFGpwAVJ
ZvMqECbdQEXYmRZCJk8I0zkOfj8EfQT8EA14yCa86um5OWXSiqnFvcsnF/sbykgW7Gc5z82jELiS
6hbdt9KRuwq3fnqILgf5AAklJHHF65yCJopNcjmOTJLgI1p7ANBBTVHu0XhgfIw8B6vVlJoEhkOs
IdZhA6BTOdyanezuQsTvO9BtpVr3ZZ7PRlVnIvOk0NHuBgbb976x23F5pHTwZO9NmCwFsIIokZNj
4TrT8OHCv8YmbG0duE/6MVUO+RTz3b1qcRXlpsMT4w8vBYzUnUhTCbAhO1lShvMNN9vqkVyjF0lu
QVOfM+hQULpuDTgHjXJDSsdM2GfUutpvL/yC9/vnHV/mKejgv5fd6tBRcG4bvrG/u30L+LdVBQ24
YNMKBZicL3o+xUN9pdKGKVD4gDSGHrbUuWxiCGm9+THXZy5m9bi2gxdJPEqcoykiXHc/MsLw4by9
l9q1AHpvu5YjskZ97ie+uhY32l5ybUouMHKC9SK14cAD240du4PLac2QUJvYTq9aRk8Ji/1CTnZ3
gaxqH/c0bxjvQ3JuPi7XZv+XqPO0YGK8MIkAwDneEwTqHpZxuv4AmkKjVLeXRwZfIagOv7TC+lnz
t/77eWN3hDTD0jA0rIoiSVreQf62X4G7JRfP/YsH4dTMlJIYXhUCr43+Bq9lJ7VrzueacV+uRMyQ
VPUBiKcHGG1yWWuZcpo9Aas0N/bp1ZEhk+w+3fsuZK4ylBMiTeJ0S8nn8kSyMdBdIaP3e37EMLpQ
l6ZmR9EThuv6rkvEaLXaDMDFSQA3Kd0VSyMb5JU4TpgGLKtW8oh4LVH1BU7zZpkFZ46Lgv91S+Kv
tqBJB4XyyeZj9EiuQ9QVG04/qWkAd7mDmMGpbqAP0Scg03e1dnYaFMZn5G4c2hb3mm4X7G3wJcGG
ml3v2E+xpuS5sBIKTpEnTZTxgzAmh6sUNaVz8v4I+axIV7h0fJwVyflL3nE3GMMVAiTNnb16fvkN
d2dGPIxhqtax1+Vex13kB3Wror47I/LbEW8MEMexQ89Mqk+CjRsXS4JR9reif4d3N68fTyqssjRh
71mSSMQbzVvsPtgbnxvG647u2Z4uNdXYDt0QmCRF9IKzyDS3oZD8nyAMaH/4OW8G36JIeI81qkHH
jQCddNknr5NHcJ7jDwXDJScNhSFgZGludmhPPgUxdVWD8Ub2b5HcSxcojERP0zWzWaoRsUQKdGVt
7Zz+r/eQJm8G+r/fvlJuVTweUF9ZKY0CFGrP3uWdIGGOcNIwHzQrHJ6tCH9iHZDtcAx0RCjkHYzo
9xLTexAnOtd2pYhEZEVhI2UdkGp3EyZoUaueK1tklETcWruIATUmZAwYBmTQdU1+yxc34UWvrc1u
koCk+KYeqviscCUA4mqF6FCGWUWb1Dc1XuNPmcquUOJ+BV33YlUKkBS5eHQq5dCJ2+h4XkZk/E+U
XuCYZnaQBpk4/CNkd2A30LczHqjJ/IVDI1m8voSPSf/hqGUEGoyEwkIZpBgB3ORJZqdOoRSv1cfX
jE3Lf3dQAHkoqPHHz+n8hJbHT07b4gHRvhq1/FyjZ7SyE6l5DVM84uU9cgTnLGPmaQ5MoaNhYRqN
qIOKDGe98iAmmzqBq/TB47+5JcEM0b/SqlmxWPw5mz9omkATGW2pL91zy+q9BcYNZr/QkxNogUB6
W3vgW6m+bSj6+gtt89hdrGFlQhs5xsIlAC3c5sZS/O/CWEpb074d8Q0cn/7N/WOI/GTh/J8S+I71
T6mLjWooVy7poo+upD0zEDaAsggNqXEd+eSESc/PPDsx/VkJwUUbrdY8Ohp47FfIhpIDt0JYulUe
jk5Y8DY6e+lIMELoGltHLitoE4aorTTIqlUHUaA5VzuH4lECbCjCdTflqitqHGf+SSDt9dob8u2k
lsyOlOVXdJqyhD8CQ0ME+IgYIG9OrxJ1BwVdipSV9lNLD1GO9oiSTE8rc7qSjyJbAOv25jvlkewB
vhTi2mQdVCKMZgLimQBJHdsHQmAOUs+QyYW/R/1UijHUpV7qE4hOLsBVMXZvx22jDIehF+Gf1ZrD
pjwuftegfd7RLvRDGTth+I4PptiSEg6lDNIuk/A9BB5KG+Qk4lFINYjUHUv5KmL/7CyeaF1w1j2M
jtMYp0ITPxSZolGQbwbN/ISeJvwrK76C2o+jjwYlGa+lDzqNS0bMpBN+bfxt8lTjV0NZbAOiSZPQ
ZGfbDZ2t+91dByhg3MbppXxfsJcowxVcMbYGNU0DcSCA5dMhrH13MC1IwVrsvEzQWqQpYCAFx+tL
pYanQXndwarhSoVkQxycaXCi4BkOGjyK0TfHVSKISvVTAY4kephcPCpZo/Kh3llDTUfAYtsZy8LZ
5qqTY2U/li/c79LwlE8k3WMFGmq4i0L10J27OSr1Lpv0Wgq0LsikKWL/bfzCGE/BXIYzLp6s1eUa
zG170F75H6uW1U7GLm7o7at+N61KoC3Bdc++NWQxtay1fmyBFmR75RNvvLWTPoVcHY7FcvXNEGzk
zSRKJNumpTSIIujmpkCCGcKrw11h/uCn8EX28Efm6Q/Cjt3whpxcPBi1gGEuXGjdRv940n689IVz
9485h9ClEEyd8mdxCjvez0d8Fk9V8OTPA4TTaZyxLduj8p9SPzb66C5yWctaQ8RWU0aMfEEHv/6I
A7XM/MAt7azt7CErwqp51pVQJme8vwbF2rUjq0ZCEV7I5E1yiVAD1nrlOQSIIajlc5qdZnjV24/X
dT4qv/KFJ8YTtZiX5YxMK9UF8ohqP5YZx5rwpXODCnET6lDk/cZvl5CVO3m47KxFOtg0oV4AhDG7
ISBSH1ewnOhHpMvm9EIt38sEtcWV6qFhy8NZkiIxjzVLBwC5/NOPF+0i5/+nbf91XTNIDriRsFRU
+bEj5eosrWKEn/2AHIrIorW+mZo5x+fRhhXGwtIfxKHnD4vPXxaTkun9CLp3GM8E68eu3qPYD7+m
fB70xyE7nw1/oL+SRqTfBj3keX7jcgO/UoHs4jCBxfeOn4W070Xn7QW/edcjfNMp6S8r58gsk5EZ
CtPiLYDEoq6ePT8WVXWduYWC/44W2dKI9vPeAMuFPs8kWAgpX2gkTMloO8v09zPL8At22SE5n/8Q
fvHFdY/Fb1zSSdO0Vru1MdWpeM6JR7TLR5sFd7wEYxHev7wjjDpy5AfVS+zp2Rh0FsHb5pk6MKRP
4+kc99c5CXA2efShygrCmmGonem12MbnsbiNx4lXQ26EZUaoN+RxGJuffI3ansXCzT8vrlsTpzbn
Q8Os0++ZH38AW0z9tN7PwwCDqUiKDlVJT2clK9QiX+9iQQ+c953TKhhvFdpZJU8BhI9DJYk+OTUd
g7qF108VUHXLSbt8hS2KmQ86E9n39yL0H3iw+V1iMwF/ZRaDMby76l5xw0fszUFnvyd2YqBgvlF0
yYYOdJY/QCCHb6j6S2lyf8Z6ShXB26PwdKCs0FUXj4aWv6e6F5LDaYTE4jaWi+/WYDPtiQa8ZKJH
eK5loraSeEA9nhw7Dq189cvle76+TSHj8nBpT0ZGZHmMo+POqu7kpvcIXB40P0aeW6NqXump4U49
3qwguRNo0re2MUIa/rid99kmz6oUuI0KSSJBDa+TPwXCL9QHTqw3c5C3m//bmVhIXBV9/H8W8Bi2
h5KwpgY1gebvzHJXLv3FebIIMQwPj8GFqLdTCCwzdrsR1VbSXaUuiGNjmEwVoTWO6fNeh/MAxCzG
XTtSP59t3DLfrC8BDDc1xQOlRQMbSsmPyJu6h7lTuE06HltvfOKUQNsLS8Sy4FvH9szUhhLnLUoo
ivQCZp0ODpvUQnLNxNKHNaPovFYjUfmsLfS4gtV+vw29wGPB6KsIstuCkkEIX9wMWeiuQygYQkE+
NflNAUvX37WJI8KppE/ysepcvyMfA20RG4JrD9q1uq8P+mAqQQ1iI7B0iEkKa8RAS56GT4x+s70S
8BmlT5tfS5Oo6mdBFo3hjoaeHskfaeAdt4h9ML3qyIGS6ybRU8xsruVpu4tme8W+X7RwXCDcunpy
ZKQL1jhCiEAOv40AT2LdHlviMzgoONEVAmRZblf7aKxuFDaeMIsmQuJG0K4NOXkYsS5f8cvljPeU
iVRLIcjjZyYi7EuBWSbx35g68xdwmad06Ln/G6v2r6mpU51teZMgXOPG3gwsz2BJsF2TPHH5tkD7
TJGiCbzmf7mfAS+pIrGYVWj0nLxGoW2f91tPUjetV5SK5A76coM9yWhVFsEWTNj1ITzqoYfrxrh1
ZHRigpIKjIRG9VU+zLdMzvUOUaqNpj0NwfU6qXKFwE5lXl0WIG2MW7u7IZbnZebeKLftyZkAQIyp
UR1pLBu5nyCPhNF05lzZ8rgVRObveLhBmgSAKz/B+0f/vXcQxSCnfGBOXibyGog0HZTCu0Y7rXAo
LeVb8lNMkUFxi3S82CWhQuA4D0in/AYFBG65KRraFQfR6GtY84WB716BxkCe5s/Dk1ck8Z7z1Jnv
DSP17ZPacZG99GqcViEbJxf4j3mDxbVf/C/VFBjG9398DM0qUYlMb54XlwXFPBBVoq3FPBJ8cPY1
Hrjqokqcmk0NTtY56P4mdHeYD2t8GVUj7rONPexeiqjFVJOdz7G+7NDzixWPIyp4zmfhaJuMWdOi
Uh/olhJLDs/CK8UdsGFatdGWFHHF7aUQ88WGv7aa18md5Oe5ZOZV2Q/4WL5LwFF9Yztx4bFb/gQd
mn0T8l1feC4hK+ZziueFGO6Djhqj5C06Z8Apgwb4ZaFHZp0w9OU13zmgbDM6pQIIvKjpa3LpUehs
o6cFjOS9U76uWHWYgHNBaaYW8yIwUObDoA0jJ/bRrOcOPBJ6QBI4qCX2k7xm8xB4WASMyZoA5ztL
h7b7pT2nwfBkOCoX6EZZIGbQC5w9Gy8P783IRJPwhOlSW6HBfExeHiHqUd/+O/4xPZp5EnnZSx7d
P04nUSjtf5z+jo+4ci43Ooz9swvFuYie5o3JNnnZLr/W4AgsJchubyOmcJNsnN4KrPJDUG5RBV+L
OtaakJXfcb6Il7iD7LrdqbxfCN/ChH+zUPGljLZ+22TQnoprbe1WEdiS1GNIL95lvNb3U/rpGdBf
PcOwO7g6/2tivtotwuySl+NVy+O6rBgcXpu05ek34gZc9tvGX7Di1R1xRNtlD3U1pJX8HIVko2B8
GCNepriOxiCFNM4zfXJyVJR2hBUfz6xPDtUgDn0qeFPwF1WcKUGbGLNsR4VHwsRtoWzN9MfPkHgh
T/xsVGdblPSV9eCJ6joHwBVBfqETWKtqdKUqDF/GE/K8Q06o+mlkMWsAczPUQk4rsbMvFsF/xUxD
jWDzevsUIomYp4kmS65yqJYWOTr5E+y/nYeK/+zQFQxSqD8Us9Sd+G0cYW67670wMyW0xc93R/FY
L42r4yGbj6z97RkPoLiqjvDY4ewp95077jcjZdTxiSyQix9xwacq2/mV2lH+pCR0OEjDiKzDSkHY
tI3FEjFbcbX/cSFYxcMhbbsHMBntG6euVhPwbo5Qhih8c6uY+2fXo3Zw34bs2H0ZAhtef9sd1M8t
wpR+WGdUPEztoaxXELOcDrqg6EuCoFOpGMRbY6kbtakfEocXbGeScADK47ras3snnaCQoJYhO2Zj
JeAEZ4NrxtZ1Ym3GOGtmprHHMA+KFJr6LIZJRq5qhOxGouXs52pThR91HOjEZKQ36KADweM/G80V
uZIfqizqbLUck80m1jl62E2Lz5YS/wwe4+uaJC+YUpRlAyPtA3JVWPE5z3kTrmaGhmDOLUPqIj3L
rNRfTxlrOOKdJYpbr8kLvZ1bpwKgkoLeVvJfcfIpenRSZ1vdsLxkR3Zvf6WoltzN5Z7hpJHzZNX2
3BqJmSt7uN0xkzmwUaoJpBTi3uopq9iLsz/WZw66n/tZHmr0RBzk9lsT8rsARb+ZuC8swAc+Ae3m
DfvHK52SfkOlmJ1t1bZkJPyrxh9+L4zYNyPSRs9O8F7UfC15to0Ywrm8ukGfXn/4vTeHj/9BtCdS
JHXE5Vyam/T1LRqJwnNcVX86c46284cBiLC824JzDK3Uf1I+GX3N7cTw3lDM0TwyVTR2uRAxJ2PS
Xc9x7Riq8BjlEXAbOoyTn7gEZhg3WFpGRIyUhFq1mcHttkcNU8v66kZYmuoGk9IQaaT6YwMCx+IM
OO4dXJm/z4LkuG/D0jkqPxa1pWE1DLJ3CUKeO+UMMQfYrUpiJiXog59AqzMEWiK/ito36o6GTXxS
qD6OB+rcwoRQN0GMbDQ3oDXXWCbfDYYVIHMD+fg+2Rcs5uk7K7MIhLmNKy3UEmqhOrHIB/Z8o0uS
s/AcNNVdPn+OnG3ZtX0vOVgQq+FJMFwN7yI59swJ7a2TNnh7VxVmvDDqtyAD8J2626e6XTQTsSZv
BzS9idch51mUcj9Esf+IwKw+QCnaJ1Hc++iuHeN2rminEdf8GyffLXda0As+iqGfcu7H9vGpngdE
Eh84TG6vLBvR31bZRXkUIksJqfkSNvtDX35d0AroCsQ7xKofdvbbyJleLv3H/Uzj9DT3TVipFRLV
zNlU24CzM+HRtwdjZrrn6jt8uC0znH6ExZEGohuOpNQKb6sEXAeJoCl+uerG60Tj/zRGLecMVBpZ
HNTTCVJu6frsHCSIw4EjREV+pnloqYCte++aoA4rx7dP3XUgWnXIy+YpVmFv+heN53w4oR+NSk1b
0+bDPW0b8M2RHg01MD5OrJoEMqkCjohH7LPBHOvWIxYAE2Q+WW4dHX5ha6pYo3A6g3NxOQFxW9nG
QXBv3SUj2ExYiAY57dL1yn9wEMYLqx77AXFTOaQ+y/dnnVEc4j4C8tpYAG2odWJuUaicB38Vkh08
UlsoZTCE5rhrp8mkUgV0UKx8mJ4TVdKjVE1ayAd99SPlNlUrepwdcFlJFsoAX65ZCBzphmWq7k59
51Xi+SGlcsTZPk9B/gAS4MahZvfYx4FzPsKTDImq1f1A5dzJCoBxI18jx6agMeZ8PLt5SENFmV7I
VQ2tIE98ltwxto7iBima9pE24UAkSaE7NyecliOJDI+tzSo/gYnee5NMf8dsffvp42ZuoWHr7Pkx
CLTsM2DkyOJi/ZSgoSvMaEjZNHVFQetmPCt0HTXz0i4f2+V7lj0C8XOGf50Ktn0Uvq04Vt+LPPVb
SodGRoulTvV7xRGI3jxqydUI3yrablh5ueZ0YrynysGeXeG8456VGkn6CSZlVHURBBKwKg9J3AkB
Nomy1L2a0ThsofLssOwwglg+sfCRDT8CbasMmu0CK6slFWjKxitxj3fr1xEexyah9ajCi/ir9f0Q
QHq/9JQdWZ7CAtAk+C7EdPxfuXsT1XXSwX9C4kq9oeyvUc/8NcFYqSvGgJfFXBEtimKvJJpK9Nok
cCd/yg1DrSiPerWUdVAMrWpV0+sTQRQqA9r0H4BLQ6uYR3N9ahbp2aocj67iNMiYMlCl0npxWFxH
4tELpchSSv4qB4KRxjZYM9MwUbBCzJ6kzpWUBMby4IEsDVebKI1sUFE3aQnKfHZd9qEcQuAEZ1LL
taIGKMADCP1h5SYC3mWEuBQUqSMOImUoVrZJ0mcjlmlMU2eo5SrmBG3GVMX1TdLHtBuB8gUljVjf
en9zOrY19s90wXTfvQVZV3YSRrwtvx33qHcr/EdJ0vWm2tu1iM5wp0Co+DIEkH/Y1cLaGEzjJCn5
cFmndQAMT7LdutE1y6SITvNPh6dVKIL76ijWkzYNbNTqd7GQOlpmpxDwcpUEQDyYo2Fb1oiSv8rg
Dvp5VNVaVpix0O5+xLhTRB3sfgpox4QXRFyPihAM1lT4Qg/0OJEn0nHXUFBBisMU/BzxF29rNUvy
2IBGb4lacMb6YQIYvQvRZQnFcvwpQsThpri4OAi8DDjTSjmtGppYZ1wsV98eOTbr8ZYoXgI0UeCN
PJvxXbjIAV4zXVF3FRJyJ1Nwtzw0GnO7iCLs7NAKIVHpxj7HAxVAIzBpbJhUhvFCYvtkLsjO7dq6
H3D42pFSCXBwIJiiGKHeQTSnK7VQllZridkL/AQGTlXCS5MWRlOxjaQzQUs4VfxnxhlB59hJ+k+c
JoXYiIk8G7QJsrHJ8gIxprpbEeYRlHudBvDQBbSpdYaSQhBqndwk3LC+fjnMXYlZCqYpZ3PhzfH1
Pa8kbhJQsZvwKOzXGWH19LNBrIVxV0Eg5oWdHPrqhNyAoagJTsne3iJdGM+pwb8+PHkmmSWYSdSG
TJZvRNC6VtW7QpgpF4gVxiHKFI5NoSKFwZSqQ6bKsuVb/nU6IELsJQjUc96PVR0t6emsSgiyu+AH
p9cBGsfm90b4LRZoe9nrtjGEC6F9GDrigckwrnS7YgI8PUw/p/gRRhn5PRf7ecus88d6QbV6bjD3
j226bc1gfV+/zG/iTlnafxd600bfxn0IpOJmrMo1JZlJt7An8s6ytEiQ3m15FDtNXv8eamLI2hwM
AIJOwj3eW9gAv2PZA/rMK+UxChzKn4xQm2xj5MtyDuCXMEfJYawnpWcRVfBTSaxax6JBB0aLczGL
Ghe2nWX90ZLXaa1+EAK52VGjbWf4BVf2ASDy4Fqf328gEjB3uoYACuVaUyM8RhxQFSR1OdldaMj7
1S2TT0cysBCN6z3KBrh7/repGR2L9UDrJ2xFagEApX8F0xxzpJvNbMqdWevJIkXJnsShzjw6dvb/
mevHTr1BC9VLnkJ7tx2h9QkY1gsLE+UVPAQml0hA7spfHiu4shDk23kkge0/RvY9WtFmDiRGEexI
gq+LtvX5jQn7FtkwPe2cSAisnxe0/9Z4bk8OJTIzRB4ZVF94fDw78XfoakK9kjMjboCctd48zkC1
mMGRrJCmd7D6/F0kvRmXO5ddJY/zG2xv7wMrcjMaw7NOBXOC5eN0iYA+DhQE7yyx4TvTpRrQrD27
0e8/P90T51RWIronO8t+2abY6VwRPpM8TKYKWxBebdgMNFhvMubDpnTmyDq1YB4CIdtaRZ9lDm6q
SRH2vVE8iSuRL90rNBnRaKpLgfNiWY0W2gQdg1uUA80QUDRVxIUFBdwVCdeL8UHBuH8+mAOjiG3Q
9EDX0uaSWjDnevRw73TPWYJCfhEubsyoglW4aUvhzi0ZBdc4XmjHOjoyl0XIi+ts61Ndp/KTf/Sv
o8gL/R3BB5d2VqLU9qN1I1lZgeesu08O+qIV2SDXYphLT1dYQeQy+zeTp9pMUs93esVRGvUKvpDS
OMJ/UMwFKcMUXcVx4TQVwdzvatLc1oMETy6KANUX8+LXRwEI3e8k+4ZAD8+49a/YqcqwfrFVAYkM
k6mNMzfhzH/aTfh8RTn3Anhox2R3NC61ZasjBM4jSxhwiuTrNhvRa0ZZrfkFLuUGCXIT/dfAea8U
Oppj8cAyLTwBfj9UVno0IbWQ0wsqSuJCSKwBgGd3MwB1f27QdpvIvY1kQhowk0AdPFOY2UIESLfl
1jwwN81g6K7t/A2iQEh5SPhpk6AfCWNRqyuBqwsNca8boy3xoaB//j4PWYf5V36ybMUJVGZkV9CE
EPj1IXiq2l8mw72T+Mj3hh/6L/4etvP43kjzAHtXhpOHKOACv1HCliW+i0ECZ1k3wK+bmrF0C7gG
UANY60egat89sLtapKsV5/xKiG6ebR/Av4c5VLOSHX+bf7juc7CFzLb1DaqtioxN9dhDikjvn2pj
LIBCelL9Wd7wQ/KN+ukgUFpzXPV0j0Dhv+pHV4S5iRlA/EV450f9nCfyW4u4+fGpyLEMRrTLgqo9
Rq+saEhcAWUxDk0Ak6hRn4oziTG5KQ1tp05W0UqS/7SS8B05r4Ql8fYELvzuxiGy7XkuZAX+TcC4
ptashwv5zoGdg7gD8y0rbVG+C36A5oTokXAVu1jil8gBFSn0va/Xt7SlmvkzmyJsnZ5vVVNmYDU9
Tr8OLFb9vHS/WRZnN450nnKsr9vjXwJXqlFkud/stN4lzUzijaJal+A6a0KAabx8W9PMylmYQECF
Q5jhhgiZfeIDW8QEpB8KAXWCSm6l1PAfZFw4XC5ZUDSr6X8RuA0KF7qiW3/e7F2iF6jpc6zjoWNS
SHLm5b6XJJXnZpePPk2dYScY5Ux1/WfWDIYGZthxe9/OTn0OuSUz0m/V/dnn6SMiMTA4M4ShV3cO
FMgBxykdty3qzkkVeuxnODzh3tv3QjJ7+NN4Z4nIHoftDiKNTxI9Wj0lwO1tCf6Ld9Ez9A7l8JCw
0WhUf4feKngqBs6AveMaxTuUJ1oKsa7ibcnxIqo0ERFilOufClbUBg8XY3SR2oaWGTkLDJZmud++
CtLhgr37WrKIaKwSxDCFlKsGBBfjazLPPkrQDHLDT2Altm6AzrrIWZCqJOns6v7fiIcoRlYFcz2e
wlqSn3mhxdj+wIuKpyagelwWLcejPHXxGC8+qWlagcnQh2VnXvUwnlibamuqkKKVkssMk5JhjQYf
lqpd/qqy75Pj6o1Rs4eO8Pfzzc8F7AkVfb0NJipljelJpEJlbuQDoqJbf3lnfuunWt7zPqyVjB39
Ykg/NNsfcVsdO5hYHEt0Z+PAKwH58nLx4q/s89qvpxFLkICYNghD40so/Pjva9ijpTE7m8rjU9VD
lZEdgeYj45IY+gQIUmqLwkRR8V+p0fCHUrOePsMKNM6LcbdtGBbSzeJ84a7tNeDkicReeFWs0xQd
JSxyJkn/t2ZyV2iCTxYjkW2o37K1keDGuiuYzx1b7IYLKn/0eDaiIejsnSV3qkSk6jPFd+AkqR38
9x/HO+MfzRzga/xOzcFmyj1tPX4pY/7Q4SmgOxEFjdFae7Ozhjq7FG5+oUe9JMlBx3gv82OyPJ7c
fteaYsWXqaoY2Yxf5EeBEzxFdmLR8aVH7ZAuO5A1jRjdBCkGj1SIVCLoqHZvmX71lq0/Dt8QfxRI
RX/xjhm0hD7NDF2f6hu78AsoOPvoRzfHQuPpJfgLd/dUGl8bxyffm/t0ZLIYorvxIZOZ1ubk2TUZ
2RUQxZ70Yud04jX8wUrYIWTChpLtf6PdXVGQRl7lwZkpkWscsj+Q8I0x0dcMG9OB2Cdy/QM26nAu
z9VS4Av7UTyl9ULUYACzYbHM7pAfECcL/X8JFyNKm5mt7Yo8O+wmT4D80zo6APp76C0RbCzhUNVm
YhkCcsBmvf9hD/fTjoePa7F4mrX3Pv6UVQQltmoFaL4v7y3wy+K8NAvDZUSKFStyoU70+ee1qyEl
M4/3OlNEie7j+lS2SMs67W3c7BzJ9xN0m2BoJfxv+ykAe+GFI7Y5lI5Ym9MdzN6Tpw5uKl8k6YHy
934MZZ1GnL5FHBYGMd2lnxGt36UhZQ1ENr9ldL/8d2WImUYmCLUCdpPEPcfqdqupMG8an3Zo+7+p
i2TGlAlddn58MpL4In4Xf36xLTdamYjFmu2hfW9PtZDnJgAMrwqUJWTjfXM24EC2Xd2UiC79Wvrn
9GNA/jqHpQgWsipma5mXwCZTqEJeHOlzJIulBEW3PxSK+gPNoP7UC2238Zbf7CClcFxFAuctFQcp
3qMpbDHdxeW0PAhobGq+McNcYgLCZCwNtXls3aTlyPInVfWLu3eJE4NiPHriD6l+ryuNapKrOyEu
iz0pqDsJyaHhoMXTKmzHbF8go7t9HVBGkXPWNIye3u1pLZLwTf93rULPheXOj0RNMFF8XwfGGYt4
6tFJhByYC7bOSNATYNAxpubqP0w39oafhuOcIBsBtif5+RI7MVt2iIyKyBF6NZTT1H8W6mSoY1zO
Ax4VGgBJnq/qsKXrcLeXdMLYYTmUgjtki/7Qg7fWLnfMh2di8w+7VYjMbZLaOk+NyAmjZkBFwhmn
Nhx4AhwfVFrWL377RDLVfzUSuI7RWAj2F/IdA/+rPYM+yFsfVuyr9Cq2Oqa/eqUnG+izD8au20gl
xniCg4gSwHGJJQUbAUp6fhadyqwSCa3qanZnLuROd46UO/ZhQs2nMfvbV+grUzfGVvnI7tWIMm10
LAql9tJtIzSP5mZkPvUlFBrVw2uB3Hu2H9zPrsXrxAxu1cc6sTmomT3wUOxjpzxl5XoZsdlZV4xC
LNKDNpInZRlVkG80ObWpuXC5ZvAk4HtEfc105vwfSGMlrFAKdJ+eaQzt3p+BE2Sk17vx4wLhaQbT
rpLFE9K0n3JAGLE18qGD32yOZlSR19HUnOJxVFxuV3aiFOrUAYWRdx+UnSY+CWBGFsTcUdLswoX1
mDZLmix2l2RbS/OxxumgMK8aE8GrrI+ZfAKTIPJaDOWCvJHhFjYgRiGytvLtuAmKS0Y+9WZk6U6r
YT3hbIURMJIo0LNXUd7pHzoWp5Hd8lRb/YPHHBtnBfD8KZXU2E9LOyEvq5OPyCWwrggZQpL3rCbe
vCZt2LQpcFnak2o20+nt9oxy0nPhTW92r/y//05CSFqs1zbTQEjdqAODYC2DdnucpgJp77QXT0Fy
SOHTVW2ET8+gRuoVNrYk23JeEVjpY9jyAkqNfNcAmBJTbRXzoi7a34Hq6cQ8+Gq7uXJyMW86AgM5
9z+/vV2nrKlAjz+ph9f1bZd+Fn8KBd2xa3+LJBj6FZ9HQx/pE1zJDc07dfr0KPCZmd7WVpF5El7z
BSiF8Mz6+sOgNd+j54SpI+7DO/dludJok3f4+gff32SbYkdlrPRsu20luuhq9g2R7swFNPPeR5Nj
1xGLbGPNW4WcaHk0lNVz3WAGNYmMaL0F4gy1wW/DFzsLAT+Rln32dC37D46GSzA5w1I5gmlRZj86
bslTHrOEvCfPnK3StWPqP6peXzP4UM+SOyYd768QCEJDVxCEUQmyvUwG+4on+PZBApXNO1cq8FUo
3t3PYznAhufKa9rLSrqXw2d2rpXp5tZQZDsTX4G1HB4kScd8niZKsvTyubMg3N2khxnDMTWncjgD
OIIrcLchYaOdDEIjK6nInRhiHG1KbQC6toVI7V3C9IT1QnXsInfotat88KgCm1CXrpQ4W9rNkdge
mn3c7U9m5L5EJCFg2lG8ntJ34ptOE6oFOu910pgLbzNB3ydwfSZaehkJ5EkySRSeMLBF3hQn
`protect end_protected
