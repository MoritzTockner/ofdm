-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iYUxRc2HQ+eMmzSfmRdp0I5h4gs3Kl0PrFGu/MeXvWN6z3kxPKAE/tCPEev3gOdFhkULKniA0Aqj
52cLbpYkF/H0lGgVe6A8dG0f8gSiH0hzOYoCHW5GWQW7Hf6GtQir21n1wlv1/zvC4I7768T+QzcF
8unoRDKIzGj1GGPUjgg4t6gG7zSOMcvRYfhsgUvF3FPkSmNkNMAOVxzq/TXBESv3rMjTdZ0Pd/l/
7KZl20cec8VcUKR+2LW2b2SYzoXIkAh2teg5mHBdvx3nawyM8mfE9UQ8aOHhfixj4pHGCJqJj7tl
FjOBRmcTMt6L7VULuLWquYCo8gLsnXApTVUIeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11952)
`protect data_block
kphg6GHTL6yIgIWJHPDg5JFiHHF90ROo7QS4RZFDgx9tNXlW4c6utU0GGuVjUVzgFrY3h/VyDzHF
D2VCZqCj0GJ9fkQXPPMDnpz6+5JU91/204+j6B3CwL2ZQ3FDNXoillrZbsFrUrohcelB2YfcWP3o
V6PhUPTdmp/7i+n7Q8WRq0paJcLe2dCRRCWIfaqGRYqRHH841KGOyebuJ2Z6oR04Q1ZeQh/fgZeY
Omm6zEvyt+8jjNRMdMQOIK+q+JfGNIvCGveTh9SmuHZ8XXzW6C+56dYHZTjALNbA9Pc4R8ubfEBi
KesD6wOgERr/SKOUnDxw7oN1rTwyEC0bcaxWpwVc9CbHxa9aseZ74eWhAoXygNAuuDhoR/0ZSWL0
uutgn0fJgTSfn733OqGr8XvnsCli/5IgbpkzKhzR/JiXP3KSeQKJhM12vHXLQ8fZojr81K2dTbwJ
yNv+O/qTWDPpwcFeQT3KgLEo6sMLSiFyRdXp1L4+R7oA5RPoBtCw39pBbRQyDnQXsCL+VbFGlxGR
t6gtvw+tbXAFKBAgsQPCENjbGrmibhi8kbfnbWBUzea35TPndqC0VE3y0UyrwCf8KAkLeDpEJ8ki
C8ZGIcENvqrV6A72sY7jk+D738g/tK60++f/OB6AHeOVXV0U6GXuKoZ4g92PAXQoS88LMyKeLxvI
hrKy1sgEGwaHHZHHV7CxRnjO/N3lfjKGm2JuWTKtgeCBfwsCpGeb2V/bBPftQDnUxbMwSaBgJSQj
b2mLZW1wnroMVMmg9IS84PWMmBSvX9wScCwrlqb9VxvH5kwoUkCexUTWn0W5/tU9pCRvLgfWCVE0
CRgDRw6OH/CiGseloz1t6j0sgctxz7O1je4jTZcfHQ9cNwPZHrUoYkrG5/okjlYr/Xr89R63Aaj+
oKv5zhkLHyXPYE/VIglRdSi9w6266RwIzKD6pA3txgMzccxKjqJhM9gYEqUbuCtuB48vIug5JXgF
SohP92vDQaoFu8Yw684dWhUdQujzWQv6s8YYx+aKEkbniSpJVvhC7CiEWVqcPMpMC4v4dIstCbTi
A0o0grQwPjK9ItGtMDce7JERX4HIJOzRZQyaO5o490bhijkD3onSntSERjW7LKVpWWuWg232C7cx
b4yHpVscRwHwyehsnMyAsoSq8htg1Nriw9N3Mp6SCX0q1CN4kDgeKZxGOGEGfUjj+2InTJ2qxOKm
tiZeoYfrTRGGGzciMA3p/1v9bz3zjh2StjjkTQF0d3UqJTsDQnkdeGqgc3VqdppHAHcHRx6yK5Ha
TZALl62j5zex2kUCvD9zfiacgc8GazLXWycHjIErom1l1BplD+/Xs/WEYCCIACyEg8hJRsVNYqqM
ZUM9cz7HjVAEdGTaOr8TMrLgihDbGGvMF1npaepw28aO6ylh9/cmsTRx0ll3rGx+4JhLm9B9fMK2
G8+GEsCfuNnBxsVemZXJ9n+WDSIJjTdjhRyPK5uwiRiFCmI3tRrmD1Y/zd9M59rzhdoaCobv+ZNB
IFhUBJe72blVjKZV49lQyx3vAxDAUu6iTHMIbTMO37i6AHhCfOkN5EJzJcxTcqFXNVo9H5smzFfv
Km8udo+D4kNWpSBduD8tUf9L6dwU1AgFLQ4SEOOP+VU7jgP6+oAUVMDx3wXIoJtB7Mi5sTpxRPSj
nHNBUQqNTiy2NopKIto+ZL95w+IY8R5j3Z23F3EXRYdMdfYyGKke/sDTXxhugTc4yUGWYsLRxPp2
GAN2Ybqt+q5JNIqW+CHNAHD8pNrmRUwGSOMshlMzykZnecfmyUma6XnUPYxlFD0H8jiJiMNDUCaJ
MlcOlevfO9e+vQk4kNtcjL+S8knC1GdsOn17uKiIWzhKXYCC1Le+X0girejkkpZUfhMGqpqLS2I5
LoipygoOt7DVlEF9e9WKe3NMeOBd02X3eFtPBFyURbYr5I78V6HI/IZ5sKYf4EoqoELRkhJ4mTB8
SVxE45th09P8LCVHtnbwy8KNLBED6OTvq1d4AmRFbIyZ7tH+B83Z+p0hHZg34UG/+7VVZE4QUcny
SdRzH3RexHdsyuhjQ7zAxjYG9w7Z1Lrs6j33Lby2j7cScUZVvcaDQ3+zjTqxL66y1shgU0Jh926V
OwrcS+ezo+0u8YigR6srSQ+gfilxZuzcWfRmofrEov47EffUUBvQmKvAOdxN1rzREEbv8mpwqALM
XmxjTqrdJyHSB6eQAWLDLW/UhrNmV3enyAEEoBqtMHADAwZZrkl7dVwWuE4yY+qD6tr6jER/xvgJ
Ek/EBuYhyTEbIGFzlyyuv2pZLkMgiTLeCJ/paen5dVWlblxbJL/jwJBVITyPgSZo2G1wrPfVlMAY
PZrKBRe2tHdP4JPwRnqDXjm0zqICYr0/VvWf6CaY4DiSrBkAPIlIYKZn1BuVuQLNtbhSNl2BmOSb
Kl9QVbopW9LSFBCoJKaNFXTXvz5EvSdoUH7W8z00Lt9DWN35XsGrbacAjJBVmjduD7czkWJzCOgQ
8WU0ZTeQoS8FPoOUb6irJsI1LT/Q9VwUeUXcXCmPrEzXN3+74nNo8qiPAwV5ysgWxhYLSKR8Fhbd
xnLJQ1HD6+xuqCPB9OBHMzF4TEKefMG8lUpjPGslW9tSUU7vHPkDU39D0bNm9bRgOYl37BlIMvdk
8sqf/Egr8ZnLZZeAL2pGo4U+pZc0pa1DohL6vpIXTi55Zosfixi/KzV+vsNSRW6UDuzogP1kbGBL
vGH79HjkjMJr24VOF1yBlR3WqRGDbgIYNhK2tRF/XlcstEqq9Ogvxb7IntnE7STWr8qRWcdSJ48o
eXMyCtu1tRngAHbM5ZhhwvNzf+aH5V596ct/EgpPkOZwmUnAa5FuKjnKww3+etFcejs5nCtxnnsM
y7d7JjcbGDD2AqBlwmhQ/hyKnedAU1t9NIYhmT9SrJAUj09Q51LBoPvF+YQCq4NMkgP+gfiEKP7k
GOzulfWT9aYHxn0msHu+dz03y3OfZUl9JPtn+M7MnOnmCopaFReZiRnAVlYGO6bGqDiDhG8E4QtD
73nUYNNXTuVps82/ReRfKr8HObteCdhhLEi2AzYe10fkzbjMK52eAhM9kx/r6PSAAXiAI0ShkKB1
DG7C1JX7syE08HE9scma9hdGG2R5KGXqn5j7GhqPzDCkpuQ9ldZ5C+3BtJH821ZqlvJ0wYbePvjq
7rFGeIhGfFuoaETZa6aeTz1Zom2uz5TFmu9khFIuSW14KIKusv26Yrl2H/EwAhiZF6g9f5S5cSNd
iOU56W2hfjbWNuPSWXaefRNUFghT4mRNrDlLDLXjh0tBQvUtPh8I7wL/VVRei7UUTD7ct/7aOnAc
CsNVvR3ELw9dzy8Gnaal0pgrAprb0lcEur7J9Br795fq6BvQyEzcn9FQK7gmE4Erd/xf4ubT21Or
vEbqhEJgXqslVCUtoUaLoZDbCWPRElafrxcdBi6+kvc3IbHayp7vr+sLFceQXbJcuP5x4oVUmwhU
CioUxnRDD6m1R4uy5P7cofj9lbinUEQx59xXhTbThP+z8EG7h2i2Lt2yHdFrhusViJqbyZg1ueTo
OD6RlslvG9/3FRte5atR9qhfpln3uaM8UZSWelyVk0qxDU4Sd07lop/xfqYbCpSXZPJK6K14Qh4t
23M77nRl0bg4j9PauDIvDdYpMabEo9b5P6rX1y7y1fM9teCeLwpbq9P+fSvCvA8YYBCC3uFNjze2
9YsZ3xD77V25C1Vpiz8KkbZz2wsVz556LDOTJJfZSO0pib6QOCWJvXOicVouLSZVJuw6wVA24jFH
2ySFgoaGvOJuXZmdzvBih/LRAp2n/l/5mnZK2IWm0NkXKBd7KWDOoUz56OojvWk+0K4EKsZ6nNVe
HzAZxgQsafORTwJTTNGVwOwlhS/oJ9EFvMlXYaFcZ721eNnfIEHfWVvXYI2GDl3+WjVw2qtzizOC
HFzNazpyONgSqZ050UcDyoWsQ/KW0lbfOxdFVTxu3o5a4N7KPruRbviJgTS8vynCMLRI82X0Wzeb
HdKAZzW6tsaTpAjmAEK5RPVx7qpEOmyYHJQL1/z2A4mBFtM+seDtRlhLl1mafde4MEVxG9EAd63h
hlWAePVPTXcrNuopHARdguK8rTz5HCo8BipOPYFRGIavgaBJG07yXWyo7OuygsKOW1KsR8gqWtgS
HWdyo4EPbEGokZW4r3iHbBq1tRVb63dndEnzvJunylLVOndTYhSC+3xOiz6088hW4+GRV+QKF5QD
j3YLN/2yK5J2+ioxFJHyQvyvW26IfgrQ1sXllz9uhmtM44I8v+ERCQNGigBQb2ibuGLXshuJ6gbs
7IgOumTJuGZ2B0v92nC/lxZ7euZVSa7PVsyr9eZrNYk6wifZApFdstNU0sRDxO3REdpUO5EBZcu9
pf3jsGuyh/k+8jXcO2tjm9mkj6Dn076ADT5GHhCgEuBFNkLRMonCfIk4Ok4AoLFOp81rK1OQGZ29
Th0r61qdpZOvtlR31uqDLYKztRYqUm8wOoGUiTkS4LkfdFr9BF0ekdcUOd0wQDTTa0F+UjhJ6iV/
sX1PO2Gj/DTohwBjIrA8Gx/p2tvqrAjMK8RymcH0y4NVwCEoo60Y54NhNuY5W/Yu0OWZy7vmseRE
UGYn6UGZ+466vDN5N/22M1Pvs/2Ngl7xMMax+OoQlEAv2ekaDyksm1EgHfnlywXH8twHxJZNAPgS
Bsj2AqYyMGLiFMQKFSrwkkAFNE2CQ111umxLPNT7teIlhw3GfEe7yDIRrP6LJScUtNpz/wY5qfKz
AQI5evOYZN2nJSt9GySSbl1sqd9pC/T0LGii5eW0e9/2IMjwIz0LaxCMoCea+MvBiZkq/58Mpef0
11OBxzP/y5SEesvJ3wGMY9+7YZr9S1J8kftd9KInHEKy9nM/UKv4oFROyfFIX8TYAeVxfzL5bBv7
2pYVrvlKnj8Rd9nXHl3rKwBtGgz7BcJsKULLbUrRQS19HZIeUzPPLva4p8ohhxT6GHpPyeWChZOW
gLvipKGvxk6jOSldTM58dCXu0zhnEuslpU82003Z/AyM0PnONniF9MPNIIU605GAu6BQIft7aF+F
pYurOfBeqHLp5HV5Na482IsZaM5jeEjkXVkuZtFvPKZQbzr38sbKseCTLTKMGeFrN5gnFQXGPf24
e1g9jKyaFPrlarxCtOve+bFaXZnYlvOo8WWRgynAlG0hF6gbYY2LyG5ekqRVpQjVoaiKLdyDRv/J
n182xhDuF4bN41BopG+XDrmrZc8/KZ19kvrq82N9o5YA1wi4dFt/Z2esfHHF7tmcDUf9ndEOEiKx
Do9OeDmmzj6EiIphueyTqy36HXBIz/FD9SnJMpd9AVkZZD/irV5k0UI2lCfHu35FlDcUUjDoXF4G
L2uYAWInyEyoazXxDMif92LijwQwiINzJYRrX6AoXOmQm2DRd5S7xBIw1Zewy21cChCcnBGGHS79
ZyerZ6G2OMUZmCptYzmVtntYmGNSNRRKHeSsUPyyLx85lrLx41pcg2ID5F7+XwdsT1R8L9bALPL/
HroyaF2AuEvjaRa0JWi++CgOfY/uujpJJ/F/UAiyTMHpTyfOgIXSXLecZAg/lzm1olA8tm1+ZN2G
jsGmOyeFcOGLPK+S263cyTUGKtg4GgYbCnDjBybCZSEBw9+DG1rbAD+dp9RQ4FNunMeKMc6ufDLk
kUfzx1kv/Ki9xsfOaUfUGv0LLExPJEnJBfr5Ik0Ycff8ev9t3n1s15lmleNMqgoWSQwfbxmjNn6L
+RIYwGU7ITHYZhEeBlWfZ8DP8TbUIKoHWIV10eCq7+/GOnUYJ4v6kBsnXM6shGhj9GNi6Y1U98we
ry0e7DZYrSN8E4xsm4i+CyX15YKpfjuy7SCwjTqfcipYp10DiuiKMUZV/mQ+j5FuVJlllRV/bpIo
LNt2PzVaBtRRnO6EMv9dX5zMfenMbt95KKsXLMatmlbInHI3xqjwApHTluElNyaygHjRY1Muj7wR
AwBIU7FGzIWIaL30a8ve5NC38PWLz9jY9czQTLm/iBVlf+IZSmhMXcjAIexX7sAlChQN0VkWSjy+
hX8Bbe//yZJu0w8tfpR2bDma6uVaD5D5IfWrp5YQHVawNoDUtp0Ic2EYyPwfrVzzG6FvOEoefju0
C4/vxV5HMT9bE5HL+DI/vTbX0fixGXgKQkE8gprNWr8qn5AbF+E6Heo9Ch5StDDT5I1g4mgQ7CBm
NkFNltASZsevLM7Yv6K4NuCRKOHbjf3bY6ZWx8EGAGZDRE6Qz4W7GiwXph/rjBjBjTuxmNWW7ZcR
UxgjeydoBeondtYa5UQCe6vbfvW5nOlmrHTQS7mQYP2ONph97/ws1O3L7lmYcsBwT3bCj0QeB5pO
2J/CQd/K8QvPGClVEzSi+e/TiD06qVieO28MMup1s37jkCTOeJOMznb/l6svuvtICm/xSeokFh+E
TTc7YrO7y07UH0rM58+nlsq+7Rti+vuihKMmd/13kjLk1mXn1DjvqQgkMg++NY9rJfMuzTvs+Ipw
LLqHaqgElFpCXEo/fF/lbivYjSGH917MjP66rJ4cD2xOEcy6XnBRakd9cPQF/6Pt3pj65HiMslCW
i0q7TaABhZrk4Pd2mjvpqtJhuF/Y6YVnG8eM/hcNlQnBp9xty83QAMggj3qXJzxBobiXAS2encoQ
wYqnJrhjJUH+Aesn5+oabqkTpHMUNF/AA3DB2qbPgiIa9ZReIpVIRLRlg85ln0zCiRchL7labGaF
jwIfrfYcdBLpELWce/pvjDehycPqrIoODhNO+BsG1QE9yj9dHovAtd6pqvcGJ1AlomVpl0aCbseC
HT59I7xrTdvJ5/SJb4i0/+vdzWDXP+cvpmHWAvtwhNPMuOpEFVQG0ctMDqgEFFn+a6WZGZQfliVj
yDRJklO4a/Xtm5YGgMJjd6xfN97BxRrhLmPIF66mbyjEQgZP6hmS59dlmbFfIMvID0cbl7TeL25+
GkXXCLzpTIc3eQE37AyT7eCXy6DNRixDRgoemppc05OrI7PwI3lf30co7ip8TGeYTQzR04b60nEC
QdE/DpbqOSAwfApBH9J8CVKZxDBNyhLmcTWsnjp8N3yOnmp+RivCP6cf6VYBUKJVSjmFfUvzZEFw
WY4kOD4PAGJSbRfwXmOh9pybIychay1cm51kBilPEwk2CkhjQgSuIMCwjgNA4MvnrSkJlJJ/3kuv
y8u33AbTnRNHlI6+/uIQlBm2FhxdCX5Z0mme6pu0ZQNqCyFJhIkgo0CJn+SIoVX4LAu2xbgfipv9
TEsFjteIlcTOPSPzMbB2zrzNNhwIVUMcBZkFwRVt2OSVUCrLfFSgrZfYHbBGd94Qslpz6PdCGoGh
uS5TxtroIijDFUnBFc//+AOQHJteH+NB9zcOfyziKvfPe2lHSUCJdGczJtCNaUI7nR7eR2Yf0kc+
o3VvzMxY8m06Ddt1kbsC3PHjwutUptox0nkFqwry+5I+1kRhvVSm/FG+LOi2q5joGlMEyHe/q3R+
NPGV1bSOueZcNugo0+R7RS8ycmMLo/sG0CNhKyai+Ss3V1o70g1yQHGrkD0np4druuIfZ7yEBEar
eYJY1viFSkzIP7claLmBSnWUmsCRwzpiNK/dbhI0OQGcyrTMevzIcxRz9gjcbamMSDQbgjq11K8N
E4sDbGN/GhOQgUhG2LK3Hw1z4jEetIPX+0si/jhpCZf0xcBugAxMsfhBS6IjjQBwQogUphl693Xz
kiPXplUc78OID6+NVd5cHaGxl8+pJlERChKYCuVerIrArE8a0dkWfiEywtfkFUD7d8O5dyFJE5z1
Edl66NZlJGpDgWO8HOpLWOmNTvpgL2ECszcGQCiYR+JGLHsbtFFI54IdruIzsmzP0w2sOamwez4u
rIo4Ss/ppY/idsK4aChx4ur542RxIp4oJwyIvlc/E0oOMLHIj7KX9Ubug9iMT+DsMr5rfDU48klV
f8iKfINx2BhYsg3gDfvFGycXM7HO2gq861vM/KHH+5QL5qWzobNsnTJuWAU8OzRVEshEyj9pSxNu
3YgNe/ASo816w2pTa6+npalryMVOKC47rQmuvIzbuAvz/rpWVDt0DAnhv+UAUP27Uu+FnaW5vq/P
VMwQqEKoTxlCkNellIAKSGHD1j5w5aTw1JgNx9LebWdrKuKRCX+yyMvbsJNHFHGrfr2HDyoTmPrz
Jbhc7X8hCy05eKZWlBfmS5Tmjydd0luXsQ42KdaA8vqPI1hV/j2Lav8SkquCKx9Sw/PbZF+0RH4m
jwK4kZG9kMykf3v/sUcFvivnB69h58j8SjStRHyFZ5Kq5p+IT2/mTFli+SgnMAGzfTNNhUhxH0BL
NCP7afptHUHkHr9RvkThxywX/OgbQh+A+BdlXqykqoIrTStL9DcWNoDJKT4Y71OVlUqCLiLq0gja
HQ/WfriLcOhxToz95Aahd3ir3kZwnzjmqWnHAyubpYOkIMumXSrCXS3O6Mtea0tBg1QpKYTtLQNE
cEUXOj9fcXeUKDoARGTEK7KNdSgiTvDtqymmRnwnyjDsh9PFG33to5EGVVbUdulgcRgJXBHRaSjN
3/J8rsVsTde0mUDfAckVQ/sjUOuI6Ad736xtqJK4WlUevrvaepTqsE0WRI2ELw676/UNo8nWobH1
Q9p7QAH6gf5zLwT3yTUq4G5liZhP/jsK8dmAgGDZVDFeFfeWDvIGS3tADXN0h8AxB/yrdeW6bTpO
mkCmZ3eCo7hisP4WnqOVeUkCzhr497doEU23olskOyMEtYgkcSfvyWlOo3UZmRACOzxeLPYWMFx2
nZM2AtF6gQzC06XHxLGryQnQ2HQzrnZlFiTkr2aOY5J0jbhQwG/Q9GUKw+o/YTwM6cpHKtXk7qSq
8nBwNyoqY92YgLoZFw5hfhABm/hBBh2FM9ZdxQK2inJDgBE90YtAR0PB8WXN026jgN6akHn5pUOt
74Xzhm0Q2zIPqx8naXhIMVZBU9HcJpuY2tE41tHkblwY/lGcD23wYTLDP5T7d+NvyOnjtlzsqkB4
mVxb4bh5ZRqU1aiIQYBYqTU7hk4pOUyoNTLoOB3KpIExLVRmMsCs6hcpzgtjKc4PW0VKuWCob1+d
FOb/muYEV+1jOimLKUdJhpq5ER3lePnLB8Ks5e8uuF0Z+5+PyvFE/HrAXAIJ56ZYe4I7CimpnDjY
0cT5FoeypsgLYZLKjyGIDVOf4g883cQldFEyldert1tWRE8GbvC9CN0Yh3SeAq2IfmkDQ4AxGSXi
K5QJ0BELlu8G4NdLOeWoWPXvldacLiq9iZKP3JHagelrCmK3mGt53o15KTXrurFtHgsyuKiteJX+
S3YD+2Xk0h1+g6VfE5LCYfdFDiM6ZJR8CNZe2ARWWY9gtf26+AqChaCdvgg0IBa/Rms/FsjYJwzX
pZlhbCQXYIlzC1se6+DCyloJxSL8SA9etzVn+861XIiA/GgKQOyTd0q0dVwJcjpwJx2+vzUQEHVr
pQHCxEOEgdPU0RQOgeRhZMTLXAccgjST/05VXWdj50aD7ICtE1uE1pkU/vO8hLKeU/p3IKVjzNtI
6DawSKnDNztiBE0m1IqDQ2uuX9Qc7ZLH2UUT0CcmbiVtQz12ajipgaWwRhO1Wh3gnqgsk/HoOMm/
ZC5srEQ7SUJ9ntcmqr33P51PHBiQTOIaV5Mre3th3DClxAJ8Cl72VJqUJI5J0A0YHQKAQK9amI25
ufg0H23en/ZERbmFCg4bC0DxRhfMgbQ0Vwg5U9D24s3Im/Z0XT+OdF+1ww9R1T3DCByNF7FxpZYc
ysBONDu5mzBn58xrrtwdqmjVOZK0hhVKqMXjdqhLad/JeWLEHzEF4bf4knWH+yOQmkL9aHTfYs2B
5Lq8rIIRjQkl//gMXNtPtvfarysX53UeO9eDmgnXVRQexG2JChng4F/CST1ujfmix8+9yM+AIv/Z
V6/V6OfLVgQsrWgw04sU58CIAkjF4EPxZCIOceztVbzj6c82Zqwlg9yeekSYIgxx4s3vH0KfDxet
49242gGwpz2h4+Va7+8ddRUhkb9vrPT79ul6HIqTuteWCjSQ1EyFx2ANF1t5HuNoGCkcSfxn7b3i
sHXYMlP6Ve/WlQAy3MvRP7dIsHlOgYce+Z9YnWWUg6lTtmYWenzQga/45+CAZGGiXi6j9OqDmaei
P3MkLLjks0GF71CDvynUqNtTmnuC3SajkPWBJhaki1VdCIwfC6/NABv5aOt6LTkHJYt6ibuC3GCD
x/V5oUtcg5YI2xpAV7mMNoaAfCzssPyeOakuxz9sP5oYPGy+3yzWeW9BsNBe5zCiOA0t1d3kGVAC
/UwfOZHtoG4bU0qUfOiKhlNts03bszeddIaF5JlR3xu382leS2GfBWhOtqG+UMdOaob7BS+reXWS
1IyDVCOcWntJTsV10AVSD4KgX7TcXVWKlBSlq9jFsnrgz6Hn7LjvMiZrDGdAeAB8EKfJHlzzWNzr
TZe+PK9ercvCec/Fw+iv441f5mq5/dmIkzFmuJutKnsraEcEN81YJSutKQKseKVJkjGoYpdfbGpb
PPNKXeVlkP2mWS+yEfxTQl2dNrHOtyHNHzyEpXTmVYt8fDJJatCnOW76g18G6ZWFDf2dfroqNCbZ
I2qV9kvohUkZPfygsd/3dZ+tBj1gNI0Frj4suKpWQJQ/sHiUc9kyghwhkBtAl0vaPsPILUntdeR9
bLxN0ip3acbKmY1Ltw1GSZxb9sbL/JchnkhnmDdwDwv7asesyxBxq0PCGeo5LmFl1PEApaQFfsB4
tDLEy19PqJ1n8fEKK9pccl9GprkRe2B11LtCLBrOWiW29T4ngEOMhQhtQ+Fg64JUh4RV39g8ouFP
zBvmpd0PEl1IrT9rR7THKbtUEc+T7azg4xvxwAkTPF2XpDGHhQZDYFB1HoELy87RMa3DSXsvN2fl
mYmdhXlr/ecoIM5A3Yaf9POJoLfuKbjkeQ05L4Y5bd4adx6UQuqzR9Dp+W5xmQgtdLzDQ+dKf/vS
E2AL4fAIjG67yW/o+q+BiXBjJ92FSukVwkIET3Gm9Phsb6N9pvkvb7zxZ2SBNnD52DbNYrGQ/Paj
uT8wbrMYLgP4IWflPjXSoReDpLUQAtx9zqWeJsUIWJSHUypemdx2IQ+vC5J/9PkSaXIomypMPf96
S5QEqgprhQXIAUJv5muSLXmEL8q4s40lu6OTNQOTkgRD9KApg2ikrlih1xSnCK4gewSd47EoMNYO
kKzNpZBU0fhOOOiFfXOYRkryk3ObzCYExjTpoDbG/T7lxnFFcklO8oN2i1EdILC1HtNDs1+KCJV7
6MfRJZpy8dPIJJsTEDTpuKv8K6JSW/XZGANKu8KoIkuaUS8kK5HlKuff6iihRtaTdUqlc8pCx3Cv
oIWzsXWfuDsWj2STgMNsulrRGBL8uFvt6N8yXKWYtlgjMenn6Ug8+8A1HR7wKLvuUCt9Ihz0pPzR
1neSbE4Z9K7oqrV/zsqyvFHuPutuZFM/mai25o78FikKZSF7h1HP7UXXgR5BveBVvra9CoauEj0n
KIuGr4ZHpXpwtrenRwJxcz/INQi6yabYlD/7knX4szbmS3c0fYzx+yIsKPh86ak2rZrKSYo4AxGN
XmfRgoXZfVbzerGtN+eFZEzLGb7k+HYEXwgDWOakDIGugfnYDGsYSNlbsju11w9FS1bCNWhRsvlB
W3rzJI+hLP7Mr7gIIdh8gAMB3t3GGSWpJiqfErg8WpZ5HrECWv/Q1P+yabqAgAutKOZNlF3Qu15u
sLThaR70hM9mj9GAD+MAYRtAsiScX9CfdQcDjcniVC5gD1YfIIpO2vvdqBRZnr11rz8PwcixC2dj
VTnuWFCQAfMyvqVe0dDscuhE6ouXqXUsR/1LMnbjQG0ZAoNlch90KuR2zQj+bzbmnJHKEmHU8TzF
8eLSGGBSWl9iRW4a2zyvM/sVcjOj7ge+wLaKEjfSLiBpX0ppCsIQCL27emFGpY3UPgXbZ4kM9aim
xvJdMipsVEBfhcHuQgtLfP99J6Iv0zTl1RD2stZbB9qfx1P11mo17wWL38aWKh2TqHJKjbJ1eD8c
7bN1zO2YzV2fhAg3CW8Ah0J/5MwSSExXms8V+Z46Trj6NfC1Zp929vBLxFOQCGv80Wx8oDH8qvAk
VVUsswut/cFMu/5YGGfBHSArRms0trHA9WntYnq+LXvn+OoDyQhNZluUZ4xrZRzTzqeEL1R4kfhQ
R4+qvk9yoQSNOlROv5aKOBiF/eIN5d5R0JD5g2Ia6t4l8k+6QbkkjUesZvvx4nL6bc7FSPXkDKRL
HG26hid+0wIHUvYGxfQpGyJjS1Tx4BYZH5Y0qglPPS/67VzKCdWFxqugL4AsAMPygYckwh6MW8JW
xyyGmxFXRNDJrpWo+wiDXy6qAmnKm9XteVBddzOitSMDNmmCVcidCHySJIE4iq/VOC8YMH3da2ZB
yhZRa1s5ycwsYijLb4+tWWqgmZdvQ0pNzqE6IRFk7mczNjnZQ0gFjGk/YhzT2GN25mQxPi8GwGnB
RYB7J78uFE4q6465mH3tvJZa4e+f36aV/LKfzHbQRKGK6bN8GN0+ptH3ZyYmXdcMGtnCOoRcGob5
RkX1z4eR/BKcZ/b0uJ35+zYHdmmYSsvsdjX0A/PD1Eb8QIC86Em34RiKAl6UZoN9yYCoxBKfnnlx
d6aGgfCaN3YzxaPL/gAftTKn/2geYg1ZkLn3L2FVtN4+OF9LPqgcDJlsTMxyl4QQ6O7uos4GhK9d
dTvRq8fAJAXa4m4ibZuetCiQbP9BSOk5JbHciPdNwc/LHF5ZFKJwztwKQl48wiLRePoNy3Z/Pgmh
l9mpkTiIsU7FdIdwGzKafsGuZv4csUADdMvXvFOToeeth7P0aZwtoxhSB+yH8JJ73oZUBVjtbJvw
Bv5jKvw9W4RU5g9dHNcVgjCqhoPg9Omy6okWJDVTXiD9Q8pCtlkmNDq/ouCoPZmBb7L0QejLI0I5
J+5AX0UKzrCOaJkYWryvliNNRTycnj1EkKfEcE01u9k1wYoLqYWec4bJnP5kbcD+npCmz2OTysRw
uVG9OyknGtnafJRAlCXyayhlJDXDpKC47vFg6VvFI2bWfrvS96wXXrBuVfrHLTtKC0dbGE4JHmSe
JPieZuMt4rInEIhGvBSXIMO+B8RTFdVPKDDoqmSBRlWP5RoGUum7vrAlKqnu12t6D5nGb32KerKQ
qzbuimykprthZ0IyGM4muqm2hndYJFqww9+r4PqgLpDhrcjjeNHVr8JGRzYcJXZNpFNqpvvmgl+E
o5aDy3rkhdbZv3ODPlif+H0Q/Zq5l8GOtGBcWSbLz6mgW2HBpBxLbUEOVnDq27YVvUOEfSTCnUan
Webg6jpY2xtijvyAvbLURvQJnIehfB2fGPgjmniNOsbB2pPjx4Q8ma3kZShNzIkE4BN4sHshiLmt
9zNRratiMtXQUrYX3dJgWnol8+SLtpdzhiGJo1mz55aDYAsk+/cuHk/eMpFEGf04v8xkrrRzYp71
y/xFdF8chehQFpQBDlm1Ic6cFR3oDszsrG4yREkRtMKi3+t3Qz8a9QPnE37plTYqogR+aq5Fd6mt
NkO1kkymowoIkX2w7Wm/izW4YnmXEfYjff8ofH3z5OX/tzSTA/biGeU0kRwNsdeS6tv8W8dQ3QOf
pidKgbtyofUEGZLCRcuuvtEWc5FrSUgfDsz9PHZ4gS6d59803MC6Oomxm/NZifVcwSE2Qx5VEPNF
OAmAkiWLRYM093iyhkXq0fvGHcwrcXB2vm2JZdMKG8kXVlJP9YUI3K32C+6XRJT+mZ2LC42eZiXW
17jcl338p8U+LT7ob+9gNFIKEYkpyKPvjZgLvp1axoCkdrLhxQ0rY/NSQZhzSavXnYwH9vkBmIeR
yihV6db7nuNusWutyzArNuyrwWa92ciWkNkeD/tM1J5m+/PcmNrIQsvYee+cFhFQvZiwRStdGGJg
J10zqBL4tztFbjY5sj5hJIfjz4VURM/tarjssNQgxvW3SXf8BvJTkS7MJpiCUqQ5JSHVO2dOEb2I
OEWH/sAfXkw7gG3w3MggJtP0YAnQPYruDje60k8lkXmop+uKAr5VJUkYPTcXl+BhnUqK9yAc7Cfz
LNC0olafKyY9Ms50AqEXp53Iqepqtu/n9mlP1htoBR5NtG2W2uYLqIJpVaYTvWwM+ep+qz6bK7sN
XXCn6yIez9GzWQ9giVbVCxCFCRoCivhjwxbhIoSVan+BcCsIeu4TrdiYUscuceTH6XinsAkFKTe4
vc4xh1KueqaMguHVGvkJnTp9XPUSrukSe4busGqv3dlZfrk+QZ2G5N23T667XiDzGMs+/JmhyOPZ
VIbQxomhVCpDnd+mjTUJbPqTJXFTRNWkxi5+Ua3u5dIl8SoIFkVyviSAnGMJtkN/0sZolJBfSUT3
OVP51UCRZ6fmmh9MhHBm2ML1uYPT3K3Xc/7AAFdGOfzJMWGvWJJLpmK/CdJKrLcnCIfeAG86hEUf
J15lNq8huzgnbMGYX6varof11bnPKsJea0H/6Wh36mw2UGRFN+OfGW5Q04IzpeUshtbMNBMFEoSe
nbNzl6XcsCgRQGv93EQKNVVnYyo9NGba4oMSmw2uKViNsSmm3D5q7yK8zsPInYwzFpJO7qeBQdpX
Tl1JSgI+z0AUUkDqqDuH2hoj4AmEWyOz5tlY4zZEeX7ZUtQ4Ay7BnW2s0kKKtGObM/3UxvgQl4MG
NjRy5UbYbtN/H/pSxA8pItOPqrMx2xJaKJjPfZAJUMVtttokB60oH7OdzztRIYOnAK77ncBfknPe
2lZkdCAZrGCy5F0XWEwee75LKZPdsFVQkwQsvJ3Lao9x37ZTgm8A1fSnpii4cVOnSA8ahfTdBS1X
DHWmxDrnr1Fu0t1tRkPba9Glj7/xo7j+OeWIM6Rm/N9+cuFWgT5tDzzhCBORKR1OMZ5eF7OevyBs
rw6r9S5XiX2XRgjqyLnmO11okDqNSr57SfUznJhMQbflaPcZd4eW0Do+iqNIFe330BI4CCEPZ1zK
J3MMstgiiuqWx3Wwn8AgOiDhgO6IiaBj+DJ1OvWqeytDY5T4ODlUGeVGYcGvM4Ynr0tShXu3/m4r
qfh2cAXMYcgGPo68O3b4MyWFKaAf9U9P46EXNTjOMoKihXznk4uv7yKIa8njNJC6U5eHbbsmPHQj
+TyelxSmet+B6722LgIyHAeqkfV6du4lLrrsaa4PZwIECntMkdmIwd2nmSA/qguhV4vwdFhcuXO0
0WHGIeJXk1DRSxRWHP6GXNTNZMnoiBQQ+OJRNd3IeoH1qZa4nRD4JN2FQtjGce3vfQcynd1F3dGh
oxb+KCU6tk4JBanKwZZiOgbas2OFMIo3HtDxlVEXsdDubp453Ep5nBSxbl6Kl7kg2Fwyedkl1NCR
GkGi7AzJzc9cPlDtE9jcVfuKy2wVpLYiBK2B8Q84F0DC9tnjemBW6juKVdoSlLDnAz5JxREXk6Q/
ygTChyyiQ12pqEZ/JzMThcw95ZC3B/r3w2jmJ2ZwnpqiL6GPslob2fDIK2051gPRDPoV3t8ThhkB
jbP/ThPsls2WaG9prOJkmK8Dfp0bR6SPXOtZWh4TCVLcEmrTd84Of7AvO7UKtebmu5+A0pd0ZB2U
qb0GvcJeQXIa/CbySgO/0pysXLFBFl+WIL3n1tyewYcEpNpLjUNxPBUuYghaKbi5OGrAEBizKXU5
jj3TQ/gTGou5igxObKlJbJT9/Fdd9e4ty578YYEt2uNFXBaTJT566uxc+HwYzL5ZvIGJ8vV+13CF
CdgsgacF0ODhtvZ9y52u92N6aEe0dqYGS8QEgeBPk0JBYHSCPth4sAIS+HtSY8YHUFNRcU1hkPY2
wEg6ChIdLqglmEZALELMr/b61I9bt/T3VbsFA6KSViQ1x5Ske1mA
`protect end_protected
