-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HFI96V8DStC2hBDzrveAh1rmbg8n0huWJh6mw+rJkLkmyNeeNdHQEuwZ8WON0vWFM999O12k/GQl
rh1S4qGArhqZNmJIqIdOGb1tr8+konxnEJgFd/G/2Ih4Su3rcgb+MplvNf9AC2t9XCV24vXy1q32
HdwLhqYaSiAs7KY9FywgkwJHuizkWq+c8nia6Rah8wYw51EQkFdQHj6Voscir4UuABhhfPKjIS8Q
UZi5x/+//pkdixTwTE9ETnwyi4LLlO+nMzqPS4yrYj16OV+Z5wWOKXHmJqg60pI1ccw3dhea64Gm
ytFfInj0IlTXxbZEJduySW02ulxwKQ0PJLe2OQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3616)
`protect data_block
LzniN9PMrjvwJxrojhYFto5akzBcCRBL3hMWuvPCDlgSQ/8d+aINkiVtflWIkNDWdsWuzR9WJYTU
f2zcF0XV8n2miRK4nBXvyOJDrMJpUKDy16p98pEpkw7leFfgidtN3J1aUttVsfTNiNW6JmADY7iu
Gp2+pANfh4Qc/4UCH6MakSHlPfRfjZvUPHRG4KKo7QEP5G7qnnQ06IWkYNbglt3i2yQHC6I3z/HN
sVeqIliANxOdUKPiOQYxm+gIIGz3eKTgee16PihLg5L4CTq2SR7fkVi6jkfY3+EBDBoNegZM47sG
IKrZrBeUc7jHwDSzeKFeGcCQCtGoggEBO2jfgTsbQoDTubgyOSrshHGNYrapVJ7MayIT9ZuNJnMK
Jhkuba0/Pq9HApjulYhSPnorluxWY/21x9Wj5UiTOHyuT5WaES99o3sXzFGBUp55KaH28yLQDDvf
WbwnCFrDJuDPz8SGCN3DYqJzFMO3BCVwKAsLft2yiyUou6oCBcRs/YS4XUIZRYd7K5IFDAEtj0Ks
BSRwPJgrsGo/cpGtKpfLr8zf+D+Zf0oQHo0rAjZ/ONO1WeAMSSRFvElw9wD5xyj3zzD5V70f+5r3
Qr53nh2r/3yxroOy162MtVn2nuj7UggPUqrAbZa9SZLGk6MEMmttkDrQGg6nAZJLpLBmTE+xjQTy
e4q9CJM+hku1q/uqgBcCQKIRnUhPF5S2GokYm8Ta6zL3B95mC6SHQ5jnfAMAAV7qRiDVq7ru/osK
DY+xMdJG0lq4yWjqNwYxaITNE1AQNxdi7cQYDIwJsmEkxfZA9bUOjTyB02CjCRrovf1bE3n9AmH1
cLue5mvJE3DoWF1twwHkIItGED+flZN/LE8T9BwOsufTHRsqhUrX4JBJNvJwEfGwXJQqBR0BF/hl
yzXfvdwE7bv/q7WuVb9o0JkOuPgzsSElJLswkJ6GJXSvr2PuYzIsYO24IHysn/9Wz9992fFnskXA
JN11HSjqhH5t9q3datyOKVFm+EHEEGz2SuzihLzq3ZdrnzK8eWTj7yRMJ9z8ucPqEtPZ86w5L9t8
HpSlMoV+7kPMpbRshAX4DzpxwOXNwQ2/vyxIdggoyr7k/V7E6iq7X3iyCr0gdpwII2pXtNmKDyRn
tYhc3tTDRCBqoRRufazDW1mkXqj3KNHQPRV6I5qQEyJQAgP+u0fvNouuWqR5wrwxZvY73gMzBlfg
KZgaZI2lNmp+XqlKWNZq8ylorLHu28DREVWB9eybnsN3dRPgG+4i/5U5B8Rr2gEpNkTp8GXN5XbD
nTqE/G/gbWTOY2ZiMDZ/k/OR+6LwtypWYWccB+1aUlebxEf5TG5PteTZyMe+AYTDFiQZkV57Ug0k
3SFxQG1+t2llbj36ccWv7YLPKQaoKZOr4qxo0KWtiGBOb8ramE2ZHTqZg2yNOXs97t4dEL4VjReI
JMjr7tJYunurePlH2ppxHLDEUfEUolcHXY/hEgWK/Z/+Fgt+CU4DUs6uwE3z4hn/llbK1Hx39uZ7
kErUK2oKqSDmPuAaVmR1Pjj4fLme+t9Y54YfXoRDPCkpSWytlyQc3htyBH3THSCwtJP/Bep95sPA
oRx0NSHAZCbvkF4HKJnLJ8Ln6qy3oz8/ea7wZGLh6Q7EXVpE0dvibDhu7BT4CDn8lVhQI2jLwJLa
DUS5jQD2FTvQ1Fbyw1606E2EsgJA7jSpUjVUxgng+9+igKJCBbUHHsQ3MzXIy19KfZgMcWJCUPeg
yOQpTeOnAW5KjsQrOSE6qO0pCFeSHkw5LGLZFI9jEIgc4nPDSKmoPvzttrWpeYjQnUN5jDZOWxpX
OnycLNeZCiu8+SkMWPuKdV1S/DgJFYHNYc4sum2xflr5pNh5FNNvFnmQPmb7bseCH5o0DHjZDCto
1WzkdRu+aRDgXcUZmH5iNUdf5w5WUe5i/RJnPopSiPWq0rKsMPYpmjbUyZxbh5Jf2EzB88iV/XMF
m9iV8OxuVbawgpx/k0I9j8i1fVHQjrXYNa9Q4i4Uau9irqdwj3vhHFFUPt41tPRbVEwMTZDzIT7f
Rm8dmI/cDxS4Cr2yzBBUwG6D72nE78BK5QrkNVa2an9PQBeFSJ5F0L0eLLLdl0iI4Eu9Kqk9wBlb
NQuQC73kXsdNxrJac+ApUmdj6ut4O/8/L9guXehgtpFPd81BPmaQ4b0FoMJZenBg9EN7N+CdB3jT
IImmxWx1BXkw3CIbLEcrfBwqjQ7vtCmztldfmC7LZsJimR4xeGs62AKgPEbilAUXuuDr/+qPnAya
OnyFjrrxsFOWV4lySAP9ZlP02l31MYKwypwuXvgeCliRT1Vh/de8rTCPhWx1HxtlpZof8wRSQTKx
OCfbO5xasa8ISq7o2NfetwUAR6n8B36Heuk0VNDrwNXEZRs/5sVWYPZlI8E5Au9QLRSHRN+62cbz
4AjEzqsI75BwjZB9hcC3l/aZg8oCgrFxeeF58SLWGmVqSKYAiVAEgoTrpa+mPFdKAz508P4S2zc1
zMle5UdzXQLjapo3MgACFBFumFKDJcK4uBQi/soNCsicGi3r7t13xZD4+ERh2oI5gXZuPSphsQmJ
uJL5LlwfZK9mOV5+OezfHJY9QnfnOZwSnxi7/+dLhWGpxKvPb7tJuJoA8wGzDbGYiOPxM3sdOeq5
LMbyxrOyGaeyGngyLB+zvTNUUSOIlb7AOWQyEdZj2dD/tpYyNENuzzY2hCuqykn9ZxeASi5YqQf7
kODnzgee06KVzk1nR/La7kIz48t1pZABZLZrU3/mDBjipTRO2fWH5yo6ZNDxzgy3pT5CM9iKSAWl
bNay9jqZkh/O2/1CTPYeU2BbR9uqoORy1NLE4TVEm2jjp7lM9RRHA/RZJOVqPas5GZiw7soyZJG0
30TU/g/Q6skIe13Day3eNdYA5zie9OUOzVlg6VadIXTw1b+66THsiiSLZssjFUtJCEDhaRJGDYxI
NBOUtwr/g9hEDRaHlb7OueKeLIM0z/VbjKLlFk5nJVgkhiycyAjzr2nu67cB/yjjQXgQG9ZKwIZS
+p7AaDeYUK0JgBshxsdjLMbqDT2m9U0M/E33OoP2qGdFm7oDm77JvmKIjcfIYiDNelZaJGags0qp
MrXTC7Ij4m1Ju2Fl/dIzWUGYm02ZsaNl3M/JMJKpePtWY+2mLJOjEUtqr1OEqROMKQqf+cQ0N+hJ
8JAZtwJDcFNJQGgLIa/E7PyZWpnMp1iER9v7E+ujqvFyXwjOdB5uD+LIVt5PmPAv8KkIBhXUxvzx
asaDSocf9EIunUjI70GDtHXhkoS6e80+Q4tH4fFogutdDzmfLZxBtk/2qyOz6HBxh+ifgDWqa5qV
Du/1yD/b5MUIxUxn30JKhS+Mj9yrPe9O0T4Hxu34nhwkVY9yF4V8pGNMkdKYBhgkpbcwGVv9+kvx
iVpPrPlNGPLhXQQJNW8uAIePvOLmhlAwd4wNCE+rXyrTiDtBCimYvHbgkdW5CajZrzfGGotXtrYo
i7qsIVBStHMQLIYhOs+eGeqaKdtcZJJ1uKgqOaML/Uf3B8+E9fmIGQg5O0PY25vOQT1myVO5JOvR
a2+nQDZneS73kT0CvdE4MVzgJiWhbM/IwXNyczFATqaQb2ufTDITMsvDk4Un5LS46u8ij8u+8GeQ
YC2tpoWFgDUh+gyPCeke8DIMj5BnqaYI8vQ5sP4lHAWGM+7GO7o6xnxx1aqQrLPg8uV3wVSzPuYW
9oED2oPK+iJdH2tuVuG/sVN5XOW/qDAN6PMmLztNrBh/lg69CfmP7ywV7idZFJ1bpkZoDQ8UOsFS
mWBsLN6kE/3yv7EGrfxLam17EH2ITA/ljCAbI8jOeY53dMkFC5pcek6ftDbqcZ6C2jnb61D1/Glo
Ey6TZA2oUe6D9seQ3U8ZJVQ3xSNH6j9oJmHyX5BAZHtGdWkkS0Ycxx1SoaoXYnZgF1zbuHUgEOuZ
Nq86ADLRbv1MmqIi5JRWyJM/YwQfkny6HoKHpWIPARJdTgkOYcskoL+jdjhm5JCkCXFfDEih2nSz
jSRcRd2Hi2ZChXwN7aSIP8MfZTbK/BeNs+PgUFo3TPw4Wbwzzst+8xykwxjio0fWk7YqZEzUitVV
qltSV6PTLYTyJHv6wzEyInM1Np4eH0B/25kLAmNEhkU7hTQm94/5MeCpOgFSL6Dz/EVVygzrUXk4
azQE32gBzYF0Jg7VIeLQ/8FSUSxYRVQbhqZsKIY0wmZbb36Kwqvvxry6NsH4lhu3a6Z2zMVV+/fs
erIaIAybfFDFgHNgcb2rqpRAdtf5BY28fJywISPoa2m5bH3xi7m8pi4HHDbYW8ify8QtOu8VNNI/
vDB2eRUQZ27Hv2ZJdefT09Ley5AzAEfJc47V5kd/3PelxpiU6iAFUSHFO+JeB5aUvn/+i54gYEUw
xiDUP2TzKjk+MooM1wiCivRFWjY12fLkI+Dr7RI2SLLtb6RL2PhJpvRaL0tZAGrDl5L8lAPhhf9L
elBKol6fptm0FuO+LSeKm+UaUDSuu7c6dlfVUlSpL5lKqekYWSHZ2UeZjRHNeFYLB1hHFFJJRIjg
N+bYf7BxoQYAHqTLcH7gdcQIFX6mf2QpkTO/EGeayhO4aKd3ZwS96PYPrIxo9YVLASGHKgG6QVEJ
VLMTw7GoGfmtOFa4YkU081SMxViOgqcYkx16u4fhSdcHtT+GQ4H1Gb5/RpSOg/0eGUFiHyv3aTln
z11gJB6sm4d+5z0+cJfzPYDyXJGNql5HPQQPep000di5Wa+Q519hivwgBU0UwO8HcXfT6/eVO7QZ
6w2bEL+4Vli00C0/DH2O+wl/pA3dTzynfA==
`protect end_protected
