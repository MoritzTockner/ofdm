-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
b0dX28j7/jI9OZFlMCbfstehUP/7UZI5QjxZI47xO0XlxqWripUmaeNDsb1y1ebn6GUmUJKYBfF7
2I6gd+aSIzhPKfDlZpRnBH88Wou77gCzcMWgl771FKYI+Ogd8Ro06kMcr1JQjxJKFVPYEeS2kyRn
bj4nHIbETXmPgxqOjOCUMvnlCFOa5NClD0Ox/RF+mZbVJIs6+mzkqOdMn+t2I0++ozPVjznrWST2
8FW1m27sTT8QVCLy0VrUVtQun694JYcgyX6V92R9ScUpaRR1NVfJhwt1ckXg6LQh7wYSUcN++17r
ky2/r7qg7a5M/eXHP4crG+eMTdZ8yCwriSsOhg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
rJG6bDpfxldtU54YzrlGU61qYyYyYAP8GxBKt4o+h0QBUJL/3PEbD+83LWKFYxdTCjI6YMUhwjCj
OhSJf6VbIslsiboWzpZakTtMEm7fK7u8pZCrxmoy+xued/QuvXZC2SB4kULIPc31Y+DJzbFdwuFD
vd2BG4r589gylWbPU2+qPuRYSLUjl9k3oTSxAEQFfg+tPRZNIUSCYhc4oHHw8C8r37tnB3uyiTFP
xjIOKFF2wD6hP8g7lL9QxFZFC5YgrpdNc/jOB5CjQ+BTa5nI6sk0nZQUPZZVF42DhzFx8ZLeaseu
CNv8WcWGNuDjnM+QaxqtodkD4Aqbhr+wve6xVwEl3w+677JotVhdsiSmIzM3h8PkQDom/QyN1k/j
0qSkRHv2BJ/NvtrDncNrfM542YUeDEzQ/IU2WC+hsOajlOxfpb0mTkwVfehJGNcFo6XS609fsebr
2RGsILDHlB46OqsQ2c6bfNs/gERdkbLp31QvGV2vBbu/KyayZBhPRB/Oha5LcqD2dO28cIJ03nkB
fn7XFrz+lrXzWleEPWOvfAVbry1nUEOS7KpKS2/qyzrvurzSPcDKvpJ9nOtUvfpHJ8GKlLsB3BYu
IoJZRog2F1LPusjB+KGQuoQ90uAtmxQtuF90zLKKM/CEq8uvVdvnXnUUAPkPtwfG5h+wK8xAoXmx
aMInO/Rg81fKHnkMosy2NXcFQrzl4y5Nw3/tQcUz7QIsPyOiitXOf0+kFY/r/bN/8Q52Xt0kPfia
5hMASM1zHjSldsntseMYLPvdlg2wdiWnA63f/nEy667tpKUfVE2MoiICzbdOpxpVLgUVi0bsCvGa
amPovxBGrnv3BR15KDU/XKOQuGuXPav1fOOVa1qvq5US+QegiKgZiyLVIc4FSI6ehzkm76XshaD8
qM9VlJlXCnq3bOBEYE3BEW7LamtvrreB5grHVRkEReC5ZxGvTDZUPBZsl1hJYFqq7ZBgeIG3YyAa
nAnp4GnAV9gsnoixbWGNDkrJ7uZXyU4Xiktw76bZ5CqTSm9YbyoYH35glgq0ku4vMnpfj+3tZoFW
ohAJU2Fd8pD7ZaRfJksu5Cff6k3pdW1z+ZEgP8TbtIwr29KuD2e7XxsRoDdx+uLWHuvxnl+MEPXV
uGPgSESLniB5O72GMbAYWWHem1ApDmWDV0k3zuUKGfuYKnS/y3cQEGNcTnLUfunqmrvOnnn0yyJn
SX2N4+I6BG6PbS60eV8lPXf5Cm3R7HTgHPnOk3OZ+T0fub5/EYCFTvyrrC4jsdzQmMth4pgNxZYw
saUtLl2LAgddbPJyxz/wbh6IeHQ7iada+EOHVLO3ed8LxouE/cxQUv2i6MSgep2fyEkyD3Rav3al
+FXtFxf/+snP52nk6hvGzFhKgw9SQD5QxKvyhixRX8wPR/UGWw5OQe22Tt99tO8nRA7JxlERUtMI
/YSFbjOumcSjsugnUBOMcXx+Myo642130/EpNeYyfCvVOTI++/66A4dXLJnSPxW0NAf8rkswm+BM
HQemlzhKWBXS5TaEOQ/wG1Ny3yLB5J49hiJGWuIi3Om1TfC3OGxckwgVfUuh1e+pIOMHkWrWUkSb
YHB0uAoJBHCcmWCM275uzuY8HOH8AOFM80sr2dJcDnylypQe6pwAT0PfCBsAW9gZ3O3Pjlr8q8o7
ZX/LXqev/u4jKdRVuyHW1BECL2zwxsZQ8Q5f/IrNWaPpmOqaEa4J15E6/wwYaVN8lGkyy5D4k80i
e6VPwYckcWB0hTOPK8ONgHVSgQj6TP2yhzYMVFUV/r2pcgRDJ6PrVD/wQ9Khrw6wZNeSxgddyq60
k1crjF8qqPScWQcL2A0qnuhzkT0ALKKwFJugW6StJ6z/uqWkv0mZhaQfiztA9LTFfXZr93ULlC2f
koPr6+FHnNgXnLpnrZNWK/i/zMX0A0dYiIgRAcwpfsWvx1qcgH2xiEStULUQNTdOce70nQWmlKoa
VMUMcJwbKVthueLdxcNlTBV4xQSOcMNoUjnCE//fMl1yudvFKStL8jpDrFVlUuUihIUtiz3iTTu7
rZHq3dP51nUQNvYOVIrAp561mS5Lnh2hzjXl9m3qT5C7bbXuDxkz1Q1E+pUH8gE7cmKTA007iQpf
NhcJ6jhyfaatguUZh0LVHmdfqM+7tZt+53ci1EnJlT+RGqLfRS8nmYsBvvpxs67/nuHCGE4EG0B4
l/Kb0URBWOSPRcqI/1AQ4S9bznN1dUk4dCODYLITUSbpGbmJo0JcG8ibS6t91YU3lD1ayWpz+F6i
/tK987XX98YHVuXE2EXvfwlL6wRPsvxqkUCYNF7mEtEQAyN6DzdLedvaqx/eLProL45hjD4baxK+
bev/b1EUXnYa2+cAdivN7MLfOLutGoChWrXpFEXW9XwqbBUey6q+9CHPUHaPnO6sQaHSOZJ+rMfm
BfRAv8neFTmw9D0WfieK52kASydJGu6/s2GCO3MqOgPg7o+M85TCJaMyZrT3P4Vb1wdHm0yyAxGt
xNN5GCLIIgVcyJVkHJZQ53G69gI1GKQcvnceMJPUvN5vLv9ZwXrQ2ZHKun/2jIEH+frPWMawphb3
OFgcB1sPvEUGdv/FfqNtQfT/kQ8YhIzkEvzLFNsrLzvHOF0itcwElkjnPZNf+WZaoGHQOJihnKFV
cxxwL21qFZCLAHQvamnJzg9EFLzFM0vY0b+PqGtx6VqEeCUz+6RoZkDf94dJV89KQ2+iRSL0bpjR
71Ts7fFcLZDPeAaLmZgMQYPbUUTFsiKeUwX1JYbsqYGx0sSq9spyGa5wYPHD1h7Q6MXLy0skazS7
cTNsbvmi+gy778gY48oD/RCURBwYtcfuLSwyLASab8QkaXH4BUWoKJ+q3+QY6/kede9zftVhoXg2
NhII1QwzDffqdywX8T7Apy+mmq75MoI0rCWCjQD9ZO+dwK67DlwGwnnbHmGA20sE8WTe7zB1OHQB
3Xmlp4yPq56ruvsyikE9qD6N23DEdS6+z4N4jYyTX1yLPgtycRqXNgpGZiSWweATbAs2qWvTtSgP
yW3RZuH9nPomhDb54iRbQtX+YRa46McZjar41xgyDTU4EU0P/TZ3r97Vovc+cT7d8eAn94iZEQf3
IDQ8r9/FontLd8aI3yVH2vQw70zXBVHcoi17jlDtUY3tw14Ji7WwnEzxul2VFMuzc5eLTYmAW/Gn
OM1pn46b6zhwwCOOEGUj62ThJxHG9xq2Nz26gJnj2yRyu2QTvioOB/m/Yxra6DxHQhcBHepSfEIT
nUfjGhyDHTjakukM8RebUZi0Tz9t3v6izKJ0RLuiSsKFz/P8WCh6C0O4a1caOKX0oVCC0HksBj/Z
/opsN9qh2tK7FGKBz3YFBsIBHiC5zionbA+iBIqq8qAxUvQIBjwOqaKIaUjxJ1uqbDRFWzJCn2cP
acD6kb4Rhb3MCiP2SXYYK2Bd8uaGVVa+Yd+zQn7HXE6K1Fx3wGJfputddl++qwY5mF9AJS14QWhs
d6bxvfJk9ebLP6hW53gECKJS3kUU+hLeRKDT4QFH5lxSCh9x11EfxRlfIqibYA5oMw1lfTJjJX5W
yulH+f4CFq8ljNQIxV1WitZtbXJF5YtgshokhTQSO9pPZxtdA3OpXjLm0CgUmEz/nnK1dEyH5m2u
2bacdCVvyBFqYDEALQcrZ3IjRYdR5+UIM1AHTKDYYnOWd2Df8aNbX0nb9pp+PdlmfnRPn7TpFxNp
AndJfOlhtVuq0g0EGyZN8xzUlFIjgu5Yndgdq8SghIyuhsu0BsRwiku/Hutzwkgk2Pd9EFXYpC6p
z5JFNMaRBmkU8IK45TjFPOQJWVuWBE0yM/R6mWFef55JGQjihPFKfeuCg9E2usFdW7rHOyvwXHAH
phIX79U9M8gATQvsaYtjxI56EHzel2RS2A9BPxMzC2dhUyeFXFAxxGPTBksqmTKk/FBGZjuMJLvM
9xpDyL4AMU3IZqlwIcNn9C9tCyrwHVNWOz/pEm/gxj8uWg2FikwCygIpXcEPalHc9ojSkjON/6Ih
DwOraa+vD8PZeRFHmaeAVfoO5P7kvGJEV5Z2p4eFAGbAaBD66yKICHJnHyFP5v7CHsvy2MAYOPLS
3X7gIFnFqfL80maSdA6VflaCL3b8y07u0JGo/UH/gNM7d6Chugf0OcW0t7c72q3DHUFtpxjoIgrl
HfsPjksheEJa7bj67AAeD4xgUJycfUrmAFpJNcF1DlCY64VdXYO5fgfzRlphuGY0Fi6N72F98n+s
KnXw7eggubGgnjmw/G7sgjQCynLwedQ7aZxMHwSExbTgTvL+QfsZPSFQT+KqYbSiU/ZrjWh5AoKL
gRxrdbrpzFBX6dMvspQ1Usf4Zq/tSt1uwLCrGt7UBmB9rpspzC/lrFE7Xmy++ZqvF6UG7dHcJHaY
gGq8j/nXstWIXta8+PcK6vDkIBa8H9jp+ZgpVoDy8rELTM2/5+qjVb15vrz2/AYEJ7auZadVFD3a
MMijUhtJIiAw9PFdP/21wPS9iSQeXeY++VpHvzZ+YptFuzPBxnFjyus1uJJ6+BOoBmk4qAx3F3u4
6N//79ctAWY0CbVLBdcbKh1RBFEpzOJLLaZpc9ClA/jXmKflgNGdxZT2gHKgdVU4U9qxZK9PL8eR
Yc8eFePyV7AbUtgmq2pP9AIwnkutA++8xjeqUmcmnMJYyzhrjNkS3nudMtLvLudtyU75GMWKQzAb
mnoZK1mG6b6AtMBiC7iQmT6gEaSjYzIzyvwhWeKDHRSqNanrBOQCCHUEQpKG5zrhRa3sHfFiaT7W
r8vDW+74xLNCEW5gXNNMpeyEUkg8ueDL5TAoCGWuE3HKHndqMMLLAMVgyj2f1O0sbhtOCf+Dq2Nm
AZLrMeg7nfltwcTx5uYEjaB03oVZDM3+SJH14UmijkthsWrFyy6fIRquBe+L595nqBkhpQ80edip
XjJMfj6Ne4TgO0lTGbJX/m+OBmgptGG0cxDW307D/gUUzBZHEb8cRl+l1tIGdoNz6XXf3VZFaVC/
f9APgiI3vV1w7Wz+F/nsNcwxvLsSyg5om6V/oP5gYLXPCtzJRpFFBEDiUQBEtQy9TxXCcw0Jo8US
gvocPpGxGZBiLYNZ5En7C9dgAQIapgLPTwz0EOkHcaVL69BdEfDuOt4w/XY0fNe96bEwhGxVX3g4
FkReCZqAtLvXt5Hxe2x8yu8tnh++1qoCP0e3laqpTvjq0/yLOcUzeYcx8lovAH0/YguWYoYLmT43
LezOxDMkyEDXsSx1cQQGDw/pEPMMnIb/k9KHYmss5kSVq28Pbjv+tvI5bLOep/W4lzU8/VyFAOtz
Z3iQMj9rKaWm6yuWNWwNRj4lHRSSxMY9caUjir/r3Lfn6t5nmUXbb2Dirky3QF1XukNLhJveYLzu
qmCONnGlFfv07U1LMmNPi0n5mwJL37lxWCLQ0ZuH0jOhLhAo3y6ETfa+teINEgGOeWzd08qIL+io
ZhWqoSpWTH6mmYxNSNym2bMkFwetO6IyaS6mKHxxkxru7OQY85yFXcA2ngumUBvwqxyVOBaHXeh/
1VYZK9Du+naJlWL5TY3W5UTPah5NDmAdn3FYcrdSyVptbWphzsftGiIedrjP73LTRwOgW28+ySUE
8AVb45wQ7mzCeZNiOfvchgatdEAfofHnQQcshXAi446M0RLRRlT+ywcIVoCNR7A7bdYash907mT/
EJlhv6o787nnLlpTF45Xb1CUHtMBVmH10+au0CZk2PgSrN458kctHdvHRqtz6xr3KH1j8lJseiKi
OHts1pphSFKaI2ucT/vbqRyT+6wxIzb1yXPKQ94K5KWonGww1WTIp9hvxn8ZV8n8UH8JaXWZAdri
NjWKFQcq0OLCta5Hnd5omcPMOXg/2rnmK31jxa2PgYSZgHKStAfHQVyMBgFgb3iJfK6PjGZ2gDrb
jDR7M8qqsaTK3cVdPEv7TftT1Q4doZcw2IIvKUCqURE0G857Hk9cYRLREGc4255c8kaT9dSQuwiU
WO68kLaTzx+Kvv5eXe/8GSBM4+sZg0IuYxYOMDrM0DyD7AJ8wcmnphDzZtT2Y1CfaQZbPd7f3+3R
rPgj2cvK8E0f3NLSc1VH8ZvzUdJx7ULHzM2gKVBFMtKUuJQ4BSuWlB01ejJUtlqCZ/nEEhyRsrj4
/isiEc8yaqtzV4DHOnO5UsUBLsLbROBWP04my6+jMnTH6D04Qqicv/jWfSlx/QwgBirf/UwKH/j6
gwivlmyTVhPxaYgpb6NOSSPOlmscx0uEAnu8DJYLhgJt1v0O57PDqeAhCEwEZorTXa9/UE/N6I37
W8Rpyg3D7fILAW0mQ3/QJrcZhSi3E9U6F/0VycVR9VgMAAX/L9tgkGdpbeH1az28sGuGrlP5y2kN
FQByPcr3yrMOh1TBH0c8rmihrgMv6UiH5SNThBmRlKJAkFVbqMyczJpT8kgT2DTp+gpJFilWAtxK
hCOQAGeuhvtdtpfsSqsTsV/COlUlxHYQ8CZtoEitbX6qT1IIo/9bvx4BPdw87iRFa4AGmG6hevnN
dLHW4bOzy7m9RBo1a8r5XKmNYBeq7RwzhH8pBUW4VrV3dTYYRVhpTwGGs8Hb7VlvJx2vPNMjbWqD
O9upSNQvG0utO5VE7xRQM9mk8nYko3QkNFJddbMFyPrOJN5yxMy3c3G5UszZz0iByVaL46Mbg1bI
ur4TH460mkGEvn8gv4JyaX++o2a/it7dcmmf8c+WjoYS0cLCQ0PHUMPURTbl4M6PrPYDotbGp/Ka
/ukRVN9Zg4BPRYYjFKa8vSqV9rAyAPDP+ex+L9IoBtDXdJyqPeQeCvyldPVcVMtkdofdWSMF8Voj
n2jV44AivgtB2+9kbYQ2Ro+nzYNf/hhuc6fUIYGMRZwI2QlhOx0DkoNBmYnRZn+0S9t5Q8F/Olcg
3ldm2sTcf6YsVXJWJDCXXpHj92CwOtdx3ILnKkK8anA3MrUsWqz3Xo+E5mo+2VM/Q6930CPiG+1v
bG6dOCJE3FtzZW5sESz5nyyqw64ybz2FZtGN9NH4GRAQ0ezH8tDvF/hBAKzd/4VkIzha8oHi+oEI
t34FGXgfaaBjLg2LvDsDKp0l25HWWJ9IT5jet1g1fOZEysWPmkfqHbX6n86z/sn8/lxnOzAJlUCR
BnUGI3Zx0B5sSbQy1H1U+mGtudCXfZGm6PnBRvpCPh1hpBVUDlpJbl2/e+lkxifmJ3NrgqMLbapR
zF+BYvZ7vq1GejZV+p90Ldd9s1C/S8pyk+Hv8NxoVEHh7yfURwrdSbZawVDUC5T7MFd3ec+2Y0Qz
rqzbzFlohpnwDHQ7MjQ80V2SSogg6q7f9Y9yOqfi8Dg7mQ8ftK7t1AIj9fmHohZuoqVyZY3B72zV
YebwEm224Bd7QZZTgDCs1KcIosFowqiUSvMLMYwVMy5pK55aYCE7SlWkp4alk4k0QbgwnbjH1Ovg
1YfgNeLijxpNAyRBx5Vby7bDHDhGIEjIV0WNwZ8aDVML16Ga/X3wW4AZ9EvRgoMPthzZTDqMYlgo
ECMvKQeBbDZ17U1/Wr0XwEYfUJbMsLaZNprbup7JAWpuO+q2fj3xurmx42gnEdBvBuLpy4H4S127
ZvNZGq0WoLODIMb3Zng89RxyXliaMKuSkEv+6+nfSQ8yUWTJSYRj2eknZCpVlt+zx5BEDDmWWgzq
LfXGX64q8+vceVpDhVDM1Luu6l7x6FjOvhq5xYuCzNadmP0zo1DvjbiIIaU9bPDHbWcpe9gwPp0I
PhUH+Cofqg8r/c8XZXNiDtEv5mqVEOckWB+CgrMQne2pv8sXrFd/vXa8W7V79sxj7kOIj6M14lh1
pVNOhXZk/9iGfu6Gr2eo9B91zzd4jdCAiV1nKX7HFN03j48lt6vdJqscepdhhOUf+ncjyl0t3meT
eH08ZkGmL7rrsG/w5gE31qZcFCp+iNINCxH45rd8khZIGvvP9NASE0EmDfBrhMwPyLJdFmjNIYV7
60Zf1KjywwjIl77WSe3T3hbp9RvtXslsSu4bdY71KbMzbn7ltDGI6rxuGVU9rvyciRIrROheh7ZZ
JglZoVodoYhmVFk7NexRWNK2IrIlRFerADAUxJob2pGT4lOyFEoV0EGL6+2MnTg5rQbcZefYrEEG
oQefEhkJV0cSPOL2pPf9POWGeyGtywKt8JHmco3n94d39MgfIITpK/2UXRN1EojNgnLtebWkQvpS
pJmM1UXNvKNmXkPDFwAepW0Pi/+v6R/TtbNVb2mi93cmMb+FbojvVRuDnn8HhCAQxS9FcAS+Meey
DfpGtXto0cl4jd0xh1bOj9mUO6GZeYGln5oM7FmGYhyTlvfoA35S/OlyUH+pZNb/nnOTMls/soLd
ySTMLmz7K0zmUATYsAgQ/UgYQFNMCigMlO2Zdmsv++XAiErd77ozciKtMlEQQ1fLkRBRaKBNh/Vv
jUxRZqd0NDprJSt5mPaBiSFqTk5OOQvd67UOTZiurumvfYQyaVtmvD6PBLDm6bliujJ8EgoHieea
f7kGDot/SckKpH8iXFTuW/3p4IKowcgZUFGptRHMTmXGZO3UI1pcMorlWzpu2jIjY9JGbPw7puBZ
IrlvSdEPyel+bOC6xNBgNXPgWf4j/RaiV/Cu2uQXSbiAqLNP8FRtUV5hWBGzsMXAN70Iz+lEr+Yv
yLYIQM57CAt5Cx3kW2JD/2gRax9hkFbFWMO1XhxLscACadBYHzisufkx0UMKfpASnskcBg8J0Zm/
lnDgGJoq+BUbQujei5ReEsg+gKBusIdd/JDZg9gaREIK/c86t2PDLOLHjYD32JQDbmMU0W06h79D
RFfJ7A1QdlMsC3DiviHrC59KArKGlZcRQOTgW4cNGgNTZS5K5E/pHvDX1+JT9pgFFSEru1zeRQPJ
WMHjx4wY3blR2leMBt6L8JNQ3yY9xPNd9c8EzFJ8mwa7pJgr+eRcH0XRBTJPifcsXF1NeJ6899tz
/qj5RETE1NAsIGEC7LzMej5Gn6nuMSWfVHWVDYKJumuBNLCqjVY884ZKUI3dOmXj6M/og3YXM2FN
d1xWd4KpFIvC0PJQAyZAayOXxIYxKTUn5HexuIu9mMUKyXU2PXnjatPuK2Z2Ut6Pt6vO+AWUQ+nQ
yqpM0/KJNiujq+JYoNWRqPC61DuUHaEQ75XrcWhhmggrY17b6xGgzu0SyNxVrTiYmQxp91QuCDLL
691MBWZKosI1iQsHmliyKtgq5IsL8ljH57iDChFUQ5Gb1dKGt9WEwGyEc23+xJyVKzGJgLItnEvX
HrPGotzUANupSKcRFatNfPS0P1aEmbPjIfLE3LGQPgB/uKX2sHsHMn/uuQm+Qfbv5IWiQH8+a8Pj
vigoIXCcqpua/e6F5GVnMgB8ZLS/sHrUxP8mJgKBZexMJiuGRbVjqs9js/KB9dfMdnToCpxEuhka
ZwNgXKlmFoXbHnN/iKN29760dT9FM4Wc+GQJKT/3rwavyD5OSkMm/TlI4h1meaerxdUZmHTq6y0I
kGkhUS6lBqlv5RlJS/f8NjODsBgDXd3SN+6O3Y8fI225sC8qnApV7ZPkcgpPT1fFMlf2sJPFrfCa
Kylr0+Y03DiUyaKmS88CIvm9jhllE6t//bStZe1dAEhN228IzXnliESGMjGiPAdsjc+bi7ZcD4uo
E11o+z0jeVpau88moO8E6VTfeZp6kR+er5zw5f2WQ+4tsD7P0JYYJ//2pKvrgwX8MvcFz+hATG9o
IFTqv5Xobz6ZstqVMLg5vN8W0XQgROnA3qG1MCMQCqX+SXc/jBi4TZRKkKvLf8QikskfHDKfyEf/
TmmwO7eeCR9Xb/YzL7d7CUjjYAxtVWgEFJLwNylA7tKqVKAlYJ7RUVpO+6EeNDBRJc6bVmmwRHp7
vpNQvNDvU3YQ86w2Ey1oqOocTdSImgTPRqt7dVUDfvwKBspREK9OgZhnRkSKLEalv26mXRWLdL0o
aVdlaT/hLyyAqM4g5QKM2qjKcSQc9Ezfeb50eLXJr20iqlHt0nAUqgq91vby8R0zUq959tPIblKj
frPrZ+w/l+sXiQ5gcUQe6MM1GXZpzycwJItR0uFGN8dY3HppSYNBUn945ogfn9ZWDVF1giuVMf+f
mdr/Ckn5LX7U661Ja3dL4HLkUIL0IVjg/KN2iQPcxerAwOgTTdlngZ+f5JmaNGsJa9X3bMJG8/BE
y11CIne1EQY+Y4f9C5eQloKlzKaBmRzo55daKbgTAYl+lI0clTsLQ1uBTVmZNkfK6dMA9XMzSDl/
XpL22r16r53cGciKvhDDwRGhM3yoOGMmzU+OgiGsNcqibEQBfceHh7xRg7S8iLVLChzY9Q9exIoF
g6ibkCrGv32hqIhWT3Y5D3zo0f23yeBgcMCco7Vchn9j9d5W9WH9nxaclYOb/bTU58X5hYeAE6A2
HXCrg58Arx2FJ16Q3lQaUBwomAaHl73UOjoemMK3RwfZfOd45qSoR1Uh/hMsoxAco0Q/x8QzKN5T
tLlYpUXsa8XGt8NZwtzWlbHGSYpoWfbXUuG81+0ALsxGNu8/zN2ql1f+5pNSbT5ySMA6YERRct5a
g3z+3bgamA/5lC+2JXfPFmKIxveEl87c4Ols54YaNJaG/F6dssxpox0OQTVad7lmQ6Af2M+DWFfF
pgXuWkCJukR3JujGQlFXLQ+bMTzDeMb/wCeaTU3VDkUEQ93pX/385g2jANw1IGCdpCqgJKJQIzc3
3dkPIEpstGnWsQLVTxssTzJ7NWnya8fR9ULoGwI45N7jAKn/KM9Rh8IbUAyY7kAbBXJRJe4zEgnf
efZ9LIERsT8dnr1oQrqsGWNANeX39MPfIKC+6eou3GRfqRJDPmbqU0MOclUsSQnrZZaG4bbyHH0Z
2lfGjXOtOqracisO4FJYuWVFky3uYrY4DFtISorjD9bCVTPhUSmwaIwoByG3YfJ+ERuwAYfzwWTQ
nLbrvKGQX3spGmjkG3ZhkuVDfcNY29cPEb+FsupkeY+hgUFxU8ngbe3CVIlFjzeq+vv1D+wZikVe
pCcgDE99kX27SpNgpmhjq761D6+lOr2AO6ei3jf953+kSsBTrtVVIUPqOa5Wtuo4uEeaPxi5wW+p
dyIYGlAk2mvQRtk7/nwIczMdaJiT+RQggZn4c1UqoxC7YcAUGfq9umNqLPt2XQe+Xo7nulN5SLmW
ftkq8EpJ/TV/xZEFUo0WwtNCBDyRFx2YZWA6zh1oAreNqyrd5Or2wNO5zvs3Cnobfn8kGLYc6cIS
/v978GHMTm156nn49FlfUNxNBumRYQ7YEBIovoN9hH7AUWjFLsfcxXVRitaNg6J8Xz1xIbRKU8Gp
HhofgwLemJ1xuFF2/0xyDG+o9vKQNb3wFqyJyng+mTfvwSIsCGo6HnFgdH+I4dQ+Vi1GKwvSASCk
5SNJ5H8IDkStKSRs6+kTaeYydrLJ8ZilFAwx5Ib6/VV3QBwboaHms1dMUFQJXu8eVhhPkoCjTfKD
otRWPJVAV0Y9RidBfSVt8qJw7Gpp1QINmruybY2EQBVatyL781hkDKT0Q9rTvUShjl1nBsDPSpR4
xUxBWcirLwux90ssN2w4bG7hiksoFkmV6IW1vQsQ/cCtPDEcGKzoL/vlRkfqYBIMjlozIh5sqEjQ
dJy7ZfpqzRuCu5kvxiR9KSXDqS6kBySdoWTFwaIYi4wM5Qa41q4qIbdMRF46XlqNTJBZRQtncewR
+6PyLtglcRPZyqXHfHKuVdfwdY8oN6AcEPRp2UAjRRPPLKiplMcmdXqQ0kdrvaODw/yrQJIIa2xM
ljvz4fdX+LAqX6RbbZsrEjGW3lRxfMfbZu16hA9JI3gAMgY7G3gB5PmY1jRu2OjBotG8mgM6htbZ
5sC2BPQvJgYYHwrgn0nKswxO5GatAF0pxDhofzH8SqslMut4b9r/zSAO0w0IEpS49yK+uCHqbGd6
PggJ/wQ5xUqbX9QBxi7z7/yNEnqsgSt6o/0Gd3UgYG2iMDuMntTYkL5iP7VuMT1VoOakRThGE7wo
LecJPKL66WTKRV8vI2ZWmiaES1kk0vLszqDPo7HTiRo5E9BbwcugFqKCGoHDQMoVoahKYh07vv/5
sQFqGG1h57Z5Mvk8miymhRq9fIldq3KeUXqZg6ov6uFklTtnlSrP6/0/m4iFfw3BsbeMOkdjP6CS
aDfAVf9UAEJEjgH1ZQbMREwowc7xZXDLGHrNDvg0jSkhWIzXQmsl4g4cjDklkwk07QG6Xn8DV9Zw
S2TWDx2pzW+aTnky/CtCbQ/7XNYoANOAEy2enoBkcrOSu5smNxxbSCtRdsed8MxeoozqyQNr3p4x
sivykL2znFXPnMibFiDXA/hunmles0RNQ9huNvtt4ZyvL1d4La6QzVE2npEbPX+5ZKV8rX2EGzLn
HM83JV7q6ulLquZ3S2M3QT5K9+1WZmFG3dMWkBhp4jRf1S0pM/ZUu0g+l1CtDxvaPgDvzfgogWfC
bw8BCJ3I/sXiWPGoe84I6TgotUTnrhubeAt6ZPBr/tlN0olfJDQQ0BgdVApGj9B/bDsoDGK8XaYX
uC/qAaMV7VWmP3tw3L5ut6ZrguZWMt2kmhgB9pEAX3fjkWJehp53gS1nJ8cCHsRihwwlBxPhN9A6
Zd0u8YfUtHUnggVhreo/wSFuJeUeUFGknsGCscQH4pskyHFGzzJkbok0FEudccdEHi6wAwcOFzbF
uMaHHKXsfiXA2CjH/6bS7rTq4leoyQv6E0iuM9/uMBmkT28liXg8FfsISTozIxxBDa/CmBg8z+7k
eT0rrk8Nq+zB6MXvyekuZmTN7vcYnApZc4lqP9iizd8nx8zAy8eT1dIpGTxJYfTHfkpiHuNEU4kz
lSWLe6xkT/0jvjljZh6/CuWnfMKkXPDXMSG8Ql/zUSWcbIeSCJYoT4rwPcCbjRh5HtJaT+jaW4KA
NT1e1mAL1CytKToZzjxFtSN+68HRMrSgIHGlTl1NPDp/YMM69PWsj3e2WlG1jtnuDSXWps5p7XWy
0n/0+7XvbIf6am+i1DjZej+AgpoTZ12YbwsppqNpqUwOBS+hIY3MUrNSN1uy4OfTt+XdvX48ZpHZ
Ic5iAfJm8ktbgM6enQXWA3P81Ro1pwWLalO/HohMUkISRLHWZBTxRU4/eisBhUGoml74yyN2DcN/
BrjVprKPqnbcepyQRDI2FjhrsAZF066g1pj3ggn4aNn7JCNOWU8tvo49HdJDxKCcFzkcdhQjlYVJ
g0Y+meAu+ZQdORnDxDNIrusexnuiFm1gcDg5A++3FLD49a0FA/ipTV4YTm+L5m93YhNZPQRkp0xD
KDOnkkq93IhHCxFAAEUifGEYjRtPx5LSIajltlMqaUMqRrdfQLpULspobQ+QmeGZpBwog407E0bp
9Xjn8SNWUzCdZGmDpmcF6QGRwQsIbIOC/j3Sgk7cbwBeMqpXoqu2gjHk4MP5DVbfiOqzTpMiN1ge
5dyyV6EHc42hfHxauwXjAvIXsYYmBsMXqkcgLtD71F0dEGDpX33RTiRGl2oguE2Ne/HENqf7bgwI
MhADM2tO0uo9ANPKWmFpp3WwCdAaJp4F4BsI1Wqs6in44vv47uaf9qi5/uFPWff94aqDVgSvs1wg
7a3xb/g3LnZugM9jOtqouL8aCinoNr5tfiu6TJguGxKkTHyCVyjJzosNriroGjUI6DLlUfwrOAeB
g9/pNpxyoKCI8a9PJ4w0Rzqzse7//72SUz3kx/+gTkL0SHoF0yKtpvYfzbnKmMQ+N9mGOR/N12jM
m2OX4i0hJvHWa2oElbVdxpxp2I69gVgOxMys31iebP9vQNm7Qk5ipxsejjBdOJvoAG6A9rs0q4W6
Mu+GNyZrplSUtFWnJNppIT7d5dzAB9O4U82rqGKNdtiekLZd4YU7BgjBwl3zmk4gXkQLQBlN1Ot3
3mmHffDKgN3cJmuD6Xo3lI8qByy5LB9puxARFqIdHf3L5eUmY+EYNTEPG1MWDGt+Isa3Zd8Oqc6s
j2q4Iah4geNq+lGU40zeKvJI+CeVb4skmS37UMsYnBkJlRds21uFHB4MJPVhuXmTbfDU+miRFYhY
RRKWviByZUzVU4Kx5diFSvTzCF/pWOlGLROc8E58YdsTynUpdwNxDvAQfJZCLzLwgqao5uJWdGn0
qeGI2gzpB5okVMKEYzYMBZ/DvDn0ygaxoZTyAQoCwoVPyREiS9W57k9+DCfRu54DFn81sdsS0zIx
Kj2k4K9lfJXFq8Ln3aXvaWNLbGYZCYbz0cDj7Re1q3D7eYJrMV/yK+i8PYSBtDABL0sbvmRKiXTU
I86EZwWx53YzZjz2CUTrRDnpJ/cRAYUtsraxKZjj3EEud6f41UqZmNZ8Y7z3+yUs8VPTuGiNmxxC
U5dwigG3L44PjL12xP08a+nnzkxEIZcBxoNcCSO9XAxz5LBrfX/7KYBhAEvfN1nMNu4+rI8tZeyS
wfqbhLlnCaPZ+vtAMZx4ctem8NfQZvmnNnKC41BW2KWNhM1FPCSFicVB8N3VZRELKVtHKiRT8X71
nSDcosz+uKjZLIXs7BasY9ix9+0JG0v5b8JjsGD3Mff3x/MOKVkzrrHWoxcPzZpP5iZkDg4t1Fj/
RyF/1tJHmU+DowXTpXraC6Dh7A6iHgDrZBROh4BlvGYWvj2to4vfycs7SlH259rulLKSlxzoC40T
6PvDI4ZhecM9hPy8OCgBuy79Fnhln21WlC2na4P6WHh0IdWhhWRQKUfPUpJ67sA2r+/O5aF3deqV
qVi9DozmzYwI7yWeYjhugALaIW7FwVMq+Z+D8i4PrqsJiHX4r5UhqDuQ7A/e40Tjfoi29+dcZ1iT
7fY7e7u5wvE0TU95l2JU06Gnkmi5Txq0lUr48jSXA477OsnSZccjwirmNY29kyJXou2eqln+qbV5
S0Tr81VGwFi0Flyj5GTY3jxNcrWHaMKSCPI8r7MngSNjr4fGSfuj0Pz4xFmGFYOM9x8nn+1+PhkT
zEvzuF2o2O210U+NmQLoTgKFeAetxLkPKyxFdzKbE64DKyukTWxm5DpJEDvNa/NBUswL9Ydg0Lnm
nqF22miE+EuYPxc0Kadis4DlBn71wjUN+Bl79dV+yo3dxWW7458Nu79QNtN7s+FilCgZAMKJ0ReL
GEnDbNiS9eOmGGFnj/ZN0QVmRoNtI8c65HdF/lvF9VmOoDJp4FltMnY6vidoYx34+MVEt/sQIVXA
kxi/qA9ZCt92zxYgtKzVZZvmmPvEtEbGHYA6f/PKcOa9sZr31NRGcB84fVmILAVtz6CuYmG7HPJw
21/sDc5GB+dfllCZ2X/7MzbXBjL7a7lBjfLkizdfMg/0XKlpCtHq3NgjgHgnbypHAE31CVxwv1JF
pxmCueoL4SKIO3hnsTjTPQ+7Y+1YE9LOXhQLNH0PmpSWFl294iCHSS1ObTltDGabW+7YKqa2wkKX
PJoHBCbfVCoxr1a05Xtr7GpgMKSZX1YhnSy6MvZbj2R63+jW48jjybgZ7irk++qwXbgBL5Kp3o8T
k6VqrBMiLDs3/mMgp57o0HU/Z145t/eEkofpplYPK7SqCq5UNvGx9KA8Xvj7kgd/1RhC5yQmyFK5
MR19IAS/iUkDXu7mGCymTQVXdRw8fcS8VrkGobgwrBPv5m0uAYISlvlmJ+S2FAJnNYfHR8Vpzb+/
/t/lwNysuQ9BeTCy4jC7OcH024NX5rJciXkOe7K0pVwvbt7clfRd7j+Yt2bZJS7Viu/ZdBCuQeAf
afu/8bymDqyIWzedAyC+ej6utaOkCAEPtvX2wN7WkHPrcQO3kzy1SRGXDaFcdoK3QJe5RoaN4f4z
5U+8eSwsuDWXCmWFrT/3MWg0DgR+1VUctkWp8iAxyFUPdSb7Ou6XNtsME0CabGXs++spv9WueXSu
OXZ2H/8qyvp5BkWgcas6OakXJqnNDiVnbu3vSNtX6xVQVuWJVgYJiGgnQQPhF0FyRA/48hZx2bXg
TXzgpkEfyOWO3CHqflt4OJGXCmCcVv01p7FXFvxwb8xhv1g0LZiev6vWl0QdBg5UkYrRzam9It0L
3z2Z0HbCQuhX0ZwdCKOlXyiuR138vcrXwodVARAf2GYW5F1C7jzA4gkSSfJFTCthaUU+OgQ/mX+M
UZATwlfWaFESLIlIfvAQfR0sGX8F5VLd0aQytrjJnkgipeOaBFoDOOUYLL1zxI5VW4NAbkpfgtix
vDDnN2ZZokyjI2oZXtaGtP/1JLO8EzI5p9LefI0tJWUUeEAE6+9MYbzr9V/yHmElxVf9mvzd8vH8
hD3IU5Pld1PBFH8qiNa9s65ngi45ZFH9VcohW4yz3FxqizKL6LUqZmFxjvING7tuY/S6jvwczhfe
nUWhjK3QWZtFvfQkiHsnczTF2cpwkl4HfTZwfWsxrajsEq2Y28+RyhmOXKutNrH1umpBzr9XLwb1
I0XfT18rUH3HCLP3DE+xm5j5QtgVV+x1PcTE6E4a2z6OCdhGyVNTMcjvMtdlrawIyAkGzU4gLqG2
8bmPGCyvG94r8A57bD/l0ylYyPeoX/sNt0GpHjfUbsU7Qz91OwTPUIGLF0CdUfu8nK/bKlsQ7eGd
oy0UvBVTDLdLAZnPwHnkqwLwpu7JV9lhQ0knpKAm1kEjphsf9AcEaK/tQMHp3U2Aaf/GQ57jic2E
AMU81js9+CT6of6BSQkp4nR5Drs/v+Jg1U+hz/xSPYXSizMG2e7VPqeZKF9CuLj7pIe/RJ76i8t3
H1a2sSihlRSRVy8FawBtYKmSdriTodTyO+MfxrI6qOETxUHc7pdtOgTbk5neqSaGJkxlShwPbhyj
cg3wXkByaGGw/jGzkhWALAkMMl8E6CP/wPSpB5eY6REHKBNfR0XmoQfqWKXNrXxtrjreG3qTGIi1
StswAHXOTM273DeW5tjBP0K0Scxjbydj9Lzw1DY5uHGZGxnkUNmnDCyKzvIGm8dZqc6X9bEQ6xMK
Fk6eH9iM7m4IxG4inokOe56pVpfG41nHdFCLrvYGM/rwKgtvYqTWxW7X8JQNrGh5Nt2edIKaVI/G
NV/GF5kshgBvFTuwm4N619SRfbbbUkkpgsC8/WwjvqfVrDsUDOY+c4RhfK1AdqUwqLb4uOEf6oTP
bmdzezk8faV+cmnMzDtFHFC0FFB0VAiT/qhBqjPSB7BHAgJSXDuqFSC5PJL7dxgDEE0V5+WOa06M
oeynWqk+XRb424aaXhkBoole4AxMrWDx17zC/FR8hSZREfKt8Gtdfm2Lgj2jNPfKfPFo1RCfAKhZ
7lY9jAHmDS2ML4cTQ0mHoT4/GkvYUguXnTGijBC/6ZU9HdMxnjgcqBjqDzDHtfUuzku/yNGXFdjP
mOZrXmBXA/Av8/9CvaQmtGb+pv/DY0ga07plRYPbjVf4s5z1AHQUgWeR1h/psrFKjSjNOAC0rc9m
uUKfDQbhorucDdP+HOg5lkbJKbLUIhvsRnXm2FJwACDqlgaGsauHIcLneW8MxZsZT/7Y+k9WYjEA
pttLiQSD00//DwoaxQq1cOvft5mR5QpDiVjYMY/luXahbKe6A6tnkR7Nnb7108O+Ehw5P23fNrj7
SwQqJTYjLyjxCMLuAQ4UfRb1vVcI25xgiIekRaKfpN2NDIWE/3r9LAAVw8I2MKuguJxmVo6f/Av9
jqhQWONailx5NqwWht5H/W3yiPV4vslPyqsUkifwyb7y37QrqTuSj3A/ADZI60S45218mt6Txb6W
sMkDo4lOMq/fmR9Qb85hxsSK526/i/VGqhtJBhKNwCtsiCzRJrBpSghyrvpEFKK8V/koyQnG8T4B
viOSnURwR2fDE6CthhWfGf/yd3hbjpR283+gpkdZxK7aC4joNbUm9cA8sSxMe18O8JIRmQfthEYI
JlOorJ1hO2aw1AJ2upQA1GNPpvoaKnvpHUbmx0wmmZd1AjB1r0rhgbq7kFJbDH/qELyu1RfiHkBz
4RFfvT9MvQ3pPFDRspNdlC+0IXwggiEgP4gF7zSB61IhjnMl27D7bZb0WRKEXMpTxXWeD7UB8SyV
06GSqNMCKF6w6yeXXSDbTZ5B6FOrBV/1htfLkehpFB5fp9LNC6MykycXqBs0IFaXEbB9seGsbD40
70Njjz7Bc/ImHi5oO8i3Z2N0syV/YMzQfbREYZX11FIX1UQT0TQkDI4tKmlTA8BCT+iPgAHTcToX
MqPUUMn0HoiswUMJU70p5E6WfaDqs9d+n/NuV6BcqgBIhApBbmG7ncWAZCbboTgjbCgNsJOljLPb
yXlaKtKJsO25LWLkFRf0lYth2Bs+yb2+aZTEna6yvBxGL2sy8r/2uoqaMZ15ZFcfufqKgWKCq8HU
7AOmwpRuCKkXCcVoSes8d11u4DlQQ6I5sC1JR9Fjd9DWVuAmBVJne6DcxVir+JAIjazZkhUIjr29
K4ThryHqi6fWVPfiPorTPKhdbOr1EsF1R9gd0Ckr4tRg85AikAz6ob3CKaPoU5KOu8kJK1vDaIIf
eQaa0SgmCIZddcgpstte/WrucYkzbsSg1SHuAhIqB12Fzne5tWAx9684TBaKrDZ+sgkVDVfum2re
Xp9OG1/+PHnAPUtGkOUZadqQK43gHU4nF1CKigSDEdM63LELN5SyZGKoFB+z1F7N6VI73N7+pjvC
PLByfKTQZTbjsXw13BreJeKx2GTW4xSVDAZ4dhxPvQzX9r4NAfm37rGHtkcJ93Hnsj+KwdbiSkBg
xwLGqT1Hus+0RUlC/oH5AHKyvEzew68ZFhmo4LN5zbWmrBEtnNwFXSu3gc8nBlsA8HYe02waEDPE
W0/fs4Xb4yvVhoufI+mO94Zf3kiCskKkAL5IjYKYaWaSvGdfWONlToPnkPJ3R8mthiFONILc5m93
rN9/0E3YsqtPdPj1rW50wHazsa5c5zdln2sMbe+TAh4MTA/4tvZhYB4Pci76bUJJa/u5/iJjmOtd
L54eseqYXNk8Nqq358kNXhY9s+hEpeKJbDUnuDJ6jS1zq+lqanDUVtQzwSBrXqswAjv5CX6bwcb9
QXN6MUzEJp5PaV3ChMPA28hIWhx8ASmGmPAODUL1bNzcn8e7w1qQbGAc62VcXtdt3EbY5DKCKxU5
oosbRWfjbvHTVsGLjiovkm6VGnkRBKXsHdcjbJbhSOdcBOBUqtXJm4iMrpkf4vtx6qOtp6uZMx+t
uvbivnchcW0IWDfU4ztSuhgnebFN8txk+PQ+evflhaNIBVGNuFrAehp18QPbDk6l9YpRrKapLt6A
Ud6P//uu/b+BopYWFRhanwno/rlLEcStg0FwmDOuTjuCkn6dt+wywKs6ZxE0sIRyY4i6gx7Tze+e
cFxHy+3/dTDUiuKgJqx0KIoKkGxjCRYQwteC+eJzfDy/p5offpLLVPgy5vjKbYG2afWqBxfL5b/1
f2JsOruul9IDmR5rTf6uKavkwezq+/QZ6qxpK3ljaDlmSD1syzf6yyOfphqtWTcaRaSsrgR6DQac
uUoV4GxzvYfcoP9a4xo1vELk5Wq5d7FowF5fW0Hy4IVHK9vwS5YHMjI3AiyLqM4Uu0wJ0BXk1Rci
0P+Jo2ksJdnG+m0kDqVEeRKx1XgkG0OI7+Kot+kTA7j+x0jItEkGyXFVr+f/LIUUX39td1pzDeSu
h0jAt0w3Ji4cU08ByD9TTDwyPjE/GFad+HjBvV1ZmsZDG3QhpwbyGBWNl1np6AGnFQvqq97v1cNX
x3zVpq3odSykSPLGaxENjvWVdEtsCXuVVaGkBBkIO23SXLXiM3OuJLfIJo54+krnclK78UsewtQi
3S8qK9hggNqJTT87yghSAzU1r9rVAzOfdF03omPUENf7585q6pwCMWQyNxSjYshMABGZc1vAjKIE
BYGQnk+cWxr7HYGwobvTRQi3afDkbvJzgl2JBthET/7gqAdPGXJO34FUNGi4YASyki8FidyCXco0
gW7JUN5+d3A1mpMQyI9l06lQ310/6gFoTQVBkTr1ok8q3h5BJinEe+8jjZaVU284K0f/VX/A2Wr2
9q8HNV1Qk8d7p22CAggdfS4N7kvo21sv+iHHUWYSq7hdrfvnqqb5KtIvYLOpsG9Pa0fKPm6fRWPq
2XrK8SnsqUJDp3I3eV6gYY8hqX8BuKTan7lX0lRPfNyZcZ2nar6Kg6EekaW1lAakNkGnO33hYIrb
3cg9vt2UFEwu3zkWRw3ygkUyArBh/E6f2s+xEYksMEp7hePTGBiJ7CunJhHPrvz2oYMN2554znqa
hFAp6n9AicNwi2sKtK2QLF/eqgNWJTmPW+RFwofXkvZlhHWPj2sc1xIDanIonD9WDuVnmfXkheiM
XGAQkftyBj4kJA072ou/4SyV6Lx1lrlsGGOmTHu19eXTFrdf27MK1eiXvj703TbAglY12/dJaMLi
t62grYcfa3uGo0DOTJL6PN6Ihsk2ob4z3I9q38JfvgF1YYn1p+u8E9IO01r8whmhOzUAnF+z6cgA
E6DkWOjIJleu8+qV3H4mUB4Oegl2xujbZTLcm+viQB9N8gtqP945X9CUBFcB3dWlYxiOL9zPqVdo
0orw7POmnyu5RqMtixWXrGvpG1XIZZKdXPzpc5q4gTT/BfCg8tvMo0Ld8L11VVzRqg2YNkSIbQkE
Q/w7A05AVontVUJjC3OUt3qLEOpORTLPPL5y2wZ5eWCZSsWPgUCuA9uxIR6KYJa/G8i9Mx8FhHbE
tEVT91P0UbqqMTeLDVxX0KD6kqs0370Ed1ojvtig9XNkMVtU9xt60ZIE5g6RN+mYCBeEXkqK6dbF
n1aZAhPZvAUCgPePCju/WNZv+72yQwvB9nQkF5W7UX28uocFI86qGoT9FKqO0HK1PiSVt6mOvCfg
mAEmwr+adZIDR6jV3HXb8lQjR0UHk9GFvGRCQV4MFv8KEKFzKvbfGSvegrzuQ4VXL448xoRQRrTW
NWjuJrbYyQPnT2KFh/seBl7ve2q5U/PsUB4PPWOEfXljQL2bT8trqAaHeTrDAij0qMLRl5WFnLkB
XGsLHKHH+Xx11iXOV/T3gLKG/oEoZNbvZsxXmWiRPRV5aN8xnwEPoqc4mR8fGtZwUMJ8WgMynWaD
JWzelT31vPpAwKFXsjZoGysj7QzGMSCY0oxqh8NDSdNQmP0iGHIZo8gLCRzS2bNRtK08KQiwDTAT
ZoXoRLEsNVnFCZZUn4adMfBFKO1FIqnEKHzmLqZzHr2jcSKP6Pd6vHZS9wDvXu8TDZ4vzvXibZKI
iob0yLoE4+WvxK7IbhHIHW2TXQo2BKpE6D/FQuZxmzIjg0QLMyB7NjbXvm5QVaEPq0qEopJqgJja
+5fzlxXYm7UXKTlqBLu9Dd/+pk4cRGxCvm1ROdIHuAfhb6ZsGliWaLBbT1IC0jMM2jCiG/wuj4hR
5iY9AlhV9juYGD7Z8sIxyHLoGJ8z2Fwry6N6uamiA1Invzg8UFpAZE0jW3haE8Q5qu5EAn2pcIW8
nyVRvVhyRUJVH+t8v1t2RGNMduFmYv5BT4kLeTYSdPrGAVHhDRXnc0S65dGJjzt8dQciK09CYQ/u
kZOqb6ewZ3mrDIp13pkzj+4CSwu2leNZIzpWEdySHSYtjJHPKeH0hVSviO2tGyJ5wpt5BspayonF
1Bz3gajY/T8gEKBWmjjwx+rifJXS1h6ubGI3nAQhWeW2hAdzFnke3aLVtZNh4gh7wxb1+3GSmi49
cqvSGhW3pVB3fNJQRmumzZSTds6332qKzsRo+voNHzi7tkyMchT5YilskUU3HjmYRAB7qPyrOv9s
agNE0a5LQ4BdRYlqU54QHOOarqqM98O8HhM7ErrsDXJu2H5p2kCgrLRUF7By7h0IyswfgkzmTvZe
1B0OhyGQQ1f+JmL01hTFp+5MqAD5gKBL88BX3V18STcGPT5F9vnHzqtAziG4CtuhF2GNn49DowQD
9QKHBERBn3mlmJiDTjxhmIFvfJ/4SfbBfTENDVMW5/lpyoNej+O+Ibh/qxnT8bJ5/3ZknA0WGEKw
VLQuVdYuHQc4OMjnQe2EdMSPnwCEUScBl2LJIyNSgcCzhOOUuLUMYx31sEC8jGwssuCww2CqaIyg
BhvR0seIvI7UmFLN25aVDBoPDH5ayG01UAXnHo1RmU4oM+KYLkILS0bQvGnB4WyMYlHJntra/g1e
XEi4WEf0zZXQ6Q5sqBZvpTwdfSoWE4uI1JPdDUR8ZC99uWtozst1qpcCAkltJv0M4Y747yF+6Sph
pn2sq9ZXIbO5IMWWHOEETiW0GJ1PPHhMj7hEjurwRLjz5AKjN6rivOFr0MGcmLf2qGoNBeT9GqqO
+COhquBDdLuPDQQ6FkbnNNZKzl2VrQzSWXv3o2mArVA9E+jc7cpuQiO7IJboNz7Aik33GkBuYPnb
eVc/g4ScH+LGenv2KzEcWmuQEgwx2TIDDW0VK4Ml5Q/pslCxPPCk39QCWGSErLETZIMbvPnofXAF
xH8oo0Om6rFZ4AznnlRiV4JvS6IS8ejCdUyRGNc1yjNGbJEhNX3LraK1RJvsJOB2n2Z7PJYPt6Qm
FWRLX7JzJHrSmKg9BWEgmpTH8qU3N1vGh1Yk8/h6XCzrBrMV0QYWdkMmM1ZTC8e1IVYFeeUlIwWz
N2pc5WKGDJ5fs1mr6IHNTfOUXIgUOkRHuI0zPM8EkxQR3tW/xAvFP5d+Qik6m+DZzyiMowBRvEzP
X3y19hDRqPy45raHvA+QMkujC0U8rboYyCVNY73/ptFyN+teKcKvQhScHhy47KS8jKaG/x6InOjp
MXB1ANvGzPqOdXXJxTxzAYcfG+467TYZL2nnbKm+27HhrABr8A16wPXalyyqoIS5zCXdh3iGkyrp
uK0CmfZmnKUQ3TYPC5cEPpM3C+hyBjwObnU6GoEkzH6Yc8TwdMcXsTwiacSelOCa/OH5dvwVJBu4
poxmW8kBd5M9d6Zley0z87eEhpr/rXTR/UoDh5q6FlalSJqx4OoKOzbIc9CgkviXWMKd/wefVKUg
eT2b7MJJqJoiiIUHWjqKZwCKrRg9zr81RJViXWr8m3rthsLNy7Xp9z0vzc8tewO9cyD5ILwct+ce
IZKVBcMuimNxwet8aeZCnOmsn+1nmNoaYS3ID8T0nY/K0HLTVqR+HmuDUYHHX9U0fcIqR4EdNiyz
2nnny0IjjHc5SixatPD4qxxkjwVI7M5+2zOGUChMbMCWp0bEXARC35yyEH2PVSl/WkNtaU1Ber1f
DOK4pMYp4CulPlyIw+ddJRL2lHjjfgUoWC32xzV1RkQj+MWf82J0lCsNFxhfPaquz2Cwf8XEjbQp
bXeCgJBZo1EhA0g7kNdMvDMbz629szQAW1tsbUn7ogtyPMICVsFmyeHloxQQSx8uCM5v0+8i20Eu
EsiH7uQ2JWqF6Lm1dne44GgfguCSeAPjZUke3yG7PLT/6PArlZl+PiLmSLkKZ0Q/x2iy8xO7Fr3J
pnPL3vW+c1eHd22xpJXOpabdDrjTi/ePW8UWs6iF++cg6D/0t48xgC+MwxsCB9zpYaw+n61C6lcO
mEdQQN/Br2+7xDJkb+c3gkOlPhDmXrejKZiqalVISoCKzzAPtXzqxNQBNtkQVUlvxVGKmsO4VM6U
PcPWBVLOD1a15cn3iwTSZWE9oyNNuE2kLODJs6lSAic+pnGJ/edp1rD31I6+NUZRcNolNSor/fPf
2LlPcHAZsGIHZGMneTq1le+GX19Laxr0Qzqfkb7mo9juUAqZ4qpzdSXhsEYTgbB/6PWUD7W9Qq76
+3W9Nx2ZDNypfItk0YxqzTkugaPy6Ar5ED2IUC0OrVl7uVKUNaS1zD1sjWPIKNowHo3O2WfqekmB
kDVpc251Iv0UzpcL+fQ+ngcM0uvOkIay/FvSs19balK0ElO6BTH+3xn9c8TvRJgr8erZycJ1RpXP
mECjEugqcHChWXFPSclCKko2Se76qdFpzsBZSOy0wXtjgsXCUcv7jEVniQxFRbdIXlacBpuxDVzq
gqiwNo8bAZd0D4uGfvQZ82VcpFEnirPyZXEO6BySUgszG+H+jb1iqi2kLMVoOWDyNitLVlba26uQ
PthlWzl8/yAHidDjGh+mDU8UvyXGfF9T6UCGoctq2Uu41qRlclV66EZILRxpzBHtsDX1xdboh+Si
ej7DfbJbYD/IYmY2GPccqw/MlDHx67OAVzk9dMhix7GOlnqKT2hUES/XOC1+ah2ienHntMorLPf3
DWEtjf8UG1/eg/NiLr9kwX+a4DZZC/tTggLEUis8VEMyUVBU8A6esOg2cFUGI/whya5A7k+w+vAQ
FOt8JM51Ou2n001rb00KozAfVaIyd5kIbi7F+GtcqI7EwpeAadBUak4y8qzAa5jSjbXVnQmg5ejB
fhfpGEHaLmgT+HmTit9ruNtSwNJK1RRuPYxRHaoqFnaUKOxwAdM6chiiC4xGSrDOwVbR8pKo0tHQ
L5SmAF/UcpLufERzhQrYWXx9u6YSJTJzZ2uaXg7nWHM+3JiC0VCebhjsF1XzhP7yKdQpfOQtsgWa
EW/PN+xfHpwJTF9QjrU49q5zT0BpId3fPr1DdFSSxEbCkBMHt3J11iaggdI98isUD4yRg11x7qQJ
2Szi3ABbP8t+Km2bGurnWD3jx4uUgXQ/431qs0WQmJzpVPSsuafAZAv0wgB+J17+aKxUDwubTL9/
wywBnbzkCzVoFIAOkJanrJIPqioxb6Y2tNWoENeflY/1sxmUxgl781EKQEPLGjHPdCw+Ynr+2KWi
mAMeXj64vCwu1E7IhhWHtuKwjysixALObDU7eaygNzh5ZL5m4EpCXberAIml12QxOQoVKA5hcnYA
7phl5nzYXBH4RGPuRvbeOlGf20TvJ0fit4z+6PD8o+ZqAv93WHhRkgdLANxCi8xJUbWqYENdZfLY
HAzQgb35YmMYcD2bive+5RH4FVxALM/0eevSFbnhnbcMwmJCNko+zNPx5ZWbNKz9Dt+rHtmlQnUE
bDN/3sCMSCwnUToT/0CQVNrojBb4idQknfYHYhVziho2ulDt2ZKl+XdlhBgL2NQhlqDomnBGSRc6
KYav9bkfUE64mMfTYOn8EQWEL3mH+QlC4Sj8Xet5YtdaMl4OMVe+6fAT7stLf6xvWbxFEpH7RRyP
MvoUVRP9q98JwGlPBOrfU2I8wZUlH8Igil7Ebjjh2TdjfFXQACYZNYHb3nI1hzNg3imtPKDM3Xr/
I8kl06zbEMxwD71A3IHqkrUzkEZ2GlPL9bDe4dD8tkxjv0JnwiGtoDcegeD6wa3pnL3ouqVTOxF5
udrxaJl8kUOT5XAH8AzVXTaLdA3gGVOOdkQITuNLG+I5u1Tk5dOeSwhCgOx8m5FovUNJA2Q7lXPO
/vnQZ2T17hdFmlYTaqp9nJCqFQMuQiMeF5nICDAa0wXEkO/4sUB6U6B//OHmiet4m++LxHgtwiXf
/Zh2qYOyCXbotIzYqGHsr1fMYc905gt0NLrKhxYKW6nvx7WtguS9ja2kKCBvxBTYZofGGYfkUKIH
G8WPyMRxgM9iUacolLtgMJ2aYfY9A0gjXtW/53X8xrmaIrMxglT48HTZPgfUpHOCfpqoRaVKw2se
B8VV6A5Rs1YIQWQ6y++iXAo7VIhbbipIjNWaPPlnM1VYCbTFS2Nn7xMNo5yKXtMaNsa7iJHdtAKL
tOvQr5L69Rbxh1ZiCyRunifhnnYvS6j7KEFF/HP5YPmlYImvevwfle06/iGfEMFbX8v3BWBp+opr
UWuKLBHLwy0YiPbVbjBsRaugOFUhanQrhFBIg46Xz2051ZwPfjMBRVD2dcXHrY4/oyqC5hQXqhfq
KUdPGTTzOPAtWH4IZR6KsK9FZodkE427s1KzFWNe6am9r/so8wNfBB3P97tchRy+M46m67b9eW3X
xa7aVsP3d2dY7ZIRS44kFON/eEnsms6et3Yetzr3W/MnXnEeCcNOaGw2WFWciWh69+uXT+otPhC4
YtURmS80WKpdS+OgVMDFsCWLlrnRCa1zNdIGR6ASXC1tRZPvsOsJ+BV7RwAQPdqKWrH5I1yHDDCW
4GGi8l3krG1jzZfw4I7Lb4oYK2IyylSKRDR4WMQX0BRocELgpNGbY/yAZxvAKIkibSwgMavl7Fpt
9zCOnB0sRrIu6k7+SpM53hQ4V8Hx9+NsqeCNKfjo1Pwqm4zUjDN89NyixtTCI7aNnCp+A+n1nHGu
e3XqmrNeRXm6GpClbpzxJ56Dcyp4H5SwVpnfoWL33KlyB5hH/WIs4VIGNqHMjfx0seLMm+D/l/8c
x6FdmybxKqyEe5qfFPYwbaGX4y1ODm7ZXo9Rch+3zSKV6YB+73HPXv9cciw0uhfunwZHLOrL0Xny
epyRfvpONyRQsKNFieSm7J/lvtw70g1I4VJ8p+JtZUG/ud9qQKL/4qtAGBTyGENse+w41wax/qh1
UH+gPANs3gVneEUYmPm+GDcbAP/5KQ/ja3rf+2XJcstbNu2jfKb4JYGKPM87U2PBZrr01f0tYsON
fn+nITIsntbaXKiShnaS6VLYhtBrovNiKPfCbwxfcSQlX20oYwN+1ehHOJVnTey8FHPbI6nh/f9G
K+p4wKRoGe+L/acBN4txZEudD7FxxHUBtCHlN8QrARK8GM1vzNNDyOzuWbgan6CtI+0QXnYapypY
A/WBWYQwcbqbpEdkciimGn2dTTqthUvPtGOwu+bSg/E0kNXKt1fPWTFaRh43PO2mP7HXfaorBvMA
X9gRnY5Ea/3Eb8uc9iXmrnhGX7DO7YyclwmPwUuesfnDSTRkzzgsL5Et/28kbj7cb8fG3mFESL0v
sEbqFz9HCt57l+8W6LxvtHxC/HwQNUvf5+lAJeEQ4DHB9d/wDcxeqPApEjgEcQ7QhVkMqX8GMBM/
LSpiGph5vf9RGWRw2We/UXqy3mbXUh80839i1OUZ0OpQ0K4evIKMErgqmw0iZdpHCiNGtxjaUZWx
wusZa3Tl+iWu57QXbuYiBBq+/VHUTvKO4alvA+MOYY0S/K5cWF4z0zeSEC/pbxwbsKUHrD6jK7Vq
+g4R6ZlN5Jr5mtwNnMovPdVu7mxQeoLRD+4yPx7Dzs/1HhT7RZKRYGoiCacmui69yKuRGS+S1Swn
LbcZcMs7gUfuaSRmlC0relQkksWaE8i+lsQb80o4xHKUhp+0e2W6h9EllssVWugkFwXh9RxIRJ9Q
iggsPz2z3LZUgEqvJ92V9Rg03MG6crJoA0dsklCwI2D5v9u6qC0iYX2Mk5nBhN5CQ89JOWQVgU+g
t83/qyEUBXCqlCq3PH0dyt8TUQ9Pm4ZvnYsdZsm3WZhGjj4eEAynra/+OREdPAGR6fEmAY5rGQWa
sWl8TySr3sAvx0vwu9vBCz7FwAAfUwWawNdVjKTRXGfI0H0N7xiO15+bHkTZ/drAIIyOGUpWmVYp
zYZ805jyvVhMeuD6HiWBcApjwuMr4M8cG2KnWo4P93788WQ6+KDKt/eA0XWZLE3APTtqNoHQglym
RMmUuK3zE/rfJ+ZyJbznwOPvjmywqgK4uzBgTKBuxyFGsqMJEyDFRm6GDdvTYKki+1RbKsC1WFC3
TR5vJ8sB+vDru5Cm98FCkcNIae3LFOevCdclyh/nKO+bpA+rvQt0Z1Nl9SkZn4aFgp0J0UM0q2rB
rOlmE4v17NHXQ4W0gv/E14ILTzg3z5BKiwuhE7C4D5lJf+6zzBJAmQJJeeQYgdjmykya2SiNkpxh
B1pVvxnTA7RkdxKhLaGjvyTK5/EbG6rl4EVW9YjXVPfFh4WkaQjiBet3X7MmbKzbqhtiXyLrT4Ch
KvxYbXaN/+u/RmwKuKrVIXMPey3fCVz28q1iP5dSNy0wI1BA7Fwqgs+vCnM+2RdG4JPSpKTri/DR
yc+NsAat4K6FYtPzb9qCkUZeS7/0Mdd+hsC5sIHQFDCoGKtrq1kgCNHGuA3LZ7OVqq/9rBnBScGc
LbUsdrKiMGvU0yIvfFU+FbUSrK8XXdCtQv8NwjTgOHusl3NNNFo2oPPsTjdxuPyIybjmm3imch4P
Bjbx6Lzmk5gfq6ouK+stYebyxLzvSyIj3ITZUX6BS0i2SVR4UouDUAnjOY1F+dkpsfwj9sVqzR0Z
ddpDj2m6ElUU7JfMef1uvly+mml5eS55eXCqaVYHfGhDD1t6hJrvISV8kUSoexaKD1AsSPV/M71w
vGv4B5G49EMIX/i12bNoce4ajBzj8WQPc/9TGwIfd7LXWKX6JxspzytNU1wJVl2l8joaOS5v+rQl
wkiCqFw1iDA/TwdvpQiGA2ilbeAWmcN6Q8WMIojA0NNn4o9ehBrj/1iLKDGRzwXE8xUcQPzOfRU9
YkiJiaM+iipgJc5vcvah9wnU2UteXp87oBfGPKDAilMg83YxRtX1grfLhxntaBmgG8QCECe1U35i
cw8PsBLVaqDB+TBzyHwdBQDG5KAhHsxLa7vSGD1coN8J8Rpylecl4t+pviZZ7BU9cnJMUE/7rsql
KpGtUY9lPSigEr4Y5+cTChZZ4I7oZyrnYvF1FiLRuPhV2jXt5ikFaqufojfOWwy0lgq3G4loCxO9
keOHIs+zBwgQKLC4faX26141fKpBQdUPDzWacSP+ExlI/Jy9Si0ut4eZjI/s9RQoZSLUSXKdP/Wn
1QuXX2KXthqJ6XIWjn+acbpvYFDCmUVGeURb+hIGiJ5Wwwb0DZaukhuE/XCbf3J6tQ8Av8Hi6A/e
3rek2V/oWcUbYf9ko+5pnTyz06kBkoGGv+zZU2veifWuzu+zyLjgC8INUQDF0iMFh0B0gSlA9zaR
8N0PKggZhbOn8NbFf4jhOhig/fiA/3AOK0lKsU8/0DTNVK8HPmjlUD1jwyPk/1xwIRhodH2PWHPc
78q5C+qIo10gI7A80/zOZVf229VTNDv7QM9oa7xXBLIxG5IHvcl//M2svhsJjcAXpuid+7qQZLbd
VVfp/wPHgBaF4T+rwxnTbFNHIJdpF6QXyY5Ly2NA0LK/C2ZisePdOTO0Gdfg9dj8oithiIdSAVgY
CsbUWKihZBY4NoJ1glb1GTG09e7/kxid5+pIlfElnnAiTJT5LKcwPgumt+EAUw37PhiFfVzgYRv3
9tOEESNmknxwfxEsrHyVkXHzih7HmNRvRR5H6KMfYeFBjtrBNxqlpThDU7HKAZAW6qg7TmZOTUUK
eotpxIuOqejpUB9wBp7p0HhIVur21Ei2tzo/22gOU53Tyt1Ig+nzcgT6BTdsoef6dwZvsV4+UkQU
nEDJCjEoOwk+HRpBrNorcjIrk4HB6d8RwUEETV9ecB0eARLI60IMyCWcGU+gsJ+EA959+k/ih5VU
hzAxqcDgpGN5fM1pzZBRNyEAuY6FirGNycUdSbHS2Tb5Allxw+zDxSXL6mJRAt8dPBHv0gnnUsBY
3FFjmOSTbSPMfOC22UwerX4Ov4PDQnAT2b02QGYuno4k/PTiMEV1Fx6kFjiS0lM+y9LCXnCTLTSD
fsMxad4SLoB41CW2Hq6j6uGf/qdXiXfGEeppUA0r2N6Rx36VNjgrzinYcD7w1E7x/bvUbar6B6LW
7c53QcuCbHFlvYl+jALwOUlsKQOftdJAMXmsHA7uzUqtxxXw7G0yib2hS1Kt1cJC82a7yP5r8fNg
TmGIt2F+wrPxPl9SetXmWGSy1xFNLFKhNVVOXo4Z3rODGtckw8LKpNsikJH5L/QwUM+1LaVh6QNC
ECti4FkvEHk6ZE4vWAC+LlUSjEE+sYya5JcKyN/lVYrR6/RQ0dzS1qFzxY44hMY64wHQf8Cb/ch0
A4tRZ6Wpajlg20ceSiE9Mxc7EY3Wc2ZhP801GpLcIcY0GmtsK9n0C2SXQ1dia1pQF9Xvn452tCrp
kjPjVZyXZ9hBGYkIMVjXJtCHK2oDp4zO2gMTv0k4ho1G/MoGG+5nn5SHWUOhEK0NLuPoGyIwOg4z
wZz5x8MknNrBrD7MP5DxFkNyuyu29MGJgQ9CITBhksGeteMjqvU9pV3JLjrZ3o56xQitaYt6l5+S
yt9P7g4DNqkf6dld5sVFL2t2tEmRS3oCRCSyyGBtyckoViNESWK+uI8GPNAJn/+KP2NIfF4g8n1E
YF8VI5X0eMn6fUTmN1HomG2ZWEbnDlcFiyZywnq2sNG1OaoEVgHxC2rMBjg51S8WSR/bG4ibtXKm
RL8QqxWLYChrh8V8D7AG7s1d4eLWNU6/w/hfkIOQXwOd2/62noo55asBS5nQsn/I7LFkRS5Ec9CG
37SXZKKe8ibyETvYnemNWruRfGOpF6BQZtCHw9j7CHaCKtxVC6UJj4mHZ0h3DwxQS4UxOzsJj/1a
rTR+gP4iVviNlhJcjPJ9cF4Z2qYABXtwWW10YhBmBo+9xlPiTf3z128RUWJH81LwLYuS3hI1Wc6W
E8CdSdnYS/ihCGp1/AjGgPRWaZVr4drEac/ZEnA97bdqrOFO8tQBKdeOcHtKPrH8uwEUT9DyK34E
mO3QMaFryYLADEwbCkOzsbQqUcyEO565pYOVN9OK3IUy1J6TD3sINMeetIJpRTr4VlHA2Lyd7oSh
ooqwObtMQsvCXiKoWv2zRGpHk2aSKowMxzLpxk2DTDYg4OLwX4O/TpPiqX5KKrwUaM8dkw/Y/JCE
iE+zkXhatWruuQjs8OGAbbJWIrw8xz6BE/N4JcFMdYuKQrQh1MMfWdjGxg4Q8X9M1R1G7L/d3srQ
Rm0klRjtKM+6WUfd5x219PAuoaYDinAlt97z1XrG08NGg6gUdHb9BAskqKopSHrFqxyhAiELls9h
kzEQpII8ljRkv12tKZnlgfsHFKNl045p30SasVUIX4Zw8+Kwk9Ircvoqycylcwu1QSMSW026dUrn
i9l04XsWkHGzC4SZFioS3NiBVRbbUGC+rpRds//8UlwScvC+e+Hi86WY4drMigMMIz6hlrMPo3ei
MDs4CAkPYbk8y3P6rufuAKt9wWqshrXOdta+aMg1pNMlifSFvP3pqkuUhkHLYiwpr8wHLlOTxsAz
t/6RjYA/GvsAKgyTAlF1GAApuBrz3lWdmH353o42495iVBpeOYFv0gjadUrA9jHBRXfp8wzOpHIl
EL3PVg54OtYmqD5zZxYD6M0JC5UEMnCfauqGx0JxNx+I+cQ8eBRTQC7fRMoc9puATwZ8C4xW8qgg
YzqUcJYZcbD2L327dhqi9fAE1l+MSD1gnPh/Iz5SC93ecBb7EvMdtA6YuVznlt6d2QAI2AVcfwzg
6gZejiebUip97Zf2f/G+g8fuqJXUBfmwxEvk8H3zaTDOmye2CtkERc1opanzeLE0KW+hJBv5me1T
jEhk6ASpNwXFOyMepL2eSWOsqZO8xEKGbHhpNWNWor89uQKPN0Elo8FFztmHYr2qavKs5hGk8NiZ
hjWeaNkEVITImic3kEcNWeBplDCoonHULv6YzjIdh0hVMQ9bj/SOICZbCKWASl2w6HKqPdI7tRdA
Ru9AK0pan/zu6G0UnVbxrOYn7qbxVSBwvDYcWrDgVaCqhBN+wHvfBIVYDaeP3uRzkH/vDondtS44
alMgg7uelvCERDre6AaeHLcLldHHPX4fQHSHNxJ2AAkpDCEqtEQ1V2GRCoy68yYaAW6Jw2UH8UjU
IlSHv/SEUeRFy+mNVFA0H7JP9ZC0KWM+tjQdSasz0DRMq8kjgekqAKaiexEQXRzEJ0PxHCbNzr4e
wRCq3Es/EFUmMMZFLTohMucxir+1n6/iGYHmbJGMgqq73qOmn7dNo1CKSPNDpyXNEckJdjRwbgn5
sUs6Y6yf9B3Kp0qwrnG1XJ044eJL35fYyssF5cgHlgjjArSldOSydZSoqhdUjY3rSgUpL5RCZrw/
uK6OhtcKDlfy0fkdznJPdHO+yMOtYh8x8eo6UeKFRRnldQtyqBqaNX84QVOa9uCiqNJFs6IqmlwZ
BjQEU8egjWfNQTsp730HiMj6J2SozOcPVG+vBM/sEwZ0R0SnL+P6rsLTr7rfXUqfdf2pB+8vtrC5
ixThHLGfUqPjjQ+j4E5zdUjJPkhl+pgAY69G945t02RO70IF7ODDB3z9UzaBhIM7uPfEgc5+BK9x
LnjWylQdqkXbW+xakqNDCEQqd1aFNZBhWZtYqUs1olQoKoUl+xAMegRQ7GyXbsZpdHIb3HuwPiJ7
I/u9sfoa7RPwoI9DHLy5A0WAh5XurBdupLDTba+KMmclKOgjjHGhX+N5zyoOXDEnxv5SZJT7N+ew
wvh3S1HMJLuFZiii/UKa7CoQsJMQDCT10J56mUkC6PwhivLmSUz6RSlNFUFS4dWP2JtCmRaazqIg
dpCRnGWlVGJIHW6rInHYG1xoucykyUDBI2dAoTTGj9h50w8xO9v2toU6yXirvFfrDMsIqqfmvnTr
piFRU5jcVBcpRWKNpNVKsCxBU/dEzfUazICsnclqndBxWy+JF/F0NEF1PwTkTyfjbjYeRr9tfvvN
vE/sxcvdYywgnyFPe5fV8f4y/rYr0XcLiNb3ykBHa7U/qwsBNLyxDYhVkbMOy9soJssXYXWtsaip
3uC2fevUgbdxc3v5YBP52mJJUHuvxCMjNPJBmRvZgZerB9oHSSqU5Yc8UPOqyd+CwJO5WpA9wEvb
7KsBaXAqk6aWwY2uZjQGnJy8wTP26c1U1vn3OKrQq9nf+LUcusT/htKGPiaLHkSMGvYUSY1g+jd4
CWjcgysars8GJ/S55NjAgVgI1LIBRSilSEiKjx83x5SD9JWh/uWlzarTMDfd8vAEeH3HRvVMbb0L
/lYM+IroPB4PgYhygF2+xLFw41MuDfZg4E8f4HLcrBi9s1bQ+VsA4Y7gLg3CGWs4GKeUfu7iTYho
rElj7P/IX30cLmSXjiFLo72k7t+adpLL/K7Gt+Gk6avGSBOBdCb6VpbtaL3hEzKT6tNWQOVUypbm
Vlm4/hnEW/B0mZvxJGN+Oep+JOfs8ZUG+0Azxg7IIqRHz4XB0abronZ0kpNTXBA1455Gg2+hgmFF
aDYpIJGWqgqeM2trNkPqpDst6lR/d/hgqOXDZsywHW90nScu2fMOoHklAHvfsJ4XrdrWRw5BGaro
tSctnlcV5JXQKIUuIZNV+zjWcl1NTgWgPkh6qbaSorRqXjV7Tl7ak8zl7XVztQz3u9/irPpZ15UG
emmooZZzlU8zfeXvhJESnIjyyxby1Xn67buPdf4Lf9u2DKMRh4LCyD/9F8mgyVrH1427GaHiNtX7
JiQrJiCCJDTFI6CE9E85A/8dMGwlkSydjaEuH41OW1THLvBs29rn3XcYvA8L/9pQlE3YRbeFvIsK
LqUEVLTyyc8ExnIDXuRta36d0tvuLDAY1yVStHye/w0t5pwsNiD1GHbnzMfdehVBkWfdfDeXtuzE
pZ5skucdeDPrtZEIz51NMSD+FZnzETofVesEk7nCE7JCWQztES+S612jOLZ+ppWZgCX2pR3/XB0U
n7aPrhTZiP3Kll3ltvKU++J1w5q1H1GynIHHCxuZhk86/NQ3huv4V189AL/BwV+6av7nGnM5i0jn
NZasZAMC8iSE42nTgkdeU0ecGH9rBtcPKMeKhZGCILvfHTdr7fKbV40ibC+PAsVpJuUVxA32PN2p
GE9ZQ4hkuyOeX/O4CDUruIwFaJDxvWp5ev/v4j3m8rWnIJPicv758bh7aEKGj5fN1eNmeVzx9/qG
GcQPqKfM6ceKNxjI9Q5Min86nCOYj0N1Riij1fUpGlHqHp6hFr1t9jT/P3MjC8JDz+JgUrJyWWCE
721vM7JOSKHBETEg7xQvu5TekVfQ6OBLLH8xSgLEO870cJqE8Su9gy551hIxRo1nyC16PVF+os0C
yZTMJLuG0duyCaH9g5Hgju3ub7/QVm7kp5jfl4PMe7oAuvf0Wp1s8FMMWswbFWVXItZdhR3a3w+g
wkaJEyAmxI350/1Ag/vr7Vz1wC8erPfxJhuv56eja/+BB1v6Kge2KqlGv+1CdLtNMgJhMTU58zzJ
DRPglKtmYn/C+FUjwbAzJAIaLUHuK5GcGb5kyGpNBD96xGaWpbZRnS/EtibVgdDqfdiwWF2Pq3r+
1Lg2jfR1388HeqJpYO10FzllEPLPXLwDKZgm/FLw/6DgZBX7E66IJZcxvZ1Bdd7VGCQfpdNAn44l
MkdXjTnbfmh+iqFMXn/rVG1T+xC4IdAQbDw2QSNFIQItMqokWcphnMOS7r3lrGISSkr38JU76i9Y
6y8ojfa2aaUqZVjYxxCE99GU9hbjL2EtP6ecA2aW5OtdOA+L9DLZtRFYAz9AKwoxWJvP9Itwwnb/
wi3kyV3caBYnEe8PK64l20TohxVz/n4TO/HXv0ykQP8jywEep+/l+bfqcQqlbUtd+FnQYXilXg+x
YqmcoZLXr+SuBNUIkwJSrqTrV3jJ1z2COla3yZXgixyYl+msIynqCIZnnk6J85Y6jxcQI2aKEIry
8Ntf3Wip9Lv8rK0Ngtbqibl87H9CCZf8sLhVjsoHTkTdtwFknJ1/6uDf1lsmbsI50HYOCy2nSDCx
tlhoceNr10O7V5Ip7JSvcdJpwDVDnybGjlhSyGxIp8ZcuLKP5oWxLHE4ffEaVPcf0dELOV3EEIGX
7EufKwlKaCT7WKWanDH2HJ9eMwmZLvwtQCUHU6FefJ3qW2aY6lOjO6QXpi/8zs132lz1ruV43/Rv
RicHHUPzLODN0Etxa3nJwIj8a0tT2NNdLLj3LjKKCdRX9Ocq+FnZdhFdfqV8qnGZZHDYMJj0KjXK
e8wMXfU2hd+ip+s32SBNB11fl70zk3yR+g2B9Ny+9XCsKQMncNH7jKBsDRkZLmgJFA00WxEOJGrV
hd9es6h6vxw6tv7JBXn8V85B9TiQYf0uuU1Ew99xgd4ntYXx+5/zjYfZAEUFQfeRoBicnWA+8JpY
HquxaEuiOZXgs9fvZSu81mFB2yWtwl69RsPDJRBPDL4UBpYE26ZgE0KUcWMRgjOSIfQhCHNSxYOe
HMyq5bO3tpGY3Z9D0EdVBAoVJ+WqxKakv7Gn+fMW4Cfdh56mFF/I3oIP6fnjBYGGIR8ou/+5c+MF
Lp1G66ILhs8UhxjKSXQKWh5OfXjeR9XDpSDPfsKKTOBstKH8ZfbSFDWMYdkD43o3/zDosLg6r1sw
J9timRIjWHFV7ufVPJTZhlIqrcVGu2Zxac6wZ2e4zsU/Zn9xA85xESAsalqz0GqYrGsMITJUgMJ6
rs2KTOHOAhCOpXYixwnNUTeNMXtVYbF0DD15ud6KoSpLqmFyJ3AnCGHXDFdq+/mNqyw3ldH7P4eo
X/N38NZP/6BCd1D5fIsCFGZl7q5SjsJkYgisIG+oFl3FRq4OxNStNjEECLQ23aifBJAcSIxUnAUk
RtjwJ8xx8AWpNj099CR/ngjQ+YOVsk+4hxq8/r4WfX0h/HzDFVkBdbA0H5w/4NU2FTwwZ+dHaPG+
EhwoP1muFiJPi2G1bJZk1SP/p8/dAb8H/C4mpsWnhFe65b0Fw2zGbG4zJjABDoiWgdg8KIds8TX4
PDIYvmp3Ba71k9MGUe1FBgcMEVt9j+eBgRJIldi7PSsw50adHIcGNBnHYjN09mRPEozH8T3g9w6V
Gh6beDFuD+qEY0R/vHlxiUz1ryg2J4KNR90wNxLNWhOBLLQu77EVRe7KlpXmEKdTdRgsEpTwdc70
DoPoX950wjuto/0s+mYxkC+WhBmsMMXNraxFzuJG+W0JlfV3Y43Z9B0K9Vjc6uEXBe4MTewK8mXf
ATSh8oxgYsnqta5edgHoDmYTEVpufiwi5ZGjyhX5n/Kv1jyZkSneWXguLdd2zU3Zad5a9AN3RiDH
hOXykhujdCJu/y74qQLKD01BoNkZMtoTIl0eQvkqmzZGXcqpsrkpujqF1csrpjhXcume1Jq+KjCM
ZEGildM4BLVgAazuke3eZXfckEz75yyyUbiNKXLWwb0n
`protect end_protected
