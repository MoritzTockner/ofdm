-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
s2Q0ygP61DChSARgYlGYETW1Qspfx1LLWjhY9h448iXHl0voRM2CdED2Tb+8UIEuv3DImNHZcbGm
grFRpzYKV7/FuHl4BlkFW35TSpEoySVTR9HZM7wiHeYbHEJIj0/XJfBCwM56ymcSlD7Wp3L9SOjb
s0Jtmk5+09BStMWt0A8p9DUp45pY0p6yvd6HMRc1Dkuj1PfZ7dojfGL6TUR/jZkxDQectOCgqnC+
dc3b26ZgdCyK8Kp/J3Ey9/P+vJXxJ35nS6HEWpEXQOd5ZMA4GnBP9sXiuadtjv6O3O4hSA16QvAU
pJ1Y54oTTTBw+jPmTFVjQ57zDCstum0folNVdQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
q5GrO8ff8tcslFTYrBV7yec/vTacsljD6YpTCCfHu9mutcHaSE+ByJftELG1+VniKcT3yPRfbVtk
tNpdMoQU/CAN/CJSu1U+kN3ON3r9QhQC8MG7l3/aasO9hHUdjv09PWZYEVU6V2RW2Cak3STjGr7U
Fk+SNCAbqvuFDZMDoBP0I3mqPvvpY5k6FEoDWpZFodl5snkSW77LBBTfFnHawG6H81/nZv8uAUN3
PijL2sHZ8/BKfCqsSpINA0Wi8+q9WowLF8sooH+Yz4DYjZtMCaZGSP9Hjnfo91a7IOPjER6NIe22
agUPjnFuTuCL6JGx3gdtO9uvkPXIAl/4RaFWaucfLSbHLPDCa8xqqIbACO4C+SAj7RV4zRmihZTg
j35uLCBBkhC7uqi6+13iWlZ1Wj0vWg8u7/UfSQF2FJlgRYqM1tO2/msmuMBvVbTGL8wS751mk3cw
miDE/NVFaKEBt+cpOug6tKVjradqcgVJp7QGb8WOGCVCRPxfruNo7A3rXjUwqJCP7s3fN0avwd7v
MWQhnvb1uTfvJsmfJ+JKIRiR2MbwK5wGJJpBdCtsq+jZ0Mu594GZQrBtNZJ06n2iEEkvIDabkyR8
J1aafk2qrNnOIVE+2hhMRx9REZJjBIXJeXZ6fvGpgYYjy3sTy4olg7EGiBN0SeE8L6A09L5RasW+
5FA9W0/ybZaDcLInYxAQhl1E6aYzmCtdn+4XhTvIZmtbZuiBI3Wg9AiFOON/mhhYUAMuHlOgsBsg
J77MUMf6s/vbwhPw7DdmtxPAbQl3GzFvm9UgNSG8hy7bRXUNB6lq4sUHPmduZ28II6qZtZk2kIk6
GUtSSs9QBL1YW2TbyF52bL8jZ487bmcxKehEzI5/UdGhx/GFI16ikTe1c5OsgaM4F/1p3u8Wu+JS
e8XWvx8pD35Iol+zWkULcklVTSNjWLKvQFuI/ITzIDZ12HQYN9CNL+4X7PQrR7Ibz3O0qElCHRy1
bmRnnwbyBW23jOzBWBlrK9I0vJC/NIE5Mo7IQVfUZ1OzwIByfWxh6C1tKRN9OTbPgyuuEErTLC67
YIFlxgrB9j6S7NoZNNWNRyET3tnb13ovCWL9rOJrRd5Rwdu4wwaKtE3OdwxOwti9yrMsJZ8rFpIg
BISJ9OjJq88bXLx0Cr9hNB0OZASIS4PDRAzo3/hq+F7P7ORLMJSLSIi2NnWIk82X+aMYxD7XNv8Q
c1rg5zq/c0xJxqJRodrukcqIM03SHudiXV3pEw0Ul6KqHy1R0gNumBP6eeXyLI2hL+E7JH5EuQuy
7SEE0dAW4nIrhdXLSlI7ryUfF3FAEt+VQu+UplihZda/C4Xza9utK5hjqYztB3XyBIMCwBcIiwOZ
Oz2KW+NNejTGagNoCuj4cWvHL/zlFCi7ETWEzWhD6EBO/2zJQ1Cf0SFHb4NC3Aqkcbsm61ZpgYGM
xU4Rws7XWy9QkdZ5qJIjnQoqPhvEpxaJNNeDPX0ugk4l32cRlGI6CwsfH2JI0tNvWm7aFTX1wh2q
zP32w4Ru4scOgrFh6dq+b205hv5Ehefi+N+b16PLq/kbo/Zt+f8iHJdhG85ND9IyJZZU8Uf+bPOW
PzjsXAsQcYLmJNcS28xUf/v9StBwMFh699pPSWxoJ0PZDMHx1Me3//jMMa34A9hopUXE8XPuPJ9l
pHhUJRUnLLdaZtUzB33UsBrU/zVtrasKWwF854NiwE844uL8+oMpufI1k1cs/8rqQ2PosWg8K6hh
rj03Ev6ibFmPHKPq9Iay6QQya9fpcBN7rCw6hdRBQubDvjyIXvR8ArNeUaRYb3MvLlR+Xg1+wgXx
u94NUe1BOFYG7uvzAYAO22fV8EYNtbrFepjY7tqioPtLMOAV2o7AvCV8nlsS2AyZ0ypgfsc4Y3si
UEqf/i5HZhxi9wncaqnTam5ue80gVp98SWFZshF/yrWP8YNvd+PXygBCe5sB+H93UNsQsrTzKhkJ
vD+Gq/ec2/cVPfQQTBsWJ/7K+9lTXLCxOq4tCK+019bXVc84OKVi0DsBuR4pwi3Gy+YMoaIjpdMw
ypFR1ZFVbJOYTNUU0B09OrY90iiPG5r8vhaY+bRR2ycqfMUQPdphQ+YPNC784BmU1nMOgmfCOnB0
2zoziflcdc+zNlJDx2hlmpL/QJfM3wSJAlATDiQTM/jhEunkFV8MJ8QYNDygWozLja/3FDESGJVi
yY3jbTVYA9utlkDL4EyZLz6Qg8YC1ZK1PAjaMAW+t2jHdowzOBZUmnOpe0xVLFFtO9weDkGSnSw0
QWk5QicFvSueIjO3liM3QKT0hWqB8RHIlbnI3hMaLklSZ2ysseVrPEzkNH7vD0xm9ryPQJxTfb3b
pM+rTG4hrJXq43gtjcWXngK7XQkKrF4AmhoByML+hFTRaTfnoKSoXA/1FMmalrOkwnadZ2h3aLHp
8JLQ/VD7jwXdzs9AT2FHdbfzabyhKPt/xTQRVzWZnALKtoCtHC/XOfvC+jzxOjpTA4+bkazk/Fcp
eOQzvsxj1oPRh+Apg4RR6n0TLLt5g5+TdcQJtKYs0QdGf1fw3ORD0CG4htvMaIFl7N7ahLcjKr5p
kgZ+vp34zaxwbTlw+PKPE5WlUcpkePBgBG8dFzLjzmOb4DTz8iUqaHhuNMsAABn9Z1pN/pUkwcBV
xkmlpEQLatkQbznWQAjWmRIXIg/+L5kpGmm7JW4wwmdn5B1TV1kOqyJB12F/k4Zr7T/yZq4LKOIN
q02gM5CSxrg6LSjUsCmO83dXfFnHQGh3AZOPST4l3RaTaKem2uoo7y6skHYN7/9fTF13UFjVcDBy
QKotWKx+7Z9+yEz6hl1le4W6u1K6Ig6GzWQwjAEhpCDF1BHZGoqli8sJcZGlXRfeM6ysV6ipVEJM
nBLrWlJ6hAwujxpqBVoGmhXKRTg5pEVha/H/SLSxtLJaM++AQmIRUk0B4WgbBDL19r7SoY7gSnWu
dlUmfwIK09ERL4JgXZx8t0OB+nBoEOniKQ6+kdxDpLC4RGiBdgueknhU15H+/YIzwPxnw2vVzbnH
xGtAOj4Uh2JMWTnVS82YwhDuT/cBeLjCOoWvVHb48mT+i8xVpMAI7OIWwRywhgN7xdiZjUx+Aczi
PJE9SzvG9twW1FHNCG1T/OneZg7dWfiteE4j4+H6JHoKIDj6hpiFZASl75eA1zWzyjRhPSN2s9BK
IFo/aYsBhtusaWsZXjmGqylNiL7y0WNt8zHjd0J8gd/UCJzwghJkK6ck/xBVgcHba1yi7eKNvvz3
RSzWd7YytTpdbmhGX6zqKDy0Xc+mnvGSl8LtNPjEBSZpUcU+R70x4r1L8Bj8TBH7KMlbbKQpE+hn
TDJUf7wbvTJY0RLa/L3y/mZrDUVyOkeKnTIPMLuCHCunk778B7Xz1GbpxZMDIbKjBTMTJ+qcr6dB
WB4ps2VkoAzakVT2PqHfNHNV0HheWwjPi1L8s5ZuU9bh2WYXMUnIh1uqBQ1oz/tZzImqO6eBtAIN
nrFg2dg7/rFW65L1CiJTU+N+ns7W5ifbpjKwHfZfeg5ZhI3VL0LVDSXCeBHgegVvqT7KN+iEmbsu
wbXmj0alnO3LlV6q0wZ5f5nJrhr5W6y0Y/r9e50a/GK4CgNaaUk76WT7z4pz4hp1mlydEgN+TPz5
9hIEeCLpbcZgpWTUkjXEw1exEea5OAEFxxRwBbKAO62Kd+CAEEBbu8/dG9iiopCqCvS9xbYzU8sP
taeU4KSRO2aT8ZN9Y9I7fgk7QbmfVrRRb3jzlP7UGOLo5a6RbNNtVZPwMgxoNnknl+Acx0rdTq4a
nCV2VSmLCEnspYykbqjJ6bmrRJbV082vOmUF0/O5aECS1147NWa11M+T6m6cZT7zkp0gt7TymjOA
bj4XLLw05dpvOonB87g2gwxSe/MoDRVS9si/s/v1VSAOaS6RYQIsSDHN/WtHoYBxIios+pD21euG
5fagh0QS/7Vyd6btk2JyYg4TPG55odqbEsuFqaopiGEuVrkHVEkZjWHK0Pky3jzUZLyxMrABgikS
3d06nTXOU+F8fjulz3D3ESXDf98z4ETuUWRg6Z3W7f1b5ohEM8xYkFeS0tjw0JjWMXCb92/YtM3o
rVkp6BLWxOY45mf7rtwUnC56Sxk4bQ/9tYqfSshQXQshQkbrhlNvmBMjmeskz3LrK/9GNehP/ker
W+ZSWFwT/7Z+H8TBHKIKJ2piM5pNixMMWakCfZPIWL6y2m4LFeVoq5GgxufrVGv+V70Ft7eqoEm8
B/BKb96LAURAS5BnpM0reJmhiF1Ip2og9E/T5WjnzyiO2VKRnFis1ncHA/zODQHW2KVBmAmw6Ebj
DJxjZP0YMF8/RntE26qVCg94t+AyMI1hCTXv6obs2kh/MzILdREivmDwgCGIE8zVB5haV+8ifEpp
I7L+lSI6oPA2VaY9pBp3uEj3TIW0owAJ9ouK6BMFvOfGsLkF0mxPiptQFlGvv76ALZ3M8Nb0QgJP
LawQs+IY9nxDI7vVEHe6lpSQtBk+orKLT75q40Na/HUYX2rXW4Yu2k4CXjmR2GePJawfnqypfBXB
bFPOI31GqiSHgFUyKvQaT6OAX7vEPXwAXyvcATXcWRalahePZdSY4iezuV2ikcnmD9IFqab/XdYK
0MfQ0DYL6BW6uvS9hwEq0x/LGCpE/DbV2qF12eLE6BWzqAnROpAQdXPm1mmocWtRdFJKaBRY+thc
1zq0xfdIfi3mYLlfcXM37DLPcz65HH23yJReAuPxcLitxA1jaPnb4+SplDSSZr2oMFhSEIIDSro3
CTOi8bP611qDvqOC+XCtFq00sdyzwqDqqwfCE8vk8/VjwrCZYeW3BCq1iUL2YMHS+LztWwmSGORz
ucEmPgLzVhe4kEzcwmqnfsSPB1XKockRJOTeBLNVYXQLs+5O5rLIo4NCfLjAQhLgvnmlWpv7IL/B
XeGTO3ieHA1qLDU9TjADE1x4Ri255FCIfc/hssPGTtf4N5hOs5yoFn8cJR9sYkxX/S2aVoLewkCl
q4qqET5/YvOW1oyUPeS+i8JBl9Xl+bMzXhR+DF89lt0Ltieafpew1sPrIRNf/59mJD3yXVdw0coO
QdoFf4q9RXUgVM45aNsaFYLnp6X2EJJSlsHqLnZfdcwUmBcBBrpEZ/ZH5Xu+6cf3qQuK++eNbKOj
vzisu7yOHh3CDQzirph8aZusBf543UfuoOTw+uSCXh47AC+bIx5FT95FEARCvKP+2dTr+k8s4g2h
RYWX7ljLzBS6sZWX6lc80gXe8xy0qln7d10f3fOp/rpcwCAAt9c1bADbGlxf279D63Tr5Z5Zi0Sx
stSHJZ87CPFu1Fx3nqJUpFPOHYlvAumS+Aq27845UNYRB7z1z3OyYi5q2dvrqvKt6MnkGTaN69u8
Vk6C7Sr3eDlMeeO82N+yV4zZon6LYefSMcA9g+5jhKfF01na2uDuBLzIv5iaTv3fJUvcNugDPOfU
o9binXmeWdES0UN0Z/uDDSJrLcIG5/61tc9Pt800dmxCdeHsIafZGrhk66MN8sSVJ4O2bEtUsoT8
caMp0Z3vSlBR/26pU2NLdVeQejNiSGjwNSiiufTw7oCuhSBcPlf65HeI7mKKBrx34jHmR1nfMHyO
ird7kPR/kBCSHs7L4csWRbwwSVd3xKml8pvY0VjLTX/hFbJyVvyfKfWwaS3JHJMm0OqOEGbSdLg4
mzu9tM8uUqldm7PpEsQEkvCJ+Olzyimpg2gcAj17VfjH1DuTrlbPX+yJ7khabDwr8SGvcX9dP0oV
fHHsJdzSHpJw3VYzOdpA/dQYhlta9tdrp/LVrLN3YP6FUINmopAUPPMMSb4ta0DDhHk9BvwoELyg
4MDROuMIUeRNoEFtZeYzARfe3D55s0JjTAaLHq9IjGSAagHWdD9WjyfparOEHWMbqPb/jICm6Wca
SHB2Z2FBr5akVPaBKh1+34+a6O2Srt+DKawI7X2ifwR2yO9vyuYFHXQ30/WziuSr3U4TNGWr2sA1
53VSXNuQIB3FiRUYKBweFV5E9b94Om9C4hlztpNPvttxs8z/S2oSWnFis1tFuLO+SubcSA9cvgwm
DyZ/Nquh6HUr9iAcPYyT7T8zGt3xcCqHVXsmE/+68/w2xeszauiHSbzJQd6/vpPtWhr+q3bur5Ms
m0nrnQMkM4kocTi0ei0+aDyHGu/yZPMcH2wJuPooUXn1S6GzIbfB7ZdIVzsLuWFFQzxuQK2INCAG
enW8BCEMHooTCxAM3315fQ5hTW16wHSimtGS2vIhSXc+39NgQaPayVLbICZwQpsQDX6BMjSd/Z5h
JUn/QvAajwBg3Ld3AOGztJif7BgWnzT/SVqWeCPR5sm0eoKIsqKf1coSS38hLbTJd00JSNJaAki/
GDrlXj+L9ZPTN63PBmk4VEEedEHxqrHwDBQSOCUoJ01EPtQUcyGuqiQYvbXLfPfKdIQSqwekSVIU
nTjiW4eSCvIuvhYpO2cBwSqtYcJTCgo46aqY/ST4HMkMfqCAJKIiQ/TFNyZ/uv4sIkoG8iMmoEmK
e0+2wSgpmK7fVnXV/cUFpyThdkwr7HLyJ3DRPe+YME71FTbuA0ILHBFNkpGzk6laX0ICPTL3YOSD
5+1LbLB8TFV9dir2uTaBFtL4RaHYbSproHTcGomB39567PVdajm3v+wyGhNDJyZs7nIZwrFBNTrO
iSZZdCqagXZXbIKcS9lOPx9UMQUvQrALricljbM5AOVtI9yfX7OVDA7CbBcVA4VKtUOoC7eQWkN1
Fs9tUgaCDEis/4KIb4T3lpq3GRqbeIJIOOEKrJ8djEcje39nNqrMaCxWdPzcCyRMe41fgbFQZmPC
gfId0nDCW90JDB+gu/eNkiiJxRE/IP9rXvWuZQpCyLE7+0piOOHrv9yVyJzk+DAStAkRf4kSjF50
Aayi3xVCIv9Ji6iia/DAQf71BXSHxhhP/t8yXyfjARZBvW9EswRXa7yskoPZCxXNb8zkp2Q3jLQo
uwk6xnpR2L4cXkvs+RVqEhyM3/Q9SsPU+/0v/vom6nUaB+bEsQXZQkNJO9TZq4/Gd4oq4bsEGvWQ
0jipFfBnK+Imj7PxTFKxDRtnrRuKbcA8EKI9M1M0O0YU4qkY6Fbn5PKoVmAfROcvpcx/u3LR+0tc
X327Stmzxwjh3bbJaOWHnXyhd1A/vv7E8d6Qht9f809ZJWQ9/Y0QrwmyhvNiO7lF33u29AVJq5xS
SnF1A4Ow6P8/Kw6eHs9afDEzxP6jhsQTFxvtq62D/ZN9K2PxL9QXySvhIZ0g0EZxTZq8HoszJ64q
HuKyKWgoMIo/Dz8CyC5gY2DKtJcsnsgrhKesvCDAnCpoDwxlqoq/fq7W9bNDxyTym6YWBuCOVg3H
K0UrjaaYrzgsI0cNEJ7mUNPd3H0RP+xx+5Prl9A/3aGuDNEAaPkkAlJnES0UpbCjcZ5ru2i4DeUg
38nm8Wy3aKC8htGrJPqah2SXlDZIknFRsrTi7EhLq8gswvnk+kbo98xa33gAPj4mU9pypgM7p7UF
r1RBWjw1tyAZvjFwaAZQ8Fl+VnVWNq40AECkez4UpEExt/0HKHJwCwtM/hy5jxA56D/JUcKSPIvS
ZiuxC1C+jfrtBdCq6iyn3l9jXgsqIF72RY5XbsTb4w4FMtaNyt3Hchcw+qiCucf6Y1e+Jwmotd8G
JHWv5u4jARNHcYNUTjJibi678Vh4A7cF2XT/6d47AkDCUFsT9Gf7w8PqK0TSOJjpiXmNIT4TKsIE
LoRxI+4dr6LDHysRBwTRI+BO7iXc6PiC6CC0oTc8o2Vl77sIlJXz0l9tOei8D+TTT9orWd9idyvP
BSmD/gOHeMduMEZ5qsEriEYOGRlYYfkz0mVVdhGZbqHGD3UViGhx7KHpMmxnf9GvGZNMKhYPXwYq
Fz65aZ7iK7Yy3iM8yVasaiiTOLn6pAD/38L6Srr2QY8K9rm3O00UD8Y0DyQFBSncBR7r1B1hOrP7
fgywSHx03c7VEus8JwyFYdtvnVoZkY/+zo8M86EHFnVZ1B1r2qHEMEPbd10WE/sgdDVq+h20DE0W
pBX2IYAgL/4IY2QZLfIsAq49iGU38KiLNiYNDfkligjy0v8xl9bQOayMDo6owZZ5L7SRl4qPfQAD
P38RAzlTuuuFucHprzNbuRjQnJZPL4RaA14mVPtCVXNLk4B7tXDRoHCYP+KSCpDJFbEt8AIq72/b
+ksrDvbQ9u7CKZidVMaPP1NuQ07Nu7KCIpv+q8gj/V3B/hPMAb6z2MLa2fvF+3ki5h+C8q0atAET
esGW3BDsN7+PIKDJdi5pWLN19kUp1qleJbTvMv3rC4RlunP8H6oQTPO/j73Mx4k9g6yI/sT/nTw0
HxjlOANrsuA4AmHCzvfVWo0ER55weDZjQwIqnQvGzRYxEfeeCW89FbEYPXz0XupdQhgaINg4+yU5
oqZRcFz0LgUcVkl6jgtiIoofrPgCfHtf4DphO4RXg5cQyVAtUu6UcpeZjGT/PiN2gyu2elhqss1v
EllnGGSZ6pAUyeJs0CZLv66MxtAKjhdxc/Ohpe5f1YV58Quev9B5VUjnqlMEHbxlJu/elXgAlvTg
f+VyLjYSAYTTkH3IQW4bT+zzFy5rQO6LikXbtXd2HWpWQz4PfzDfeBhtAAqhIuqUlw6cb1Lf42y6
JQg2GzPQAPRmDelbU2hQafNn2k5/Y4VkLfJcJZHDs/I5LLzEXoLxATAFvdFNSgf2gFr6WWlIxqGu
SL8xa1ULy5tDswkpArtNBrZvo4QNGwscMMQqNAsQJZ8uSeu4Wo0+WLQA2GlV9D8fDsXdnLEIhusx
ufpKj3/95FVp4Ygi8f3ojdN6rrTfSIKmyN/OAoMx/hl5CtsnGv3A42CCrtmL622uw5H3MiHG4zpq
BuzJA93tPF90uO6qcwMrBiyNl3XbSrelIqVesiZfURn3VYE78Fl6nBDkCm4LEAWgvSa+NBiJKUy6
i8JpWcuVN0zEV4ogfS7GuDUykqKDJhtDwN+VX3TNHxlR2MLysuZTmLWx5qZRPXZUTF0QbSl1AEQr
grsRLfniQ/eaRHHDlY6aJWWsPgJXdlJ8kWjBSZ56n4QnbkPJksLZG+ZRN70v2Bok2bgUngCRaYMN
dYhL7e2TNhVhIOgv6ES/RTYpynS5cjtKg2yqbr+f8+/E/+AY2XKMB30xhBnyAk3bHA19PCFTq5kC
maNyVw9boBIM+37XOTgnNutLpfF3Ny+qviYeEC0wyF0a1+tu0SJvag5l8bfcj3ssi0vAPZDOV0ch
SOkx8Yt2lPOVprPetck0cO/hBoJ1QWGrWNgQjTaYiEiZ4mZCfsqiwT09QUZ0IEjfmMWYhke1jBSl
qVYMTX4egJepI7rJx8HGWkjQ/04rPwswuJsi1TW6Wb8tSkEJ9ck35Loi66rXFsCGO9/ITVFl8HIX
/jc52tpkr7KIdFgUescrZrnR1AmjHr6dyT/DlLqije37XqV+xIwrJzaYkIlORImyjhpQVdKVWLZE
C+IExPxW6KG0wLx4QFNsZgluKfk2VZb57CzJA6RrcyGhpZGj5LuMN4IK20VKnJcaBwDJ2e5vNFDU
dNSDJRrk4YwPsJtxJ1ayjX6KK5eH0Lf9s2bbDMB8Aoa1j/o0vtJFz5xbuaG0nm5xnU7wHuJRlHxd
iBqvGz+ZeopCwPLfxkHNdMquJ2ddDPrpHlmyjWX9g6o7QWL1Dxmr0hrJ8uWAybNuPDawcUrG10Yf
r/dz1vsL9aOABu665kQtaMr91+52e3SVfIMjPluytZCn5NzqsKForDaZJVh3AlJxj0xdy/0FtWIY
jTKKZmK87Qkxbe6JKE4g+Ql4Q0+Ixn02ZXqau3KAhSfsjPNL4Al5Xt61jugDEfK6P120c27OLPlk
+qYinT+wCWHQ8O1CxXNbfWcUgbLHpubw5ujpQbkH8vg37yFWuOtrHFQ+BJxY6pT56icZJ0ht957v
jvTzXq+LHC13q/g3UCchoNVP+CEuxsQu71jDE1UJUtGvugR1J5B3CDQZpJi968o+05eUR+BwuMcO
5X5APHk/+44b18Y1u6dOGWIiZqCk9G+5q/8Hz6ynKo43MrVaI8jVHOdncCl25nDZChUL9J1ZFu+K
ZREJ1cT3nguSBgE85oPKSgW28Py5RnUq3eLfJJf5Uww2pBR/pA3VMZtZUfM4HrPFo57e4GuEygrQ
+ZjibVZlX8CuRtabd2LcuY61BwlT5seipes2oY8UHYa8o5ZQMl4+xHOgqVr/5ztQDnUpVQpgmr1F
5/zACdN1mQhbskxMh8U02I2irRjOxMAwIZVLAQFvHQCzAeTXAK9dmVG4CNK2Hp5uxeLCcS3KIupw
KWYm+a5ZzNoYzX6SH4bORb2IIRLF7zTgfe4fv9Qys3QK/61GdASBRfXr2myhhWsOfCSWgF0Fwy2X
i/uMYjDnBwFj+cFCJjlkGvp2rKv7bikZO4jJ03gSvbiizslDIoa4Z3P2N9sVqwjmLWRf8aXzhfw5
EUcJriniYsZ1+0jLb3sZQuwZykvDqxT2TlgbAOvqIgelj++bteycDbRrTvHPmWgRroYF26XBeO3z
cFWApT+C0+QbggbLgLSc2asrOHvvvm4Lbjoxf/aFj2KT5hDUzBUnhZ1f6lVQelLfWd9g7PRsQw7w
L8rUcEdWR7Zy8M5FYxPf6NUyG/5MKFSYR2ZDVpdTLIt2ntVs3TbgzzQy65BUS3yqyBigYP9VxrM2
/L6oSb4juNRrcUoblJ+jytB0er7lpLJ6eq0F0c2nEZSPGxkfGI6JNpuo0F22aq1PNriA/ZqW+Uc3
udAGi55Rls8npDqXbJpWkouJVTGMTy0alQSVNxq0hWzyq+e346z6ubz1IE9V4WaP1dWNQ6TJx3Y7
oZ+0Tgb9fsECi+gn7imiMYGx//kPrjsDoSZZVrouQo+A3a7Zr9GsHpMMm6TluMrx+6LyAdeENCR1
UWE9Eer1N3qugpB32P0JnF/4rlTNPzjypB5K7izcrexHvUYo4NzympXUdXSSkHmLNoMv3mba44eM
R3c5aCXxnr4ppC1oc78bcExTaR//Bocu9WmhoDS/Ez9mwD3/mXRIA5Xj6fdulXMMcCI0OosLixY/
vtweGrbz0ssbDowXKFtYh2G/enWkZEt+nkKX8VilHEqhFXHaHOg7PLhcOesLEJnQrI+QydDdgiUS
dan1o6A97TpxZTIX5tEa6++EGTgyQaNeptr6xHMWmxbHROukMqdJ2pug6zPLAycETTDRcqYxtDPR
/ZiC7J6AKpjhKDepo042z36TkyKJGryOO1OtfyC4Yh6GX0cs1iJ7QrI5YdOkuocK//aQomZp3axA
7dr95OsjLzc3fzjQ2Ca6WH9FNrK+he4idXQN8XwYpLQfLq61X87jy41yV2K9xc1eccCgexotpL4+
4Vu/6LIo0mX/eqgnmnCYp2csPkwfA+cQwK+uBtV1zVEDtbMAUe26+XBAbZTvV0tVomN4dN4JeYfW
cmREgtmG/Vg4GlXzgkTVITXzF+Y7ROY/vkMvGWGm+tMTtTdEqR1EZSxN6hI6BjK3QSjNnzUeEPI3
twXitK6rArUgGoNSjip2ch7socd+8Rw8pcTYHcKjUDNHVU0gUdj9uMwqyfg3OusnHdGxUY7ywyLZ
oL+FonzpzSMZM0P1YS5o1mt5OHgNOvobYzJYapiUK03Fo0tjAZvwPIhP0XaoXP1s7o9pjYFHQH+p
Y/3vS+meafF566UVQu5kXnTRT5rGmA9d5eOIKOHOzd2V7MSk+5FOmoxUuadEI/RGmh6mzc8TyEix
NWRDsTNi67CaDiwEveWuSabdsyBT3fibaPZK9/ZvhBqUFBph9p0FFOewVpX5k6CL5Um0QapK2Jy4
BmCCp2/1BrmBGO/nBlDWEv2gCC+9eqQaA+RVLOsDq4nAmEdi+CRSxIxtzoadoo1xLw1dRW1/1tFo
fVr5iQ3QIKA6Oe2ga0IykrfLLsSaBriEjWcJGQ/XprsonnAGgwcd73Lm6HMfIOeA8gdzqCttrZpT
Ub/CyHRZ6Fqfzswq6eH16XqStoKUcPFOYg+BhQQluO9awIiYufO3jJMsYZl1gD5DeYbPRnduuBSy
OxVjTsKRMu9HjtO0z6FdtL/mYRgSXsh9qVJ5OkKekvjEdznLZ9MX6DYVkbylKUt+e+sQgP+1sOJz
yBB9TOFU9WglwXPSJETCqm6n8u1namIyojmO4UEUxujIBJzmNe+Ob4HLyIUs9nHGB56p/IJ60wxA
ghVZfgSRK8GuaBuTgn2yE3kEgdJ7xAFdBByvJC8nUs6Ot6+Zfyo2k3mFUDFPpYvmKw7Oo2fvwlI8
oebOgdheqbzmMWYNAxB0i00VEPHk6THsTS+9LPiqZsyquMNq9H3nmhg7L2tGyaBHuGUeaNpiox7z
7QHezPzGnyF7OVqDvGHTVljVsk6FNqoBjDKl01YKzTkoevlahUef0PDsIZIruKtyG+vLau45tcSb
GAFvVH7tgMOG3oYnsrO+3P9/YCOa0x428Gg56PqvxraFMjEjOVMhi3Vmx801SHlOCK6mtYnRXKr2
UeNf/uXF/7nJpkdsebHVhnteOUg2kMSUnOzbvWBQpLdpfj4VTIpc21OPSYOyTtmP0zt05xwP8i/b
rXXJHd/6v6lJCT6iisTp7K9dGUxKP7SVtb5TKHs0bhrZ4c+sJKFZ7YHF2B6nV9adbq5c8znZW1xF
yQ8Erbj0eK1ZDcVl49Y+J8CMNovV47difLv5NviE+aY2pxF9YrUKXJ3Rm8L6TQWk4kW5x1135nA7
EEYfjXKpTSu/dWL8B5+N6J2/iLr3UW9dl1+gQuRYeEP6Csa7fOQ/cs3Oi85rNDfliqdnP3H6fA2Y
+H6vESGj/wPWsS7XVoTFo4mvr+fka68qFJ6kB53DVHj45SZFLxz/Be/TIdbyqOC+CwpFZC8JF8D/
nmqMihK3/tYUlU9suIGYKBudmKi1YMBhPXNH1IZR8+HqIh7yKXlfkJzNI5t3qG5GT6l9L2qyPNBY
cdJQn6+PMNTr3NxWyboIM81o8f4OAuyPnKHSZyA0ur2o1U4uz1ueVF8bbNVgsYmyDYyDMAaQhOoT
RsdNt0AUIQPF8I2tlAirHDHhhfjZiGPI9Yh2pM6vPGZmxVQztRQ9NJPzppgdrxshC80hhUsUcQ/7
jOXn37MfhxHfEwTGuPWT88ijovrRziEBKfzNYpyE3g4huc4FPt4i/m2yXUq/svA34FB+pNa3OyQ3
3hzrBkA5DCjqVIcX+wRaoZDx9zsS/V7EBYC8d+AisGgN56uZTdCqWNJt3gF61sKIb+dVTxCmkuNw
e5dO874eNwJcFG0WTkpjKE9bahA3FL5eb+Y4GQlypP4LFBX5zM4cLlFScUVDHuU54AHwpSXK+T/v
OTXJsQlXC7J3DT19HEM4d1HRR67uNPCTsMpLsM7GmGOkDmrf9Ak4QvvmPZEUXjNVqvDYnbrwm0D4
dPKDIL2Ky3Jv3KTkxQYJ7JNk4oGPu6yqf4AyWJbOC0WTjhHdkiduiCU2pIjpM1jNigR82/izoXU/
PS86UOlUEDSuXRDUVUtSRPTFQONc7AcN4a0w7n4gwQVSVAcMbW0g+dJLuWgY2yr2EwYGJbr5ONta
LfQ04nZraUTg7bHhtb38OsvVFbU+1ZtvTBIVTUsw1FbaxuTaAbUbvSoRE627lhZRY6Gzp+snEByV
GNNLTNXaTvUYFAbbBxfH37Eg4A7OAGY+DZtdRDYT937CDSdkT9EM9SShZu5jrM1wjS5o5ENLb70i
5NZHctwpqBAZuWABRdpsjtuGtqjRtE7D5a1RGblQ9fWhQDb8/C9M2JaGCvFgTwqhXLZ3W0YFK3dW
LH8M1UnS5MXwxx3aDHvdKw+3Lrs1C7AP36+BGgPgQ/3MiT+mobAIcK3zYnVIpNpfCHc54sgs7C/a
jEunv7t11hVf9yFfX9qNmbX5Am2sq+Dqo9PohXKfU5cLr/wSPhkQdA+PC71TU7M1frHbT7Q00496
HJJ8ksfMxePnrBbCvcyDDxgEaDLQ9DebhadSzS/dUh+QLi5+UwWWmtlb9qUBAZ9aShPjvuAhlUcu
hvIywj4wk2Oau9Bt+PEoHclcaS50Wh4e3jiZk9m+mwzcQCjHcXkuW7DFfER8SSA=
`protect end_protected
