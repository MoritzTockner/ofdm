-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dU3Cw8CmZMf7cw8PrqUxRVKt77lmcr7UQMCQ4QQSr/VrZEq8WJ7+BPXYCZGwbSfq4NOh2Pe4m0di
74dRd0HTx14ZAnZ9TRFuS8CkqFHT1QMMJGmzkFy5aqNPBg1gfwfh93DWGUTmeSNJ4NyYO6wFuClY
0TqFYosWWjzhxwe8/sstgN6uKGOzwe5Y+H1lyFaQF0nENBq1W2vuLDiwj3ej/Ht9cF5LwP2iaGD8
09uYnCwHUX3cD7QjjZptRWvdL3Wz0WUhxHa1vkvdECZ8lEO20qhCa4KJwc3n8MMxfOzO/vLGe2RX
TfZ7uPIgyhkgVBSaDm4BCkTS4jeMQOWLXz8/1A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
qeppsdyofw+dxwSlFvhN+8jgnM2pvrtMAX1MetoVXPibkt5COEqG85E4gG570pnitXk0v3PMvTHH
DhdRjsnOj34gsOBh4jXJIC0mQeuIGEn/cfKDLE0WKi45XhIoXBGGeM4KOZdqUS38bkPqKEQ6gv16
4VRPwqqxDr6bKDAGM/B739VoCYfCw7tMILEzLMulBcmHSMY/lWjHMtYyKbAfWQ0PtbRzfNO8mEmM
aPn4YUTwaIc1WlyWhTCBR4jEgIhxk+e1XgGRnGjZJpiMeMxS7Khqsa20p3JcYzNkmfhMbWa0BzIj
aWde14KCoxW5m+Q+Wk7IvS1e7M4ElzPJoEEpB5XHac+/0qcCcLua1B2Ys5y2kXTpEpbKCYn3k0Je
smiwyPd71I61Brv93XfHoW42XyNl7dUy5bXUACTYogtIG/CthCEki+ypGymfKxwpuylNX2eI5FPe
WEli5/UbxXQUURm4WCq1cIM5GR7oX+sfeIEuEs1vtENuYC5o+kqiKAm7jC1PVNBM1lfNvzsWYPBA
nwh+6tWKn647WjrHi+I4wKo2CnDz7ZrkB8XrA7k361NGNV9jrjwTbARUGjcEJPdDkCFCAVaPowQk
1UuJ0fPIR3emPuznQhCnGR2dAfC3Gfvq4ipL2Q8mo/gqnBUo7fW6saSZQy5YXp0/4/vo+cG6n9pw
Vs9YCTuA0FjEhMGgv1bJHSj1VxImI8BXuF0VqkO3OqQ5VzZAtlFPvNIfHGTl/xFPNL3PIFKUlIb/
XAS9UKJV50NbtUjn70BzdA8JrxfAJbPc9NbFP4DH5JWT1qkXAKTXm+wLW7DatUqZipc0fYivy343
/UT4nreSGXYDVwc6HgdGL/b5U5yE8ruc+hzmdSNs/4UigtBitssRUfrr4gmhEiClPA/bXf9+LmDm
MQ9/+6vmtblZRJ3e70ybRf+grEUnn3XLpSkvYGoLnq2y3pkxtjHEU9dB+zt3e2R1w/rgUnAbblMe
4tUoDKSknMbnU82sS1ZdtQdp8kS/8hnxx18Dzs3GId/ZA8EbGxigBdEygBu1Ya3+vVhcE5pQ+MXb
5u85Cbb78lXvqdfT/92f0j8bI7K4Ky/z3tHLJVaIraUqrrlHWIysyvl8RT/9m32oz9reWynSJPAS
hyPOn7QE2ZQULfhOiueZ5S5R3gdrDcTGuXYvbXleHLuPuS2Y3cwzevF6XFpklyRkh+DR84HrIGlY
Zcs90LLYiXe5xuXK6zWk4YAZ9YAesatR7ukVKS12ayxgHl61l6Gokj5LVtIPvYKxPF8hKnWrgkEn
JCL8npGeBOQLtrtGKi9sBjE/5vRfwE6t2WRZVqaAewnD7xtRvKHrgivP5h1iBkKIGshkAezhBefg
Prvkr2wm84PH17WF2UXjj5CuAo32mRXbEZhGzolhRZx94+bnb/jaGos6EHlIJFv4MsCHhPOYzoOU
NG7FQqJWcyzOsz89kTO9/RTBegTj0OL1oEIAcpXpWYvRhSen/lmStCT6AbEydj3aFcRxpUcSd4Md
Ze9UkqiXIic1bYIClonBNwuWFh77Llmg/9oHsBOdEyQXYu4mAk+ovxELGyMJIWHj2C44k2Y8WTb1
8Jyvy5aEj5YvvDmW6PC5DkWKEriCWvbFw9c1mxzCQw8lNoLSbbobWqimb2YD3sHXjwGIRXlWg0Qi
sgKkhOoMN+Fa5vnd2uRKRIkGQjhRe0yPkcEGlA+/j/LVjGeJ312ZwM8IFkY8W7p4OFHxam0tSNki
tx88VJcwNBp1tF3qQrCIZFwUz90z5/IFnN/qbao9ndgEy450laylrfpdcun2lcoaXJ3owsVUrHGK
nsQ8fcId8I7DhNTD/ZV1Wo9RSxHQABc++aewdr9tELw8NOC+xPSQCshZjSN+Hu7sD3VjDhd0xJ4m
SJPSB+fXCqqYEFse2GFQhHL41H1rKQBm1hPqS2uKXJtA4qoVFlTfEG12Ir4KNi7JfCzfuh0+5u8B
qpwj279oEMHxpOws3UV/6D9gfFZM3F9lmc1f1QyBJ1nf8kfDBhUV+vgn0MxO69PPBvYWCHTLSrx0
sx0stpwyszucnGF6ZCEItPopyvU76Ie+G9B9n3dBvX6IVjIEhCQEbd7RpKl45B1M4soPl5U+1QwL
WJgWDmdrAy3tix6zWIew9gxuLcS1qYHd+jQChUS5eb2VNQickIfGac69EY7urSVPTAAAM9taxTf4
aJbrJ1QaD1oGWIiCwPWZK1AJb3Su3abMSeVNFCFKXslpwO0bqMHAeQWLrhrOD6CzkJSx12aS0a9+
kG3M2DQPwJyiIDRzt2Y2I1RoRXnF8Ak5vBxqXcQ+pRrzl1ch1YjLH6Ytk+8ROonEY0DVd6VI8clj
3lfPWkAeEBiU5Rrfu0HWVlNeRx96Lrs7LFKeJpuZU856QPGfIcEXavQw5Ke7wxZCHtPh1E1lt4nL
p1IV2ylAuNOKh23yoJ3CZXh3RUZqRKVmTIy5xOfI2LH9hFqBolH/v6tWqniwPMyUdrjsIXsQfmF9
7ZiwOksTzY9O7us2MmTdZr3XGW1YvHai/fSDN+obJEX9xNDV78//xqcXTeS3yl2UoL9U9sj8v7L4
fZlhO2kNgAPi4LGzD02iWz5ysQVWHVkgwOZMwlVzLsfxwMynCvugjYy+jnrW6fdTPSb9TkU7qrb7
pFM47T9GIUE5wiHLWhweUvfHXU45GrJwVCOHojf0/IcmOXCnBJ/LMiFDqLvyi8IHvkg0nwmSKvUp
w0VZ8Uvb8mBJajILi4n+OlXqbREd/LGXKVSHw3Vvf4aEaS5IfF375ZxTpRqAnxviqNuqR+M1K+TG
mQ6bu9b4HrzDl1jHHJuKMBBBPsM560zT+vB9RS2OEw0dlE93uubuTqfPP2nkHsng3IYLwRK4U65X
W50lTs3M29PGPg8/NupUMcnL4dxrsnhpxUK6BjIje6za1NPSNhgIo+xMz4WGLDMFavPVcud2HE31
KIcC1zS0TeTKm72lHYO/wyJVOvBHl9bbbuKQ5o6YBJekLBbENKiXergaUkngziWthPu6RNm4xN4g
xVukTUGjZMY/GZIwNj74muNQ/6BIE6xfso6zw8MytSou1/NECzBzX+vUKGKlnI8WQ+Uz1gwBFyPL
engoQFlKfpm406MCajutvcMpowuJZ9tcs8bxaXJAStyTiBaX0aEx0Y76x36fd6mAqojM4w26aMQz
Dg5qrdxHI75v++za5EH9ks4AW9qMBmnfeYS5BdfMOgW5Fb1Cr6zmZazCuztQ3h8g0leQrkgz8hTq
slbP5pkdAtB6UNc+nZ9q0F0YEPkLjmzJbc6k9EAJTmtMpJzeSMSKNT5JEkNt3Cu9C14zgcCnAMF3
6PgRMBr6NTQ4MwWa1vB4A3HyXspa0je50QJjdvY4tLRRTUTk+Yov0EqASVfnWZE2Kw0ta43kxvOW
/QQWUL3y0/1LWJqtxspdkwQQ5ocuwR+I58xlucWT77Pj0kKYtee1QFTTc3ywCXmyHVzv3vvRKIR/
nmOAPMbsNVw0TpapLWK2DJGxLUNCArUNGeqzLksv2JOwPKvFbjZx35TxnA0vJad6aIPicCijCHn0
pNzyda+OB6yWp7v/RsK0XypkuLS46oA5p6iNcpizYhCW3BfEIsg08yC84JbR5qzzBrCPthHfevax
6QDCHDrEYByXZs0PbD2i24CATRRP2Bjqd85ikKW5vnrvY83VxAVUe30CtqfCoqbi5lyncHJzSr7E
nEsfT5WRb15iAQ7Qy974niJEPZrVGHZ05kOQh/kPYNcMR6KhBC26Ef00X4Od1XmdX8S/6NTrUOE9
gej/omTtBhX+dAzhZEL2GeYo8uEsXTT3n9v91MTar0dcivBDNvltoI8qs4FyHHQcZzMCRNDo+eHj
54jUCuhcvf0fQyMmdBM1IWYd6a8qByf++QLOB7cEvT1QNmKYGZ7o+Q3Y2cPGv9CVI/W3YFi5mAYF
g7m+c7yMHJ78WgW13m0KTOLCHSF3TgxctatLXi+qMpEjyzNWD7NZ036mEF5e2qGQQQt8ZvjHHUJg
G5dsw032vqeYSgT7luyU7qOgeUQ+SE5YH3HE1kf8i97Iy0ddeEyrpa/JUukqgZNYUnvRgaCsIzr2
iAZmPjGk+B5Ctyany0GewWjgNPXVjxPrzFo/Y6w34srQPk04AHVVV63EIq5iN4UuO90gwZvi6W/o
gHHqhuQyxr/bOzLlST2ntvVie3rium9C0eT3FbJ70vHfvorn55JzWqgLhkSnw7r7q7PigSuIDcrn
V7HzmnwyiCOA28dfzDH0ikiSGi2YImb5PBwa/IhA1tcC1sm/UbMpoDj3asX7/HNkWndPjfebKDpT
MgEutW0jQJ8DG1LwGzEW45JBIYro+2HqBDsjFg4xnM25Xekuw+cTLkgm+QK1G/fN4U5vqn0yKO+2
MQwEJ0Ms0eyr4HdXX2gaSsooZD6iHnASv18hslpSPm3oGoJZusl5rqatbNSWqvcuOZsi6BcRmVgK
XzV5W7g6JlSvVu6QiWNql2QaYV0o5HlghS865iUHFNqCNRYOs6fqwWuY4s/5nXK/uuTfO4unIYbd
3U6RPkOfRWXr2NiSwhvDcDjzWQ4Kckpj+9fNBPh7v1PRx5NQLXedFISEWMB4W7wpGl5KL2bTxBv2
cyTmQS3NPvECP8M0ItBo5V1gJv63O51eWFK/pgqUxl45H8ASYRhLqmev7s8Q2vXp98ABwx7U54Sn
Ons+kZWMg9COxcpxKy4/GQ0tM1dlZuW45PRZepqu0p1vaG9NL7QaRKWufWWTeCgYEBQ+LO8+lJ/3
JuE0/BRCRI212KjXB9beAj0+9cW2l3pvf/c7Zv5ndhUDZRCPKoDs/k8Trv/UlS/c72vgYWZyISXf
mixKCcOxSab39mYI+wSd4IKg3S3m/G0QptNM1bFpnz5w34ElH6y5Bh6pmPwM3AhOzPxs7LLzwjJJ
qCr2r7WjByXha9AaKpqEF1o+y0dR+tIu7MMWZc/dfDiqTn8lmbMwLbe9/3jDvseo4WDtUitL0J39
x2KFrP8hIXYw5T376boDWqDT1I9+BNYJRneKVreyQuoRF6qRpWqMKBe9O8/1SjvZngoxWxzU4rMG
rsUYeS9zvfoMDk03Idwo/HFTBHuABKyhAiBslIwIHtDdcwq4DZLLUxv122Lt50H3yhCJPPh5mkNH
TStnqsXwiheiUa4LS8lpQtnUK5hBZS/tawD/DhGudSD/NqM3iLXIZaOg8Z5VxUa/deieCm1lfFBE
BG1lnX/JkaaOhZh467PZCpDoVfWE4svkx3Hx4pioKlEkjA0lIaZaZ6xxbk2Swj7uqogu6mgjErqc
D8aO+PGMmP5we79D6ELCyh+Y9dVnd24p1bBOeMFP8W6HuStTRmXDN1/KLDSjcBmouq/L7DsJV3/f
IxRmh8EG4KdwCA2oq8KcYCZL/zr5ojiuc/eSkZqFANacEzMGvGwkWVfffqLgVVwFA4hL6OcRjrBw
M9Le5hZGyHeyTNc7iCdCw2YVWiiE4nIhAdBozSXSPrzgMSKvmjmYaY2YsUdIWLobOwcffV9qN4pm
dAIz6IZC3wIWhozyeqAj0Q4H8zYGtXb+u6RxBKw5d387uiWzHJHzJJLl/a7CbJZw59HDz6P6SM/O
2RJwpAvJ4ySmMPO4l1Cf2xQTsBPKLz3oXQr5+HmsZciMdPo8GeQmI98KHQUGf1pyWE9fQkDGWlyQ
g/hpGAgxwFwkxBMy8JOi47hOA4Nk4NQNHKzDJuij6CTC0vGm0gomBnY13RNyUzApjN90f4YjcZlX
4LqZ+RctrmmU4ukfk+L6G7iyFA50m1YHdPtn+VTSGowaA5wVO1Y4GPdsP2AmXCS5+1Vij7xiq5C6
fgF/6McqdF9yjzIBZTv4M8lqtce1II1e5yhzQEI2vTJdYSodS+BYPNhDugSR1YvL+qF4BWxObFEg
u3v0A6CGKkdKmZYEBMJV/ukCcSx6vn5SRZ0ahG1IkAfCkfqKN9Y/6Upl54kzyi8nb9UlYUPAJXtF
LIOfZ/0b2nK1JYq5dwQqhgLr56CFK4rbZYkAOZuXqzRSvX6eS1IW233ePHN5ZDE5biSrSkIfrPrq
YA5cRpD+x0I6fvcK1hrjlMXCXoZka4kfTN1EBjhwYjZwZzyipHb5S/wDxq6f/gCphnuuz4XHUokI
rxkkYFF2T7ylSO/pydre/E8Y8eqhNnvkAn2SLmtvlxw1tWS+z7LcNmFcJXKqJiO5x/Ri+N2QLzVW
3dj8kVya0rH22M3j5E//YpYCLXTU43D94U3P0mYmBDpAoFshocy/7EHOY4h9sILxFfKoYa9RwRqc
qACUv73H1hI4TKM0mnogOYZQl04CZY6OvZ+wRJbOnG+RQv/9J6lMP0Rjq4mOqIwooeKB8iOigx/p
tz4YQWB2aaxT4Em3Zc9Wc9BRwRxS2t2z4I93ftvLFZtGo0U2OY/APp7uxbb9kDJ5SB+52gILDcK6
7vCLEJwqWHP/tu2129xeHj5CsthtTBZhBnomLbAudePoIrkL0fRcjMGzyiLkfscmK+b6oIP5Tu4V
CUAx+hhPJZd4+nv42iibYQtFYwmn51dZptuo34HvlMlmekoS1sZmY3fz14DY+hNgnndtj4ZAKaVE
vnxjVbKsNlFTPIObdzj+/1SW6lZNKt1AqXsSg6eWdHaptt2KaOpZtmrbaSm+JnZ4PMDxYVsMLSlO
gPzELD0/0hg0NtaMGBO+BBCNdjHzh98oz3+VVzCNoImopqw6d4zXCxfeCtDMIpv6XaeEl7nZkDkq
zIKuXxZ9lMaJy03gtwSeODPj/326XHq7nQ5P1WZ8QUQRdw8a1ho7YNrnEx/R00Q2JRK/p6Z8c+u6
xVxsbicoH2CsKczjrJKk0CiWGvMN5T8LlCEJ14NW/jebrdWp+zTRoaUlU7jRz06pQXoEGLimPkcr
7Xdhn8Ri+XqQAQaCl0BIf1B2NnPiGvnCvDbpv7njBNvDxkfAbn5y9TSoWIq88K7tefyZM8AbNSVP
kzT16iKRCtoMfk66yzo3AGDsRpDigWdnCJcbgjoJque3vw/N3G0u2WohaJm4P3pt6obqhcH9TmUB
Qu3iQiWRQKBnHuaMOgh8DY6NtEd++hcev3scVUtcVUQWoUOQ9MXGFujd9yrStTLi+zCsfNZwPM90
3apfu6uirD9u/qc8a0aCwQlA73DoCPgiCzZC7xRWpAlnKYueDvOG2bZ3M9mQDtFtgPVv7bxgiEYA
1SU46wBmrKiJ4l7KK1unl7pp//nstbM2Xup6D1HACfuvVGGyVv+wLjxK3xijd+4q5r5CnxSjsDEV
F1yBXts5f9gA4JeZP4mfQO68F0QqAcsIevehRecr289U7LTL+LF6IA9LHAPVlxBE6L8cH4mQ4gcm
GEPyNjhFhV6+TyThs9SfbVqaUlp4jrBWH4hixs5Oi+5C0tmhI+TmHV3nN6fGseq8CkN55WuFqS8m
BRmJzlpOWD+zhGDinv4RIP5M7swITO5l0PsprUUxwTNxi1p8YlcjTLWWo6aIQujI1A+hK02xRSNa
EfRAd+c48QlzMyiihSI9QlJqmy90ocP6l6Q+yrMHbMhEVBlYvNorHkd+h6hX4RDWklviQ2wLom3+
Bv6z/33cBM85pzuEnKZ/txTRj5+9tRRSk+iBLbri8087DVoAzBS4BbaSBQAro+7vTqJS4GTsbOYg
8S2cKIgdcONH1ONg/45eTsOYD3nLC1Cz9AcCfEznDBTadlkgcmfSql3LIoUbhs0dR8cjYsIKvOup
AZ5suk6XrH98zHUlMGl1whB8DID8NW3TcY19LiAlnuJOTTNR8SuAYs29eYcgKLrFaSv1JwjEXhEC
2WYS50/MM1Y31WN/1hXLMumDlzdFCjSmqEjxJiaNOWXMRIntg8rMx7FUXYg6dRoGEVKPJRSh4z9D
u6hnnmd+WOAMSfoKVxISi7u0e4ZKqZjweHO+vnptPu8XFAT/iFRr8j61nYOqVW+0+JPfjG1okbsg
Xa6YGl8SAGkkHcoWV0Q5+ai2mC9CPRAL+wKVLc6e5gAsEWXDtqic/th5sDhpD9D7sCHyd+DYelpE
X/ezQDjUCQs3J/VfkAwqHx/uSY842sCCj/ifrDb3wWeTkoDQHn0cY3cGFeiDBMV8zv8ZyVov9Ejg
5rRzMfqheRRzfsDTp6Z2v37fpeTfKQP36tGVV0TiQtQG0iERbAFIMiLUuV9OSEXVv7Ufl1TykU23
IiikwxmH3umw+wCcfKtnAuFnSuNw6fPoFB4XpYSfCtkXFHqzUtePpf6BDrKLDQLjQOkjYnYuhfDE
b6FqgtatF0X9ewV80ZrwPUsxDX+JbTccIWz6HA6n2MJUi+7eyBOx4lmvnb7KZLferBzwkh58/i7L
SBblYEtEysVs9husnAzyGnlvPFOSBKJ+U1oddjuqpyeSBZAsXZLTSkczwrmuBF6Z/2dLZEgteUN2
CDHu/uXOqzipqIFV1AbvKyLt/weAhAkvSuFPbmVPLjvwPhJD/zBPd8qAUIhGMfRipVKAQdryw09H
CMf3Q2GBZP3RysWCZTNy+UBnB78Qo9YTglU4RUgl2ucOfYS+XmWeJxdS4NRpWQ63i+h1j5oBoA6b
VKFTlvGtVgA8uzwebmFXOmr4vZW+D+xneKnYuhbgx26UdSM6dwdNtTJLubmQNoSSQui96PLWkJgh
8JVwZLlECmo87fD7WJ/YI4oxM1FK3VFstNe4wnryd969CNU+zxDea5vZzWXv5KU2WR3SVJstb3/j
9KbgtHO2JtMUW0aHXeR7dyxg4XN9mVb/XM/CtvBK9a7bkfwx8i/qEJcsQgEtwRf2AOI/UTPN5vxG
6sOxetUd0ENYx5SrYhERDVz1Fu4s2tQGXkwgsd2j84H3QCtDywvYnqx/RgUOkTU4lnTZGiygH6tY
grweYdSJg/pajW7UAqNbnQv78gaBtTfAssmw9lCiPNgZ6rAuJGwlZcU4xgxbjVE8SHM5/3//x/Ai
aTR2NAd2+08ayB/KIPO37YAtseBv7d43+a7UXkVtXqVkjwQJueUGsnTMfl3EsEvfPKxUfctsOD+t
PGf2mpTBtF11F9TyIMPa8jW1yGynbysbFrLI4f4opM7CftdCXN8FNkGoWM8ph0Y8479dQ5/58mG2
sk/lp6ImGnb+RrteDDFBPcFvlVwldwEBPrHh1WX7OaQTAbOTRo7JQvqixc8jIH9uC1CeyPyRwSM7
PCj0erAjLVHSfJpjUxNLRLf1ltXekh+bK+2dTseOrb99B2LvFrdAND7jZC/VHgy3e2wCocH+4qt0
FAJ2l0S2axjah9ErFzcrd8eWplNf1pSmWvuAWQcxI7awa1ACIzj4f1ua8lPb1d3CSDTl7ASH0j4p
Kvr4QQBMii5DxPw4Qh/NZVSym5bMJUlqxPiqeh7RDic7AWi/Kobgd57P6JnIeKDLZFuH21Tb98OU
iO5720YMZHvGpsqoKJudJ9RlsDjahMFl1nS1H8QBLZX0o1pMX4pS611/OL5GqcBFAbeTgkrgVty/
Sr4jQI54a/ygxxq/BwL1m67Zc8N0s3hjC2K1TzaDyoig1CpmDAtg83GIU0qjslj/CNWxdiLP5N6k
Sr7jlBI0lv5/aODFbGOse/hRD3fmZiSUsqJuzn0xpWlNu0sXbvyH/APBKcmMZ4w2uAnMkqB6T8cn
A2fAX3gFgcX+cQd5PPTrk2u5x+fTLpPHcnc8i5L01i7NCr3BtPSK4idaYPZGRK9z9zA3lf+c9P5+
4u9Y1Es82BF2pjBgL8VE124qomLcKuSY0oP6WqsuE8FuIOy3A7eAopPeOZvz+0yl7BU6mMuAx59R
/rWaHQAVqtZPO5ZkWa+oqGUxnWDrSsC5EUUYdwRZi/sEIyswFEnrQB6C0mDONlSv6scBohnwM3Y3
wmTY1bM+9cvrwbrHRXPOXHXHrm5qIfhYJSrOs8r/Rd402jrV61ed1hloNzr+4Cv+rCxM3A1ybWIz
/cEUkaY4RfyVif8ThyRoFv04Zbk8N6dYMn/L53WJoEmkaM45xeCGIe2b1BRibk76HscUsaYxSy4U
N9fSf8wPIZz3VQmnLlcp4WLSBxy/vwC4IKmOPex6izlZbDQKqhWjVpgTzjmYJrA6VKOObFOewhmX
RrfE2VmsRKuCOIYFAR12kuC2gDREIf0gzSzsbiGbfT5oi6QyE67pmtZJAvvkKtjNDFNiF7gREc4/
+pRbx2bTzSa71P2XjgIdljmTh4nPhhEf8DpL+AMpC7Vvzk5PEpIBYcyssHvKrgBskTUgejOZXaFL
qpyyxLkthJF0mEzRGBq0UWE+C8U1mJ3JbUVkptGMhanPxoLq5zqZdW5tF+uKZgsZlnJNpp0IcNg8
zpDNDv9Q0w4+PKp2/50G5X2sSxGWZ6HwjvGGZ95dQ1xqXMSQxw/ypB+xxtVXY5e+BB09PcKUR7r0
bs02oXZ2Du7dJ/kwHI49TDkmviIbItGnamR4yvWQ9O408fcB+x7apwOUgIJXipacjXm0cHYmbSV7
YyAAMsbJmqM8kVs68VUro6cj4QdaR8TmrG2utLq8Y9GN8DDFPZpFxK/0NcGePQNQa4quQ3GkQ+vk
hw873HdyeWMHnHOB7hwRKCzkokgfJIPDdM+Vx8TIhZmlhxlmTf1/mEdLOXyHPHsVIlrm+pv7gImg
hHiMYXBLvQ7xxhJ5uJaYIgP971AZc7RfY4ELhQepTF6lV9hQfcnjmVoPF9DsJy7YvJOQLcGRlfGr
Xng3sdrcRfI0kRFmMty0axnqX9i+SidPVrzqPEkrIQsSiuLp+hWrFF6olq3zmUPUotfDJDN5AG67
qh15ZyNUkAACja6WnrwCXeSmFYrbvnK3uMNKnS024OOh8pLbTsxwQbIS57m2b3WrPUOi1iH4rkYV
MIzOJp6ZTkoi1IV7wAPxb1znp8r6DyF/qbnrV2kNpYeH+tl4UH+PYCUzy2SPQeRPBSV00s/pW8aB
xhuit3ST+yUw0O+SlRcO4s+z8fzzqI3B5So5UfjIMQK6nncz+wQ/6RGm8X/2CZmRRUKf7bgrMtFz
9axpqY2UXXU5rYjvrR/Kep0obBTBvooQIlafW0uDsuz/iqWiPABd9MY/CqHO0oeZOVpduEh2IS8y
EQDBZEz3XdzQZqexx7EJHhPd5+muCAg55qvgCEtLleEI1cx8i1VRcxDtQ9cuM+or4cDy950SB/wX
dVwC1NTQSx0+B88VBS2rH10xoU1+zzV+jLEzze+EwRqMBUkIT7S9WbHRgeqPKMjqbqamLXwDMM4C
O6n7O3S4MR69IPm9tlgDVlGjSSEoNaadfjmx44+qPvtraiQIBg5/rCMkfWU+EYZ6nn5RnZUWH98/
9uuEvspGA2BZMMSxC4y9ei2IkM9eSY88VdUBl6mPUcoJTsosEyZAfzAcuI1mvIarrB3BoHktGowt
qxTlp6PQEkjUvCSuewfgvl0q2i05eLj0OZfL3DVYIrNNw9TmNwmf7AwGgwKnncmskuyulo4gUzzy
dxhz29hU0vr0CdK1B7xYj+xJwfvAkZ8KSwo83ZobzTGNuNtuGabg4uSxj16J6HF2gJOMT7JA12K/
cTSvB/Ko6n5B2lj/haKDCTZ/bS+eUEPh1Cw2Mm8IodDzmXN9oA5QHKE36mmzT9mAvlrEHHYzXfKX
SFSNWu0XGcn8aWa0RLSnRXft8Be9dpvZi4QsccIRKT98aQ/a5l11a801KTB1FdOBTeraTAHe3XAp
fif2/V4WPnaRU8vws51pezjlqdFEkxkulk8ZNW5K3nOXH2nng01HxCJ/j9hxyiNp8a827zNC1cEU
XWHucxODPGkhl93v9BznVZtEpqiKeH6mbfn7koOUfY+n+vRyy/iOgYSNC5G4ZlHLmzKg+BzJ7KS+
Ph8Hu5MZELHM3O+zlvablTDp4mcCvfSL6MhAYWzLM7GtD7xWng0fbnZ+h36jdsCkpHRhQAjqvbcr
uBT6spDun4n+3Toa/rcXPL24JO0ZGJM/V6ZG/zx2SAZw4lkRN4wBSkANrMjmBflfa2VFPX04fBsq
ikAlOyXHksIkHTihqBQ/mf5sKJldrB8qRxy0xm6/dVdJI9fK6KLi+HycxTwyA6gpTlcPJ9At8aWp
i0NiJ96pfM3tHnxv5CRLpbx3AifSXL5i62svX2X8WHenLciP/J5pWB1cV8iZisofuAhAuHDaOiw4
6Joc94RI85pOCZHTqHcLOyPIENHvteD44bpWuJs6xIIkw5AB7+A91hctt5ckSthdEc/ajKyPWI/6
FQBqReAkTz4pyN1mlTwQIvHloYIb4kTxIUjLh9H7JWKhhrDVSNFaJmFB0Gk57wjkplZbw80yQkfO
qlffT61fHhBP2q2MaCBwmhnF3430ncDvC2GByprEiP8IAMAejK8VXqhtodGkQQy2trqMGi3QFn5j
2pirXd+NzuxO2AUmd0hR9+/eR8KuR5BgoGmi+jH6sZplamxNISsJ5plBhwHQC/MnKicyZkFdIIz8
byn1Z9GT06V87tLczgqLOkz+ZJWyDexLUGeAmRRDbdccqUiixsUkOpFrZxQlmmUrqro4Y6hYnr1S
tu1dbo5tgx5+jwZHtpGNo0UOylTKqI1FKO9m8DH4CE3iOb3RlwPLs4oiDewgII0sf5eWKd5uUZht
iWKThn55UeIIF+Sob6Y83Y7ZRMcdz6quJtDGYcDZQva8sZTGbVlL+ZUyPiQErBoI6j6pxSCWF1xL
RXH9mtlvJvu3azKS8dk0jKzhKk6d0hyQfRglkrFBbnrxP9zySAYSilrPOw61pKyTHPKt1UYThe6k
waq1wBe0z2JOqev2NB76WgP5+3ndoICNL45APt7FRHXjRus1bnlZ8X+MswpA8WCWidrcuq/plcY8
oex7bwlPdWMgTy4m3DKpsTWW5+AYfpUDSZ//4zcHB/ZAbGjSjhiv01aYy4lnANj+CfRQl3cpemLc
nKnb7RL+ge5PPQ+5h3tbei7iLGFnxbmkrdjJnVeCDgBl1DGpbJat880Yrbjl6bbg1sYrW7OpSv8Z
+i7ZzarTa5WINk2tC36IAQw/iLj9U0MO9MxDBErzsR3mrBzZ6sOf43LHgaUN57c+FamwFLx6SuTU
mbN5MUyy8bfmlhD3CudzHE8Pu2S05i8NBWCzgzmPBKzUHf8HM1efcX6n6yFwHCbYNxeO4oIRh3dp
+fFq/f9ED0yyebNtcWAtbdIqE0sD+udsjYhmNJ2v0UniU3Oz1TVX0wbCgOsbTGflumzaRtwJNKKs
cr/MojttKIauKIIglNCZ9RTRZo+vstqg08zxHl6NqJW0ux8FqDZ8Xw1oOMtm/7b2xFvI5/t0H8DP
4cPtvy/U3KzsNMX//fZs0n1g5Wypp+lGDilbdXAazNWf1BvRUmjPyrdOnFgaMLc0jIYE98DpuL/0
Rp8+rnQ08oidKcX0ZH3iBwD1UNZDCcvQdlzklhHVeyIXZkDS1JnlZAF/Ozft9t3+0g++gwtTZmlw
TnTht/wrJkzVkBMDPPc9vO7CdoirBaB0BF7459sknjXlrGZydCPwAf5FpXGjCTf+750fcEelfT8Q
ajYxLJXPC+wR2xc9LlW7ZmisNeRqxcWm8yee2u8WUUF2YV7Y9FH8Urc8KbHaj+yjb8ZWc0RBAefG
epTZu447L8BWd3/OGQPRSoPS0OOnWfy0CbfAxQGGwQumB9ffzjMmU5EsKJ/b2Sse+8NZXY0VDIOd
fUHnWB5EBmoJWvafz4s+N+CicA8k6VfUvOEIZ1oeZCgvYpHO2utuwyHNawGQMwpXMHs3F2K/4OhU
AHu/D6kCikY+Rzo4i9ufjiGyMvVMgs7klAWpXWCcVUBOkFJBVEEhrLwWJNN/7sss34C52h+GP2wB
E+aEHwv5Z+u5ehAgGZVzAKBksfvIYQJtesgUZq8KCKUu0fKpSTzCvbPJjeVHUoC35NF933heyCDX
FNhL9KsnaKSWMF/0RUNiSbqqnV/2xX3/HmBAct88iF0x4AWc0UImGMjM0q48VMuzgksAvapD/GIw
uzzc40/DR9TNQqb5Uan8RwZ4cnjIq8yYvtb8rJFDEm2shBu7Ft/ARJ405Yd4NpbcxhfpHAqZu1q9
RxfOSPta7xI6kcF8d0wsT/TNjvSatqCTGg1l9oMq1UF6sAhycc7cRVFZ+voNeBiuhClRp0co1mwI
MNyq/idZfOwxcdmQt3zAzNvyuzCVL98BoPPiUpnCULkVI50M70mH20G6W2Bm/SwkzH+ezWZWxjvk
416FwekS8OvR+nGhl+c5ujIOEgSDb609NdMLUKd/6te5drMXZmx2xFIzNUfz3ZKDzRGim/Rnx3l9
k/BMHw0nTDKtYRXu4Nk2H7wPm9Z7wiM+vUmcERcRoX2mN+aB8wxRH9xw3RbgGNoBNpgXAR0Af27s
Q5BZGH97Y5U+Ucaqe5FJkAIBF1y2/USgD8NhXc2OD8DsTvhSh6brmQJJJf405YBPrwtYBVCvK++M
MosW8d//bbsxJb9yLffPzneLVuig82KNJaqTAGBy7qhAasIno/gR9gNW1/R+JPY3tinUBnyGAe7j
nbeitkV8Hfn6cYkKIC6lpGM2zbn0McynpEhDmg5H12rNGdXCigg8qL0kYnhDPho5f/yzo6ELDD41
qa+9gyIRoiuZhiQU7uQR3MMWE5oZGMmJy1Jn96gzMU2d4S2P/WQgUkTfrwmuvFFLPwhseq6ORKuQ
KaTx97Y/+CloM6CAzS1oV12/4IJIGOj7pzzwQDlEYyEVa3xmMJzTv6wkR1KYJMz/04rwb1Bqif+0
1qJvBxt7z/SYOsbQ7eVw8RwMG8BbDJw/yhsv+dTWW1PAx749W0oNh0/B4MU/Zs6zqKVFATjsrvtw
wmW42BDyyMlQBY/zZ7xYnJPaAKmXktEHCquxn9IMF/HQUVWMBSwnn6Cql1n6WyGoo9qrRfM6oI90
0+kZwPQXaaWT8ZcwrYzxLKThpVxnFm2DLi5/Y61Yf+iF+oMcRqbdwLmSFhR+xHjND2s8hYU+D7Ns
ny8MpKmWduINfpSv3tYOxtf3cVrAnuelF9eXjG72N34eDuVdfgxrlcJZLHXUvdx8eNQt4fuRM8Po
IQc6AaMNyX/XbryST/F7jACe5lSdzMiQKUknq83EGmuCyGPbqH9iaTXh8Qxh1OERaAz+o5ttRe6A
KoltQJ7KoqiWqz2+/fYJxYyUZM3SVo9hNN33zsIS55l9zbiq8X0DMNYpn84rN14K/qxtCanxtdeB
VuPIFhfLSvedxVyKz1kzCtCW36xYNFaFB3OJgAQ/VHKe5D+fiHMG1GZobAC8zF1RW3TLQt6rVbxl
4GKUnSbHPAAcRsgKHgMpix/P3r8m4lRRRHeHDjmBstpJ33DsjYNgMH/C6ymrX5kSjZhcczRzyRLh
oKt9IteKh+dOx2MBaStjq1aS3rMGeIrImuIrzHHgTVJSkbVqW7xZSiOSPRyyX/7WsZD9s2VLv5xK
uelMxwB46ZZfucNGQ9q8xGYLJYDMsuXGBRWPbRBs0JOX910BT4TMPMBHKwHT/pwrlkK4JbUm+tP7
f69sRJOg10bBvdhkfK37nOQ6O0UJtPE1a2M8xNj4cNUqAWBIIXCHB1HGc6oCRWlvkn7OHYrA0VUo
BztHqtQeGMBCocSQsfkX2/8Sw3MzsCZo6PDpmi4dxYltY6JHGXjtwVvzkS+n34d47chMYeLgkTTu
VKShg271AmKwSX+5HPb6d9gR8h8Boa9OvvMNFCPg38aiLpjlV0AM3Rq9or0wu10WqHfc589f1GzN
dA+wn4qA61x0auZ/o6P9GBc+0fmjkWKZqDjIjVA8RdaH1/bdK6zxyAJsyVCleeSfnw1mQmT8JUqU
xU/0p42IXkZ1X1k/2OWl5pCAnA1ox/VwlhcL2DjsZaqvFj1Kj+DB9EhOMQgrFWklCVQx29zKMPT/
V0Ri/FruYcK5UcfmPvPNl+ZWLvMiat4DpRfRC+o0eS2pSToxFctl9pz8bzEt1khXgth/YHuTfaFC
jBYbeqUyNEaiLy8+ndCq/xKPrd9zDxPYHFfVCIwrxKhhQusQCZx3YMig27qH07h5W7HXkzuRqFKn
0bbMIAvbXFPQlHvG33HCKtiU9XOdmHcPJDOAYCJrFf782kRro+NZ3/fVEHj4axq7c7ntQNOlJFup
iCUoOASK0bhafF2Vh4WqeY5X3PIkMM0KHbPm0qRUGItEiuwQx/3pN857n4b5Vd6w8AQ/npgwQP9M
pYhAEDzaJI+ZizfZlJYvJLetKDoKcj6kxCuob6Qw42OO+f4V4hZcNCjE3TwuFiHjM5zED3GOD2MP
C51y6d7KLd0uUAMptlDYf2zAMjCq2mHrWiC/AZyEJsWU38GqFu3vVko1wqpUTobQvNdbG5+OD8M3
l+tTshAZ8WEHQnyJedZ+7gR1bFeo2vnwu/NAz2JXc4adTg95VH82lxQTwF83RqI8l1CY/Jv+/yBx
CWRF0CoeuNl59WJiX1w+FuEb3ln3FYDkK+RNj2hUkzX6dzb1gXoNyRvQt7svj9ql9Jxs5nbUDUHQ
/p6ZDMnfblumw1pmuc9yKXyr294JrOsO92xEtGAqUcv2Jm2EuK9L1NVl108CPl7y9YL3z/APCWXG
8u6zZtBGHUTh9o7YGUW5/T3byy3yOhiOd+ZJ8lSX9wbEFDEOlm2teXSZAxHT0v4cfSM8dCvXCqKk
HVfQWVmO9QT3rsdwdOZB3U8giDT+iGfZT/RMntPk6ufT87on1u41zVcFJ+ifLC2IrlA3yf4e86Cy
jZs38BTqF6+k618fSsMWw41nRaEnvrTWpjp5Drecvy/qWDq+35ZjxMoAsRin/te+LtUKNfWo7qQo
hugdAien7+Aq/b30q+mNBuh8uiXcO7wJnovTg7eeLtxwRP3XeM/lTrPWzFCxNwUhU14d56cnIDg6
dBHffFvq9DqXrb+RGRJHcwu2I3rLIueBg9vpDN3K7DsstU91XgOX75LrkVRBLlbMHrKfxB+mPrG4
Y+OuRI2sJT+zn73GhN5gPSOwzbonhAc8YNzbJmjYbMPm/c5TR6N64pN2JskrBZwBTPgNxd5+qRPP
xS5N+qK3ppUOY1dfcSeHXmS7RtcsKNusZ0sAUIq7D5NV1wMjZH3pBleFdOzfXmlfdSiJHiXsAn8y
a82V6+MLul7yw6/fGXT0PY4x6qfDiAOLPiL0JvC+2ICP3Jl0qeVVbBTsZvJacv31cuNiDnc2RSlW
/vdFvySHSr+i2Q5bQJnRphKRCmgUoyUayhrvgnDixdld8eIsaeG0xYL5AwgkOreE6ZgcHoj9xw0K
YiMabeWr5nP+a/mdMmzt/ioiC3Auq4Pdmdtn6hFrq0zSFhvPSgmx4xYFfsZ72mdOA0lRX+Z7pztV
9h1LyOpSqX9BhVsaT0Xqb/kjinFQi2m/I0HGIyyMoGlwyT4U0AqKYsi4yfyqoEXYmJRCQRjqmySd
8MD/1Ojksu+XwC0KMzzgwfK3vPbySjLxRQyYIqWBBcvKgRreuvAY+Qm22eopTRYNlHHZZGo6M1IH
AHhBgTo7U6L4fjC0ajvRTwV8Rp9DOgZ/d8bskBYWoH0Ebw8/mlknBSuzRpYiAqegAOwHeYwhOHin
pdkII1jeXJkxiV3x9JId2Gq0l5QRAxFUos+V23XAFnA6e051HoL2+ICPDYf147r79bdjoZA04vmz
lx9hozKCgHY2L2X0DYzfGdjWsUY7RmMJ59K2ZkqqjqUWuwCR1wRkuwqU8tTXZkFMPb+v8+G9HaE3
SKujsCE0AIzOR+oS/LvusTszui8tD0tlWGnZPdKJohpPEkj6HL2Rr5BtDrBDRdOT4qDJSsn6px9D
nPJAT+QGn836VNWeZtsPNnAlh1Qq/Qscip+5EUQIgQ+NXVxtlB5jvlSf48S2vSOl8NFPNnlZERnG
NF+bsV+7mlG/EDwFgs5z604e5ZVL30G0A+AgV9XAkI/+pl6WUtQD18WOdoTivE9JCsAiDveoEq+a
+ZnHiDsNKWMnke1JeZBZV+Q6zAZf+2sjwIrpwUqaBkBPO2zP2A9qPjLGzwEcEBxq3IiJz4Fcljpo
ZDDvpn4ucMihvQUYaT7Kr0EG0ZG0CLEMi4wnnKBxXswk8H9QjlnnxT8GA36UhE1XH9/cNzIxtKW2
whyPjfwlA2q8rhINOVvIsdUHVhgFW7X0ySDPi3pGMApHKotI4NjOfSs+D4rvd4MobdUtCDyiRxjv
Y9GeiBIQR50q9ePJ66F5meKf3kayxEfau2dI1Os82MSXDWPhtRE8dvYPmCXRRVwKN51jhOkl9tbz
hwErdrLayLtAQQGLiJYEAssF+CzUaJ5FU2qLTTBEQltjrMqVjV+FDLTdFXGmgn3DoEuHZ8vxAH6C
zgNc7FzKCX4lnFUIS1VMisnSsPSuvj1AIdER84bqAlhMvLDQb7Sw4gvrx5Ve0TMtJW/UK+WBZRA2
X2r2eVMXoIOvbBc6PTCPO5ajgpDFSgMJQFJwAnAk7ZO3gYZ/xvpICRgoGMScxJ14HN1rH4tJU1gO
/pOXeppHK887QHKYi2EOANxwPKJYQSECn0XVq0dhiJbnE4sLSTaHuSuYxtWyR3xwtRH3NnDHck7W
tmQDumjOf9RLYKkR+kOqYEwBIF+xEl5+rObpDML0YA4ydVovkekQ/3156r8PcCZXsC9apvI2HCNh
GeEeh5F18Ol4H4B3UObjOu3olLSkhA1jG6ficMLQ4da1fPeI/i/kF7NAfqLF3nVuaBOgkUsEWvjC
e1IUfaEUnbjsP05eROXfFNVYcs62/Bv8JkDEq/ljSD/Uj/tPE/F0aYf6WdToZhSQzxLeZ6LzJ+zJ
YRm40nBfWFupJE+kU2U1kIlaQQ8IqF5hAvRmLuyUIioLhkDAgzFdknTGX5GctdIUb5IxQ5YUJcV/
5SqeZr2CsAL7p8VtUTj1vze/OCYOpW1gzAI04Z6WvJNDRVYzoAkHAAV/rMBMQuoiioDIgOQYV2St
UWcn7tFySQvQIcQZEa3JdJCMtMBRSzkXAyrxymZkcqdMfz0XkkE+khp856Ilws4lFZUBfF7p5vNT
I1q3aVqfiWUHwtPw0wk1GKBBiSH7T9omPw/7czhmJ70NfZgXjzzg28NFi9L8SVunhLQt70Q/jM3q
XWY68/cbsGXLOPzaQS4Vw/SlmVD4upLGw5EKbGuPooGwCNs8nzL/fv9HsVjACmRU6dXvjI3/v7fP
99ydxzvhIxy74qQ3yehzsatGCCeecDKwqM4jytcSYRptz5j0Y4cX6+d9DkmS2bUol7Lio1W/KYDS
ci3YEbZojNcKVvi+n4AikQmiyt+fThjhx7Dm0HREm7EeBizqEPx5Z/hKP/TUu6y3+4dqNFvPP1co
k9lQ/ADPumpNfYKnS0YSurZjmYUBJFCOxQkQEWSnccC6ZuHc2Ub9vjRO+tbxftLctSwJRHyJ1osE
WbA3+l1NOdDGU75j8EMb7ii5JA3fqpXRTELcOcoucJmBn2l5kNzAwzrlxUnRiTgDj2kcDyCLFYeB
XClFBGqUce2cH+vZJevN4DEy9cJonoNoj8NGEMymD00KMcWyUEJrgUetDIyKr3cO79+on/t17wqd
RroiHGA93Q==
`protect end_protected
