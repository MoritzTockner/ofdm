-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
l8yhtKFCHHX4d+aAl8XvjXK/pt6/FlBNYTOdXLYzQrwpL0c5Sld7V/7v4G9OFM5+Kq1CXKRiq4mA
YY7ukyXhosqLUqYM1L/aKRxsGoddB8n3QTcPdvlMFsv5UuIBQsGcVcmXAHoLengs0/8sxlTVf9rR
pSkys+WiNZ9CLYS8X8F+oq4n9sdU+6eKLDd6FgbJUm3bBmvf8hXfSXFe+m4ZtRj7Wozn9rG5rmUM
YD6Atji8d67tB1y0tau5AyLojChItxTkWRmmwTOHuOAyWXd2qIvFBz7BSkFHn8QFPU4FsNkpLluH
Qi7Sxv21VadIsayq3JaYR54Ik6ttnAaGiAXoPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
Yjv7Xe0EJBZnXVRuuF+xVsyiTy90Q3MPstJMHp0hcSnGuERCVdoEztUJ/G7Dpu4QffgNxP9dgbA9
tPR5sARCcAwgahYImHZk82dv29mzfJsyX1sLq/mIHJG4iQSRqLXLyLjGa1N06zwpW2r3g3D4eZ3U
zZr4f8WxdIKJj5QdNREWlo8GQyr0BxFLA4IGkhAupgKwn28xdnx6et0yYl5l8Y71a8Bc5MNP9GEY
f/f3tyCq9sKz4DFqh+qta1OZjl0sv3eThSXiQmwrob5KSr0BFZtFlHUdvsDI9Wx+ljw7qq6zWLqc
sdELGtLfNhJffEYpzT0JZ7hSXLZML0yC2IIWuQ5XIKcPqKQMr5oZDWJIV2cnG9eMZoLafR2/M1Yk
6++NQ0E7TC7xSB6qU19IK0RZimpgy7o2e56rxxrqvuyEQekGCviY7wMTkgyo4Ddjawz0UBHd1nmp
hXJIDik2zjjzverzzN1csniT9steGt/SLQ5RKNnW1738Fm9EUS9XLsN5kgx20DSGW2sN4u+tuFOb
FPKMNCbd5UwbsOHgQlj4aP3uDGfxzENy6y7Jz6b8OKOBixXOWCXD9wFFu/6RxE67FQd37fUAGYjg
VGLHrd9gSPnixLvWEKJTAuSalFPPm0XXMKPg1WeonK1jMXCAPlf4TElZAA7XGGptepRnmAEjKAKZ
sDKc8IA8ZGAt59GeRxMGXUUCEUl+n4Skj0kT85s1rlovTDpx2DJRAlMw800V8flR10ERxUFYvkRp
N6X5kp6hKve7gFUMb6Kov1Y2yJjZFmcBzmk62HYI9VcvdHhUlX97pXz/UQyiRpOLzJsZpdksM5nT
cIPvyw3miBZojYqOBRPevhuiNqnFRRCCLfBa980NYpAygdfLsPhZztib0eQj5ymxfyjHXTEROu3A
FcIfux5G68QqzmxYrtD06Jz/EZY0gfCjxCacONOrM8f5gSqXPUHsqxu9EKBDlywSY1a/eLLIx/3q
w96/KerZgQWOi3Zl5bJldaS/9rQpyjIIHqoos0OZPBYf57PiUGPakn6LjKHoZgiQJw+6JKjJ0bI0
YzM/wf36F5/P+mhIgEq3D+cq6JDVQ9542y+ZyFetB2yGOld42bqikEwFrFuxA0vJ8uEpgoO2EDEk
8HG85UBw6V5KSQPQ03fqSnTTQSoJ2UXMAmly4TyUhJGhC0yhYLtZsYTbuAjmBTKWQq2jr1AeKZwD
n9L76gU5BDz6ZTLoCBo9iHAwb8zHKGtE6kZqmALpjCu/GNuDNHQhRItgEHzAS0jS4IXINhJSvd67
lIT4yKtq1mPlOvDHDDH2dmHcM4Spnx7KqW+X4EE/ZqOmNSiVAswsk08gSxhwiPV7Dt15k748cwEJ
3qbvA35IjDidVAHJy/p2N7LVH73LhSiAvi2x9lrDgSFSzfq93dJ/rIepq8y7B1yX+FtynJTojoFH
fLWIpQ2plUyZYFNlLc67LVEeFvPc310fJq+xURvL6jTx5P0fekuIAwcBjUVKJK0PtbwatCYXj4qR
8V4hdZfxbgSjAkJMi38rmn24t2zNfVTO3eDKYK4G27i0zDVseWYmuqln/8M7ZVYSgIuQkCvq9H4H
49cPUcPBLTxfiR720aHuv7T8FcYiEowIY8Q6O4iQAPxTVCQscXXN9wi19OluDC0mzZzY+/bS7QV5
ekr2fNZ6SqH4EiKUKZkylX85mZU0SDB5qwzEEWWOYsuLjxc58dj3D17wUuGDhstq8UM9fL2sGDs4
Y8W1G0RU81vsORzgZ+p501/UbCgcKSXIBFuJMpKV4YYxfjh3JD3tzC12nu6l/MvalDkkPkMMtNvS
w0F+oBl4dHY0MX3eq4ZHrpZbSQ+O31UobGLQFcFm3Nl0QiHQ8dQ+OdbtX9nSEeMh8pvNJ+28DvRj
EEgBDW7O4IZzgnj2jptXUpiKFyZgjfjeEMMT+32xQMUWApHQJ3svL9ArQzHj7NrGUHY8VMHDczY7
vhqDyAvDbABRHGZG9m4ukWO7jBzrtZ24cxj1OSlWAc5cEUtopZn6saI/v8ubfbLHwfgkntoqyuwz
m+NYqVRKpBSmOlq1k1FwH0vSl/KuT+Flka54wDQ2BTBSRqquywv7INFsvaAdoFE5NWEYRmcY4GuB
olIHFNV0pcUY5rZHrkG7R8e3obZNccK6kZV0cyE7y0AmmlCckh440k+DRQOjK7nQpMwX7CfuCSX9
OLj5AfaDzweVufZ94fBFZxYfOzXaRnfdePoG00BaMRGYPZQBAfRKl4Wz+cjTgZ03UnxSpBhJUz61
hir9z59BNLSY/AqU++C3au7LsycUkIwUvijTu71QiDwvsqUWViLVZpURZtbwTi9hwLfcPyNY8HHr
I7qDbgqL84a35b8Uq1uJ78LrDW2UytW75pTSBi8vZAZKUA8Kzs/6Gmns/vQE97YupvoCR2ZqrKQA
Op9N864lKaRMkaFrl/blpGWRWVmac6F5ZgOefNHTeBb6F2C9By3kfBoL+eE/Gj5OofJ4AUQEhIVw
mH11mc/QKug/BPy6bslh4C+LaAVge0kUiCA9Hfg0EyeAny+5WSjhTTrQXPpDT3bFlH8ryIREQZE/
LZMVHH/rSEBPSK/329cv40lWaS8UW+qVgI0+15f/MXxvA+LEq3HgBiNC9MpyqUgZzu72sX4tTm7p
cFuyxvWjTWF191ZNdCkDhfYX1VgfmQYL06wD8/yWQ3eJM7tpOo9OcwleSjO4RGqqH4A1NvYH4Lv7
ZhFuEh4hJibE2ib1hoXVTcVRKgUJM9lf6KEohX98wOPY20p5g0iVHRLygXSzfw23uuPeLktDcrRO
/BrVQLSFzBp1suWQevQrzCOuhPCUdBrsK0UQyJ/x27qPQX2MX/ZXxGvKAYxuP7Ef/SepGUqkSuto
z+SCruw8IshNJYNVSBlEnwvuB5OqifwkPPBS+Nirg9O/KLJ1CmIKSwuTs9/ZIAnVPFS2dtpojOoB
43b4ijfr5oK9Ka92sQPPxFGng+ZiqOKfYZPhOE7ijsb6qLmsFQm1XXKmkiQWRulxSq0A8/8Rp8t+
nXXYDNz94uCUp7j2OW5p3O0iAJiC3SrifTRf7ojH21xpG/q3sFnoBTO8jpLxO0uRyG/VPuW0pVIN
6xgaJBIJd7I+pgIZ2Uk9g37GIn2zgHnBkULS0C0qsWrtBXJ/GwLBttkBaViYf5XSIOO3qhxdg2EU
G9rZZ/HVPsh2vC+1pOrb8mWFZ2XH4CpIzq6FAWyOV1mDS6aIz1HL7hFIV2WW2YzCWq1lazqsUs46
SzxfLUnCPKXdxSkh6RuQsxmsDf1WKGj668LAeHU91hAoA7aMvseQUnFVWTuATJ/OGq9sP7EDH3Qf
8Vsfbkad4jaE8/hI58bfQvOs+Cepmnd3hEj/C+HlX29dV3UMCnaOxVV6qlZ7xYj/0OLP+2ws6tzC
L3KHashv7pFdVvdUhYyn0J+xFCYy7QWC0RftdEqLhMcf1ZsrLU/NWm/As59xZe5om/Oi/AtmdoQd
yIMXwLkY+psgnGO9L/ABtrqNJjy0uZ/7NmxWad9Y+7SBwRqHNaxHLYl9zoKhncpxan7GXdyrrE7w
onveyhis4ZeuJ3quWUOndEMjf3kvemMuiplu5uN6EM5dKxpkgUqdpqDL36qn02ASaGfeQruQ19HD
I9YXoI+d227t4qhkpnZuGfIOkMGfk2//n1xFn0zrJXiBLqcP00t3MUV4SkkGPW/5/NraJfoebDAI
5Pg8RFTmhbPsQ6JkwgCB2GbGdZct2MR5rXHh8WelxqekeA3f4qCM2Xdzm678oIOTLxy/npBGbhu5
9q5ECpVuAT368CnO0Uqd1IxQwBzt6+X4IN3MWsll3FEZioTsSgrHOKWAPkbg5o3dsE7o5VtuRabs
Sihq41BsmtrZOfc1te/Mj9LDtNFIBDIzorMvU5QyVQ2ujzkh+z28QHBu49mrpz1SInVZShZ0B1g0
Sg9H2/Zi65mHea3youYbhRNK0HC1BjUeL6LnROoLWLsHhuRbq1REesJQzDRsGPwxlyRtAV0FG+il
oqhW9aWxxglYtfyAF6utUjoZgTDBfjD9lQqkI+pC4VfPkp0Rc/MKUs5vgBvMAejRAnWPdc9K/yJA
iUp6LaFchfxlEjHS0LsHjOTFf+J5ErFXKVhh4odC1zpJoHaLv67VIuXINITaToiF1gYETMhI8/Xh
IAhZAOBFG/eWIhved+OE+1DbNCMLyD5nbgiQNOnPBTXpqj6sdGpxyTd+8qi3DWl7X1HOUXNmT5zl
Njv4jQ7dFDaQv6OMJC1ONtb7ddOPEAJwee1RDVGzwjLW4F1CGlXhfj0s8i0VD/USeQ8AsrktruUi
r4YVnv3Jnyn3+F8mQ6fgneQGY/FuBZWQqr/zY0hdWLHsB0IfgmEpBvrie8w/mfWiXSU/eyuAEYPh
Z7opFmG7oP1slWrNfef3Wvd+3abtN3ouGUkNJSis+ZJ8/96SphW7cdIC0uQqZCDSZ8bml3WdZhoL
wW6i6MbpuhfS00Zw53pniythO4pI9WBp1+hnwlyperDE+U+aWLldxPyQ+EpAApcyfAnuHXPkTGzy
6tZ1EIlt3nQGeiVh5JlBOHduin0GgCNBg3i20SeQQmHIX9lYTtpc0niJD7rk7MnDVHV4vgKPnefM
6ngUyXyfopba+aymHLMsTIAtYiVaCtuQfeeI/I5tF4M6eAJHA6GVPMYscY4ysyhpP2hKkKXoCOzR
bVVWxsXf+kEeUpjWPTlTLqH5q73o4Y2bIgf9p1PHmVZRId32laXvX5G5Z1jl62DXhO3/4OmkyuRL
Z++IT/pXeXg39No5NBKYY2jRYbkDc2i6DyXCp7LZ+cT8IVHI0qvKBmGtuM5KcH6x/yCrNpg5ynas
ZoB3WmVmc4N6SAO/3W7gcyWh3X4sNYkkWgePt2Ker3KssvCvOPkLvc8GnMMfB30N+AlG6y7vS2YA
nL3IijC4MC/wp2Ed/F45L7v3Nfpk27b14Oz25M7SQ2sSYxYxIeIKPuW8PbWekD+r3B/TVUYCjiMC
WoUDQCgkNe4aPkXfr2Sppse7PLEAh3ecqt8UKchzsIWriSEKkhh+amV7+DmMxT3D00RQUt2kiRGj
GKo8rC0VBgbIAmgZea72UTWPZsMf6b1aiMKE4g0AV4Wx41cGk4KnYaYmrHDdt5kd2NvfjYAlunVl
M5fve9D+3XTaTHZ7z5lsuPUj5u2ePSau2IYTczsAp0kqdQokHuNXilbP4784JOeHB8bpkCbU+igz
S5zwfGqNtFEFvYGf7kwx8Z3QAdVpqOcRXqpDmkhOqhBVPRv7aJ9Txeo+/WALg0SDoBZt1UpY+E1f
KBjLmgYGwWk8UcUHTMURH4OFAhfFRTXXZK+N5aNlD0rmUqoEZa7mps+Noc2WA5mmix2ALXfh3sNz
vn4WWVyWE5FsI7GBMfXHGY1c81hP9lfX3ZQNxDlSFLTeYb63ben21ZvV6fSOSMwOH7ZvUE/IV0qa
wjpKRYFboo+WztmoQZD0k442woHCsr6e7UEIEkDbtVm0weZcxiXjJzn/NVfMyH7W+Q5RuKhhHNdO
YqGRwt4AuRSbuAECBWMhppIc1uhTp2nMG9lzcRniOzCH5z3v2XF7vZcVtFWFuhIvbO1B5zLrMi9I
tJ6T1qnFIDubDoMkR1eRpEy2nJfuOmg0/h4uvbDHT3Fl2l0d52eTBbgitKTOcm7npET4nqG7SkaC
m7gTM+uHqOnVYbW15H3WO88gbLuYkCYuPKXROyAIXz8S12Z82ITLqeyQOQIU1TELLKEUsznOG9MZ
r050O3kAXwnkhd/U6pRKqovxRXYb/8hyot14jaGS1n3JvfU0A0ascXgV2WYP8m0YOZyi5WgwsiFd
bDVmZJJk5IyBd28G8TfHdpG+RIEtZ7JMyf2XcWfJfClEaIGZhTp5ckTkSYIQYejlBHPJd/qSgU0p
iPfF6ol+k+qSoWT/Db/EApnD3Uqk1NGTPHLneV/lWCFKeXuG+gPi9o+jnKfNIXIYtr0E5IlO4D38
eirlwOr0G0YzLZHH5VV1rxt3KdAyIDklMFHlPfm/97v+Kf4w2Ek8l9Cq4aoFeR3l4R84FFFjAoMu
DLFVQG4VMdershy48Kmhk9IGuzTx33KpA8GVKE2FetDD+YWY7xF7E5kV73Z+NzkgpFswbHJm5Hju
g0szPjGrtC4fu8DyRAQjMQI2yAo+w/EDMkAoUdJvGip31fA5Znb5z2+dtqURhfzDMtkQ6wV1uDcc
jK4HD6vNp+0cEQphcavRD9Oh0zakyxZ10ropg/6jaFb7bGzqECVs7XX17YzFyq9Bmo0pPwT4Oeu2
FepCHaJzsY6dc3MGGoayCCkWQcDWkv2EQubmvvb79EEKNXWI9O7W/umPP8Eq7UBuvNYuHWdvglrH
+r0NcTCD6ZSqMbPCaDdRPcEFVJqyi4uw/a7xQVKSwLGZGyamDgDyU2OGtF+0/4bdyxZpJdhbjLlA
Xbn9Szv8IQrJ1GaHxgyBQETUJjMTwBpHlNDW83UmlBoN2an4pkdnKVe1QOPf7Nk7fcFyeHJsUPGn
zgRuMrHZTPulahSAs3bwwK61g4D76hXs58iVk2Xp7TrwYDcqdsMYZVi6GTEyv6p0tLCw7CDFyAsW
ED0u2vWKFnS3MWlXODdrzWbBiQ6Fi36U//5Etb9OyioNS/F8b55fU1Tce2aSFBr1hkwQ3K69AfpK
oILwG+ta42aO7z/4EPDR6cLNcrA6cD6cBAm/55XCKJawZKYDwXg3+tN4/CNaJ3llznHOdf+kAG19
dCKPu/qOgq6pzhH32bn/rmSE6ofiRcF5bKNxzK2YrHnFVaoeo0qP21BcpI2M97Yeozm2znpM/Cw9
HrJdu4lOXbUSOSGEvogy2i5LJuSAXZpvTDA4Zb8BDji4XTvqD9nNtpCRj1HYqcwRqkpEq5q4O9Vr
1kbLmT1IEIxH4mQQ079H9+xkKbs406Ju6JoCoTU1HPhFu++eiXmwppCr2lcf7v0VD+Bkp9x8uBxP
iop5hoZlWeLG3yLZCjAFzR9qQwbeXwGWmNdAYH5Adkh0gTxLApB5eGDHlOG+xZhEnd0ZRnSI+NFx
9idzkX8Eo5kablTBOKXyjVLVsC5SaPkucKnRdO7qs9BVeSEPQ/ma15t8xy0a8cIuEzXnITDI/ZFR
I/OjTwlSKLtb2kR2g6GTr7ZSmIN8BZl+hV8wDIWFrsh75G1ke0K/CShMgmMwV+0WDmNyEVUdsIHq
YSK2VCvfwmk1uneu8dFutwJvqfAO4R9WbPMs6IZKjIZ/94WRzkKeI/Il+ZArpLLEFhyMmEiKXE1Z
OlZb0jUBcKeR96XgNlRiJNnCn9p4fe7PM01CG+wQhSElbGCEssU5tawUGd7bO1EZZRccb7OJO37Q
ING8dAX9mkfCk1qgJR4tCDqrcy4Df8BMtqDcNZ90XGr1BJu3ARDsAvyHVNdv6OKDfWek7VBVjfjV
22ESt9MtGX85H5VA3lIXOTxRE2jlyMfcZ3jObvstaTPv7ef4wfzSMn0C6cEIQQp9//IOGGYijKuO
smr1QjoJaSJ9WL/bTR+2SuU4s+q5LLjJAxsv+ao+rPhs2y/F2C9gbN1f5rUJC0MCVeCnctIemvqR
RlUTKkTrnAy/uMbdCTcJivDF702+bf5KRxpXba/SSnKqHS8c6qHoO57oKhZh2bwWuaAv2WUgakGm
ihUniO4v+Owke9ZPPlLS8vUUX7So/zJ25Km3b9LTKjo50qYtklYy0Njof9MpC1wn7i1DOWmp9Nq1
Zt7S4SxX5SBohYiYebUgqUYaW8tF+fg00jcA6+Ryhl7mZKmq7kY2XPhgL389CqlVc+aIEopZOspr
27hGk/xFC36tgsf8nMCLTRY7BvElYs3ifc2fG5qC7hkj64dVR+Nc1tDSC5HhPpoYaYGOnHRmVaa4
nVd2+KY7MKU85unqCe30c6xH3HzQQR0i4xwJ4T3zdKDG8XYQk3pdgb4shj9F/qiLBUs8sleanXdA
BSzruqJ/DvHOBnn7dBJKHYg05Q8cyN6OeE0tjmS5FykgwMi4qP4ZoauNyxHVKpqcPiwIZ86I0vsY
1CH7Nt/8qbo9C8UVoxOxjRWdjlcBtKcySytzNaB6Jvozz8nR5PeilNuaTW5YB+i4P2IP3E7ZjcWm
CUMtsaO6o4xI+5VubPZt9t48yGP0uxuLcsEEqEDqNeVe+DsWXIxL+9ETJ8n2c95BZG6x4y2qX193
VQ+OiVG+oxztchyl/VAos2fbflV4q6c2wqkUSO5NcD4bjERl312PMJqyiBDL5mP0sh843bjv070u
0OuRZYqubO3H3MZxl6W4pa1QIFAgdKIHXA8U/pC8A5RpQY5HC86y9U+56oMplnFE9pVFcHEE322U
tIAIJxDjtxNltmQZp+L7PDx4f81CLb5+i/PxWjcBz0WDAShB7dI7AGgeh6XPCDvtqi04ZYSDNk6T
p6oyCwJNI/GZiGKuq7jFyqMZ/GsXBY6wddq9fz2wmAeZptYwEIJaBBkC77uVzGSDXiEn5JL7hvy2
Od3A78qIbsciJRXjSy2ksf/kMxchXEeNFgtyoqarRc5+0KF6S/Y5Byph6iAsOTqC7w8Dddc5tNA6
BhPqgserO3zO0aNYEuVWNJgQutGUQW0HemGSVWph4x8h5+giXQg+TkPJbQgVsbyU5HZxF1Ag43tA
QICqzXlXz5QkZLos+oLoXXpml56Swkj/QKyCxOjJQSV0TV6fYqDMCprwjt6KI5qFPoYEu/Viz1RD
NfsnHEW1+DumdG/z+/Rppd4fyg9XgRcmsHGZ8+WJF4i1fObrdfwBSIID9NJTWZXHePiUi2BvpImR
hWXtmvhK0Vx2j7umrW+cBCnZIuG2aJwNptld+76KVkVOIc/WNpQKrPSj9CoZMoq1/fmLrbKUaSYB
bMTrmZC0X7M9R9yJSUMqjAwKbarb7aNaKiel9H6MEEWCvuxLzt+B3qNWsxbdX7pamcFXuy1w3wPt
ZCPswEHmd8gtOic5ctikBfwR/uJz0bdzITlT1aScXeUZx3feP9jviiYbZghIYaAapiFnVeXAdvD3
0/gIQSdnVZYHrtMlCumqQW1wmP72gOwXS35Ogd4hyuiJdxfUPlPX0a/TmBFYedx7eXbmdF5PGZeg
LnfDht8gr9etyBxSCLJKCSKtv3A1V3HTOT2oxaOtVA3AybZ/QYV8W0/TR8nWHqjv+CsfDtAlGrKh
m5Kyn2w/JwhasWKadcdUvcX53caDpAVrz4xOMkHa0F1lODS9SNBZxON83Ep+7YoOsrEoWcrovCps
+7fcVpQy3OQLiF7yfZ0ryirvq4Dej41WyggHsCRMG/rNUPxKo1jv0SlclPdIyjOusC9m5IpTVtSa
TAzYKT2St2Px9ciRVdTM7gSSqWXmZWEf3iZgMMFKBeYo8UZhSQBhtxxPmwcRWatJPdVzIFmrjv3h
P2Y2DAcY9vmu0ns2rL/XMMX2l/tpziUvvHVafs6TU9fVUfOkOK7rnEqPklU17jvGDtFpaN2k5f2o
qpCZIOFLXnaR/h8/A8bWsjXRbp9XjGfDJCPCe0G/0Yavk8ipUWsfGNruvtVPyYNC9eujsdLAMA1w
vAPRtIyBWbdgl8H/dFYhnRWI22k2DEWW3dCZe80tbEbUqtwp43ZdHAEZAinHzUdmxZwHPBFil8kT
HpfLbnTJMTGCnZHjF9HWVL05AzM6cotwj/I+96vHlGYgzfpUzur3T6NQIYnHegewwGYdZ1PfvuQz
2vfAc0MhuwzFaD33Sp7G3DIRdBeKckn5ehu0+UG54j3X2EqLkdoTIuDflt1TRnbjb+krR27+tn+M
RShK//IAYo7EkHDN2rusYvO0pp4H+ebt2JNPGx6TX5gsss4edTvrBy7ipTkqMTpuDWYB2ghkfDPN
gZevyG47FIcbInRVycYgFoFlzoQsxvaNOp+AiZNVCSfsrAiqrQtCYVdkhbWCTWYxCtEIYKnrFlGb
wW/vV4qB6eyYLim/lV+Zh9eIjaKcV/YZtreGwKA9PPSU0sYWQC5UOV0Qa9JdewDb93BsCdNVaCDL
aMZ/v2IsPDzHlwk8Oo6x3cEAMrpk5ZCtvNeiLJDSBMQlqHW7xmMBJ5vqvFW9KZX70dx0Jp446bUo
QKCONfxspFxBACyPKBt821+belwFUYKnm3+QOX79N8PaMzGg/9j6XCnIYm7r46QZexInYIAxERIQ
ad7S/ToOQU9oMhTvtOdai8Dgv/LXAHytYZ5aOdWT9cXmOt5UTg2DO7yhuG8qijwLkmOVy0tmgklW
fQdebHjpv1+DLzru5H8gZ6DLxIw68iY/aY/AWoOVHhquaA+xtE3LlQpwdUxGbss467nbD8YAOTah
d/MjhaO0WlFm4Aja+zQG5dkdm0Ge1M2xBcdoMEKE/7RjEkNCE6bjYLdkea39/WpGVftGHgK53ku8
h49VwgMxeClnqS/x3swT9MMzYrmA1K0MEShKz8ck7jNNYGAvzsjthfkIPzdNjcjhoCfpyHStObcj
odhf/nZ7Q5/ZFUP7bRo2UvNIXKDge74fBfK6Gt7IOHd0+Xy0FC1ESw6ohY2hKulptEbIAk0Q9rGp
A9f3MVB+Wjr4bou3KvL0bNevmJ9/1H/ruC9cOtYPReaPJK7gGR3u/yp4H1GjiC3uOIiFz2KDBTHo
QiTV7k0Y0Q4YdU80PS3APW/bABGkrAFoxnqX3of700am5vLm7HefUkTIn215KhjSkZmX64ESFrVF
NaIteuZKFJmLzzh1CHwh3D55cbYLq/QTM9Yv7iUwmrDWvNPx5OFKb2QGLO4Y2U7PjH+QGK+0W15w
3MPDNIQ/QbdNoMThaTQWpJPhfTwhpKJk85jppUS3CH8PNw54tMcF8orQQB75ftMG+ZNl0TtpTzF9
dcm1/QmHA9RaEl4xeZ4WkHEDgpnJtdaZJj8NapJte+/70qkW7YH+4pN6bHsx9+S6eCYmOfPcPKP+
ZN3CFiXdU/TyLPB6EjpIChOriK6+qOwTJT232gtu3b4e+hZ9d/jNQkDcdRwX5V4xRRnw//p8WmLR
WkowuNJjTFL9g+ogUSyFDlDTixFUc9ICc5xgrYJaQYbHtv+/RJHXv5SG0vT+whpjTuE923SIXmF/
qSJke6u+xcUYFX52sqgQwW0GXNEDtZ1CYXEb/mZWhguwtRZ3z8mqA7Pmc3mYsa7yehhZuJi1Eb7+
WX3x/TYPs7iU9ZCwp7NRJ7jA1+fIvTeRpfS1HwC6g8gofuoTBbQfY3j6/FhkOEUMoJN7jHB0jWnn
uVRiQ4X8OXdmeitGWltn7gg6bTDgOoZMC+NVrv4SgQUu8EcZvxq1FbHQlMW7cWJuJLQgVCOw7Bcl
8zmQhu4Wl/rv+/DJ5BTyGpInzHdV3MWEpMIA8k+KgDgcPqNP/OUi3nHxQQNmjOIvNaXwE72BdGVY
4RojXpFGWHc0Hhzv8GESpd7skaSctBn2jbrs6+LrewcwWBp8PDZsRISvJv1IwhNWg1f5D7Egn0Ob
lbTu7uVlLGKMHXJKryH3Vq8gxqrEjGB3rIoK35Y8EUbVE/dw30CWAHk135+Lpv83ExZHJA5+qcxn
v6nbCnZ57HF6dxh6jH5ASa4gSERSOIerJMAiFmUhssyQtdpGBlQmRcu7VoltgkMN23SRNMjrtkiI
Bn9tfewLYRmBvlAsRtij//5p6/3pdioUIqB5Wvf5QWF+W7feruJNWqt3KHyz91y1pPE9sBVAc/Vi
ICx2gWQSmOJ59N/qa/yesMKlVW/R4GftUKjAhHIR/DLZG7YarKvMDtND+b8IhnMoTNULzjahgB2E
s3zydS6hNBGe+Uf/5db/3Os/6KqZhbC3gVqXJheSxjOQT7EfOK3A+hyGSQXfhbdIyk+o13geM0Jo
Hipx0AB/48EsuH4ig0Xn0AtJeSN1Dy6kiIyUn9L+gcFct28cMDtAoGQ5rlcbVgDDVIn2p+txT3jc
lMRefIez2h0ydlbKxZUZwPi4SvCREVI0nxs8kcHcaWf8gtFSp4CwiTstVFiB5x1IPs0qIHkTkRiN
ZzUiXexMaV844NpMr9teYw3YCH/H4G8V5fHPrKDDjEjnyPGswz6oVL6iDqmBzXKxSDwQSnycj3YF
S6+BnIk2FB3QYo2OERMIgQWKDTaB8rMr+fa7NEvSW4paI1ARg9qTuCJ0POMWOUw+Gh1EWzcZAkog
Hwddd5COzeS/oXCnOQGgArSSd+ym1b5Y5QicCPFxVzv/COB4YKVcJbldM8ZbJTfnAnu3cOahj1Ep
FCB+WvfKQJP8ZMCzobuvYqGq9xN3mvtnJz9IGQcKrwjxsQU1DgKGGw1p4+QOLBjqHBdybgBocTbP
WeILRI++DDD4zLS9wVHbM2u63TePXrdX5l4gcRTyO53556YxJ3v+ukmQ9d3oPE8IViX2xRv9GgMd
lEwmkv0CYUSAJJCixbTfoEEN4XuBPbxsfheh8knxIIAHvEUIizk+W4KzcQQF5ak7AcxHtEoCWfNj
eG4rRg5+OJFoFxjbbTV7gRAzjlsabU4Ld2UPxH107vwsLT/dsnPAzfmLja/q/+HWdArtWnnBn5Tu
aCX0vsf3FlG8P34z/cV6Vxh6PlC3yJo5ODlfvGFx0RdK9JG7cKBShS4112C33uuirumeF4F7lFQ6
AJK9dVWkia+Q4DjVcqkN1RE3S4c3EI1FM82kmiw8ZCyJGYN25QZjA5SwzgGoT5Zaovl33sJbtxyv
DsMeJuc0/IMCnpvcJ8LJLkQ4eh4Un2Dt1EnqJlUx0IUsJMopCNqnShmulZoFBlhsO3cDQHtPbJhc
vqIQKUKbEA3vI/zNV94SpOVGM+3xlqAH27RHreGRp0uU+vFi4I9pTT/Dyfj6cxb/ABGpTbfeVNAN
WHYIldg7sLZi3wDEklo3MBYv6YlxylsJuDh3lmeVTYIuOXOsm1PIRWwwytXHdj9XACUVMBX4106q
cSe7nkCvFfMAosRdrqGb3Yr1i4UqTCF/xYqqaWnU9Lr9HRWsym+G4pBDrO0Q9TachfrqU0jHdfVl
twyHZrE5siYLet6QQy0RVoKw0yjCJWNKFI0FqSJ5wn51GyC69zD1N/BQ8D5WBRGw13JsqIoJW1+9
YpGaVZbPe+sN6EmrkktYmupvj+Pkr5i3lXyNC3aecviabM6jr45anuhdLY/4acGplT/+M4OmjqOi
JWeHt7AYIvY7TMHxtlyWTO+KEM6fONOdT14BFm/PIzBdDsW6MfJ8HKki/o4BgNT+Qkd9AT4m2xjn
VB4haoUCs5+MIeVH/FjqlXNN4BpiB/ZlDfAVRsLjcHtUGPzOPYTrg2w7xLdt0O9DKaOwsTFiswDq
qD+lvkE3eXOpffRgoCLo440Kx7UZCZRtdQgPAg9qX7LLDXYTVIX5K8zhy4lQn5huzsMIf3PMxHIf
ebXOlTgO5BhHbgNM6ZqxTUhHu/Hkmf7pXqPrP+Tjoj+862LDzgnKpz35h7XZB1/r+DrdPFsbMScV
x6uKRHdW6No2Y1miscVyoyagHL/CdG98FXfOMd2uzZ5G1ta5ALyO4FwrhJbkLdyNeYePcXHUVw06
a7swcTYnAdeYGZZWmFgS5afhOga8LI/74l8B7Jdqt3HUs5VfcDE7QbH+mX5B9YCYICQSuHp8E0xX
kBqMsW02e/5o6Dh5/kcv/nHGmFD7gfuwxt+q002q87YD0mPVJxDz1nZ7n3/cI7FjVi6jhCQmhqYb
PUTWdTl7K+29Of7Nkkru3K/z2OV216Oo3G7azsBxVKh6+NywUO52lW158KvoNFLwJdWjtXm72YWf
zdwYGik19a88e/DdWxJd4pVyJ+bXVl/FUFHI8YgfYJ7vxbv3W8p9Vt8liFY3DdSqIoN5GTfWRJTy
b6hKNZxSdGZ5KvgEYqwp1FuEqLfSpBz0bHsal4QVbffw5YVZjLDVk9eaujjXRptA6mb+wCWl4Dez
eoRAS/p09jorm0UkA8j1TlPGzaJR8aVyb4Rkdt7FXxhnmLevRbSZ9dIJctnDjlavlxeJAcaomBSG
mKlmkA9Zd93r8ooGrNbccDVD7iQoEOfot8DJFGRJFXWrO1YV/LX+OoxxsE1HrFZcLBVMvxt9mXvL
R4tegumvSVPlBhTipDd0zaoTC7jUZ5C38t8bD287vPzomc0BkHfsJ0TghxNVxVxABkFydcWpTM9Z
HJtLGKP9
`protect end_protected
