-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tcpTP91Xsgnu6ytdLPxoepvV8srKDvGo27VX+JJJbImmG0yn64IhHuHBbaIGpB3AjNnMZhNj+IHU
IeKNBQQcW3t7jtoDzlcNFFl3VKIwcYuecMIPsGMQFXd+L38WnmZnzi97SHqagU/N2uPB8e4gDlVd
jAXmZsqk2Xj1CRD7DmFEDuNEsfJhxfbHxcPFf98GFgi1EFImKH4PgJDvK+BeqSWq4Iqgl54vVn+x
LMmyjTuXyxnTYno0t/jDOXiF0G3cl5fENFGqTdZUtkSzvmijMy7cXEdNK38nidMnsyN8ZuUpoAdD
zfKyC4JnN1u4e8u1y7ChBPjLqXGK1guedZPMMA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
gnm0fHPcK8tid8I901YopqW5fVJVuc5IbggxxbJ5A6eo/cRTb4AzG6oXHPMDrCQ5JVsGFoo+Oj5e
+TOFLCgXYmGXrGP6Lm/LP7Km8LYTNzY7BQD78lcjJBf9+5FFK0Zmkphv74IxMOSbwj4a/nS1uvSK
uI/FB4oLmYsPc4+6PWWaoGD9wcd7ejabl4snEMJtZnirFM92N/iwttiqrG2XeyJ2QftHAhtcmRKW
KRV9VIGrlHIGi5Sbd88/bep18gxj25a5G58WpmPAFCiDznstsWAmSfat8hvrNSoiYZW7SEWFiyEP
xuDWt3crkRQxBMcgBh/RHgJCmZdHz52M2R2HSL3DDVjz2DtukZC7dK0+z0Pzsytx1ubSzf/S8Uc2
we0z3jlu5w2EbYMuTEGlaURCk07oCAYf9o22fhA84kIaJ7zilC/FsA+SwTYEG/fau2D9DkI8/tl2
GrbKub8mJY1OHd5jLOC4a8xQG/TEe/EH5PE0QZy/4fQXAieqN7Gxh/vs5Gg65/yE4qxn560NlElu
8NDSmxUYp9aPFnHwqUQgG5kN+D17bpE1U8NSnZ1iF9cPVap+PCBUgh7gztSENbWZ6Okg83kWBFiT
EruyD+bTPRUAkR/esfvWw8rpS+iEmwS9Um1cSrWaU5xPryQ9xzWdFJUqWeZKmqI4Tm5vvJGIItYT
jEJzb6eHRTq/2iLwzziQSCwh7TyPkPKJRXS+aQlrJvgcQ++JVDNC+8nHlT3daoEZagAVPO6WI8zJ
Spl21vwh+jTHc1y1lmnypWolMHQar2YvdqE2fP2t2I5/eLTB8ZkreyR3WApIAqtiWFw3q0MSwdis
xIacmX0iM9XLCItIJ+lEYIJQUSX7ZGWgu/ZgH/GtTN2bo7BoseuJhTS3pGeqpb0mO/xrmmX+q1G8
wdOXURK44JRDlz7xXKGz+wGEbEt+g/hOo6ekc8ckU4k0F1UTv/17Te15w1xc4n4n1CYJ5JjF7Aod
xoGOPK2Y1EETQvcOJImU9ACa+ceKgRFAe27pUl4erGMTd3hPHTXZKpgsvO75+zdBMi7kDjjlulse
11e8lDbi6ljI8Dqbgo5EUj9gLrtvGNn3ePnK5tpHpzaX3RWIVr91JqQnlbgpx3XZ6nASAYUdM24X
b1cuaZGmcu6jK8ivBlmsgAVQPZrO4FzFkIuk6GUt13h14KA0MV36hdSZ3mmy+nmGia94DX/lZlJV
MVYlY3+qdyETLHr2G7ZkWZnai42e/187/kohIfsKeNqE0nDx4HuMUh0WElfldQSfHQZBiN7b6qxL
1Pr+Yb3At0wS++z7i35uIHaELRj5IXSYHWXWMt+S6aS+8kTMq+Ic1CEDagqT+wsyfm6y49QtK3YK
8M8aY/xfPpILUZ5dcHu7JhfxaU1hvUVFnu++drG+Xxwq8npuidrxoTay8g0i+AXOuSxB3q0jFNu6
3riVvnSEwOARNUcgAmXI69VzxFcJfGQ5w/PZlsN4OJqwr6r7jhiSbp94mDil4OsbTfYsz7nrUoOT
h3zaWVBkvaUr8njZlJzT4ccv2w2v96gNHo96Y1b7Qy1hMgYyZ+T+hwLEwwSfTBA9s67X/QeJcnm9
nuh3Gxg4j690/TMmhJ+0OP0yKiriE1HM4rNAfURKZJwCMu8DkdQoUWdM/bdUyhsOmK5+ag2wJl6k
Lxj7kxc1EM+NlM+iY98Ut1fhWHjbDRNfzsKVxj5uRAcApSVRMCjxcRqzTpZpzHY0TaA/nSIdZhfD
gWVKwANqzy/e8HEzqu3f1ejAaiZXH+2ZWeCSpVvhExEXJo7S+prECGiISSMftWi7jSAOXRcy+sMd
d0111JtK4fvmur/4Rj4ANISgpzGrAjQGdElHT/vOcXXxAfJf2fp7j6TDrZvvrRAR9VhLceZOZRDY
yLbGoyffKlQmsbuTY79YBiSjnfUCPJlFBjLYLr/TUHja2EjK27tH3AgN/0f7UWcxkJ68nYNxomAI
8thO4RdtM+cke8iThq2Stc09qRmQMXsvmnYbUPE0IWXwdydIiLmNj1zHl4tPUCJjCblFWHtwaoi7
UQZ19T5342pxmdB/HdniMLdhIyDeM8PfNS+IzcWds+cEJs9KCWx/QvUYDHeeRjowN9hI2OwF69qV
Cke/whJUerbIzSIUzHaQ0ySk/UghKBNVYPLY1Xhsop1pP4saQOT2QuaSork8nzpDjyzsB+YOIX6a
tCTcTF+2OT0SfK4KUYGrGjvzgrYRrfDRUz/Ha/2SDbTsxdI4XUy027xet3yJKg1MQUTIlIidTPOm
m9T/DyiL81UHzbhxj1sKHgbp7PmjTdvzY0Tm5MkKsKxtcAyDBs0hNGNOaX5ywtNmijLjiI13+eGe
hGa4sVr2ot9rt26jRW8G+yUnYQ2oLpFxM5SBl1BL+NENwq4u80JtS6DLTNXXdDS7E2VsW7F1BUd3
v5oWLASuiN/6dl+y7LCY7R+H31Lga+oyyKOuGIZsTN+ovm0ej797ojdrh/re/oApekpG/rW//y6Y
2ma74MDMFlyhJoLjqEjhU6fy+cSCynOE25YpODiKr/RYs1eO/UZtDQHlnwyKeyHh/rxwvnHRfxK5
o/+vZQ8ffy88HZnbRJgSqcK+dNNa10Rg5QgzW1U0xnieHNGF6JJ5cLCm+9YC+Pi3X+plnOPWTI14
/a+mOYXI5zh+aUQNhUrX4T+yjh5ybucpM3NB4RTMCWPHWGDy9YTn/xOr0ZyuAphtzNCbB2ZERR4j
AARpmaiUyul62j27MTWKBdFYBad8stYTCIKgFE5ZovAoF4DNV+iS/tfD4p5TKtL4/e6wz22axBNr
Q1zKz3Swu6B6AmZwo4emhs1NvVBn6iwbDxBtyYTdr2LGYdv/BFiGP8Ba87ylcks76PQT0jd5cS3R
O57Z4CdyEhSwJvArQq7OGUETygLwrbTvWwFkhZNfh8msEmBNkfmy0NIxb5BsWJSP0/3qwtbt6ujB
dI2WtjmZsh0676m7t5+sDsCj88s7tNN5C/nxbrBO2pnDny2LV78P0218siao6C6Ucv8huRkz+4zQ
5CA0OBG/grBmt8vNIDxxPsJhDR1HX4RMUMPwbAY8Umzs9QH3qVF9tdrqua3JRmwYjwkmEdboj+Ku
eY9Aj374m1/52INhiJ5xP+xtze8J+nxYrW/yPodoRpCjoRtOid1UMJl9RVxArRKwB9Zdl3CqsZcB
qzbGTJn1ZiUmJFrDUa5ooKcL+Nj6ZBGIZXeN2Ns5jgK3gsEmikesKFGTs1n6osl/6Z82mPA0yEPj
tDHwqK00/yyVNkCxrLGlBevSylODMq/8I9jp0pBt8x6Lpxn/sZyfl1aTj9nz5PspJavBFGKok0+Z
LUcnU2MH7hh5HTBkOeVGag5UKzfO49mg9W8eMWIWLJsJBy4CfqXDW2rvlFgt57EVNzZjbWfugzgw
ubYPNGM1WzOrWPnPLbno6YlVuq0lRTAP85QkYN1aylYwHkq7ikccIpESeHqKBwca7WpuCAmHWI4T
9q88txPEW3KEPpYStuDdspHz9H85opCeoSj9LiJLt544K0yQqA6s31CJZ5Y+4NNJfe9SoDFVpmlV
S0TZzIw0d/HIZLVgEqF3XVHzg0cqqxzV9CqpnULK6eBXrQpFGWiPFi0v5WLHAofxh1UkMrNChbQn
LuL+cGmw+MReiCUBG0ugiaoBOYKVyAHGtk0KpC2bGq9Bd6J3wIgR5sh/neIaBt5udKQ661rBGeo0
hhVG5nGK+n7bP7rwlOVJXOZ9mF9effHhO+ORr7sX+4WbgitW8hfV3+IG8FsjLPjx5pb3QPYmnToI
jxvcaYKLPyKNi3q1dpwBtH/OcqoCCWmV+iXPhPvoRIJZvtkKr9dUnSWhAQLTWlWw7AmuaGnE2qfG
/8U9xhJ2lXTjiY4VAvUUFBw76bprYIqbz1AmbLq8uxqMb4cDQJ8fr1mBIK97pNLudZbbAcnCK9iR
E4idLJLSwsGgqrAzeNDKuK3KqwkYmMs2ufE5cabUHJjxDnE0qHU4gGJtMx6nRix6NIz/Ppy8wYee
8bXdHkkQd0RReDNlq5p02a+Tzjh/WbVrpwzs9tBP8xuKkdCXs6RQdIvZubpblLwXVhHGAkeiW6uS
3bicUApM5zT2rFLwn+3eiN6+/QMYZXfgN2yNKt4vtX+LAodg+4Fl8LtMmk+wx6QBR6SewATCUP6S
7mqDtZDU1JoF7HiKXOmRT7ADHAHMEf4IYqegEwTuth5/TspipgB8beKLxxPVKPA5EkQIwa+4nOUd
6spyStVYmdX1soldPpxnpfG69ztAxkV77MuJYrlugxkB2WY7JoaUiUB8972HfJSwsydDUbhQP/gE
X+ki/7l+p87uVB5UFlsNDPwF1lMzHZltsfZBut6/lkGveXyoawJP5mU+FDbdRtJBLJEoD1HEiK/g
ODcO4q7N6k03U7u77xAJ+i3Mfnn3UkY3BnvgDzJJsXtXM9VFsoFgv07zrXYhVpm/wMBtSEjoDqim
Y4YieDrbpTcDwK1Qireg/wVDMpjOhUxL4IhWYeex9hc7U+N0RoYF9pssDCiTWUq027WiYgibLgTT
G1PMujjO6K1k++hNamTA9F4YTqRitv98pzKxAEDRih4fSK8hpAb8dtfXSehw8ushTNGqI7BvriOX
x55USHXBg99lFehfO7wk+3UdIYqYrxaEYy+ZnW+WMEBJUGDiDeVG0GwMFDj4evFXxxuEeTV0MslC
29xOQ6G62O5OUmjsGXwPYZuKB7YNkT0fEH8qZDeAk7SLp5MIGJbLBjG8RhJwHJz/PkULokeqcXJz
WRbX8u2t14UHt6Vw0c3V7z9ib/jPaFzmbvVwKhQPj30pZJHIuChNxtkbiWq97qK3rw9VJm1AaBnE
Kd2abUsYZ0JflQh6iAd1+sG3SIOXFp5d7bMZLQ2wKvnvXPPn+qZdEKC7UKy4XqGQIGrVCxBMcu73
QeCHG7cgF93cZffy7r23fPus+OC0axV77l0Iy83b02GEJR4jf0xdApTttLs9oypLyK0qgLa3FFQl
xgRiTEcNqfocg640RsLP01ZR9Fpjo+khzrJgynD5t8revKKFVTIz9+UlolB7wIVckMTLYjyoWYPd
K86DngjrPDW+RC4FUAhDCol6eEXvKPUB07Y6prniL+G/WiwdfMbPNTbTDSf2GDbwWDa9AjqiQrON
bPPI+gtxM6g/g/ZnkNlKFNltYl61i3oG8gtsAdenYpwXEA9OA0u8GJtpW7MP2jw5A2uA1SdvsBak
mFn1q5Ox8ezPdgmjdE/w/iFXpR1prUXiEKni+ToTzCS5mGFWxIixKQ1v4KWaJUkoNp9xUfqOKc6H
MHyfHCo0vvT9674c/vlsdoTc066Pkj443aRt2wJgAnbmYavYvq7+iIHmVd0uGs9rzxEelr2Wd47A
E08NmIo9pZiQLI5V869P2NSndRZZ9LwXipzayITyvBsuEgUs22/0s0Kb+iyfRO2B8/Qs5ep+Glsh
cmraHvKXzI1JMqbIy5Sxoxv06ckP0TD1R3Lr+ZRfnY5AX1ywGuDaWEWOOkhfiGhnT9kA6eiHYx1Q
0413NkbO8RaTq76veozXDIvGMJQEiprSA1y3U6jqIuztz0TtNOahkM0gw27MFzSX5h5FyW3Ocsbg
dwwvpO8ZCizApPpSyDDIOe0SRV/cd3rKZ71pgZZ7Hgm3q4XevHpkpDjBgCrpl1VMsK4ktRSS74zE
abNoPx72xKiPSvkpXB71064P5bKL8iL3UG5+dZhWPt7AF1fG8DEJnUbIceIGSLmblJsE4Qg2ilJz
6zw+PJeyLJCqR4qY70JWLUKUN7c+vHXivxnrI66TI6HxCZIePl5hiWqlKkpPtANxrJS0I8Hgr/Y1
WzbjmflCEO//aYu/+Q/h358MTtnVhNNZWEWS02hjEdZC4hud7G4C/ikil/CDt9n+7NVszpktQpkb
9PruqBhxJFfSrORjVbEIt/RGE/vtxlag8lTZPfe3j91GYRjV0IgguF8c3DlhQyOyR2zw4DdsVJLL
VWkWHOHldXpi8t42HnQLh8D22NxWj41+wHOsLLDrmArAgnewvY/5PzWbdF69NgfeQvZwREgFcJE2
Zi6D3Pwfo5knjCXYl81lzErcxH9WMqJ/t4Ps/2wtoFq1kxhjJizxru3EMAIc6dyJVAS834/kkzv1
00MKq1upE0D2Wm9WbIYDbYtT4xwgvMliWL96Hl+9AkrFoqtLKNLy4MyTNeKNUqFpDxASD5lStEra
br1Ox3Yoq5Y1azQLxmZxg6CI8AtsnLxlWEYS5Ejz2r4BIaOlMAXglSVd/E+Ntmb6CU3p3bG2Y3JW
d9lIMvbozFBUxJ8qzz4baProBvk0K+IUy9lF1I/hqii8kxRzrhEyVTznu/zGPZta9X4uQXPAI+lE
priNhCoCQx/rtpAtLklEnQ5+UhYyP9ZhM36Do4sfYiCnhN1pD7Orc0VCw0BXRQBHarSxWt5QfKRM
pdC2CIfsuJk1P3MFMqlYk1wBNsVqVvnRvOQ9UMWdoSxGxqJFj7oGB3+LT4IkjtKrXU4z6xrRtZ2b
920wNZ8TuIOE4skukpTChtBQ0HdEpnd3U35NEXeMxHML8vurCxjDZrmJPed2gGb7gU0x/WiXSOJe
iYXvgZ/nFNzs3s7WzrxaLUMQOyyh2OvPZm1lt7Z870JNENqxQjo9djWRhzAZOCkMg251JxBHOJJL
eVIVSE/Y6t+mOcp6ZMCnmkU8cqLmbXhNtZVIfJ9QEy7go8wy+2fnGGU2YoA7ndNX6gTbGG1meVnR
L0y0kpFvkjyXi0/63ezqjU+Zl0asMRPWNhdb4Kd0qeIosO0v09Ro8aSub2Tfve/J77witwujJ5Se
f6YYvvAg4JV3qnzp/Wxy2BlahRrsJakeI5czp8+9kdGVoOQf1U0QYk9jL1joKYfnOmyngLfEB2iE
sxrk6wIrk8KzoyBKrAIWYeLcoamtcMZAEJN3uXdJTnExNAOiku/86ACL2yjlxlVYzRQwMyX7rB6s
xgYeA3PEt+f40Eu9PQ/e265HDFYMc4mO8eJT5Qm4fMEWXY2SrFezDJiUxANVyWVzhAbMjmqDObpN
u7x9K6IkAuA4HMJUjliQtJXyoUMoQmqdz/xwLmjk9LAFAhJj9a3Hr2xQLLevLqqzbtPOwqoBGYpn
5lDWcxwlyOGe0sdFKijVN/hb6PAKgtK3l28VkSv6WEZS4236LRrZ/aMiywGWTZGE3CYZH0WewZ+j
mZpr12m4JiISQEhkIJvJvsQzc/pDD6B2YvM76qAszdmWfv6PSKrHgmHV9UGN4Q0w2RjCc8U59pqA
u6i+EvlXPQhwrYxC/rLX4DdHErt95FCZhYbBU2L4L7SWOEju6g+W6craRPZcbg+As17jHBq/ObGj
aVpC/EOmC2037EJnO7MJi7fhDJLyRIDipF+3LhZUL2kLn9kk5XJ7I+xAzfmIKgW7dOSStUT8x1Ji
vNTOAYfXLvq5CfwO8OgzYGysD5zAoUyGC/npXOfXJUUax1I0iLqk7zOsJceJP05lpC1Vys9r/aa3
RQbTZG2LxufLXL2+DOE2P7b8y3LgguSBXlLXYgA8Rwndwd+JOd5AVK5l+3h4ZdaXYbrGTe8Y6GHn
Y+DRIrWmzp2QR/MlH1T797luj0GI43JDNP1AdswZIxO8ACJ671kva0WxC2C2zJIDo+TTu///Hjst
0n5vZkqW1VNcQqj23RMNF94a0iwbF9X3s0SGXTiXW0Yo+o4XCuWqHRxCz6SYbnmjQTliBMEXifsG
g9u3PMLyk3rQ2KrteTWuwkVBE2EQlae6FC/ULVRvqx7zcrbFhbO0WC+YgdWZeuxNlkRwKqf3vqwI
NgWM/+K7+Zb3SiRailWevY1kj7PKGHU3YjO0yHUl/8zajKteudEphcwZ0CFuzXkSFDLLqn2/hLqP
XPaYrJvPhibfG1yAYzs7JkEWuXFSnf9WztwolvuwOmzotF9OmlZCniNFDTJqaIQ8C5+gI9voDFkc
FvCYU+8G4zYQ2i1bWqZRClK8VGzsLVTD3i5GOsOetwkwLgPp/y43F4ejAQLeEV5NrWtupiYIHqsN
qB8o1opB6gfOUnn8zsKinH5UMK3u9oQwP+Nv8QJ8hhf59Q+Jf/ntQw+7iNIbfW/p2PKNhs3iYpHG
J4r9oY0VjbUntU8pzXprBat1Xj9a4k/kt37gB42WPEt9tTI+Oj4FU8kxJkt1H73AOG1YW3qy9wp7
l6gINnHPgfmkgYdfawg3gQj/kwE1d44eQFxWc709PNBdIwTWyIsEzZ3zDbBr6En1GjSRCCZ+XUHK
J+Sf/+D3p7GfME7+23Ern4AzjVfpwTuzNvgrEpEBNfjVE07ZGeMsM44fP5+Il4tfTKTFL9ts83wp
jw9UyikG9Rlq/eFnb6PecoFbQG4kL6jKXMXNHKqfB4wHNg1gt5LqhEoJ783EeVOdbpr5o/9RKfzm
QrJJba01SH4D01/8/zg4Wu/CmMJti8GQ9Y7DBgdT28kkzhvMI+51n/ll1DmNYoGKDVkc16aRzVx9
hX3x2WBYn745qt/1DhrK05gyMzpv7EYA5kfpseYL/pIvb1cVsUrkLP75rdLjHcy988LHgucSql3B
Gw2abmowRwWvV6d/MAk/F8ZtTqhJliLk3RQXyzolSttDATHaJpfBiJR/Of1j0W8tYlN8ME8DJ26x
aZVQQmlr6Im9bcd3Aqsc/ItWIziSZ+MdTD8wW1DZ2fFcQXQomktGKqIUJAvcibxrLgWAZOlfehLs
p7M2AEAedHFqBbbeQgQ1R+HIJ3IMCJ6ezK9NfH4icAY7WgKG2Q2TqGIxnK5EMJpbYl/CZP/J1fGd
gDcmVJdkifmDauXgA65+wQ0J1Gtq+ll0LY/A80RKqYG9AhbD7+b9m2q4i4E4hWmZf42iApCRlzFY
NvSJLFcOg58nBGba81TqsX81NWghASFd7Z5ttqgzhvfIq23Wn/KX31sFG369cIuBfQODNB3GOp8J
Sn7NNs/Op7x3NBuTK0yEXXymiPa88xNuI1EtcBk6sjZ8Sx/ZADkvzWpqi6R5EmxZCllJPgzzYZr6
Dl0M0RCxa2TobC7y/JG6gIJz3GJtkJd2e444JiFfQiPY0oobs8xEwMpfx5AOOsv/Jm8DPrYzTZiL
3SALU7SGp/JTi4qQ8BLSjZFOYxrNjFJ2CG7TF66bg80bySlocyXlPvfrO7LJnEB4bNY6H5aTxSy7
neMTY0XFbZSP2SG4/KDzgkLKJoJttH544wvRucD5STmhmt7O7aMGNesGX7Zb9HG+0KGvP9my3/aT
dneId/v1kjgtQKhoqiKVyJCsle6Tm+qUuoAJK2Z1MwJ1tAa88E1zozdBgYivVy2NMQkopZ4lgoMX
VjCyHRYfEor7eNXXn3OKDlQluXHfEsM1U9yOZ6OjehamaF8nk56A/qMzqiiv38cJw2LB309X97PV
bKdBGMkLfyBtSLJxjYaHIYyj5mE+bVNpN0P7+vagbmZ/nQhyYxJZqf+LAXXFtAWs8TcRsAxEhCNy
oUi6kP8R7gR/Rk7NcvhYJVTJbJ2Y6IiMGmTGlKGN6bYB60DZr+N0vH8GMioEtF5faw3mThSEfGFA
EZfbcPSmmHFZZqGBmA97r3RTotStuQ4AxEaJvmk77GPHEmynDaIbczujjQCqmSS3qR0/VzXPm5KH
iX2CMvOVsATVVm7WTZj1zFM5JYQ/fAWsX9+uIsfobFjk8yWWKQnTX0MMsauOnT3kc8Jp0vI8HkcN
dsHLCWXBMEjYGdYVq6ULBwW2tnZMs6fRMRtW9soGhtsoBN8LZKfG9ja6t71njyYwkVgQxGj95Uab
pw14WJMD9RoRt4VUAgg0Zs+Y00yiuFNSYJPovbh+oHBFHlFL+rEPCqEiuKSeGmbG7jxIoWE6ln9z
+EcmnD5+mLhnFp+qnIsqBnM1gc96B4aYdJgXcazZff/eC+RQCpmoqyREDEp+7cTxdGhFZu6hqA7G
EZ4d+5PjjwK8FXi2f3GS113oek5FgMrSN9pSmwQ+++x3BjXUu6p3d9KUZiV/2lBk4k2CsXZUMtwr
ByME1L8njk9lMPM0+n2Q3rqR1xgzE8rp28d+jg/GBUPluQNOLwBkn16OgVYlfuCNx0PV60UoYfNB
fY+o/sCmMXSfmy63coxLuKKpfsEuSbuJESeD8Bz4Ste6BrFU/lbBETPmxSSwxORTCx1X3t6rtJT6
Qit6AXqC971HdqRRvRCIrm8TGma2g5yDK7TdZelQCB43FmDe4budSG0noEz0BD1O43qRiPvKCy+1
pkEzaRKfDxZR0k+NuZ6pQweSFBypmnYj2a94kEiuXRAWKxweSt/9FVvDwx9gmBuFXqmM05P7XeiE
jcDbIFG+aO3RdLK33Vhyi+lx2NMFKxYf9vvbFBESoiADHukc7X9MYPjtDtgwdIJwaFIWbo7TGdd7
E+/g9mDjpsZpJXsQUMXoEc+/oqgk383SlASuUIl8pKaHS07OJkAt3ZvXw9FIbNTxgGzbKRwtAgp5
pcf0Xr0ZKieDuMkOjdErUu2cGWCSm9ej3RlAquHMFKQqB1jt3SuEQxH//aTVANKYcC979XmYkud0
FTCFP378lbknlRdwb4C7J8f+1uf8o4lS2Xhz6Nu3AITCj+gHz6KryH54uU/kZVKy9HtTNO2OXaNH
tGFCGRO2ENbr2xygebS1Xavfjr7xC5t6vWaGHEwmdz5Q6+lvQcI8fpG85yFi9j6n4llILVN8rV/q
BASYfj4hWHWlogRQO73QbK54a/PKbXBIVUJB8rZ0ehO20SZOHbei2Hj6lrgq6jfJqMNHH3hGEWww
zffvTOQCdlfH8iWI2HAlLkLyQWBrgJHhjO5Jq0eGa4e5OaoC9uT5FvO+l3F9oevkt4A3Z0iK0+3Y
fA/62vYd3+xfSjXUnJdqRo2ASrzliMYZMgty6S9kn/1e9vyf6nL4Am0AwzyKKl4WGBkvxB3y9TkL
JkJpQgMpuNE1DmvOlqUIX9EUdoIkRVHXt5TDFkmD9hFOwFF3o9s7waVhze+6Me0sh9xlZd0tb6iH
dGD/hPtgzC5Lj8XeF1LCXqhxH9v5Gd+tgXLVeWiF5dFqbKUvl650hbC8RIGfbWPuY67dRMPpP4gO
AmvHy7mxkDQWijrZiQNgFcFZ2ehu22RvMXFM5291Qk7Be1lVbN2gBkT0GbJElYY5Taoa65uWCXSw
XcgfI0KHox2T0GIhoVORa4/dN06N4+aw8dMjL4n1WKCQ8OqfWNnsnkXxS2RavlPcXgQF1GDlzzOA
akqCZxVQZZj2jODxoCUekcwS1skDcyrN/cPHbndtAa4udFeaFu49YWa+edDHowKarPqOHWem9EhI
/qIebPC4rlTecIVBOyEwVVh/fcV/Ea9WUYU5icc7JyUTbgJgDJ6ZSW5KHMReWKejhYNnEiwM4Off
/PwpNYsEBHN8b602nXoyuXYGAa9PGEp+KtX7g5qpLM47n92yVUFrMVHSQgWxc6IEf2f8Dn6W/x4T
Qbrj6z27sK1ad/3z9+8lDRBazZtdBla0zh97FFiH2JCbwOaaPpZFIanzdFHxcg52/wwLc/7/RRqB
wPXdk8VA4kr20WQ2iKYAsoPDE08lmsXGda8OFmOJt5W9AIm0iUAxxm6zhXcX5Q7hSq3MDU3MtRvG
PN+NWYUewDYpKCsfN2mdQobWhB7krmp4GAci8YPfvwdF0GffsrXnYwtn2uF+bA5xmqqrnMdQ04PI
HAwJYY1kz8FAfXDDwpl67FUy97jS1r58f0nvaDCGNH3KMclus0xP4m71v7AT6jWvvBOOBsIeW00E
+DPwlHeayfJ8Ql7dv8c7EdXJhYxFcHEs3s+B5L0OseFEmyrHjZef8E6RqKK84mvwfONls+90MpS4
ZnIIaVlU0nfShyrJl98IgFLp/9seDkT0BzaJhq5TaGNTy5Ys57yRFLs5BlDWT3rjJhPfXcpRH318
QXEHYbKIbVwxQ9EcR2kJZWm9AGqk/DyIinvyYb1whAZsYjFQxUrK/BifXEudIuFP8oUeVvHmIKH7
m3392tCU1ZPuvsN6b0pCMexzMrmmqJcDlu0pUUtsf4OUcKqNl0VHc8urtDZ91wRk5utaFZuYlmNA
AK2OJ2e86a+YR8vxm5fIsIr3ySzq3es2Jzpn02tyGy1UI8Cc7x2op8JIHtmewpca+lqcJBJRvIrG
GAxQryLMt6b1ajXyDpAyB0303IyidQlMADr69TQWQISy6gZCK5Onr+4t8oLFgtn+FIEp7yOmNetv
3+UpXlDTwjGu6uMKZ5aG0A84SgeyVo19cdDrVxtWG+JerrClXd4XR079PdApgHLPq7nfKtAnPR1y
EgDDYX/HYL8jkaG9GIdyKNtTvsqPYBMpn6WxvMlVXinu59xOk/z5ASbmIqDnwYZidPh2vuSCZtLF
IlHjK7rIkSQnPIUFyimGbR+Qrw/h/Ipk7GulnR1MeiKc0kepESLaLLfZ7jbxhI6s+FdSoRUYHLTF
REDsiU4HE9ra2Y1zaq+Izqa5q72tMmGl+bJ8/2/D1Fo7lgdogAOHvVnDS2d2Gf8qtVi2BWW9W8WC
uRBL0u3H/TSdCdgDIs/VlvoaS+Ea3/O8lQiGb2G9jbadOgyF3gTq/i2Jgr5cwf7AipdFYYiQIwPc
l2ZTKAfr0SW8Dh0zlDII/SvhoStwkg4LL3uNvvrPPH28mXGT7CTjPOFk0D+6PRhVOXV/l9FrIJ9F
5Ob4sBQqDYDKqDaR0ZnseqsVEtm3DW/GMpGHe6X1x3buQ4rk+c6ewnFlt+5t+Kc9OXgheeVXurAG
JwShdi+f3v9yATk7iG4Qwd2BWsD7VCG31Q6cWwFUC2hkyj5IrLD0/6xuaWRcoMrqpZI12TX3nLa7
cLB0m/XUnPov0mdyJ3QgKmZBFdwQCHJ6zh7rSyt4QL9m18uRrIC0F+x2628cKWINesD/+Yh9QaAX
k7wRSbLvr2TIABYrP7fc6lJZRMLbhQ==
`protect end_protected
