-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KinNNmRgLTTDx+iaU2Y6Fd8HOvRPSP/qg2DO7SRgR4pEKwObAzm6ge9h0rX4Ncty0s5/vrU33DlY
93bF6lgSxrdcbCEBfJaMtVh9pg6Eji/D1+lko9g9+JrzW+grhDj4Josn+4yoGmAZeMoK8pLSAHhh
VgMMjP85cjqegkxmU53CEjKbyzWaUDag3TXo2DFtyQKvA3qsPBadqZgOZky6NXMZHRCNxcV8xK98
4TDY0IH7ILpW8YpZZ3cNXZW6P2pt0g5Rm3PK5h1qij0Ex5Xeotb+gCqYJPmv47ZfPqYRddGY8Z3f
Q8z0JzrCYoW8YVAZszuLTbxf/tioVRoaNOPmOg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
1FGqATb8UaYjEHUy90xaPIT/5L1y0FHiieBu0sZiatB6hpeWfClTjKYqjxpNopfpB1gnPFblYPsp
0dXDBixuUmiz1hruYy9sA3wKLpZ/tZZR9t4RNQXHBO3iTzWJvCfRpBMGgGqtDsxV5B+iY5A12YSn
Q2EfdqtenIp6WlSZVHAD03Ss/eKk/Se1x4g3r5bB0NoJXCDUXoFGVnF+roy+GfIKPUzeQ/Gh6XlT
UtF+yQ419O5zuBjGTrQI11Pr0Q03nMnn/BhVvy0GKZoY8wfRjIGytM6ZHDtB8DnccqAa3gDSF8CB
tYG6PrF0CQaPTawuUFeocuhAA4Mqos/upN7KeeBSImfGPo/tCR0uF8r/do5IjrnFY2c6hY0/wM3J
l4JdPdEL20ZwapxomHhuFLCkdTjbJa5BKFJruElblclV2f74Mz5WYXUc8fBkhb2e04zsVyqQDgvL
qAdSZ3EvNPCjXfXkYJfV2khFdi7AxPtTMxUyUgVdBJqs7/DUonrZx8NEaZ/QTmqwaTZqWT7sVjKG
kfX0nmg7FiKeWmeb+JgztSyGx7noPUqzAnFXukNTliMNwOFFgRLoOI+eKugBadL4mFgIYUfXYCF/
E9CMx/IJofBEpr2zyatuKElHbRgGPoYmCIfRlSLPEHDnQOf1LUgjK6pXYsj2KvEhtUFMmTI2HdrQ
jNZE5pjZ5R1Cig1sA1bTVJwgjLcQtB/zRMPeZM0nodTylK9Lg1gmpX3YYxob3QQ76sobg6AZQplV
u/V0QxJQt8zR6Qx3exs2yIDW6bd+5q4vsBJTOv1/ZlZQAN3Y4DKD2KYkzTkpOHXzMhawgX5E0aSF
Rm4MnhwOknVSINzKVFO2ESbapCy0hPsbuTEIfPEgrKi6M8io8DRAXil9EzY/0TCcG8FqMDEXrZ/j
YZGugeXFUI/0PRIdyEGg26IW50uSvOl0c1P3S/v721N4t+HqqoCNzxK5+qBJh9kCda2+r41lks5q
xAde2Tcjd+fRVyH1gFkOt8v3Nei6w9r4/dmDfgRQ7iyJ2spGYmNolxgROJdW9iDZcehI74pI/Wct
eg6J6qtncTv0pWnclWd1rsAqWbjX9LuCs+7jofAOXJCi8jkMbDU1fdwdK+kMA2dVgCCTqxYKndXv
ptj0rxBNGbi21phAuOvssXsyy2gp0Omsd/gCrK3Pp+2+1iRkyWJSvEClsa4yQdOzzK3R3pU+m7TA
wDmkXE+57ItWN44lj+H2EpFuGd0WI43MsoDfakGK/oP9r+YadEEHoUueMOZocls2KFwI2bBo0FGg
rrB2WSy7BwvDBQfsXH6V9kLk0iWwEHR5twf/wzngqDRDLRY58IDh5vHItGCQhb0cvEl6KE9LiGin
FUR8gSFX3H5x0J7TV4JDKq7umPqKMh7fLU5uwnQ2/2OjycgahlWcyBOdjcpJxagH6QakP+qvLsso
XxsOPOO5W9UL5uVlEqMUIiZto4cZrlWh9hQy7bGGIe2p4qDaZSvj3iY9E2d4rZVMpAUGsA6zKWuy
MbaHP0/dDLC6sBva5Y3yjYEKcYlI2I6fQGNcLrNzRmeoboEH4j3ZiOcZ2Z34TOcTxODf74tMbw4V
Op1ytjCuh7X+8K/dfkE0l+c5uuxYtiID/tmuCEtl66goZLu462X86nasQfCRpbTXFHEBw46T3Q0S
M78aM5NusvNal49XrvRpipLeHP3FAd7PpKNbV5dgD5ClthnnvFc1M5yszvKh1iR3+S178Oof5L7P
zZkQ8/3xu732TPcZh9PPjD30S8lqoRmIrlIv8L5a2i/IBfX+YlUs9Uggf1w9DT3SGeMol6dlzUUK
3ZFySs2v7WpgJdIonAQH/aDgD/dm8XTJmq5xLzROx/ZMvnljyjouIL09dRDJt5q43VoJ6mm6DSsS
vWcOYkb6hbWYfNGJhX65Xb45vhT15SXjQ/ZpvloOFpfoKh0TT9yvgflQFjvTD+5m10665kStvts9
wkBMeG1ZT/I5Uz2FRmCM8KrcpAMpck9pUqs+1gpqy4VTGAhZi2ergXNYKU8jaH+Qn7bkBRycfgGY
ZX+7WUEUJbqzVJJxPEa3H5giF/hIp2ivX9AYV5cjUFGmyy5ugFT6PHKulpnr3ejCt6nLDzN48Es4
GOQwDojGokmz7Mc+IqRMBfK4kLCWPsGn6NAHSN4idsoQ37NMHDv2N2GuMW830Gw3S1G42eriX6qJ
lAEU55xfpi8Sf967eb6Co7OWRF7Npc2lzCOIuqHsMgjy+fcAkpYPVlPWxVqNKPUCcZd/5Hvp920h
yjB9b1acCeasabS7YrHIprwNftH3KcWluciW/mfoS2IiSE75Cq5GylkMTqIe3nPY3vTJdPRuC9+7
rLapMbMag4bHsvS8jNy4z7P7fDshGxE8e9Sd8aElw4+FO+c2SFPM8YzWJn4P1kUusZ//q8imfOQr
OVcdOyK5uQdm68MttKS67b6rjClRyMdSNSZH3d4UA24WSUuGvutyepEn1e5X9bfEGqKGWsfJP5Wi
BBKctz2SzPtl0safBaqnAyPlC0r56z1KJ/LtaWTt6cknoE2OsTNVzHc+CkyWbBuDEGWVzL9YErW5
JeTJEEvW6QZHnRXFstqEfRKP+tOA4PKdJnvtInvFlztWMTEGHNSdib/1CI0vWClRDsPXLM0hxWyU
e/yAm2EUbnVcAARHoVPTdIo93FAz8Gul7i1j56a42MwGgGMOq6UM6F4keuGkaQyrs+xL6c0lk7K8
4az2aWy7F4somHaAHw17YMjSVXFqKqgnR7nie39aGdseaq60d9F0ZJy7MKuqU8JEOpdUI7MRE+or
lHhduY5hScjZJDKaZ2xL2ab74O5lrxSYs0GIc+Zl/xyr8Y/9jk0lVIzUb5Ro3WN03ABdCuIjDeHe
V2aLyBZxmqGyrvdJ3aNq3GgiDa3MOwqWZXLo7PPHVOqzm81zKtIl//QpaG1JHAKoysAIL4r0sr2d
ip55AWeW4/O8DgL7v/VFbtT7WR9bg/FR7NodfQLNiTIReJx+5/xRSVYUf8HnEzhF0qG7a63ZAjVK
i53oG4H7pWwJwTUncu2i/E8G8pyPDu7s6beHzrmVB0EzrsoDrf4Ym/BTWtofycTnruZKgb9/qwEH
c+4YxDUCiWZo5SEgUGBtRsq/qO+seLHQ4CNhmFWKFSsewCn4lEUeTmuYqC8NoQB8VyhSDYTN5FPA
EJI4nd3d9/kqaKMS1YjjO6T9Ov/Y63Ob3OqwAG0UFi9hpXhVMusCYobPXCz6AB35o5QwtoRBaBCy
Cjwxhy83p99cCO095sBgTwtF6T63eLS4XmdEtk9p6zdCkBsNgKfhhmfFANWquc2ju4IRhAUMIBPx
+hzfN/Z6m6CxkoImIsYCR8nnSrgeuALQQn3CLD3G+BqW9t/yl/wOw1DoBo9ZNn4lN4rOrBrmPAvk
ZfcavluHvIM737TJafo8cWGy3si5FEgQ+wNXN0qEQlTq9btqp3Ljpd8qJCmz2zXinjzK5QO8p7lv
adQSb3FWKwhxKAESCCHD1zmnxO2jYK4UEybrZheXsPRaPspfOVfhq/0swb5PAU+eIIdcaj4UqBoK
cKTc8e+MfLtRfo/2s1KdCLv/3SEUimApGfWTvXS2TzzXH6N1wXlWvHEtaRVr8P3THbFGIU54LWsd
BUGKq1Ttorygj5bK9InpBmVdspcPREkxmhUj70csHduGmeZeXk55SnvZ11WuieNbJG9s8TeY1sOD
ZDo66ujkoE1oYaycmzTzQhNSdiWlPjM6FuKQnw+EGwokMmYafGmIZx0T/9x2EwCZ7W2ua3gy41xP
roHPEC9v0cN9HiLG9e3pc24x7tVb+FgbhvtSrYZsquxdBYg4ErfqPlMeUKAD2itnDrhAoi14NnfT
6/J6I9BbShXrs/pxfiN6dV71gY1bt8dc2+kCRgkm5w1sQaq0+dTsE96gsuPHGxNbyNdDc3eB82A2
tcn18MOl4tAJCXH3TQGuIgsj3Q7d9sctNOC362nRlZlZPcZSojIQXzRIFcGATyg9ufh3OagbnsfW
gBUE8tAtXjXyVk/QYK2NetaXks/d1TennF9I2Sb0oObpelk0qwAA2RFV6VCBEoe9Qe6HlnxvcsiS
an2m+PbNyikVFZy0Ffk+Xysqfg5IAlU7n3wggFNr7MlNw7lzKMy3wkRGGJUgkoOdLc3qm6wktnpL
aYrbcnwKKdT7/t59QfZQhZTnL/yE7qIGQLyiXwdcTqjTREynRWb7/SvcOVoeDFkO6h4BH0Ymy6bx
eRXel4fF3Du8jcmQ8IsjWVssZeDCD7HFKkP1YHuPD+FI+EkUYmBN3l3SoUWjhmOPSokDckKu8roS
O0d4+uL5tIPDg4kavUHr4r4QBjYQuDLPvSmRKXws3Cmq9GCXWJJGf2LL4w94avtJUKj0pnSG2evI
fhGhMefH3hWfd3esYxyhqeknWx4QGC+XfIOkGN/QvGezeNzT3R5gW5bUSZlRIy3/DWHUXgSQGruh
nHZSx6zJ1YYyC4IMUIYNwa+GVW9VNNmRWfzjvcrlGbYNyNES2sVfHO2RuUXgBTOCAYGgV5p3lWrD
SccfjsIVmWwl18qTEi154CKizMurRnbb2o4JNLx7BHs4z6G/WRYbfzOcvbPzj2N2tQG5yJVK+P6c
2joyBYwWyMbyRw4GLQo/rJ/SMs6QYfAn9BhWmC0i8YlK/807iCxIjUAu7y0ntd9jJHcuCVPe5r+W
wO2E4JmrSbTYzZZ6hcILmfxEYT/hQYU4zTNM/s5ooTWVrsriOM+OGn78hk4srnYDHQ5hAiwYoAfh
kXlAotvpo9lfdVFPzFqR5FJSG1eGjeRTz3MqI+XEDbh0vyg3G/A2bsI0M4mbHHXEWxnxxBY9DwcB
+tMeONbL8zY+nfKm8OwU1FSQYeWnVsMbq2j5LQP/bYFEzKkGbsl+tn1t2hXTmP867NSRv+uTby47
MDT99SUWa0JpRe+I5oe97728n9N5phbPZ0kKZer+kcj707KEk7XvCMBzzHLpA/YuYnnADRH0ec53
64uLcm29BiPLTrKMMcPMOZTaaJfjvAPb430QsijRkpegOr8hGe4syLRt+9QLlSnwQHUyqTzfCd6Z
LGvDi9WG0MuVXHsa7zKzqxr8xeDL2TV2aXbCmmB1dVUBkqjUCMAWT1OU4cUmFnW3amHiAPEn35Zq
T86v77tds9feDy+QrlqXiNjXhvVvIbkuNB9O3/+atWnqILWSSGyMhVLoN30gaA22ZNqw9cmdb000
UmzK1BN6UdBE1c7CvDayrbjfVicBRSdyEOSPUon5O2V5p7CqF72wuo3XBcyWQWEAk0AfwxbnpkTL
ZOruaWQp+VcZxtZV56S//Ju34cDfMhldKkSMObJ15i61EstqalsZ/HtkhkTIxxUrE7f6qBv9NjCG
vCA+SI76FPtQsod7H1aZv79VimN+rltnOsWTqkclbL86+7wfEHY/VY/wYpglsLGTIeHqpnKuABB3
ZdIfq3hffNVzNiufi4KvHNIHjsfqOutImlc0MI1bSg+bnvFD13gjN1vROHz1PCmyGaJgkyOvSVMo
irM3F5iRUIPNWkNASF1jX6ztepvJM9Oz/xCgn9OLFLgJw6nyyu6ra5DBzsRas6aqY1N3uxtqWIIv
LrnQ63a23pA4g+BC/7+b0e4hzvbl5neDgV+XIu4bb/BpNaHnE+lo0I9w/bcQWn9GCzH/ApI+5nRh
gTs+9XGnicp8FyErlez0w5OnRSylP7OSlZD4acIxBS4ctQ6H3YEgYw5M/H9T2chMdTPb7He1WfLN
i++eCMe0j1qcYvE74LmFrO2DW1y8h0CnDLTek/J9D928NsHMdNqnffRg/TJBmnRD4B0OV+R2FxtQ
tr4soBmwHCWSmkM7QMEsaXwa0dLxDEi3ABpxjdCAwvQMRJtxlfPq1s5w0iCHm93dYxHv86JbhbWy
W6zUQd247VjJzhd8LJaBUGMTpKj6V37q9zj3owkxFF/cZQUQuorlG53PLAOQ6DXTrAv6gRknujIf
jYvf7cao8PQerg/tFYB7dv/ZX74Zg3vAFX/jF6xYnl4vqE8ENXW3Epe9OmfEEBpOdGFHu3TqKoZ8
BWAESGplLigvQORstmJkY/hLltJdAb3neNPkndUTp0UE4xCpfwVj+14YVEobvdMpMk2lGRfDYYko
aAezZYBiXbAHINWP2tGV4fd6pURLdJ0GfjRJRNF/QjF38gxM2mgbho4Kx71DRZxhT7aKQCe28QZv
3uVGHMGn9SvtcL3RdjV0iLMHSJx1qsj6DcAQFkUuXyi/pDNol7j/ttXTFZqUhdTp7IFxB1Cea7az
hZs/Utp1O4DsvabhQ8M4HrVJpmFhWrD2Eo/Zd3PKqQ/Rt4sCWzrz9MfTaLF4C8NYP8W9HUCRk8Gr
4OXhOcmVEzyArKAjKMxLkyZKtqeukCoKM3kEDXsgsWot+IY21zWouSkUWun3+jMXjsbcCTnZ48CP
VS8OsYaePZlM/uVQJO5y3ENnGMxHiqxT2ow9upn70kkxH/oIst9BREhl1YLYaZkuAXYOITwtnLLe
H85e3l6AAjl+2fwZLJYWMLum6VqbP3gigXUT85fopgKsfoaSOZqSxMg+UKeKTbGWOKQ5Po7+F2na
Zxa16V8nY2XTdzdScV4eNJ47Dep6E9EAh4KMxE5mF1vbieTar09N3EZ94SLoPOhET6a8lesrK4sX
rSNLLeml31/Foir7jvpQjy+QPogm2NOoemxt0DGY5pXzFPpZttGC5G7mrEodcj07zcdZOhvue11p
JsAkwvz+LJs9NnWm5G0gztUVBrAAqCzgqfGmN3FXPkzZ+o0Q/FO8JH7CEg0v2kofysxlk7rluW18
WU1CvXwuq1hxo90m8cd52vytUXZFSxlOlQOCvLnkcIgk6FGKP9o7s0JsZlC85oA31k6MM7spqtOW
YNZKnxka8YliwxEzOGcCuN4F50byaNVx7JhcpZqrIqcRmsMZoE7GLJ0mxQtleCuhnrX/h7WHwmyz
kFduUFBqD6fy8W3PXWZqdrwzdeM7DBcn/drmyAZpuAKS2zfMFDehJveZM4pQ48OFFB4WYdsf78Dy
PKIHXuBoK6UWwG8LxtxX67dVEyvAed0bFEGpb8EOcAod72YjUo/N/tgE6zPottw7O6MN1fyjBKk9
1jeYCJGPo+33AXK4RaIjHCbsDItgtKpoMnuRbyvYG0GyAJ85NpSr0H3aRLLSkn3tq5L5d0lCJY4H
cEknhoDkgWzYMolyxmm4UO130chG3LhMKIiaNdWOmTVv73dkdVYSP+io0HDXogMvUZDOjc/xiSWt
wUkRK8lc31AuGwWJzMqM5xw8TtwogvxHLwdOpc1YvAH9Aeef4VW9934DRbArZVSuD2LYaiShPfuA
fcq78+GVV/9I4upemzX2gJJtF4tKtDZO0+ZRHieH2Q9VszzFB21wv4IrOgjOo7VPw2e0OVJi/71W
emCX7Kzp9djVWPaU77MvWpDqJtGpCbR0mLGws6Hrrz/SrapTQ0Zzd23jOxboiCjzbcxo+rQYvO5Q
zpUcGecfrlSiOcsQdwK3wkTSe7x2GApo3LKCm69wNxVbXv39EJ8/0VHFy3nob/YNosIdlROp80ve
epMHcYvFx07gTGebpBNNroPF3dLajzxWp9fJ/viPQ9vOkLgSlaeJ+443nKk6oi74I15rPFNgsEjL
te9h6zCbpURjGtIJatq9Sj0MVSuXEZCVBy5bBg/Z0jwMYSAjD3Na9UQZhcrTr61/UZjzyDIpSEj2
nhEucDVg9dyrc6qWiF35zYJxfnKYJl6OyaoZaN7GJyKhbXT1OoVvEITWchn0hPdZVRFM2UMFmS3b
edTEclslMl5mtF4mkPo0Dgmww/8xPxGp8N02Hd8jEam5Hl7Nety7jLJo4ArIpLXImfyaMFbjH0Kq
QhoSMfOQhAp+c+KIsFjXFwqi7Wyqtc8CZme1iA4+dsN0gFOjAdQYOnmTkdbDWzqb2M8p8bUSLU4X
JhITu/8Fa+GdcIN9IPJr3aDumRZP1bZ4UqKbNZ8aT90WMn6YvSujoiyOe5ZwFNgBlGkSS3iESl9N
t1e7kg5VXptwmzzKJ7IHY040fAtkAfq3eNXiJF3TPJ55oQA7GsBDe+snPZRUvHjhf2JOqdzq7CSg
5l/zRXAGoES8rcTMAxDdMnOdGzVsZ/6UcIoE6DB6+bDcyxmr8s7PBV9uYYPLEFS1aKBiA/1nJc1i
cDtaGLZUxV7ggpCiUmWz08KNLARnCRsINk1BiYlUzsszBoqpVWN5lHfOgi6eztzbfxmqiFv0w9xA
PpeRvjpqO8Fkeaxp8+GJkYyWXaWJW8DqjOAqoHJYxAG5Okfi/AXYpB55rgISGqxFcbjew4zzcVFh
BDQe2mSv07006k+FAdnR6RAMoz/kShu/GkoRbxFQ2ZM38KrHPXd/xkw9m1Nfseu3+30NH1LL+p0T
KxCKOWqNrsjBVgrwTzj4xnUS/TBVuGFIkFJk4PLsZxlVLCPXtI2kFtH8YpHoAoBMBbx6CZ7QaPpA
mzdeIzKLP79z47UWnHzmGLXyN0Sz+GPSHKv1LKgmYL6/+sRHttDTYDC0x9D057I3LeloiF7oAsuR
MwhaqsKw+NijpnAWVnsZaLGqoCIpUUVYJHZDaDdtzNbr+BEDBHARIeVI7RLK0nUU8zdrYfTUDdLb
Ef445ngu8QlUAgDOMJM/WkQjjDqrccqKEtfuCQChhIehbhYbWZYLHRvqXMAVMKgzwVvKqOOrNXZb
7PMabWAAacrdYCvKEJtb1hZt5zFfDgu6wvm/2cZecHGR3usolvErEzeE9lOWRNDYakwXS1zQZ7FD
KRqyaiyhF9DjDP7GUeird6LpVSftGUqoRhXehMDbc3oSQwE3tqm046J6T4ogr8LrJZxnM5cRLLFl
16DyCfjTD/klkRWUAiOBDXijsFITma9ygyV8lFM+l5RbEINyqwuLap+DLP8C0wIr62s5cevLBQ2N
BboZbgaMSna7u84ccwceoxK1fhYX27tw6GrjaQSw/39D5q7Ci5mtrcEB2ytnZd+4i2ieOTuotu+9
mkvsAA39wIzmidwbQ8t2D4HLJaeQaObDFVBrzfSpYIRpxBN19YhOHPEzd5DhOZiOVKwwHQHDMCiU
9guSYFngfQXkIAFX4CW8xGpurKoWr9nStaZjNdgOW5ECe42m0Cjn6rNgAfPGBsA6fZYOPJ3A8pl9
TYQfugp+MoFQAoGT+sbfANEevnmhufWVJv2VmOWybqD5w48oykPOcvz0YX+/e/ZSr81ugIsehzio
By7hl0wnXE8yb9Hp3SoMkcQAXPr/+PmLzD9d7762qAIPFo9ykVz/fRlVGUiY1vk6/xu+qfx3KSVw
YjWBz2cYjWGZiAEs9glesPukMDDqis+THSaEFpMRXMI0h31JaOsjqGQbIYFsYlStAU2IwundQ3wk
u7ESUme6b6ZOLH88rwJI8ZUCOTlqTgZldNdOPo9l9E0XusavaTidImPk9Asi+IySktiIpViABE98
IVpuJRCs1x88t8RAsjeMnZT4ONc/FxUCHB92n0WGDkfRAFecp7r6HfxLKEmruhUFJAqr8VR6Awzy
rlpWPyQDnDbGRLFq/0tdlmEs2yg7e5/61NQlNNt/G6trWm0MMk4NxihcYIOyNGGQ048K9LrjCkNb
41lX8rilvNpfGzcRHvLwyawepJVr0QwQn5TlJgbh2unRxZ2ZvOs9bSrq7eK5C1A3lHXoOktcClet
EdiLh7xMoWntGKFB1RLwZJFajl9XMq0GSjPWre+yEIpt1npRsZchRvSyYaXZKy5a6S22rqj7Qx/e
G5CeqxQCB3jEWs/w5pgBRIUfpGQtpBvDbiCZWW9MyiY7J8a0DToEW8Sj9OVjsRXTH+2R5ZhnRn3g
zsGV8JfMrzCWm1Esk5ikVlPS5Uyi4dvc+4MwsX+N0rVSZQw9kmvm8oQJK7cylM7MqE0s2k5QnXyG
6hnL2fJaAqAylVerHQQt7tsDR8KNo3F7V010uE0fAQ1Q+Qw2gyLm6p75PltdK6/eprC7eZL0U0IN
QylEqVuSeP+PEr5+dVSOLDCRU/b7dZXiiy38qCHhU+RgeRe6wL9m3Wb3nXhP0nnkQYy0LbNfQBmo
qsnZcbWWBqBmcy/wc0zj4nIuK91g56HzD/BBjN7e1fylXe7oeYU5EWhKzVnUABjTwh3BNqIiXEQo
iHz1rGHyyrIFiC1RYLMxub6SIRPF7NZLLj88e22JMT58Um5/gDHa/0wniq7HAxHpNiOeix4ueIyr
2mPVOsXRlYAj0SQK3SrMTk1mERhf+zhQ7jAbTL3ftOggAmhKRWVOaX0HYX8ZghoyshLCcvbdkoUv
aNlwRJGm8gk6K2q6FnqK4QqSTamgB0MPaZH8It2Guwr9RZgV+DfU+Mk3RwQ4Zz6Pc4t5UMH8ZQks
2HHqczEaTh8vG5TqjPQQv2ItA70FEAFThi+zrltzJnAvTuUdy4LMSI4XKyGBDM+H6Zrsjd3R90oa
gqj0czStmsVGebxzKYQNZCAAwV6Wzd2G2vg0/qTo1A6yX1sZLpeCrSonnBzcn3WjVEKCin/SR5nh
PPt0Z6Uq/qFCkUIKdeWJsf/wOzRVpt6EMd1GYP95s7NJqJ6Hd2pnPUE6fwoBwxzO7+oN97hujl4Q
9luEhSVTRC0vBVd2x+ZS3QOhZVmpW4BFaBKfGfh5Vzda8ad4PlDDRbEi9NxuiEWgklSLuk8Y0QuM
wWFl2UKwS4+K2xWNhD2cRAhk0g5+u0O4r2JUXN4xA4xlFCmyAHckGDBE/9rzEKmSR0O4hHy4qf5i
UjrinNXfhe8J2Sn1LqWFkPENCRzAwyPtvEOSUnl1APuAtAOtm2CjVyhqtC8EVYBTgucBBe+XmMr5
aNyn5wvr7T8sTgXb6BtVsQ35DZkLAGuABz1Os7+LqzR5xLcmGe7++lcdclNeVQU7is7qJkI5To4G
m55ZraORsqj9W+k/9ACGKHO/SRpr+J35iqTssDVMULeIwtlMNlvvfitG0QxEht2GxW70QuUwC6QQ
2EdlazCFnLc2e7LkEUbQL64TlklZzQTEi/EHqaRMOPtRAd53HAqvmZhURA7xCjVJsTCLTSM6W0SQ
lAt+KyMIyElFt39v7BtA01Hvhn+9fAtY3MTe38mwNkN5MeVCRsAdgA5enAf2+nnjpULJ4/7teyvw
04ZmhSobAIw8385pgptOTvlDSomhfXNCseExNE/lqVkZ9U8ctWcVWBNLPXxI1YN48DWUxVe5CZr+
FzFvqVeMkJdhBvtl6x7CpKjDbRfbN2T9VAavZiHkhHMWeHZtkIABp3oH2VixSdxHh4lFnpI6uEFi
wA/D2p7OaIk00ThP2NnyIEiExIDCVlH35hJXgLIbU09MT9ltcrDe2afqjAC+H+M9d7IhlOs8OqZp
IMROSOzGphRvHIsNLgnQwIGUgDGuqQXdHPM4hBVnTw87yR8WGYbOmLeNSvgJ9eQGuX9iQOKKKnTX
TeFa5QDo9bmwHrxIIbrYyXL+0NIWNplM0DEkm4S4KU8b1rUKT6s2S2PaEwFWk0B/aAIYB/kzhGOp
zNVKJ8rZlN5XH4S+OuFT6m2XHsKoNlkQNDCx9yKx4UBlLX3OPlznUOdkanhRkwX7w2CJPa5vshVC
UPZ99Zjo8FBWtizAbiC30gyhU2kFoePZpLTZ/T4Nuh3PMqz74MtZaWxn9kj4wNcQS6ilHIw8Q8iV
NXpgKq/OYVl77kplqI2RwALRczwMZ0qnRts01aPwTW68l5mMXaD46taIf2X+qKvLYWKvPXrKrzru
jH7mKKwyiDyZptKrbhcxebzwRyqkLuOG93B/TTWyCYdPJhjULSjqP0SEYIByuRQoW1G1yQs8NRJp
pmkNiMSNhvRm2Om5YUfdtsnIWFvADJ4bHRT2bLdGhVv2x4m28YPlCHV42W+x2pVBXL1OTS0TOBRZ
vR2RSO2yyUIg2mALcotf7V3Ml5V058ZdsZ8WCY0OQnrPf0uhoyOCa3dAbRPyn67dWR7pdzDSlxVE
zLdz5byOU2DPGT6nUX4+3CqI0hgzm/BD1creGxzFb63PgipyCujQJZhwJ+lO2caddCrC6t47SUzf
92U4NTCccou0dTfDorPx1lZLLLyklZMvon0oQCcT2mU90p5WVZ8x19nMR+uhhEB7Z4/POB9kkcaK
wQsm6ymMJLW0K4ChFZYE5yzy1jFUuldf7PmrlhPVt3Ln9hT4WhxNQmu1SR7ngDK5GK1aNcPu/g4j
K0A1Md0+dchEfC/jBfKqbCaO+/K0IO+uQu4mxDVdGWuRJINv+Krg6uq8C9ODiqHwlcJdhqLwyG5V
zSJMaDEAOaSHp0X8i3MU9J+HdHeFGxrA8s7cWXZw7WdONof1UZPrYbUCVu6uQGTzyCpP+Gsh4cKk
YOvYJ4dyYRZGoPLpZ3oTl3Lhanx9WkAbHJ2Iyw/MmbzapRzJ+l54V9IrCYocBiXyntrydqcCfy/l
gE4iUEAxT6G9eeO6xW/G75lXJIHyIOxiQYnVTAhJY7ljfLk59VcgVhpgaIbpqd42w+q70hc0kbuD
1ohVRCD7I3zefFgocpRToHDhp6sTf8ViWVSsgxmI5YA+ZoVi7Te/5PoaztEGhSqP/fawbo+ufYQE
6rL2k/AV0t5ONSc40UCi8cAP51LTNjLc+/HWq4NsoEw0xPV1SYLb9Moh+dTXvIjfC8sU+ujoPlV8
Vk2xgHeAndn/ZPo65PArE2K1By/nFr1u4mt0sLxq5rP/iKZatCdB6y2NISprUsiaC5JkY1sVCaL5
1DYFjpPZiHODmkLnPXcWWnPYZQzyRj1Eeu1pqaTOpi6YBopiLXEQxwre6tfcXSaX25hWMEVw9JRD
hyWwNHS75z4tH6fhNGeXftAqEUD4bhxeFDgl0mZw7oGS/UtnEoSai+UYMC4AnsZOqTZP8al8AILb
hFEg8ng1crwJHGyaFskkMX2N2Wn+11xBm0FY3YMVXcsp5zS9WpZ3nGduHQ6ZM+TjV68nspzx7o7D
HZg/22HBxoLz8RPNelBtp+azlpKTngTAxvxgZ8KrxRwZaUKezqUn/Hsn7OsgIz/2ZXqQKYfjK/UV
T2unjXVPaQa6jCzkLIMDIM8OMzVl6ZSkagE6E4NhCUA/IowUYjTIywm6+mLLxj4y3aycw8v+Jpep
23gh75TfNLRugWPfz6E6PkAsnScGIZ/mukSJwcMYZanFhq/FCS041yH2vwMe5AUAE/NrFtHGF1sw
Of8JF6VONeIWX/vKao1rk9EXJg5qwgodr8gXMGy55TDNkO28xivHjTWT7RmNh3Koun89maHj/5DR
cptqFhUgTDktCKR/73jo1Y+HL9ezOyfkgNgogCvTvWA8tHE5mwQBB6y7GoUUdwSed3acF/RXXzTL
ihPgjG6PRSrWSGXWVzgbtGscFCxkU2Yg68kEzjYfygvSyA/M7DkCRM73pz6lxFVV6pjdtLvRnxmO
mGiDtPUqOvdXljl/gMyt3aX9WLBKbqlysJQPv4lzJNXZpdqqMlUZUlVRitWX8mrbVbe01ETzjBoJ
NYLSKlrfrXyUcvydY5xGmwUUHUPiAHazoHdfvDYm1Kd7tsFhliqA7d1bnxEEn2VqLnIq/3QHnBka
ab9Mv8BQc3YcRWGcR2WIJoSHfoNTsQvDwGn0z1AQeuFDBbHVIMtBOUb5aG8FXJkN/2EjvV/6n2+H
CmhP1mDYAn+qoFA0myRUpLF23FSOz2ndxVN1pj/U+R3/8pSfl5MzA3fG28twucZeI6ZPQOw44Ts9
rOhnwi9uzLoSl3M9s9jkKGLI5hT2Lo3h/IEWady2g7Nw5Q4wq3Uw5HJFJVPbxXuT8GxUhIaJEmmB
VeFIu19CNltoWNH3mZxH1yuYNOfxTcg5UwFESQUWR7nrBSlOJRFcvVxt+BEALipa+eHhNw144Bvo
aaDsq6Uxb/SoCcp0RLFrurryc2oKearitA4LJBQNg7ZrVa5irGYj1ucG4OZBV84Og+Y41J1fjW3E
r1GVOUOxi0P+tDCbg/bM5ynwESHRwZRc2tnBM7kq9dY5F1csx0NhRtz21NpP4LYDkKqTYLzWAXEB
832DJurJx3RP1ci5kqBNHxmfpmFbm1x72P1DYJft+5ipk3K+KHUcANcyK7ozhSqLdJdtPYjfb558
8/FRaPCffPYf8ZKIXGLKprlROthRVAl5E/pXGZhpEB3lhW0ko6evVBB474Pa9txMQbmvGjAhnCS3
azpPqNYCqRh8dfb5GDembQSgKAgkepcwacYeKCCyX1zPluSFOpySsWa3l85/6nj1WjGNXKwTcWon
YHJkRZA6NC2WjpGShe+EeS0/2kZxchRtYPXrbTlvRKDlTwYZU8rVU6lQUUajpQFMGSo/tkFWr6tz
DUzWMdDFZiRX/LXXQYjY6rNl7/1ZRsvZAMqfu8Mv7OOU0JbcQjAzgOEyibq1KqhGuXvfQL/nEwA7
c4qTc1Ojejiysb2U47YMh0f5pPJF571sVh8z1f+pdGquDtyWKeV3Zkds0KdD4MwCsM0Cku+/zVBr
GZ/+hSp/ULjwYdyY5GOFs8uacvrr4MVEtca2qSLfGZdKoUbPxTnuG+cS5BczXLudF4Gbo76Z8ztx
b7Vu0A5Y/814rsyvd+qqbYuBTsn09SQ95wZWBJNH8WN7knVxfYcjPtzW8sP4IJpeflCEIMpoBuc6
zWcJaTcZiTxC4qHyvKJ9ePS++y5z6hHI1Ke0laQygunr9PFBE07b/PWAX4JkafqyaFxM93TjZkV8
HERR7rTmWxRFXdEIUPV3ULnYMZ14dO4FeKizHxD64kbCxt3ouAqKH1gfNFOiK7JbGRFvimdffqn0
TnQ+fT6x4doyTXZaqkbzEgNOBPb+vUGMvlsxhp9lqVfNfKovCJdlbM8e2/S1NWhZv2PeHHnSh+4h
0zTNVMH87TBKlYi3P31Ongyk77w/jiEWb3qDdrxlaKyDpRoulioDM1tVA+5vrLvWFb0rlS8WI+SV
i+PoxFJD2kDxYX2flh866YNWzifr6J/oJTjHNMX+Oi9+LNOexln2bwUV+1Fqy3IleRhKBJsLA2BZ
Qy+LPZuKZb0IVTlyGX6Dg/swBiTeNBERq7vFjxoAqRei8sGwvhe28GeVDhyjLny3VUxOuJJTo0fC
TwdyI6rOmC1w9Ij/ZyDWPeO5+i+lt7X4V0MYhNjhdXvXnUMqFGBMVoWm0YORIoRJsmp3lYtoOIlz
+vrIGt4Siy07A+PZmGbX4iVmJoKVtA4HBD4pXse/lpujy8L+9M93kzGLnojZmyzsRICCQURIReHa
GpXKG4AfkjKMBum5T6OvRH2EukuM0oN+Fa04KuxVZFHqv095Nn3qkFZ8pp0/uX0NLsPcwkdeXhzh
xv/sHvXmM4w+RBvA19veVfMCfdxZm+EqeJ2kxQjADUbnG0f6U6vKvm3Q4doJG2E/EN9+EezEVRVW
7G2XS9LMgjSBkIdXITFRvvpp2bR1Rm1shM7zFnEz+ofMaUE/OJwjcmj8JWDtEOD4VqJlpfVrBqZU
xEaxC6hW4wpzxoXY7o/SsQn8YdqX4qVWFy677lVap2PTNnmbXRFQZf+6dgVQujFPRhNw/TqGrfTP
XA5gUrjCaGYq86dHBJfxh0RfjRbkqbgCaye26I3tx4+Biu5XbL1WtzVTnm1WxLhxN70ExSGaocpS
AXIKxwmS59BSxsqhGD70n8ucKQDlD8UQtjUCZDIlte0lPPMbyVsL9ndque/1wL3vYYFVlcXaP6PJ
GkYOlW9bZHZ5iPZvq6smwr0rSK5sFoNYA5w1TBElf2dsRcpu5Vrhx1YxyIX27/mJzt1Pzts9XSRu
SdUsKGfOnqOXH9TbaWZWKZrQovnbscw0PfzbAWkhehY=
`protect end_protected
