-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e51R3r27nWx3C/o/bxF0sex1M5dADsss6TQlv2CQD8u2eU2oWEm6l/+0FnroUgTf5hiBUsLr26wA
26jDx+Cog2G/y0f3//hazT7udqrIRZsbjXPZv8gL3p6I5Vy8syGuPsJfwrFvqFeWer1mzbQECx7K
CiBhHu67QRyrxT/jmm5tvK2llmZ/zJ4uaiOaJh71xmBc7GKB7A02dYMlcsA0BBK+whQCzS9x+eqf
1f2MmNe5xguEBejGpPsmmN7WSV/wiH+WRyzT9uclwQl/nLrG2Dqgt3E8kZob7ixo02QyNBtrHhmN
zVQC31FmDa++gtaBFdg2e5ZZ6iUCIjm6MYYWxQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
3UcKyA9aLgH+Q2r/nx96/1kQHQ90OoRjmI02yupCd0cLyGjB0XbF3hfMJt39JOc/YUexTBOFMREZ
sFjIc39uJ+P5XnY72BbxKhjQ1J1uXomclnqjc2s9Mg9hswmKFhkWR0/vR41/0a0IMC7CVvgk78Kf
M/LjRYtmtX+Yj0q+i7Lj49qNTNIv8Fu56wPBcAaB3BPo1jQuQjvLGHJ/YuVwItNNSdFduOYw/qhS
wdoSqe9JXRUBYZ0ZNc7bqqLW7jHap6eoZO4zCxBBWu3ugorPD0hYR9+mrWx98XGLG6mhLIdxnpVg
53fTosCDfp91sCHQhvxgGsV8+DOn0keTFZ07bm91jm8sEvenBjAm+Cy71asH+x82ZNNmZcSSuwTB
rPPC+GZCB9GxBfR9u1yLWXMiYHgJYoiphTfBLASg5BjoQQRebAgy8r3ntHcgyf/Z6I5gCcuvNS47
ucLo3U4H4sMUF1aLh2DbDZStgOPgX0E/k1uTzJm7TSRjNnBMG0PrE+MLKLorRMhoZ+t79l2VyZO6
rKxV+Vjgli3JLLuzQQ1tK3brdPhU9iExJcU0EIuskFT9C3aia/X70pgCPdoS9InSV8LmJV4Vfp4A
agm5ojbM31BPje24PbNHxVYMcTjrEcWtI5OoZkWfHDIP0T3p9jAn8Fm6Lym4Kx3LGnOBiM5foB5S
o/+uMGka69HCMvRSR072jIDc4n/jSB2sdlxhaXu4BnztlKekFGZZlJuUrziz66B5zQJMsWRTJeRb
LZVyErq7stGQq+kJcQ1xn4szbXY50F3FfxfD5Qo6m+bIM5/isCZt1UZVliMKGe11GBtS+w1xIOSt
izkyLNGc82Tn9qjlwcfM1JTPM3Ml7DtZaacg8cuNjl0AgoIgK3UQX+3mRV7oTeJ0Oy6R6C5drIbz
Hpni7c16ELMj2tvwiSx1bNrw9HOJ8fKydrtlaaejYaJwlznyCvFkdtOP/JI0vg9NAct4f5qMRH5h
J4EGztFB5xexVMM4kAno125pmLxycNB1QM6B0mRe9ViTevU3bRynslxZSXkRUAZlar6G1XV4364s
3THHBQkgGmWnB6U2JYRLwLEjtUqxagAU/C1LFiCZ0CpRUv6r73IopXXnhIp1twFuL3x4VStucyLn
7kZcAh0zjg8bzoNjlI0F1cYgIeINspC2PP2SuCjmlMSO567Mlx3hG+9X+QK9qdZleL1QAt3PBxS9
QfgRpETmr8zFfhZvDtnRvdjSb9vvP2ZxyIXbyUfDJdO/UgRr3NPp6Sbkuc6rkQbDNoZzXvikuk34
gSzhfkdgRrCS2y3l7Kn/6XisDuAnIzTvK8TtRd9q4pH8OjdwD2fQGOZ2I/vC1KKaSKsW/VBJVCX7
VvgVhgUOr7cR/Pk9dDrCH7cPscF2fbldyQrt6Qkz7wz+rYEhMcDR4S4dv8GJSP+c38h/nGs8KLWP
ck06wN+AvexS2DeYoUMAcIxO03buP7PFz+P2XUrfAfu5Iy+pIlZd7OsKWf7+rdhxfl7nXCBmI9JW
EKBv0SHby8V6U41luRx4r+CWXh11/XmlkGG2SUTmCQOrIHUhh7Jul81wT3Z61FvcWWQgN7W0/2mP
jcix+MV5LiPoDGjp1QDiemGQDwBI+Hw+etfYDGO3Vk1bw/7wtybBgMHxRoJTR7O9mj03lcPsoUC3
8XyZz0cR1fYY6VjqPcl1ZgkhETASt5KuEliyDZdNqetC1rl5Pf1MtZYey7+4LHuCoiP0MZIxrVlX
oT0wGX9cAWvj7B0aTD4hIEt4YCFf2rZfH8f768bLgB2r+rJ4WoiuMlaEEJumAqkrjJ3rMeJhSy6h
EJpp5ULVUU+Pit37tohC19KLeBVjn8qehi1CeuIVtVsaFTdnD87YrbBq5WS+GD5fz9Q8j3Vf5NLO
H9qZpEHZEuqAs+4xa1FHoH8dp8WmMssdl7PRoo3NPHUZwzsYbTBIq8mrExQ/U/z0UBTS/aW3wTtq
r7pLMPDh4k+qPcrwGQX/3ityz5NsZnJLyKuJYhff/ef9Fk40o5LVoaC+/OqTqAYYYjIZMsVj/MqB
QEqY6qE3pgQF0p649UQmRuVsCNK7kE7ysz9FETOFGO/j/Kyi48YH6vo0q9evk1ToOlkPiCJPv9gU
YfwcwNKfFbDmDWuCvEG834bga4PpL7ldTzMX44zkgaENJ9MAuygL9MNg338ZUgdE0lZ0d5s3KrBh
7CPIIEV6AhR0POvwT4n3LAa61DnrvXVCjiBSqxZnSj0NGvysxdYD3scwAZSVJNsO7qbHFmVb9HIT
PbVw7Z7p9CJM2DV7EDX5YcC7CwCf3xfLddZDsff6mo0gOjRcD8cMqUzOjh69QWcRkTCWIwZjH219
+mMwomHohdWJP/Hz55NZOccalIejz+K4/vLU2XeAcIt+TAKcPdsDzRJwW8JsAk56IhqH/lj38czt
0w3O6A1S0W55JrIhwzYsJlLVwi29G77Xd3wj6TniFn/M1v3IMXFGmBjXU4mDFxT8jJSQOgmxt87a
5aoPWtmsj4bpMHRbzAGHcX9N8QtviSBmobX0XgwZLApgVfJVRwF7F/VrOhQcrTJAfg2h324BraMK
isixm+Zxun4ErP3fXfb0W5cfvNxJbfI0eIe3PDZvbdPRrdQeV6to3J6Q3Bu/oTFIAG+aWsa48dgL
UHMno44mvHdCjA2FLRE6DRWYJP7waGZlQXHA2WHg4aMUlvaXpw5xcxdik20mgxeM1b3h2o2e7aj0
DOo4joe4e7FzGIBlTwtUMoXNlTMv55x8q+YoaCRhyEK+iZPbv0PbHrW2Qm332dqnkZdWOCSlLxOy
l9cbbyD+C44t7MpTgg0YMH+z91vWIpLQ325kFgY491d90zR52uF63wYm/aY9B5ZXpmlqW4CIzoO7
P2AY7/UWj668kJRRvYeMIghkpwikTsVmJqU7H9V/+G9pNUnNlFgeQWkqrFgrePM3gQAuWVQTVFvT
alS02otVqeOTXjqLzPvB4rtVeMA6ebU/olW50EHOUYydSE+v3rqj7ovX/hlol12BcAi+q9AEPDwd
lFFKdFoZOvv9tD48RTNGIvvV1D+2ARUg2miwoDy9MhFyUtruKqPtty0f13UhrapAfDI9ubijSZoM
xuf+QChFj2twr5bszONWKaImpbq3z6T+uLT9vrwM6xDsoDFbQP1InZuLbPKRivjDL1gnpxg8lzTR
oH9TBDZZi60oChvN+dhbJ1iyX1+KJaJH2nD8/+VpWHAzWwphwuZex1ZORS6OdB2UNcNxrKXMcx4n
fHW32vY8npjyWmBVrwCbe2XIkCaspxi2HZdxzPbb3AlTAgV57sh5uPClVshBmgpVMd9NIb7TxH+I
fhp0ppFYuB7GCysKCBh7nmFSazjj/WUZ+I00dgDKEOX52WbilrbK+XFdibUJpUjVt8CyyEA9fkP1
J4wD57o2k1hbc1ODAW+la/z+1LfA7X03YGejGDmXjOM5azPj3sy4e98xMWRZpNcUNQVRl3QlrTUq
I5IgkdH883sf6AnWG6ngq/pgv/4sE7xgssnsisAZ8VYOdKvlWYJK3x0wvWkk+ocPQqGzi3MeJZ0K
t1b2BhwVbmKcgTDaNtex5Yg/Yq4y1BdeZgCwarQcDF00gZwryGphLNVlHctB5rvMg8Odo1aEmWSO
KlUbvgkjx4Dql84zMVmJvZ+/O1JWqygYH2LkhEodeMIfd3E8IqaO6LOUAo0wc58OaO4QuUcfk9m/
f8Ghn9FoMpYmGPHXs3ClDpVG2DjtNASTP7PODBb8VxwyFXaujFNKp2v/vQsTwDHEgt0k7uYrGm+Z
VJruH4mk36fzET30MmwGJx6XrBV/GeNti/npO24f0jCwW4v8BnwEkUx1CNvtj5kqsm0gJaC9aNlH
DR+z8chg3UUEh3doGQrKDCxAod5f19x6aXmmh+XGQQxry7XsdYgzBciRYd85E0vwkzN35I7xLizT
W07MbE6sPMItrVXTObLlZH44V1ALmvWG/g0ynkkclHUHSM0H1tfxhjt75i/MP1tubaEdwHd7G+1J
ieb5yvepKmYyEcZktFh5pLpUoQNTcP1oh7Jo7d6k+GIFKJg9dwNhM4+AYHAED+8y393wkBV8IVtB
F92S74Eb7MCth2wNDjQ+EutvOrtOlUSzZi4wWkC6RM0+msMwCBQy4lLO/1mXJKxzRl1h+r0DCWX2
8reF7qsQZBvcflOUUXbqscNx9YjNCEq2SoemNU/rg8OTjSuQAPfabd/1bIzyPcnA6x5AeffKIsy7
JSBbYtFSQcWuAuXWpwfztvE8oKlu4cEGx3vg8Vvi9+ThkjvmUqyHHQrYWHrGMlTryKTDqVTuzfsH
C9F3Rf0u0wo2zQ0wFDkHVtJA6Nuf97RcGqPoMBWzaWYvVoOyPmYOKWg8RtToaJ4BSJwTUQPVfMYb
85eN1JOsxqGgQ51LBZmbPEQo30WlQfy0YUyBy02DY4SYMIXd07BTcM6AE6QcTLOIiEdtg4tATtFO
JMEoeRwotwIDZsYY6zGKJwimscKl6uXKY4chqhbbS+FaqFXyAHQ/cP1Yau1VTm2ODPSSgJUodZ8V
bcgTrHDJxjsLDRDJaSWN4ipVuf6DNMwrY5xpZEMn1oyOFBYnN40+RvokO19CMGwAu1Q0vA4SXdTP
TdOjcZGTOgPNDlyL5qfiLTdcCR1HYGSchQ0PWozWNm82oYpZ/ydacpBRlRNLMnybGdlMtklLqPeH
d/q5sBL+/TciEA6zfCz+FTVdWkbg79EIAUyG5eofSB0LVEpQiPI4/74r2tNQqyH5DzlD1cLTywkJ
xOtW6+MIW966Uw09ktyuQvcT8noOQ5cg4hs4hoqrkVTZjtNOhFsAswWy7LzZSiu+ZA+GX5BDn9mU
zUOptQ31QXvyeyAa54k+DgF0TB2k4fHhZCaq9IY600vxZeOCMGheKxczjbXNPcvU5WE8Nmg9dSQL
T26IGIskkItJLpJ/75DJgPGWOX8gypovTXMxR8XfuBkg7Ae6h6/yXsmnX8hToYw/OXUnKbFMdzvQ
EWMS3ENtOJK083oWv+rcK4EeOU0ycASVSNwlL1ekNnYALyFh6Yfap5yrNl3McQg3q+nC5xxlB3Fh
B8WjZbDvQYR+zZuQsyDMK2atE71g9Z4UAjB7Qf7aB7ME0vEYQQIOdxaBZJj5jcrnbjZ6/KBIvvTy
IFjWXEXCiIw7kT018xOjYXvnKbsatOCWQ3DWgDAEzTiam5BG+ujHU3mgkG9X2HrI4SwOw/gPvj8y
dMoNIzVQujyHuAlSukz+pRuN3L97JiOXZg1eWdZqziK8GbknD5sSyd3ZVAzd2BNz0Ifl2M20CRKQ
um7wb8BFcJ8o1i55gjOsawvNyxJC2TRBUUEXX+iPqjFYBYjszljuF9cu8ImORkKXQXSHt4TKx3Sw
hC3s6kPJzCU5j0NefFFo8ZDixzvt8aGqqRaqs4DD1Pf4bEZfo+05cz/Hh2UjjDqOn1Jdzw9UkhjL
Ey18DsEH3J54rf5fM0hFfFFZMsSV+R7be75n9c0nJ2WmDSAKddHsfF2kWZunhlISjSuPbgYbO3RJ
vURwpeoAUxAdk9aQIOK6Rsic9Shikmz5MrcWQYz2FNFH3LWXOPe0g2MaNofeSnF8026fNFxgcXr1
H5wg0kJ92Y1hYxJ5ptj8UMsKl26fEQMviNSjaGnF5XiE+ZItM0xfCJuWOLHETm7v8Bn3KB+mRhse
xUBeM147YYxQ4eG/j/r1WGxFcIc3LFPRX5fCzkdNepRJrHWO5e1ax0YJxhCb6x9QB4kCm4mC6NKl
FBQdW3LQiTcLoiai2VobwDtTkutlAoFjNLoomm6bsejjKjOEq8uX4dvfeJMiKAs+lx4jJyrqIcxy
gaWj82szWS1NEWsIZ8BHAKd5rnXerLRq53etDfjOf4DKyBiJFExAZL3Qn46eWl+G+Ch5unfpw0nA
80FXiugrkt2GmOWpw+am8V+MRkLaaID+r2sBDWLEeND2UaeEHU0WLVtRlcFscL/LARqZYfYtKLFb
9TeECCToBCBAG+4hAyZbF+hiUs7HF/4PbXY9o9LToN+pgaUtphImxpg3ti9YwcRADkqk6SnGnKYi
LhwFH4XgnJyvAdJEBKN0u3NPebKu9wldioyjaMbswX6Je5ghMBKo1mF194Au96aJuOTMSyKge62x
mtxCvYXG6bW8azNcD/16+uW/CPRL/7MZvz4EPmvd7PRjsnD4qzXmRv2cGHyMqbB1Qx63xtFbwIgZ
bpKjzRlyH9c+46mIHgNsAQWT5KJdmgFrkw9GfqXP7gYkQXHCjotsJl8dJZzz1ruwBB7GHLaQDZzD
YiVuf6ImpGQbr1mr4bLG8sBXFAqbQay3RPM76ifQSxnYuP6wmS7V+XGTiB3yQ8HvN9+u8+WSxm7E
U/Uy9Vx4ryfATjGVOGRZE4dU+N63MWfVu0Rhyn9InJ9bWiWAfQQ/2wWqJMFoY6aORS4tKXkC53G5
7uLExUgOVv/v80RmT2gaQMNEhit2/PD8KlzQHVUFJmwXb7u2M8G3owy1ZSoVCuvQC1CUFC3KEkya
4AABOCZubHw8OYNqV+1eUMslw6JyUW2btpGDP3DYOtLS8Tc9CtAtuBD7vPLaM5gPi1ktjjN5HFVI
6lMKFeVY6QasllM8CTQsqrS7XgNAV7s+C18lIbJmyfl+ox2SKtW7/8CM0RcNl+LNHAycixp1YWgQ
6wlYSTPDiRLoV2McpFxG2dr4jWmrUDfF/IB9ljGkpnXp6jglV/aUevksSaRetLYIVAEO6HoQomyg
qHkIok619al0+zVZOUNCRaNhsX/NuQQh2RkhruqgHikDXmKopzgU3Qa3928zjQmg+BBQn52X/mgn
V6t3SeUJDPNsbiFtUZnMg1RGK6kuaYg+mzUqeOnmE4HchmuTk56xldHRzj7wxPAFeycnSnZ3u6FX
OSt30fVX/yhiqhfhAiMT8qGka7UAXBH5I2VlGEF4FnIMr9srFeTvy9ZuIcmzHn2N9rQ6c41Th9+t
0KC2D6GMSbgxC8uh1jifK/SIiskxg/IxwKvEJ+4xNgcXb2mZyX4wB0ELvigzdXho0h8AfozVDs4K
tt+B4OR6UNny6wFFqNJFivQYtVC28arChCfEvZ21LC8fSFEZTsqhA1jk0T62SecgUgpX+IhnsfsY
MZaNflfkENE9mCWC60QTyqjjVqPStAdHSVf+m7q5j+7nNpCDY+0KaCrp3yq52u2DTZjcjNK55B/a
BqZd9SNheWDea3CUYX+Wjy8NhmD82LmSvmnmTfeyQbfPXDyoQ1uIA6PZMIvVo+y0Iu58xR+fGFFy
L02UzLjNLfVzfyiYLOuxE7I/XA3EZnQA/ChOYntHc8eF7b47RbuTuZwTBrJsxT8KoVzFrZGhKGnZ
vGoseuc0M8/PHFh23Isgyuf3mwR1m6CgPcp7YPPwFcQBzuD2dLFR1DSQMKLXNCz6lyl8ZfeplonO
PTtEgG+tLE1HZP9Y/uL6RIAua98AVNJJisLKgv0rbuXNS3jtCQx+me9qlfiyECInPGBG+GIA7W4X
4oEt32saZ0Ts/WRlzmEuwlPLVeJfc9asA3Olm7hQBnaOSroGayuILyn+jLLOjO+k6l0IdQeUJmlH
iGrh8a2dHG/qWJNQxGfhysWAmZCW5+rpMmJ3OWg0TTf9TrOmw8bvf4bjHTV2XI8AtJG7NosFGGhL
FlR24Hf+iDHzS3+F2LMvm21aSuwg70esA+MhXjIWg4V4jqCQ33KDweKxqTP1MNSTEdwV4UBnBul/
Vz71KnhGiwqwz7VQ0y0R72lUxESNtliKfMz6YJamyAXMBse3wppKCqqc5An/PVifGHeiWjuIEIKh
mDYaX/4Hx+dereLVd6Emd9dGuzBKAfmLPvnnK3FtybgoGbl96dxR0EIqxcg81xdq1sdhd4c6ZhM8
hDEL4M4pI42YMnyq6SJ9MpH8toEXmHm8G+8nLPjGIj7uC/kYCU4xHi0AtlZa5ZZd+JRV7IpmMev4
jMmwKenanCJtoW+HA0ySgrZJZz2XTF7+hxJkvs5ijT2N3XYJlLUhlo75bMSPUrmaF8eCf24DnT0B
qsikVUO9Fd01yH3TlrkiQYPqxCdRlNh/qRIH3hgvKQRBJSyraIuGVqtSo9YeM/PnpLjBJPJNUKQF
axxF92tHgQd2uuw9UjECUXp1GeGhK1KWkmkgabOPk8sPS77I7mNPdTnUuYGPCHqRfMFUBRt12TnH
GpiQj6TL2uMQlhXMEFmv8O4aDQsgRGNv7hDEyZVJ+HWb1OdNVf+5eD6C0lwxF1DCKF9nEwI7R0Al
BiVj992YlDGDMV4X2XwYkNrVPROakzBS9hnNGd1ZRwcFXwnszimsAixFchoKg2go9tCbVSkmo3/7
Nr9sSEVspaioqs3Id99Fxc7V8d6mFaust9ipVCyRaLR9muzszVOZ3kFxtEdLsN5jy8DTk9Mebm9L
kCfDDMH0jG1soN0lvUrmM8w2ncB8zuHSE80fxAqJUD1/f0d9g2qHq2yv+6InPKUp8IEb7kQpCkdp
6Xhgjub6Gpa4jMnvJR5KJtNu0wOWPl3flHrG9vKhobP0G/sCtEDkCx88aDT7M6rCvyrE8vAYoLbt
+hKQ/5tPXMywjS/JZYEhnNnwXhTIvGiLae36OkzBu7sRjBkmCYXglKV+cu3/lsehMpA8xPYFwMk5
ShP4SM1ac13mNLslYfs628Vv0TnEe5s3qFBDtRMU4FqMtfLdqnZCWFUlcenZRRFQ3TALyf+S2/Bq
99C2dOkqmurCB9XEGSvPidpKoIjMQnWY5ecqCHZEw9SgMGPV0zk2KOjYHJvg1UDpSxbvbXrMJyWB
aoR2LJZNWG2HjaNad8Tp2p4TExg4SJP29vlcsOkrOJ/000/fqodyWu81l6TN2GUxPL9KicBKZyjk
Wh82quT/S73l8CDPVSsYwiUEvME7HqLtvQQP6B4BFU2Wiwegrw93SwkP5nNbUzibnln05iBZjjgy
QllK+U9DN5t1BipnHKTyESXo0r4j79aE6WN5SaA2GOnUvITJ3gwQNG4lluOmKbnlTenqJNRFYLSp
HDeUze0o8gGjkJ0+Y99WGVsj0J/3eLwGuu8sJNnxE2+czUD7tLTGQkrpis+yisKgtDzrcWQDhCnW
2t9DgyTn43PumyokK5cPBHrVO6TjPl2XXkRw2u1ICRovyuxjRRnF1e0xusV4BaC/yyssK50jtxgR
iAaVubu37KEIDRHY4bEGbMeGf0Z5JzMh8kwwgO4yXYLRmg1GoCdVU3jbXNsb8GiSDvj9EqWU06TB
8wT+INa0zbG23FZH3kFtbAEEdia4N4GV3Qj4utL+ryj8EP2NuxvSVhWbdhcqR0LoO3SlPhzcGZmy
LCam0XP0J+LL7ejPxf5P0AlWseUrNj+Gw48vcP4m+fW9dr3Iwyfz3aPbW0HZZsYu2N3PgbjXdvHm
2jIqHQGL0vLFy+kf3fvYYqbfwe4mN/rikQaW2u6n8ZQaq7SWdyT7AeSIQ3ig38ncVwb5Vfy+ixS2
EAVanh2vXS81D7fJnEQvBgf/meY6RkYTYIEORnnxb6q1XUJrR4aoJFSuiHzfGgQ8E0hrBRJU1XYd
3kehJGRGCi0AHq0LJy50oJL7Iu3LgRhuinS63f2cjJZmnJfXlSYqw2Y0ts03S8uvSzi1nkoeDKPR
tiAxoGoYEu5Iqap6hJqxPA4p98bHvgX52j31O25aEh4WqNg9r7LthnBHyFb0N2H4rxvdsXrQczoK
eA+9C+EcbVl2RbJ2qg3nXrFtxbv+27k+Yaj+/l9bW2+In1JO+JDaJdOthfWzd+vSfLISB3MOo9/z
92lwL+o4bkZWkRwl0U+VTlLCEIKt490UvtcJu2b2VQqVC1jbrPbzjCsKTglHpPnkh2s+OMjvT1ma
AiVdRiQ16jzBQ+l45+s4t7F//MZEFzwwujomzQKBl9jAp1J9tpa1NuEN+L4MkMJNK2373RCl+mai
pwkUBc8+DT74Nl6xbgeVAQDjQXWfmXhgQpSWwGDgpWzQa+rJwIGbCKmmu3lm75ZPHngOWgM=
`protect end_protected
