-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M3/WtiEUOqVm2mDEUlqXn2eeoH/mME7Wh8akpWWwf3cxBdngF0IRMECKPWUyChGXL6kF/+m4LVA7
QNd7c3ws4SJay1qyjtwqmYnS7xibFLaWsVu75GuOMkR6AkWvPT28meJoXZcZlgCkiWu1s9iiL7r6
/2Cy/gkf4oq18ugS+yHbHYdnLaIOGgWi8MRDbBcfhf0m/Fhhrw2kXyq1ZRaQDDRiZ2D5HWuzl/Y6
DGxNmOtkbpZeZiwvsX5GiU8UTwxh14Xw2qWJEeBAtdVAEwP6roRqeyAASox1eY3bek8YtmVaFnRX
Ss7HJZ3071abfGWMveA4RvbSpYaFyp2OLzPZcw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23888)
`protect data_block
feCEHK+CT5ZI/CvRBvyzPK54NjzSgVw+ZGIAAcydRRWEOLD/uwtswn4ZfeOYBP2JULdpGQMeV98+
fDrhQlZjsdIp5b+Ed3HCkYHszIkjryvRY1VSG9Vzv3hoj6OY284XSdG7oldx3lcIIPtR+SAxdAWC
GmDJDiSzfqpCJUVY7tvPvi7ruYM7vP23CDrdrbkEJaWXOmo3RCXF07zNHu1cf+n4fXNpBo5IG/9G
bArxO7vAOPzExc5+0nP8hQ7Zc8VXG4GrAqXXs4wTRzT80o1FBU0NzY7/NBzzyrlRYtq6TNuKg1CV
cu5XuXdE+F6GkJHEKf92gDgE7yY7Jg6CC6sgU/OCeXCTcuiaetkKmUyrwF7RxKQTSu1FfX86Mksn
L2Fu9nuvpR4MQ3+dlwqsEGvu5gHNN0bgEfY/NkkXgMTar9LgSbayKmH2CWK6vTOlQ1vUWfmONeIR
N/Do/aNFly2aItBTuNxrSki99j9ZyP+xx7Tjn9OabgUddTP4sSg3wpf2HXmbLDlL9jRc9d+XdRkS
UTKkwAQPJkcEgYjF4jp+QUFoQWDeCCtMXAEZebgLGSeOfg8VrZpleK1HIgYEwOyJ7jswbMzfOsP/
mUOANSvICIWDjjnD7037IZ0uII0BGAuR9UZeqMZC9sJzBruSVdMZkz466McYyhJS32dHwXnSWpST
bLuLZFOZ/VRlpJW/WuX1vOiz+wwqabTvCy5sB7ffHXl5j/7FJlLFbkPQzmh6aXfvBmz1XQK35vh6
Ua1qRBPB8k7b2LF6/6q0ddf8oU3TyrB/h3UJqrWazd4sw1WJEMp0dWKoeYKNYCip+Lz8BPFT6kNE
22oEAIXYRXTS7SYKJp3qAQ5JmbYMJeyp40a1B2jo+GmXvAxTEXXaery46mjQLdFK2J+xdGVXzt5n
W24/gMY5sx3dJDxXy7xulPhTa81at+lpToQiRmnTmLNux4eqCCwR38K4ARYGetd61WexjzCeluEF
q1j2N2QpKo2vxPH7YUOHYFYI236I9NlSj6unPpYK1tL5r0ZOzPP6H4VZAl+2/09f1lVOGrekz99b
nQ9TtEaxOvRDge9fjbS+GUpBrcHawH93GYYQ6XCCRKFVArrJt1u63SwR8iOTOTyiZkSYtUYRmVb3
9+SuGUKDOC39nyIwAfDFfYNVb6YcgOv0rQxow2RCWkxicTE8hOdKW7gr9fkmddmx8QgYIMtop6ti
MAp+glS88c+mmBRhIXnSlcGk8Iba1ESZrtcpJllOEx/99Z2YT0NAfgG2T/V1oCv5v94jBhVUmrAy
6qmPmIFaQFJkOunfJ+BuPjhmClXf2v4jG1v7FZhP4WyzhlkfQeyE9El0q+PKLUB4ZrrG4iTymnPH
qe7tHK3Mui42USesC25U8clkDL7Gb1oGoofsi8vAVK7x7iZL4HRFD/p7wYmstcvn+y7xoY0rsutB
9puLeBM+ERM+yYJfrj98knmvoniiEHvUYDoeOS0L6mnqJ0hSv2khSH6DS5OAqWXoaI3Zv7PorYAo
teBFiHNrBwSLYVaHQ/flKCgEDO8aQsWmO+lXxJsQcyZLqyGnc8gD8Lh2qcL4pKbjRxKr+IKmn64a
qgSIIHd2kqz5QCbVcnmyLUtwEtiFYSqrYC3x4XvLT7t8Rnm078Nm8tquuj+eWt1+o9VmThBv+mBh
EERlFykc18x4ZdZ3hYlGfJ9T6PDhqeOafF6DMlcHHH0a82XZDOhKe9LoYeOJ1GN+NIoVF5SHtHa4
FtHUqV0WSTlHQuVF2+Ped8pOZ/YCSvKZJl03fmWlvlNPWLEIB2JvKGEzx78Cr/1jMZ2h75N96M2o
bwblXN35TjhPhv07hUXg7vOaBBMREs6U4XXuyDQUFptx7nYy9R+CZSbiUejaEzXGbmrvna5Ue0b3
RqsMS0SksEzfH7d7TDzyA81Uxqd5LmxrkyFaX3pxff2FqCle5+VEPhgm6Lv0KyTSO0HrX1fGyEko
Uh1UxEUNcya2WRh9f0r0ULMqdXrLFTcQgc7UPO8zviBumEyRLgzaNkx8YG8Hzoj0QGaDVatz5Owz
I+dQ3N4ll07fTz0aLjixicYV3D8mN0UYsNvLGId3lOkoXa1tqrOWOUMty96XtI5CtkHrPfgehASg
gq6hQDJb8JQG43h7JckSo6EwVDdf5o3FSq3fHda+c5jko5sYMjI09XdTkdqGXlTEqVwBbMeT+yW9
1LenGciLydSv1J+Dlo/1jgF2DTp+hHRKwYVOK850izfAAiPAA4+KkbykbXilLNihzKvjcJjZL1Ed
holx1NaVTkJhjqveRtlYgxx6PgrXBtTCo51zKotzpCcLwbhh45BsexmjkrKoke53IzUFIy127es4
HEMDiAGGYqe5zgmyo/zVcSuI/54t6mfsllgCZD8Gwb3qxHIVkYisEHdDsxhxGKt3hXfaKzM2KrvZ
29DM/aEUOX9RCfQB5Bg1woX3ReV02ummcOYjDQY5EABOqC4/5oxHf1g3zTUqslBjzSQl/VDzdPR8
A4OSpdvl96lOckvs2E4G+xjYan+eRls1kf0k5eLaNByJtw8WrR4OwpHQ6YYxyLP2Ir7R/DI6yKYJ
F0O7VX5MGjRVMpnVfdUlZONJQorye209QEKJu9qPtegURyXK8zrJ99jMAU8D04IuXUjRtOmHHzh5
Yrp5mn9gf+YVGdTdI8Sj70xDQF5CnKE3tKilgHbUjJWQ7ua9sRwGvHKU0m3HrvYnYjA3/YE7+Kyd
N3uP2HRRIGF9EC3ppWt7On09ZeE+WTs+oXkmNle2HL7RUe4yW+J/jljHtRZksJgaXx5nTXXS+g4f
90Je7vPj7/rcyE1607zytNn8zSTXnYBuktafpOZae6JZWMH4yqTdcNZjq6PPxYMGWJJBPnsbf2Wp
WH3IBXAoyHrLXuavc8layaAaWqiKszWmk5WmWg4u8JnhUAvrzJoft95mfD6XrS55BeK4mDY0WpUy
CGTuIwa0WUtqD0wv+24jJY7d/GbIjM9abHqi25XsR2EeDk5IO8HyuxgamgLlSXg8B2DM0uzIV3iw
+I13UQJ1Uuaf0IVl7ZA/frCKed5NdkiTQCSmnFDWUWqkKhnSJfe06IedxB65lzAskYd3jmAhxmmi
5HvKgsfOFL9vW3kL7Nh918Lz9YcsOvXrfkv4x2CrU84XhY/chy19cP02CN7B0+leDhob7DVNUqRP
YhEjsulEK77+fUnzBmigXCANgk5ia1Qm9NIhsMgLr1qujrkhSSnl8lVw2uupl167rhuJfH+8KFWA
TFeBmDqC4toCpzbpNbqD4HrUBpJyR2urv2N5tlcWrb9S9GIUKCwtdgMRyKy28jL88169g7oJ8Xsf
iRa26R/UVQEaRi+0Bbr4fpLerxkjpQIR2YnVwBe0QkGU86/QjZ6gIdx8Zh/zYStmj7WEM7TFK30k
OjU94zWIwqpb0Rd9ZwKYPj3TRavrH5JyXRXX8XEWq/T/bHXebgeUADAFNLC2b7f7ZWU5GzBt2bH4
A3RtRP2RPLacLOaRChwbtd91u5FFPjT+e2dOIxuxtIkjHWZ5Lh0GtVC1CiB7z0byJnxLA3C103hv
sTCiMz+bKm5fAEBT7TdseaEanv4vWyXyqiEjDk3UplC6LLr2Af7BKHM+fmJKPV6HgLzBGygpSPeD
+GQQ4YaKwr4Qwixyz9+cw/C/Ni29qnl7ir8qgfVDT0c74+JJiQzEgSpbIRrh2NElVqYvKggL3mEF
mHeJRI0HJeLADw8CRcfEbIwfs6UpnUJGv15XjzAZwNGmRWxYsKyO8k9okTIu4QMexEK3FvQFBpIq
twLvEJwrPlTHYun6GGSRvxJxOTUO/8MTnd7Vr9NfOLnv42xM/3vRlJ38YwNgYElOI24J3kg4m91T
KFV8Aw1yV4K+5ncpd1einxOYwDHiH9Cen25MhGThkzC8CsI5EIs0mmh8dJdbOwypvHpwQFTsXVkG
AjxTjSORFlzg3gbbHWNXCdxe6tCpE1nFs6wU50pmwtpf5QwUSMRNgIW3l4qJbs+0jJaw4yrpJysY
2R2std1b3uzjJO2Ilr3nmPht/gKi8AbKsG0K520rvqv7cU+gbt6ZTIABLuEOpw2uAuclm/zPKEOK
l8d50MCJneKTjT/Ch8CiIZKF7cH+naETWkHkxoqWBcXY8iM9UJZ8dIdIR406pc52+Xkd4nJo8CYy
JyGocdopVNmwDI6JYrAtID3uzmEIjvbfPDVbcqNvM2LZ7VD2BlnUvIGUi1E+OG9HSYONncuypH3T
f3QYD9ZE4Hsr2Ja2ADzyGpH5XZ6yd6/vwxzl1GHBBjreIA+4gFUANAgmtqQx3kDtc4AGX6QiOv4N
aXGACXmyy6oluKNDWTi5ff7sbirAqGdnUWaF5zOx2Ayrr3Xb3UoxCxkVXRRSFwDRqEegiv7vm5kw
ZtnFMgMMMFw1jSXKdeQD1t1+12MmQ58zr0JocR0dbiWi4fdpjuujKFlyqPpOBW9yEbkHFkZ/dswP
s9BSNmkFwhPOwFJ6XoaA4KvVu8zeHsH/GAJnzr9DV9JbiWiPYcqpu/WbXw40k1RvLYU4E03cFrVq
VWAPW5kB4K/NgWlquk3W3EIZZN4cBLib1HLAKn3/tA7vfqmj/+iNePtTAFPDQTxqtCfRmABqWlYR
MurtEvDwnEC1RBYyA+FK0AY0niG9HymOvABglSyMp0/fxjlZ0PHblVPb4bJJSGFxwZ3cZNvK0Emh
KBT26SZE42lGKcLUCCQnc7Dnet7xNmkw8eL5l+eqzOe2HtnfGh/NITW8c0NHVsQVH9Cbq6Kpu+6D
3LSNSmvcZAsT44lFjThQZNJ7YrlnndBVUfpTkLzT3kPANt88EUNYbJfaucjO8KWLMUk13h8K6O6T
grsqIRERLmFkaiJLBKUruBI6Ww+JB8bk7dvIRxWhZGOlbhvCuFevHMuUamCaJRe95Oa4/980aoRl
83ZaKNEh2/1Cl8M3xmT/AGKrtTyaFY72i1a5nWvntWFH9WqUcL8eL43j2G8mJ3ra63oUONHmspI9
K66ypYhC10jMz3l4lPnvXsve6LDjOMGRqDkoOW/3U+Sj2UfdjsTVWogvJPqILD2RPRpmH6fBw0p2
jVQHLBzqY2st5FZd/UiRTQIDj4o1a71U5xnjAXqyVUBiRRDmcgqbsmfLFkYyqZOZE6uGlba7LiLG
OYMLjMFThUSIQmKdM93+In7p6bYMSZSnyQYgVT4GSSL+EZAFyVq+lm6LTesB665FVerilPwK8NhV
a+DjIRAy4FGaTBByrYAno6WCRwbwwPLBUG1ps7NR1iH+eDPGAu8lmClWtQxvjIW8t0qcDAqMYY6J
QDb53EcCGnIjJTPVzmxxSvhpeCXYyYv+5raoP3KhuSh0y3kVOLLLodIQgUkaUvirW/Vdqfom3Uvk
0wd+jBxwjq8PiBVT9LnhCrDkH3hOtPJv1/nw6gA4LfURd3xi+1C7xbA1uwTmVk5yrOYBYRyXoMbU
2/JZr1y4xFj3CXzdgRh1OUjwfOEjg48OwWxBgF50r4zluVZP8hO9k4rabNdnrmeq9mXWIvHt0bTs
s3dRtBRHp8a8jCEkDThtcvDb2vr5NDjlck8/H0KBVO1dghbpgElDbDB4vKe4JcewjvwP/GcF2oFe
ioDIWd4kGgm6i1AhMHMiMruAVOL+d4PaXXm40yy3SDdbqcDwS1ve1lY6NGvzOOm1Jyf2ps1nvJBG
TuUhkXfBZHgg0/TqEXB1+oHlnIRHAdBfiTQL2L7ASwTejRAAq8E1/hSkGwLDMM4eVasGSRhL3KAn
lo+SOrJYPqMzX9cfmiJrQJmfFSX/qAfjAaxxZ03k1hG0z3O8Pbeg1kBHHKmGakCGXPpyQdJdmAvk
9GCGT6UUtd7y6XWrn0Qp2CbS8mAfQHPdIOX8vvlqLhZbz7xN69FFYtZntdrZ0Vu3Ya3SVRE/Eltn
BV3YKLdkB9KG77y0PmPbQ8kSocLZ0EqSU15XVF21ukfPrl3NW+7mDRxEeSMTCBzGjz+EQQYuyE8n
EM0K92AiHnrfIdgHvhtTjWteV+ylWvtaWalWACEMbxW3LUnlo/KwPcUCSDGd+I6tc2Ig8f0S5xut
crJnEhlmX6FGVkOVyAO37b9SHgjSy+9nRbSe1z5RGCNdbkysyC5uCurbuhcPyE1cE5iItl9Eh9XE
VGZdtzlFwnbsrJALONlreKqARFxuehvAES32F7pJYQ4Z1D6OP3Z72urRgoFKUKuKtZNxq8aerG2H
aj14ahcTK4JkhrOKp1AL5y6phP4M6UwoEpjaFtwSfH4QV2kOZ9vwT1A0fALYPQB4nN+XQQbOAWho
/o16jlS+DDbOJDMCwi/G3gj6ucCVf5ZQ7fvYNjoN4Zm0I5s2PnlxEKFGrMiMIkBaeJaWICaEEMrr
ZKFVS45a5rLUUI+UbSfzjrUdfnsrp6CVUjPUtGO9f5+nsbc6fausSb/iGQrj4ZSPJmKdJguMDk3v
ECQ9AvoING5YaPocv4eTWD5mV7QHR+G7/5vlJB0THz6rWFUx/Q7FuJbfCy1X8ckxqwt98vCkGbTr
+8F+XYbUIqGq9LulCmHQbfT/RmGqKOPYYaQx1kJvxUSk9+9ohHDu9meO63dwZ3QhzQrMfh1lXLuV
fi8Lulx+A4NsIasOnWd3urJC2Vsw/NonTdDW0wfMK2bMigkl6qmzWXu37BtykdC0BO2ilIOfoLX8
ra6l1Wa4DiKOTtsaNKDrYWPoqa8E58avz7qh5oFKdOaDfNzaJ5kXoDJJrJHpFV57TCVRxUMhb+bz
OHyT/mG+f+ohA0Ykd6ufRGRcFT2SYS+6j6mJ+KASKEAxmnSTc7SbPGJwd4oPr0oDmkUim146SqRW
dWMA4nBnVJJ44EeTFsCeYw3c82fFMZjnNzl8VUt+XhTA5B5HNA2ZNyfsMPlP+1m6ErH7S+A0fDYd
vlhXsHOgI4TgWLajmMqglMCfP441Tia1hW+fSNyZc/S52rK+8jtMyH6bSswBkWpYQ6lpVn/bPZ5w
qWEoKOrFV3x4CEwG3Jt6GN8HD26MdMUFRq/8ren/aZFiQZfnJD/H6FZe7JwnmAjz3RuuUTSo3hWk
zBGBBAT8/+rj0ZSxbBwyDQ7fjSJpSfdNnN2IaRgx83fYRWirbkGCWKDNWJNIusmH2JQC6FJep+pf
wRZRSoTMbVZ+LpnjrU//bHSbqNi8rBOMo0d/bppueQQS2QxS+YmWgJBw2HnLqkIjeYL14UzWIFuq
Sch7+F3e8PUgXhh5gWzyBryKWhSjb8YzUbXdPn8iT9KvQW450tGwB/824NibPfafDd5pTM7X33HR
WmS7GjkKIj2r99DrUFYS4mNDHFFkXBnyvh3YiyoKDmrVmOTfPIRQiNABKaZhyY3TE5ifSFjAPg+6
xHi8437P41oD6Dlai1hajdhIOOWipeOoAzQ2YtplV6b5s4RwYEZcFV/gJPKjUkYI3sMTED1pbiqx
ZMkeHwQ9Dt2stbvAtCYGU0vmSyGBYb8hupVBs0+Y7ZEF/DFGBvYJ5PE5FzZv/a4gGD1gqEe85hRg
N1qWulg7Xv25gdCRh+F2eLiqdMhHSbOoMlRn/S87HVlclDdPFLfSmUK40Lzk/TOsk1g5H6lW6Ukf
3UAYr9GvN9lFItMpyFIDv/LXwr7lTkUTFxC1zhJn2to5fft87WVd7mWHRVxWOu53MlWRziso89dP
w16sm6IwUojsM9605rticHOFD6bA5KOPlrudULg2svM7kOfx6SGAJYgTD3tE31eIeN5ooBjAF5ND
e5/mIelIsOXTB9W2FNh+Y3W1WskvMzgi1Vf9qrjoYb0i8RxPXqG4IGCv1kQ57i9Pvdc0Yh7xfbO9
GFf5laO6mudhxCeXiccZGKaSwgnCm91Fro0XV1vRV1+n0Vfolto8rf76j9JR/snVsl8NmDimgSF9
sBKdsxGWlJXwsOIvtcGP/20oq2Fu+AeeOiemKAKdVFE2mEqUINjaZdB/Hq8ZHl/w533YX3VL2UC3
kplXwCSxRKuc0YdWXtmk0+llFz+LJg3QzCK7kw5SdYgvDHS11kZzeL48VJ7RxsIC3e6szVVw4tb5
SYJVrEs84tJ0qd2l/RqPhVO6k5cYvf4isf36wu1rEQ8t40b0EGMiz2/UR+DL3Azia8R4EQJ/AHFj
TVzJls9eKwiHS8Cu7Z9wX+3ErRdFp0ta4Ojb/DOoT+kdidt6a4Npo/gfwH/PvtJYfy9ivn6aBF/v
mpMpnoaYiCkIrnIkp72gcVu6YYludNypdPaQ4Wx1vnocu9Pkp7BAiiokON5F6MTGOrOrSzBCG986
3dh20KU3lH6p0FYIE7QEguzmpDa9UuIxun99L7LRq33IyULC4t7eqtagDu9G2tj5KXjHB9NrPpUk
RTl75i4mzn+Qq5iOuqhxqyy0twQUX9jlTYDzWqobq9RXCNHlNl/r2M8igAPPPR//TjW9yR8ZL+It
aZxI7g246Du6Hq3ZanPraJ9cNlHsyUH5Md1lIV8hWkGkOSd9I48MgDg8igv6VrNzIBN6wVWrKH5l
3ObYYSec6rG6hJDHWYCev/C9D3UqCSAhWotGXLWtvfeTyNr3z8Mw4qggPSV9IJwwy1T301nygBkh
fDsSwKv/8ifI+IScjGHeXkszZUlDoNbewQz0zY2PNYZVw3G4VX4DnespIVPJjRzlmDZkuKFi8WtO
7U2Wu8Hwkwv6rm8eWeAQG5+YHz5s47T+ry4XoOmdbnPjwPnIFGIgpD4tHYdMSh3Vjp33gRm6LFQ9
U35KannpsyJN7Q+pcXakKFKf+bKP4dk0o5MoeNaknwDjgjmA/5vOgk4jTo5tZMiODr21jpkJvkwT
YeRv45cEVAfa6nmyL2ZyAq0Jq6hPfr86jX8n3rOGYt0KHBNN2WJlmzi25iPltLR+b6/W2XL/T6Gp
BxlJ2ZHvzmgrh+AUgbjGly8Q1UnK7/A7VEnyWVgSMNVVNi//hl1DjESCJ+YBJ3EDxLsPNFH35F1h
lZYQAkGIIbjaAPFc4mzw9dy4fbiu9GDHC5ZGvfBiK1RGYVQTAgzJAODnI417DTNuqS3+gDt/IAuB
fmICGXnSwYKZWUZphlBm2RHjs6TAL1+E0kSKQBn0l3ZnNPRMyx0Cr23IWouf6CnnDn9Wq92Yax3W
gEiF8jokIaX+LNdKU9YQpLykDApBSWALDpHDcPXRghYNGGmFgPoU8/+/uJCUrgoNNo0fR+lTvmIf
1p38BpvkiXPyK7VCLqDGN2QOI2imjVKLstaaSs7CQ+XJAkxgXX89Fc2ZtuL5gfoEIJyfRaESOKXT
2W/CFRRK3grpy+NqNIijfM6K0awOH/AL0qeJEFj0CcgxAFPyYW8xvsfLS45/0F6AV/AqYDiwlkhE
o3V/AqmzpHspOwaj0ZFDdwdPq1kD43uzBr+EZmmTXli28qdMR9/6UarXHh0V7XT/cSEZbKajuavA
0CcpiKaW1BdyqRhulTZ3svcDWWIoTw0FxHFaJuDBtLr6y0yrJ1eEVouolhURjOuQraemjtRuBIJf
UsJ1yXwt3nLWK/EHNz1+n+NN1Txiol/yNH1FoxY5BBs9/W5O4qhOmGlanDW4kO3QolHAxiskweq9
THbn8dUINdDPlaa7HIO+G6loTirMAkQKTL1E2Q+q0m1TLQMHXAauaKnlnYkHumVBo98XNaTk4xQw
hp1vY+r+aQNoZyjQaecCGXzhZ+gAskSVrkYOouXVM06qpkt/WYxVQ87P6IXP8VX/onKivVQcdqXu
ftv6zYmNO3TBDsy9eTVm+ySMPRD/CvqLSK+amhEvM5ZDKQTITLH384dA6a0sycUF8vDr5c4T35DR
gbJMz5W6ZzomiDbR0WueUkbpugwPF7g7sGYjcGtwwxjSPhnX3NPQClHYEDsXFbwciffY3VJi4HjV
eIKubV6F8vsxlpHAzQPlYVlR4E6EV+rEqrmZQbSC6F/IEP7gguuEaiIoKkOf40VmQzUxDKoR/MTQ
Gmrdckxze28gRuQjGegRH+msCttzN6/7EAYbWHocv9eB2uLn8kBLy9dPjEwew2kK3ZcPQrQLCiqY
bb7OxJnwPL8AEJyiMpE5pTzeOSFowyZocAD8d2ArTWoshfNjDHnU8sdAf7oW9GQfL5gjdnd4PoIg
DilkGpT8D4W73EfCSyPBZRcFzrS3ijH/3cEXrOOD/YSd7xKqNEEfs36IXQmqzZ7fZ/SWnKgUxDZk
zXt55AJscgqSjMYjbl83P7Rkm62sTbXc67UxwXE4m2xjcUHr/MheRGk4TES/psDWEsruhPj8FQT2
ixf1uXJoOmcS5z5sNqtKnKqNTpcbgGkUEdNDUvQHfmTdIjG2KCIe4jMs5h5wTjh0EEE4Be8evo63
ubECYNZCOMhxRkSwQE89UI28nrHtnoHnYhwURUTSVYZrV2OXxf90ZZlvELSn9S6dOJUKBBGkFJP+
Nh/FoU9mifsmU//VlMAEbq4vxz5GRCqVAvuLrtK7GgrsySLlEVe9QefJ0syX5YqC6OrOt6R/9YXY
6hszonMjJ+efMv38YZgof3p5aSqYI5DYe9Ispn7efrKjIQEhKbB/339w3Ewm9HrUz3A7veWlO7Lc
h5toeyL1gCSCZNI7gEaAkwgQKzvXGKOXLCMtYMtNgsfF36JMeDMTNaCV1YQIrDB27iMDlqkcYOSK
4VrONbfaPYCrcboinZfO5JFQUimBy+9n2JMd+apEMBgS8063UJ8YwJ1lZwBVhOdlK0mn4aEd7hLf
RgldqUVs4GxD84ODC2toyBPQiA2DZpEF+0scwAOf9a9gsscZxcXG6ROXsZn81P6ro3KH+OYmJzjA
ggdKBo1lxO73cYUv3F0z6SDrL3g3XBSqyvT7sAPsIvVim5HDN4qrUMOxvY9HbyWnjWrEncCBVvp5
Qcat715v3niHnEIXLi9C0QwPN8QrJiF5mV02ytgcd/VxgsGEVa2ksWd2xhaqqy6lKTUnAwpbowm+
XoS0g2LScSxVLg9HIGkYIKcpbUMqNWpNgjJhofXjuqqZvls/eEWfsmYj/lf9ht3LEcEKsYfu7Dhf
5KpIzKsd7gnoeo47IsnHDOWVC0vzKm536qnUiWKr7qz9v2xnUH7Keel2JvdQRqYOwVKD6mxZr2y5
jYPpevKXFUDwTK9uKOU0nc9x5DYBAcxNOzbIO8kTAUn/6Ct7qkVBltfrbmDx4nw2tbb1eSK8mcRE
/Zd14LnkS67NZQ1b2uJ/0jXB2QZraYdqPjYBbcfm/Iocul+6QDd9qY8cxy66aumcGM3ckUa59c50
i36UOjZ+ro3sGJVFkW8mmrrbH+TlKWMKDjjuEkQcxacXy8hN9qqG7L1A66f22Wl2zt8BN+NMBI6T
Mk8C30gYpTKq9sklpvr5ckdHcw69Cxi0F8o85mEILzrjbTgkfSvz7ZFJyTlxzvykRctEhISwljA/
5gC7zD2BfLSEI8/WWQ1re/CX+x9PTL9VCOv51RNQ66+ohPICD/3d59fG4x3qJyaDKBapzc0+vqyZ
Y80qsVDzbr7C2t73QAc1WXijGejUOXoAqFOjN7nzu7Oaf4IXaoQXs51naNSH/9mPDqG9q50N2BNn
AvtPy6/5uSPGtJBrl/WHlOM8BUF4AYNzTa/ArzsNysH0Ig9U+K/izRV6sENot+PbfQhrj7mx4VoX
VDGCdZZEps820Q4n/LDOC027womZHpU9YKyDnmkstWJI54PjVQcm35An+gQ7ukxmTdqmX67/7i0S
snP6jG2xQvgt92gWrYpHOx5aP7MBFNCJYV217dGO+f4owjyhk/e8BSivBaPtL2brRYXwRoli81eW
td7P7FBCJ0MJksInltAzi2+wO39nZRgekVcr1KDPBtgRqA+XjLdCVkIA9mgQpL6UGH4SSOJMyLC/
gemOxNdVFj+7E5nk47QTdPjKlkb+TqY22UN1edym5d9eTz34stjTyF+VD/bfRldkZy4L74pwPhG2
1rlSUm9OV+jAu5Hfx1TqIvXx90bwDvXG0TbjjFEvOBQVO47jeizq3O/9FpCLARnaJuc7iVjujydT
VLucAZ3Jt1k2f4o+Y3udrPwkfIfRCt3XYubt74/+pjBsMbYUOscr6aBpwh6s/KKj4xV+tMD930x3
pDwPGutcpz/P80kKBoR8PUAS5uX2XpKxwZYqOt1d6gJyVpF0EffBxzXgqU7e1ThM4oYRC3JQLqnr
b9Falf0AVsK1f3oqJiYMfPq9phdCyNoLfax5+GQX/CHchV1ShXXFFxkm57jNvDKmLgZivRhQoA37
9jBLZeHrZq4LDV87YJQwTq8CE9sxkjJYUYue1/6wPXazyRHm5uxlWCaVq2DOIFIh2jcykkHSs7fN
WrHc3ve12LkG8qUUG33IZSx4zptelFtAduAHb5MCX1bDhwjVY8c+cYVrXfDKhCE3ZfohVI8gkdED
0Dp/nJNLX1uWA2bPiIa9MC/WHPMM20eq9vhO36A0qF+9kYtAztLf65kLsmTWItmwASRisxJtR8F/
FyJGrlhkRKt6yI33CjvfJJdWQrwhpV7DXQFMMcPZ6yxbPffNinEUNgNJElLkSOJzmcJgX7BNtUr2
rtIhyhZWbHTQKiIqFZxipmD7MsLBcm+nBStYtjS15hOQUGGOjrLVvHDkVfwFdozUqr2zEAEBMOxK
K//IlT8q2u8J4H1OC/9inHr70KrN21WdF38BqsjDDRhsVL5DNv7Z4D3m6FCWaOeO0dUhq0qU8xxQ
7fSf/ywTfR3wsRqw7FVmylCPsoqGeEXprm8P5NLLPtc9RCmzfMu9K1R87xCBKF5gZLCbef/kGJ9h
7M8h0GwHaddN1LKBerz2wgNJF1BS9+Cho7ojYn456uND21fpWAGNl/c+Z8d4Q3uF6jcTGOmuGl7Z
9DACZrabc2D+Q5BXsuUv3Idipfjqvh/ubRxZ7Z8D+Xn5Wq0AImkxuExJ1HS1s34xmD7lzvwV2ijP
4HP3E2bagKzYeemmG0erPT0kEAR7KJTMzrjsrlW5nwgBywaBNF2CXs+SLz65yrswrFy5kZO5UEol
Oou9+3RN/w0Hvuvtu8SYvIqjbf+Q1B3PuXA8cH7zT24gGJ39UDpGrJjNrBcB337i8mhx7xOpGAvI
s5SODnvMgS4jkrX2buiJaPUD+I9P98FAfbSsM0Yhr2CdP2aIsGqdqgMyvjgq23dgghoLYXG74u4a
maOyJgwvC7pmWvC1qg1dAyd0imlZuPDKcyRcp6EKpQPSo/dBtCCGupOL1XX9lK4i/dvsZLFVRoUR
UIOu4pwwYgPMwKPi7nzi1uSc9jSSxgt4ABjOgRopwMOrdWI/aPR006NENdY87PGn/Lzw6B1v8ow1
nGBfloy3UzYrOQ70G6QshNjNnJhYj7L00t73lyx431lnZ+l35vnVPSF5eTFjE16jhJQ8Y44+npKg
Kvu2IKudNZVUJQp7AerjkPFgqiprUnX2LPKqufuNaY8xApmHNHKGn6dQ8Hg1bo5Wr2aByyVjFAWV
8ikRN0x7Ix5OUV6WdTdSOLZNYk8bvw4MUx/eVANDLjFadLwlp9Yyk6w1itD4MrcxgkVBMNmpxAGE
R364VTY+HpxjY2xZxxLJnOuwJ/0/auIlrLGuh4PMR7J1gBURqhLOyAC8xgGgCNxGWLTwxoR1nkS/
JfmxClioWTtVps5dEtlVUVmLtpF5hRu8Yoc54cTnAGA2U8Q9DvjtIU6hULTFTKWf9psowIFKNmTM
5BzfEPze5ddRAEngIlnLRtwCxcUoWVfDt6V5jssbudgwysNrGAvenSwoKC0DhkZOcMi69d9F4eVi
14LyeKDk33317/D2aKSSuojbdwG9ZhD+LrnzO7B2wxaJyxHmO//Y4KzOEsX1MoBL9qYPXCpYQqx1
GoLOPgp2T/KfNrdzcvqO3V8nR3rz1JFr96FPHxLagVohBB5JHj9uTh2a+PkwbT5cafE+vMJOCmFJ
d22lkeOLN89WJx0dxEH7DgINPEEnQ/ImNSdMAdHdgxKJvUIM6nJdq71MvGyb4PtnvzA/R5G8amIy
+z1Hs057bj0ozuzA6HBiEEE57pme7bauwQzlL14No15Eqty0mLVfLrtH+2yShrXlFXQ5tuoCTCu7
R3Mk5lwXQEDrCInYadaxo7uv4Hr2WTZy8r/jAupGk/z85go5QdYau5OVtnkZosIeH/waCvEOEXHa
oECacDOE6LwhYBrEIuDCKhgkbHADfBO5fgXuS5J2Q5IS2uEAvoSWkwdB+jDgeYbGYfRb5MVKM8yc
J0mKEhGoxIW+YL/xRU8IS4tbedSL+DXw5zz0PVyAQAu5IYngSOsGDL6oaNu5LuvlCSHsmoY9jdMz
PedCK43xUgbv4ekxY+hLf5WhtXFoyWPQ9rNbdiNUrm4ckVcPxLUu5kApblHgUWETmYIujO6NCDDq
uFnitXmdwuCjntdOuJwpBjePelU1RI9COvd2WTXYuM6/0xIpLB6FbTxDJ0Jb5sDKZWt/0oq5z3yv
tOISnFl83KYmzrmH9r2cMZ4r1QARiTFO6dEPqDPmJjAHWrX2FCmFw/cYgS9BL9za1eP/6Hvnk5nl
UXr+gCEHhY/AuORpyTUoIxyLpzvarWdNBQBKgETOjQAQqm6NSLp1zbTNNFMrCzqBVwpkuBAtKSDJ
FeNdoj0LuobHTA5HLJ1VWWUomml79U+s7pZ8OHe11PdWRNXZdUbFMJyN1PxzRb/oNwZNE/RR3SDZ
pFf070DnEZrbss8MkVgWWwfHbRO47O2Lexa8H3QJ5B+8PaEw5sH0K6E6GJyiRt8PYFnweAVLH7Fi
8GAkoyzKpMf+MfhPCU2EOvibBWylICfOkLZD5Gzu86it+59caH9i/jFf53GN8YeMV7tNJ2of7kET
s5WjZCW/B6vwJC98D5vxsip271ZLC5qSkM6jtqU053X/NCY9m91kFDr0Tj+TCNuQ1E5Vh+Ym2kgC
eo+TvmVzalqqJMQy8zC9D6+W/KxQz2DZfU81TrK1H2pxDPnX+GUs3zdxJaffJYb8zQvCLyRpInIq
yKNcyk69658Ib2n5Frpg3gXbgktNg0J+6gTSLu9COZKp86920MeolNxwS4ikXXcEZRTeZMdgrEgG
jHTaWBgBhLdIwwVBaFYg/aXaPqfpBBQ1NPpVpAa7QgN23JVZxp+04trGMt+Fu83P+VnSba9TOIX1
3cxL+yUwR0Ab6C8drek7pu9cva/G5G7NwRb1zQSgzlMTotRMwlgfH5P34Y/VuIEWg66Sjby4lQhv
r06Zet0FoHmTvGEo+skBFW0Iau1zXHE7fPQZfjLZCDHWmoFjz6kip0tpidgSO6JnD/pIOuloufT2
vsuHodPf8+MOn5ehAehDjCra611pQw3EYk7RwmzBCMoguI8S5fvJpX43O52WJmgxpMauAh9lCZ3n
NETmt5OSuJwKMkre7goabEEJ6t8JrniE8uizf/ubIsSaS+PVA/lDe4aN1uP+heIwK6QYxEejkJKx
QJR+1wytEaxdFFjT4f9LqkcsEhME7lizRCbDDm3I4GulcasWhVBIKuo/ZRkSPX639RCJlYOmQV8S
9MYlU4FxOMJLyneUUd2AdPmt8+rJxL9izwxbGUCsyD27cjhmWcn4+pM2aVHK3cC/GSCWYMIBVjDW
C49FRpgrWJALaWGPeUr1UoIFJWYV6/bUlyVmXpdyHCFV3MXARqpZOgXaXP2jKNwyjRVGdt6POJxo
0oD67IP2Benwj7UzIWeZ601+2233lr0mueXUbVIbcDxeusjJWTR/az+puSfjkF8nOFWNZ471eMk4
lkSwOghwQz6QeDVYAW4D7T5n3OsQ4+QbfEKQcP0USHKmSsSLURz80RTXsH0o/mkwsh/981Wm4seP
GoOFnFc3gjm94ZzVkRSg9QwmPRyP6GcwUXJejILj43pbZr+dzlmN3DWYMfhXG7tSV1s1QGAx3UDI
swn1dKdX+IPxnXB86bpZYrMOmhWE59IgiLyqoPuhcklPb8yv/3KeR0mF8IKl+RujgfMgtFAAAxZc
goI4nwYAyOZ5avjDj5i4ISz7T9lvoL071DYREVG/vOAlutnJbKePfqcaREZrTyI5L/GAKE0BDOVn
TQoONqD6DTNlUz5cs1ZvSD2/nDAJCcGX5U60lbKp5tJN2XloM68Ube+oFf7nmJVBECTqmvy36VEb
mt/KHj2Qsbody8nCqnKLVoBw6ORll8MlEivVZzJlu5IT6pPjDiI4Yxrb1JSumYT+Y9isA7rI9NkV
WsszllZLKIivw411ib4djGsN7lW+XKIKkSn2FKdI8mI+4AdqUe3jHp/J2a4kC7ItALdwwJ3RRk5a
O8QXTUxIAsNfjwzqyjyH+FtnIncv06AZhFd3JpAM9G+ydexhgTeOYCNqwtj8Z517IUlGdzai4quS
DZb5VT29aKSMd/t29lqRPH5E55G8U88XPHH9z+THQRuwBtoxwFGCmbBMrNP5rFMi0gU9hXq5vZxY
Dpp3uGfd1y0ssUyTtkP145XmCfe8sd9KbEDqiKAUqJ4xNDcU3w4yZYjzpnPexpmn4eluMZGwZWbf
kQiSHOZQUJ96iS0EyvkYbUzOhOainIFJXd0koySZ3KLb8kFiXEMLQu4BHpTnX6/DriRGuAmqEZbS
dxmPzRig8vH8mLjrTTgEHMfuVKsBOSituxaQR1XbmsYJ/jlzcDajBqyQnUvj1DvXxHeDsUjuA2Bf
3/2NQXvV/eF0kmeycRE67XZ0ctP4KWw5LgRzfe3XbLFft1ybsLvUjFh4YYAU8fYd0TEw5aaoEJkT
q4vIDr5aVT95//xazctyTyiMRVwzHqdmCc088zjWqZyEpFV6KzPIWbyZsAZPaSs0IXPXNj+Muzyw
nlUr9ph8BLqhTaFRg8RBT91QOxJIirHZt+QYVciRjBFHyS9r5Khyw74eNNTv/TpQI57sLO4UPxYk
72Kp6v1+Afgi7YYxZXujIu+nlKBqVS7UQn4dYGPq72pnwjKJn956t6/YmG/zV2P2JKQyCrULFKDz
kDCvAyh0VtXasL540Hcmtv5UTj5OWG3kJA8rZ5q0NYmd9UF6IyVmoTKJTDFxwgzE0CKo5fKOixpP
LZlLbFdYXkTKV2BCe7z3KHCHVjXtcQsiMMBZlnQUK709G7SLcMAaBnVP6FGIQUBm0WDcLfs4q/1+
qQJeZoVQj6VxQlkNdoPpmmBd0G/c9t6I3jUqU3K+2YV84r1gqK+7XqV2MpWqGuDvwzP8X2ldeuzb
ZzNcIxoy22J7v2ELLOg9+Yw+/HZbCq4degko26o/8cgIgZiMjmfz5uv7TWaSz0gcf7QZHGm+GNl7
6FGA7TWN9Z43uhtJjeijRLVsaQhB0Ry+cznR/JynEgaXg/9o//lst/EDnQLwW3Z7xmiSrAyFF9b+
6ieJvPi1Kwkyht7hYGaIC3TLHlQ4hqKK/cjw8Q3DWzZ9Ebyl/ffRdvxHYftinML03FeQN9JRDNgq
qIlgwwrHP9HX0xLHB0lKUnU1k+Of+jp8fGSJU0A9TfmNKPA6pNMoKbWodjwESU02W9uQvAU1eiw/
t/FAhxoQNhxm79A4qqYIIxuIQiwkGTQ05Pyy8KaeFbzYuGc4dDG69PvNXjIBxw20sFdF0kfbE1L0
Cye4DaZ0ludm/UUxa+caCrekzPwvtK4T0dah4sd0r5jufBrP+QiBrpAiuavIik0BfLogp3cvhgVK
LW3h2EDGOvcIP7pNsNul8fZ+xMUdMH8SMhazQInPG8k+AoG++bqdDcnSJ60JmzK1plhaOwBlrB+v
3y4Txu7xWuxgcSWdk+L2KNcPZi6+z28iOb/Vmm4EeGeHthYVvR7E5z07amcaeehsLz30v931Mn2n
JjOQ+l3RO/sKGSY7dXiqOzZBxR5sf9zCuaDLGz//L66tJSuCbRZMkT9eollm9KkvlB0tyRrK4KBl
bWwc1MYjRqnP4gGI/rRTy5c/EA3XkXkDyY6Wxr7etxRt4Xhsy7Lr+rAHckEITQfi8sAYI33fI1Z0
MAh0ilQnUXPHx9Ctk090k77IASDJ/i+xwv5F+Qyo5w/j01Z7xIroqjFvE2rQI5VRyKZznb4e60lT
IyknPcjs4Il7KulArrcNYxDqmNKnaeOKLFl4KrXnZpJbRKfcLG0iYCSMP6TgGTYpTFpJFboo+jrr
zPpKRWkMi7u3WzRTxETh+L4vuR1FpeFTZcCLssU6v5rpcMf+w1odo7Ru7KH8zLkblN78+PM74MDy
WYQbv27CLxW8AbwVYEYWbPfaA0Zlrtck0W3nd/XKO3G2J9LBakxyz9+LIbput/ERszVUCONv1uka
sibAQ15F1cl3lymN8q1juQlmOihYCfIaK2712n5ErU9DlynVo35VS1vRYtH72nmO7SvRoXd5bHBw
ElvrE+Bkwj0Q/3jDb8OIuEJ2KI4dUMruOPeF9Tn7RrJHzTaleINaZDYztbh0RE0P7Pc3PiGVwJh4
LjFLi7MPMwKwlYLJ3bW9hIuhDxGj6XUsm8IfQvmrVPSNAd5+1IjjzXZE1TtrIlbSsx040c85iWiQ
j86suya9eizxogbEJ9WHGCAue9IPNsx7AZjv/hbbxgbOOjpn1CUCgv7mqK91whOVBrQpl8KKB20b
i0aO/bvqnbWwtmgMWGcZf9Pp6z5txEmAoQ8fWyTLmFs94Ny2PRuqsmCARXc8NWneu6AGbsBKST0D
xrUZIzOMawPuDjH+XdQSu+OIv2LU4B3Vsd8e31wqqrl7wLJfqoEMQR+OAidZpZlTkmpUuFP79yoY
ToKrRQD8jJ+R9wabATEexEvR0pLbuRao+zK1Ldm41bXnbFBTYgObsmIYQ8Mglv+8DcsX6/I3qCOD
6eccP2pm7jvut/wPas7KmO/2CCF4Q77Uy0+hs0UJNEMCaaVjOiTxnLf4sQ1rzl+xUU6D0hhdQ/Zc
gb7DzC1HPPXDhB+ZhBtrVWIrC66Ii8TbzzwfaLG+mMwKamyNyn6TEL+FpNBLlqmVXXoSRGv8k/U7
QUdjW8RBJFmXDbDi6ApPWsUXlmauo+KiBlg8sJSzxVyOeOfUBLkwxVnwk4pNB2hGluKv05A+eypU
mT+BAzk9WFEQvE0xAfIl/ff95ePVsqK8F+KAn/e3bO2+BRJ5yEK9V2ciokWfdyuuvnFzf/5wqQy2
Gmv456yZhWoqfuhA1WuSYjHYWh5Tq3VFBjiLYMeY/YZC9O3/5YlfMaUctGXvNUu4Rh0qZVzklfc+
jA3cHVokXCmeCjUfb8fOsKMqKG2FTEuUgJLc96IpBWJ2I39DZ7nQmMBA5Zv4N7t37uHeds1Dbr6q
BIlswvbY48ahtX/Kh923fxRnsxcO0K11CzQGqIPpF03NgS7NuGPHtNFE3CvnBAJaTtbKG35q/f0K
S7u2JDhSB/vebjz5N8QUL3ndG7aX/MQoVIt/QBaLVGAI6tyLIMCFcK7EdAMrU+aNc3duRWmBD+ta
FnsiRNKUREiEWP4I8dH3B3sygKJDwqGFMBGcPcNkxm4qTrSpClU/+I/NN76j2ZZzpY0aQOV8Tebv
XSl/np7kDzztIeQixrGtFa1dHLCgNtoBNFOPHKTXyGGWUrjg5gP3afsBGqwWBUHTgO2HQOlJLtiF
77AZrlmW3+3vumUypVytDAmE7/jz7dqRDCVD2gykzOxqj5rDD2/gCcVePkVI9ChmEqdoMPXnMc9U
+eBKSMiNSJCYRuCLKqoOZTrb1sWqLKXZ9roxx0CbufWOeT+9vWRYSiC4mCrRb8SWMxhexD2sXivU
BQ44o0CGH8K1U8ok/G6LZcU8Ulhty8X2u3ecuw/g3/4AZV9SQqZL9pyHk27XuHNPx+FNWZionSFG
fiDMJ7zwDIcMzTNGvmwzg0eE6yxhEff3ojBMZMhsUqhxk1gG+oVeF671jPsIfkxySgCit1OqKf86
x1R1AIe3qUKjQiWtE/N0O/Z5q3An5X6EgEHHmeSg0tSQsBkOnfgME26jwZ4ABSs7Q9P1uGJdEt3+
Ev5cfDYRtCRQXM+NA9EYXzsD+mSRGNdCSkZDEZpFgEcvf21DObCttwByk6xrycyzs7Rtw+HrtYY1
1DdRRZhD6J33BYSmVjO0V7u2Sery5ewqKcniQkGgHD2VnU6FVpJ93t83MoPCEBBAf6hd/JSKxK0W
5V8WG82l8LrI+5pJ7Bnidwjli0T8F2dLGozmRIP37K7wSobx1vlaF0K50ViVRvJf69vn87sDuVn8
dxKsG4iropaONGCSajIWqsH0VfQ8p4b8HElZ7BkJomPmpXqOfSIipRteCcwZ4hSMky8IgVQfYtap
Ox+qZCVrhyPuIsOlbt3fBSsRIzfuiOvI2n8h5/9Y+BJnfF83AtHephpkd8fzEQyMtpNI61Rn1Z0x
ppvFJbfcKyxFEJwlDZf1ThPHt4ssfvLKGl993DB5JB3+Zz9+HC/M9wTKOtcsq3OVbatHERNrJEcW
d5ceykRWKAXdpYIrZYpj8mRXEkSf9NBord8px11RTQMdA6B7JDicRuJv9YTYcg1pxhpjb+htHt5B
DxaNJ32TJuGzqQkp6DWKI+ondwIL632JK/ip2iLIOGZz5mFnlDg1llcugYBU9CU+icwL9feyK9eX
wCrBIO7ed3u3O7xmVGDTc5nDwELT711hgTcTn9wMGNNVed0vE+q2f+TvnXVFig0oh6QO25OkrpBN
6MC8CUMCPYL0Q0ZcTJgEuYTOt6hvwqV9V6c5tfjnVtzjsPA1DzT4YfA/U9V4U+OvGL1PP9sufpSP
ySzoOeU6JCjoDEZD0MXWce3AUUO8gKFIVLbncKQgI/qzC6bcYMti0+7R0YXUfHoQS8RJ3vjl+lav
vrdzCenqfcmc4u5pH0sziBkdN520F7Mc5Wwx401U1GqvD75nWmQql/V2GQwrS/BRSVXPotcSnBpx
ot5iv5bEHfumHNMdO5dE50AnWJBwz+m4E2w7qh7S5oE1djctlabTd+6DGJEtC6lh/KRh7u/C3wNP
hxsmHkbFMJpIDeocSnC9pF4cJqa8Q1y6aD8+TUXvFIheJznNp34ckHZohM87blbYUpwF1y0wcLwY
ZK85Kj4VuMYp1Z34g5d1a8NxdPUw1+w2FYzGGlAmYHxPBppPMMUsuXdEI1RAd8Ty2ZIL2TRcdFLp
fOXH0Ip8lzZWDRbsDqGq9uJhPP+gjSuNN+ECMiVsq14YkbtEtQ9RqtfeXLJ2c7kmh39QE0X1N/G6
E6S0JKij0HcH4H/htVzvRJiXJ6Q+hJ6Wk5Ta6IJV3uz1IXO6Quqv/0nZNX/ilHNADOeAzaT2oBNp
8/ea/KaT8F1giTmxbX/uZQBtCtRM+NEldfxjClQGJ/G2DABdMFSRAdDt6obz8Ogggjw07v9Irud2
w9kfk2I6/cdn6A84wjYs9hNkOhe3cLpnAsldLbLQWDF3EE29fvZz5M/sTCRXz37GvCXnN4h/ODZL
tb7Z86IQ7m/5HM0ZdFSmTT2THo2zJCez5ycDckiu+nLCocuK6HEF5hp64G2NklhKOm4htdy1LSTi
OkCK/DYZrHrAx832+ZL1IxLv+r8+vq+jztoBRfbGCU2aLnmPbWT1c9sxcYk4NxtrRBw1iPpfQgse
cyPDo+sUI54yGsPt4acmn00oY7OhsuBlO0Mrq8XQjAziF8Y5/GESVjhQ1Z7ayeY/5XY5dHA3PxyP
HYhgnbtJU5p8NUd6RqyE2ooULx5f5ryp0szNQmO3O4HDJRL2QAK+BTAfa3FYGDes33djDbNcBk1X
GPY4Bt6COwbyAUg+uYTBGx3ogf+Re8Tnw1sBd8wPwt9CXic1e3cLGoZY3bPqeqpqumSdg88IbHDU
yevcnSQTqoJgrolJfrJ0vb/W6jV9qvNhEh2kwIOeABT02/c7daIKaHV5rXVsLJZNcguKZB7t6mAf
KLAm0is9tbtT48EHbDNgRMH09mf85Vq3DTnWPeAMTcHycr5CMj+NOp8EFhzRT/97jkse7IyXzM8W
+YVT6n918m7XlDOanU2OBpq0kzDkm6cqcuS72O3Vm0ZM1gou4VCWabWnommdCckrL8JaYtteycM8
hCUWACGV+NB+J3pkUq44dwEXFD3FpPLAgnueUvTtmqkg4mMKd22vEfh6Qpq02m9JeqbNkpTRqbTH
d+x49YxxqDd20NJTAinsKt5Cs4xmoXtsvKW/UoNQxZNlCtarWQozMIhVgSP+AxcnGx5gyO9UnIPH
gDRnwbNzR5PK+bK8OF/v/ZJmStmvmsB4rGeeCV2liQWFqXjsXfYCpCPd3v+4VV+Sz/+eLQ/1Q1Wh
wMsXCrsP1hBC/f16ore8ylGPIkREIqDq0V8jsca9N2Rk2W0JZBFJtY22xdBgTY+vOpbdP6NV/h0J
zyMmYvK8UjlDbBp6lbg158FlGkwnJqAwrS5dhR+502vXWuvQmfNFSY0ProG7ql6Bue/L8ZIpvVDr
vSgOza7qEjpbpmlHK6XzypLDSx68aatb2DoD2TJcAr0oD4Vxpj46MTN+tsS7+OwY5Gjy+Xe32/Vj
8/sveT/hjPb2YYOTn97PudFFNRg50v26hzP7c4L4uH6xJqSE6ZPfROPq1WiIdWIxx+zlEktdgOi2
VQ1rVzdTHhXcv+rO5QyynJyzVpwpEN1sdknc1fMqs6Zij6Zn0RAxNkW+vxj6saz8gG0CphHOMg63
K+bhA74dy7VDfH4rRgWdnOMZR5pixIA9ghheoOYZMShlHArEA6YTPNY1PSw6W3KX6z5+qESMyzps
qzg2MGu7fQw+m1my2huefQFZP7ZdCLlIKYz4uqk4YrjSX7FxWzl+XcPpWy60+idRIEX3GV37Npgc
ALUGpN5aHm0sPzFopXT12KSx5oZ9hKp36LVhaU2yjBP4BLY1Qus05WSY2tC9+aOEcf0htzUAb4es
2o3tYZa4ICZ1ppkWHnVRPW6DaRKmarHwNlqI3FBlD3O5gYU1r/UPHo7IDbIjg4GaQNCXGbbdMerp
sE6RbFEkYJbCCCcp19vJAyIipSjV8nSdT5ZvXMhQmh7FFkM6gVTnHGOoZ9tqok+3OfS5KMmG6oaZ
CdIbZDRhSIK9ItvudLcS8SL/ju9489HAtPOvCiWq5CwG9yMAwucubw1AOL+l6/LGBijjMBaEFoTp
CFOAaIiqSicepKirgm0LXe0jb9eSP4M2EA/1/QODpe8sAK5HgjeIBAkzAhJCS+X9DowNDKd4P1D8
QxjAU+y2+qs6xGqapdbSlIxLWByqPE3cvOPmfwimIfZ1LFiw5R6a0tcURDgCPlY7zLP0wN1GY/m9
5alcqwjSzsFhOtg0a1IHI9Xh/MtzTR06BHXMDMYfSkSlnz+eUngbslGH+3hH9B5v60BR9CVshLSq
vdqzNEWlpCKQRC/jlimKTptgsfggpxOwWpqVgEdbBB4KIX3jk64n40hv7SGWZWVK++JHShgtY2X5
YTwFPh3svVxScKE9Q28qJVGwbr+VloP+nLMTKNEyhsqrm1I0qfqwaICATMgS440TfVnGFBW26fba
i3tGZT+kNg12VMSUnHzl5NDTBC1O66J6HTKzmYTQkSEtIUwZzuMUP1Acj2z5vZMoIpGriK0VZ1dW
UJ+xdWlPVB+ijtesbaNO8hAPE2RA+2BH8Ko5Hx/ZblE1us1vl/YWm0jgbQMgOwM2zxsaok4pIQtm
c+GCkaYhbZYOj36kh3R2/SKjllbPHGs7VQ1pVb+Hc8BLwv0GhOWrrcpCgNVsl65P9mcqtIMHOpPM
4GIfarE8Ads3eXT6PVZmYTYpwladC+/InzsR2I+qDp6D/uUrqNAmKcYeDEnOVdKd7Clk0Pa0HrqN
wmgC13cYgXYZRPYPzHPQ1I5chi5/iGEl+MhZAPYK1jnigieKGrgJV8DdcbFrMPyCUThFvK6CrXFK
BkdXeV5g0kKK0PA9hneBmMEY7TiJJ9yo/vXI2FKPpYldnebkJlCDwJV86fh+ShAw+dBYnbaWQZKe
ZWrOyagBE8AZGWgKBgLoJPkmFsmJAutNCqt0Y32l88p54T6J9Cehf/atSFX5dyRXQbsLHmQcQPIv
m23VI2f5z1pQIDcCIrsPzGRB52ampuasMpj25t4hQfgtQ39LrlWJFVAC753naGRhnT/zdp2J/1Vd
ndfke3pEZtk82sUihr5wJy1f6d+pSVaUZ6/Bv9gN9jcPxhDOffLtd/UsZhle+oBka1nbO+nCJvCC
nnOTmo9Xh+Lwee6Y4naXvczVo2s8PQ+EIXD2M7M/maq2MgNts1IgDujksV2IJfGv7DijXIl8D/wc
GYg5gur5SwzKvkaZk8Gvpb3fUBG0gra+VsEM/9Y99JrWVCWthoq5RvYPkI+loOPaSwjkaexqmdB6
h1+qqddY4qw8Bj1E0o2ZdXl8x4VnDKIUM6qJ4LrvbO3HIKxsihogYcsJp4/biPO3mzlpTHCw2Tuk
i+76EOIY5ySkMEj7oIDw+TkmOP/nXHuX8jlqJKmI1okdBvxn2c+3r/SG6OjCpewBPwC6097CFS96
tRM/MBnwLcaazKItt9e377vn/qdVhUY2A0yEeJPX5CcHur97NNALaEQ5QR2JHTtr1Os3sehtjrVg
vG4bHjyK/4r2rvnFbxZXAJYRlLRmLk6dXHpq3mPRwNmjw+gq0PEU36ATzY5o4w3OOXIpKpO20klA
VR9q1vsQ5OSe04keSRmzuTrMskYlmAENRPerzb2oFBbSf/cdsf586gMD6zP9C6RPZCl+gGZXtATV
NpeBavPJ1GP7a4awa6AikpvwaFnVlnSWR4hndjh00Sluyn5dqmYq9G0pgtPKf6n2OtuTYOYIZr60
Yo1lS1Zd5BZlG8fP0G4RTne+OP4E3ExKb0NyNsrzum/wqqmppwsxu0RoizqvsoLODPZVCdtSJeH/
Sz21Cb7S9av05Mcg0PbOuhSZXDpF8fojFBGuuoYdRhpM2Hjy7uV18rGxFn6lIaAmOr9vSkgL/YgU
xTQKYWQKuQLruQ6dDjl+1oPA/Y2WFZmrVGieLSIKl4z/awlHhzKRPHnHHJEAdDFAXdncYgVnoRya
AwE+6QsecowtlbkNwp5SF+7cXuuSFQLfAOIE1TBUGVg3nhKpg81q9IVYL7ef4XrPBOOgRTyhLH7G
FWAbEOZI24rNFpmklDfEU218vnpDnLSeLwdvQUl24ziy5TgaQ6L8TTTkop24nx/hZhA9TAhvtdUX
Q1g6YOYmeqWCf6A8Jvxyld34zHLYHciSHh0P0p0TWpHmEd5jVNRA9eLNaa12gsvyOrOiBGvBBADX
fThcUE59tfuZ9AIiANMYoDUwlq1Lyx4oXFhbfncBN2WBeJNcQAkFG/hxBPeHS861GFFDCdafCleX
fNDB5tRiBvapsi7IQYw0z3MsainQ/xesenrCBL9nvBzr3MHNiw/MkRMaizgq49bHrrxaO9dd5hLy
cpXsSfxlK3cIA6Z4xpKGNnQXy96fRS9ekJOeteVLBvzXiUYuiuTnqVMstSYn7XumIBLs1oJ5Nh0I
hIRsOaEVn98J1jHFlkzTgcqOybdxFtjKPUAGOpeWFQyzCq6vlyLcK5WG/1nH7UXJEVFhT380D8ll
WSafVDlTbxmzGwFLxhzDWpBqBcf3k/lXBqUb1cFmAGkRv/2gw3ew9g1SRSVw1m9x7/feJl4okfpj
g343X0Iov/xLvRd02ijwIi7EiHBMY5BKG0nxsRZ5vhCst6NqgJeHZIjbPy/+WUE8CEINRk7/I4sx
lQuPvB6MxGYnuQ2rlxAwQZS+Vq8EguSoyJYIIcIk3fmrfv1xwDlWCu1r8OI3VYpIimkndP6p7lqc
0jDuG7ID+jJ24hbjaXJ08bQ8iGELI0X5qkR8+znr/86IB2BYE2dNRLv+nnTyHcdP4bDQ/yZ/on+h
dSN1i7+tRaWj1Tf5wg6YFiSQXngnSbcjkeRIrneMAeizPZk2eK4eWmqRc9HJAR5XSbq/RJIoH7T2
eYrDz7y8PZrkd8l/e7eoyMBivsEMbq6u0MnJudRo5pttdLbQQjkAOaEG2zwS9JYCjSxeqS2+B1An
VwRH+HMiEv+61sPI3dsDi5Oe505PvPd8lIE3Wugiz/7/UG8WQ83c15HfpO+QSb4swq28kOgDpTqE
GhJScqoiCLiSFD2SAMengtMU0MN70kj0olLtKCr+xpcVd8W7EIUtKYNNCaO5J3Ca+dE3D7gyXBRx
HTkWKe99MHpOsgh0KEIm/JWzNGcFTfbngxeqdPPACVJB/kAbV2A4pucd4ewbyRwVFZIcTaUFxrWp
OY+TQGiu02OOyZPzhtzcSScxdNFJo1G1wAWJaxMdoKLxpuFpZlL4WMYRzL4PMhk21qz1xldSeZRq
/msNGMFb1RoZWOp/zdIc75leAIyrH7X1Dufqk1roNTxQlYOYodmejNKga6JFE58E6FiTdLWpkUvR
5T668BPipqZTxWLdInhIyIF5FNAWHmEqOk9DPDWHuz4OutQT0j9BEVXgrjqMZXHqMVJhkKvAeuBm
hnsbypuNTNb6ljl2teIxFofJmGhmk1o/NnelfpK7epAIQd7PPqqP6VknwVxPOIKx/r/f11oE1j47
IAMGTqQAMG8o+zzQCbH94gf9Rv8Lofg0d8ALHdV4GwLb2VpaNvpLyCtUbiIrx6yGdIRfqDyXBCmt
xNFfMP9sIBumOzFZM+NoNX0iGcX2Idl00m3inlkN+Qo1IzPXuXq6UDedOCPFZj0f9or47dXY3ZL2
xkeYfM68VBUApMA+90+1j8jeb5WKRRH0zSuAGkpGUmegj8IegMohryYR+Y4gNXP44yKhncpw/jHE
AGSwKrn9ddVNtvu+M1X4T/f/ZQqpfB+PmXgC3jKkjJINEq2QvXV3s5z0/iKx1mvhHUJju8bqVhdO
SVQKxl5uZMFunF0gS7qbqRs3TwG/aQLQTZVqQ6fgpR9UcMMDyOrPIAZlP25S2CKEi4qeUe7LRQxq
Nw7zAnRAMJc5hKxSeuUzQjcloCNBJpX4NHz0u0i/ahllnbccr5103cOoYU4lsSoLlhWk4zvTjtGv
S92ngHIOrdYGwZp/UfQkdFEUMkNWE/u+58yP/v05i+X1xsF0pO5zAc8bp2Nd89IbnuRmDjjbevnv
EoD6c5zr+B/sRk6+kFqox/1ObsY8+XD0/irMMtU/UwVb5prR/tSSgBAjZLwguyBe30NyTeaPKXwQ
8ban3+kAb59tV++Tv9PiwsE04WhqvCve+xivdjpRw7Zr8aYR+9nhzbCnZ1XZe86gjsPkGPCTSV6a
kVsFfvhszTcOlL8BUDe0DI6iE6uPXhMbhEaWFohJEZIpuNCjjj6hPRCh/w+hXBMPB5EuNFbnkR+7
S1Upy6mvliRkWFQW9aP8GwEsAgYLsohzbehsCKqrXpOLVNJoikzItYZe7UkJ9ZzPPXPq3kUav3lC
sSt5LoNvKXPrcyoUsVRi56BL1ihPxYeExBTxOP/0JiWUa8IMkMbwLW6LSJGWaHpUcT3IJNMl5u+D
V+cHnpc9O0Z21oprujLdNXwRY/JwLW1IfPVLVatULEGuN9mo5UUiTRjvvZYrnzSR7JGBQovFCpJh
QyxIwHoVdK0namdPkvY84FCAEVql9w4vj7mkreu9c/CY8fmCqpFmpSUoASWXR4IcIpslXxp5Fynh
oU1+JKQEFPSPmsNUutqQiofciO/3wbaFUM5lQN9c9sU1OOMLrQio4yPa+sUMcLwhU+Wqo2nN9A9P
Ro/E7NEBOTm2N1A1b/M29YtFy85HzJ/RmStMOIxlZkTvsf0SGfzJQ7PIfXoBsadvg973hf+p0zAb
mEFH5olCA2PGuZ52SEb4fTPskUPnOWKLPOlS4aed0Zh004nzIQ9gxn88LYI06rVaW8ocZud95lEk
q4o9jbmuAwc0fbK4cnpdQml9hbOzD8JBBP0lpgPXFATiaoPaT+nrYD1hJ5Fi5FVHHweuxxQakm9S
GUpDe2qA7VyDTFGfZi2+S8hCQW1LiLZL2Etc3U3QvVCGxR86j3CxRVQyjACfWx201wzy+qVuLLPx
SxmMoNooZvCc3rjYlrYzY8hncPp2nK2I9TTwxv9bi8IwoiHUFA7BWq5NOPtVjjXT1+iTfymXEKUJ
bvvDkEEE15op5JirztFlKywmKI0ShWRu9t9BkGKjC/qO+7hcqWYXxMH6FnGsJ5QT6N2pesBpOPk7
0gZ3G40K9rWnaJJuSdZYrsTBWQPYsjGP0gqqsvCDhvb3MnB9PTCSMYUvVqOEpUyRYocdln9RLuEx
8Nu3CrjB6kkORCbuKabvpK045m1kJHkzHJHH9moU4ybPAkfJUfSHgWY8j4it9LyUHOT0Ckwah6hx
041K8OxGo0F09Fz9awi45Bg/+CZvYMwRbv2e2rEJFe5RPHzl5MmF6yIkVzJklqqGOkPkzQMnu+75
ScGBtzN87JWuhhugalT3J88ImDXk9XP/S3bl9rQQxWCZu8wzvuH+1FEL1rJVOjOOzQyqSTwZcLQA
KnUK85ddYYz8wNKTkZQ4kKNcOguwlZMknm3Mh0rEsneGWJCcCAUrnBnMOXnHCK0zjKstyncGHJPo
db0E5Ynpih2YZNRBBg1sML/1fUn53ZddBOYMzQ3/bZhYcxyT12KLPI25/WXGxNNw/ukWmHedaiOM
xGyF5M3ZX9t00JjCtDmnzrkhf12sKoHhBELnHV1/eIRV6ani8BNWfVnNS3O5TDAFlpAMgNDzo6Po
kQqWzj1ISNJa1H4EurvFWcE5nhZ0wUv+u8MYEQAQWbIU023eSuK9tsYJ8iRghg7J8iO5lqYHwElm
Lz40xn2D46AiZ0J/1ezfyAki18vCpE6ZDaXpbw4Xb161ifQnLI07667DRFD9BF80KUfaL6HsAG3D
TDhozcqR8NccgTr1ZMjPvLo1OgbMEPCZ/oD8RVb0rhBXzxJI2pH9EYxVhQkIYa/cfFHNoxoGUYXb
Wz2HrNWCZWsWYUFIiLV2DfMQRMkJfpz3jHs+7AT0l4WHXDfMzUwphHQryFg623jOWXOH4km84UQN
CC2wwVvqwx6VbypxsuUclIEYOsPgsYkoMLZOaLPizfLCYmW5cQKGYF0+tNktPgSFkA7eTAutag04
mqzef4Utno6JsB2msDut87NssmNuyBSBVYRddpSJimSTdROigHLYGowHvYOvSiA2jwxn28CyfAxa
CbTwQp9QYovF5Uyb2cfSGBvVxRPLZ8NfgmsNxZ1vhfEcmuMebllnMqxGOSd6BRX0V7bpJdt8RgDZ
UfWYSj+x55FsWk2Hqs90EKH1Ospx5UaoUIET4kRfSVx4xTU+K2vUNFigB46e9hOpHveRV+oUsu0z
xNGVZMHq6HmWX4Devr+Tm9k/srjjrvnV2XCkqgOfmAp531djr+2TvbV9ko/86DtC388x9CbN6kLS
Y/wycgf5va1QKoXBRSJd5yBaQSNz4Rv7MV1Y+P6v90iD/HoGgOFag+qJNC9g/RtIfcJ5G041Z4DH
x2I2nBlv6HB5+exfczUI4XWPHXQs+iIqaGtyrDDXu0L8c1pKYtSNH65gZVQIEzCca+nwD2SuaakO
zepUtSgO9HjuuzAXx8HoD9wqrcGc0hd2qaJvZLR7UchsrkSFMxNW2uITO04CPcwpkGAeK6dzfb2N
TA+HhcZ5WArNFuXnILWAf/7AgwuxptA+gwC8WxHSfHZ0OGXuWRBOO7Ah6Xyv2ErXoSjwVflQowfv
Z2DaIV2qFRmNjn00Cx2qwIkJfwNbpWdKi4FKjyF+Hxlg6kvNhdJbHS/VZYv3+GEDvqy/SZeWyZrU
6cublbXsHmAS+K7iMHNir7dn0SYDrDGECrjD1jv6ztEj3V+uZWSkHr2VfIlUwzLlK3l4XndiiiZn
ST71mUATlafx/hOR6ZHZFA/d4Hhcl8gnwvE7lMfw3wb4AZBV2xfWJDRhGtEfPqZCLO8tmFfd3Khj
jU6Lp+Nejv+x8hg6nF/Qk+c9gk+MZWibN9XFVcAwx6nzTxmI0YEECScgeTJjj7GMfb6iLWcII0FI
lVRZRDHgSZ4YvNnRmSXRHp2iEwuKbsYmVO98xDN1dz9l22qIj55il13FdMOjicf/T2CG3b0Azz3q
vt/AaCIX13vQDMxSsIaOsW+g7Yj579eORxYY4VwpeyOe8mOb+63KMAc031NdgCfvG/wE8DO0wkVA
oWBGLVX4tSBIl77YRYmu4+rTeqOWzGkQGpS2UJc+AfB2vKPc2vxpMp5PaQFAs0yXWT/A0wBLbqDO
Kax6SaxDsIaN8EtYNRKcTCstxgujlLpQJCi/bIjAvnnXsdD6/cVo7SlrkvGMDvqi+Ah68wkWbyi6
VgbOKYR8ZI0fb/D+6F4DcUN0sDZVBkavNRivHXLT23A3yBna/x95ZNMW4nb7V5AMHb/cPqKttUH+
h/1K+ub1VI2RNmDUUgyrgRg5vPabIY1EQVIcIi3KhGkR1fDsrIcrDibAkjhP1NkeKTQ1bwQfby5c
NPRoW/mUn7zSetZm9cCC0Slc4FyIgZtz2n4yBsnCKQ9D+dB0oZ3Upq1jkxBtJRHk/l+xrTdQpuZo
wjxLb7iv7zQIGt8YvLQAMajQbugn54nTPJ8YcF0LoWFLOlbUP3tpalKhmPkSd/zB/pmflX+vDhD9
dloKTQske37OBsL7LuX1QHBWuBwpv1pMqp4PVh7yP+qIL5/Y/JCnaazeglpPudjLLiUaw0WhcnAX
sMmt9WzXU4AOmsjldRAtTHbEZkoJpSzSF+oEd+DGKbQyLGG8VgE/bOwzxhAIECSEFZtvrzgXuFBJ
M5GObO88z7gelFYnV82vIKNQZWtgg5CWMQVgnExzjELlAOJhW23/Ogp99uwYfb5c7W7imelaY88k
XEqgkCu9qnijv/3kIVc+chERCHXuuBfeANRTDgkLT28nYlSqgSexEj1zD7AIu48EgCNxzYEynP11
MoZSFz2ruVKZAnpsIbO6AMmw7Y+wcXDtncdNw9s95oAuYVmKR5owY8Z7b0jCrCJoT16Rj24w9QbL
/R8ajEYDCsnB+MGJeN7tTX3O9c0+D/2+g39TVBmaGqBUCHF3W+uo3JvL5SRw/ghnG0lCc5R/bUV8
UsEB4bGBgZv1b0VQ7F14CUGymY6EMFnKmxApBT62/SFJ5IYnd85PeFEqJRFq1dXNJCcSzp/9sGC1
E1vaOSUZHCMB4Sl1jiw6HpsgOVEQZwVy/8/vriDu3vCGu8xp3u5ZmmxXqzSzwaEKfc2Te+T+bCnV
TdrFV4kL6g+yOxs9KGi8WGJNjyv2DRhxcN5VHC6WS8PeZl+WSAUADlUeRn43iPj6sN7vABK1WkMj
10wPGpbnUJKSyVWBC80TrQXETjVec9/RL5TwFWLnNAS4MmuzbNSuXtzPfQiETymgvGOSI9+39YyV
5mjgR500g4Ac09tiMVZZdpcA9tLw1VvMDXJBpUNSV7A9ArrN0OO2b9bt1pEV3gTBa4tmfAxmbhMs
6mwy0+wWq/R2E8O0o/nYa029+CJfPtHat93ftgKqzJJyEPBlVcnG+E/9Vr0aO+29ys2/kvkQav9N
pAys4VoxhgOrrN9UWRI2yVWCiBAuOzzMz+y8QVhzbCGxMqhp2k7In6MUKBnh3SexxCR5c461IpFT
RbDPJvr0H1pJ5TnZbDDZ81LX588eways2GjgNqe4phHqhaQp9jKqTSOrmRJuR0tnNxTC+Dr4yYpg
7+sQi+R6oYgOJSPEdKYC1rRsscW+KgCiDmdNoYh36Mb3BYYvQnEYR4VTvXoPvysGMKiHPmhWEcC7
juhQ8RhraaJ/8h5ncnH5At2xoe6LsWx/XWbRJv8VSfvFqvTUTycV/ymm305aQYy4pf3AQ1CUkJi3
HMcQ50t65Dk4gDpemhUbaxI7VkOnAlfpnu5yHHStw6v23srRuPEpSk8todTH72I73ONTFZ07oPAU
DrqjIER+IaJU/6P2Mk3PpUyUWkkaZg/OKJx8pFlWHZxriGllzypBQC3uqH6dVOHcaFTAN68ytqOb
dfhdJxc=
`protect end_protected
