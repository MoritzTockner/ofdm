-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
waUy8KgdvsJpGD1K2OcFtyQt2g8r/PKqqi9+1DAW7KQYkKArUIqdJJW8mnz9i8/IcEx1nEXS2wq3
BZgJVptZ1t28KBpMYJMrKrEQhQiDHLUQR17QfS78eLacdRMoaTyoGXAX4PzEBQdakv9j1o01uMMi
MPzhLr/2qbBxbnrwCRJeMhDh06rNhm1LR89LrcBU6q+UBKGx0cDqtOpb8IjsBKck1q0TlwmBLq6M
5ps0YkyHreyyw45jBC1osDHKwqTt176iYBjE0IivlDa5Pk8NpHZKsh7x+02vAN9aml15EmU7IOPq
mhoxVuTuvuqjpW/r0pos/mH6cJD/FeqHc6zdKQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
toJfNHT3qIzqr+z86etOTdteLHjNeb6z/QDIbr2j07MXvX2ESTVhgOrXPdFGAYFG+EMj3Cl1GWgc
Rf9ndYNuM9X5zMbLttqt5nH5AE5hrcORr1B9M5TK0KopgQ3tNvsvCyLlOn0fCaqjA9MGwQLuQvrH
eqEMAKlMQistNn3Ds+Mh66tosZI69FJpHwLq2NW3mAHhSGWnl0ZTEBhKS80PFcZqIibbI2MG03GT
OS0/ximSauFFvIXsWZ+aLz8gjJwfHqcrrs0gMzFF4td2uJ4h8zZjHWfTO6dOjZtYzMG2eDI9FfV7
TB81frfGkgZ3UCev6RdKeVQFFTJ+9oCwvF8sfE2E8ndd+sLLVWD+a1bvSHqA3sxEX7JfUppwhYFW
ocqF+JksxLu3jqKbkt0evIAXXb5ygEyG16/QiCa5TPjgplRj9PpK32vi3ovs5MquxHBAHj5ReNPz
d6gvzz68FlBTCw9WHqARn1VuJqg+HoQFmNDpVrwkXv12OcPad+lVoVfuYH0NnadUFV4LUD5rqnXe
WbTMJ2An5/2THtEmniqYQ5aTY6VNDpfWM8uU7EDtTeU97/plBwfpmDHySLA2wHvdJEBZjwzOoyA8
17hDPZqb73rLPvhBl4vc2hExRDK0C/Pe5TQ/3rlr+yhnhD5F1TbjJJybyyZf56eYowaDOlrdC/Tn
vzvs9MSipRWU1BacWlZqJs7Adxw8MVGx+rUuMEju7FsrN5v+HQW42kL1B1LWdpsNpjJ/fb3+ADMs
8h7BjsXhozEDcw9UHlvqapqIhdlhuwZIcaTljTfZEprgo+u+q5bGWAzlut3lU/a99FTPose2jk/x
lM1ph3TPnyb4tiqfdhPr2whYE7bUO8rW+DFnBayG7LhgZB1K6cgYSUn7cgxKjfX0cQytTEMcTifR
Ob/KEKuaBccrhyd6xgsUzt6+JfGkRa7FAmZQGonLXX7KOpogUZKy7/P4NHovmWhq/lIk1kr6rJ3J
KtY/SVFfeRK5THtbGWw4oWkw0qo8tuST9/x6JCfvVkpxXlitM3vbml3MHPBvwEuOYqq5X1wExIog
F2eHD6sROxBdxkQTgwEAm1nvkuZoFXwKZ7DtwQG1HI+Own01UEmENcADGdN4g1eUb2SKflqaRBAi
nvp8WB49Suii6ol7mOATMif8YM1b3xDhde95D0lu3WomxyRMmlXHJqsSuBCEhQSIgs4/21Q0tsiE
gELk44Chsygx/qppfSgqkR9WCMu2UnKSeounB7hUiJMk0YbBYrGE/qwIsXhHj5N4YCWWrKsovLPY
AD/z96mJfVdTzhJf6X5m2nMzAZKT/7ubg0zXypP81JvRh0+4GMNBzypU75or3moH+0WCLOSPgtP3
6ab2AdMjIVr3CXmG2Hbn0KfqK4fCgFArzBGynjmcKJRKRxx8dpe1DxECD9qEco8JIIJs4P3H8Ns9
obPzLeIZWYBYHZLHgwk0FoqE8S0nktFmTGIHI+C0j8rnOIJe0SWxEAnlY1jot0C+oceE4ECZTNGJ
tAs1y07Pk23JW5yk+cAFVgZ03t4+hva2lXB01vmmWaYr7MtPwHUqv+ujW7wm5q62OeztmE4B1cIu
FMB00ENAr4UJixEwVmrKPHLY3FOsNLAUlaBzsl1fNjqD30HEJv9r6BolJ8BsLQyLAGiI6P3PbHVM
0iFcyfD2MHe/0VMC6FHVN24dftay8fSd59Bq61ue/RFjVUIVQX09MWH/Duoz87kl+3NoivEgqCzP
vucmeCjnNZ5Yt7SJJBmFbhEIp+LJMBh8xYFEyuLBVSK0YAYlP9Mfo150cnqn88/5YD3e/fdShe+E
duAXN8bI0gq8oTGtY21S2cSPXFwEB4L4oo1hxAU2BH9T1ahif6XnuLdUBJavRhLo/YlhpbPxh5h4
a8xNM5N/kl3jKbXtQH5LTAuiBb9wupKt4LM+8H2xYF14TjemVQxrnMb1jX6hwmN2RDYIXC5XhXm0
pU3gph5rb6kAI2/VNezfdQn43Xp607yskjHx3TPw9+bRE462ECmJXgHIGmyzguQyLnvwhLirXYMF
KpffWEoQU7VrWEtAIFRXaNZPh0zaQV4/YOpx6CjmyaXUDpcDFD8CZ30ja83kd/ffRY9wMdtRQrjE
TdzSnfBspnmsoqscpdcDt/WcU0CYU8IvuB+mBBOK86+/lyjbw8T5DvCOD9hfble3LAYmiAezOzfu
dRqQH4BjKRCHgcp2XHW2/ryZSwuN+/jBAUICZ6bmkp16RoNJkAK79DzQ8IJejnrigLmmCaz5dRp0
9XsaoWIVtNebVtovXSivxGM0mTG+SvwfBsp2uz++DQQnzVTyAnvMqG3RyJPWl+oLvLmbJ+jVN75K
S3Zs48xLRwVqmjG/TwwqXutChhFzzV9vb0843sfO07aJ0BzdhB6DxwEt1zVDiA1lSJrhI+ulkRM3
/5zp97CSWjdHVkLLbues6dTXHOi5gDhp1CBIiFCb6bxgvXQ/hR1/PocPWZp9TNaRU3hrTkMeaOKe
4D48BRql4LYG0fUozjlTRXpPafDOTo6JqZ6SgN6vVe/5oHQc8PhZSRHchlJH5Ea2wFRjWoFJOBW0
cV2tklRT4ekHakymiEL2gg8D3ruJa/p66toaJX25vq2W62ZBBAwfHdRWPkzZ7nIHzLxCVxGxlCUr
inYRyn10/GX//s8SsbiUmkLejpHYbE9PiqF6WIRndoX5XVfaceP5vrXyj9MyaqsfMjW2b4VJ39nH
4EbHRPZ1Z4/Xpk8pXhyZLNZ7DGGOU6hHWDjpTNNbwoa/2kQS3NxnP+rA3SuxN0JyB1G8h6IjUG67
JmtR9djAb1SEIQkE6RXnOW/gHi6IX/ogIe70d7vDr9oIlJ7x66BH7sw6VTaG1puAZE6IiftssPQH
WJn/WpvnOeeerpVmf8d5ajLwMgl3PmfyXKBsRGP6G9Dhmwoyh0Rg097MbK0gNZwZL/oFHPfmr7Xf
x517WMihMoYoI0oU8P5hh2GVwAk8bkRUsT/0krcxLNwWh7jEtQO1t5qWXOkZfWFTeGU0fM102us9
NQfvDG3pEXoEPNU4XRV2ymlxt3Ik7Zk1VsNWFW/V5rBqeIOkgMr0jaMuTWMDZgTZiUw4aWyG8wRJ
lRTq2ysHIidMD9ZTnS583x6uFLiRwO1tTsB2K79u3pWPiuFCxuncAo0cNhU+jLiq7q1grK0XNhEc
hLRMzh8REpdqYRAXhLxECCkGGKMduMzIS4EZPC4Xmm8NrlwxHW2vO50LrL9Ck/d1sDKbCFSWXk5Q
egLqcE1SBzpBDJWtkmrmU7gTsUQsZhQTUqgTjGsyQmmJih8rnxMIzxMWFcLDMOa5WwXes/i7F2jI
7a9WbXKyXRzm3hOvawedpxAheMsD1vhiVQ/Q3B2aTMPA4GtxCRQMjFwTT6F44+2RwUatogyBuibG
bBSVXFVbBN48B/UQHero5NQgtL9CA6FOw3pxEtcQIL+Mn6M+kb97JhmFOuX5EeoOevGwRMZJv3oF
sibgTj+7jvn3SIHtbN2qIB50a0wt9+K09ZfXdKtUHdijLSUxgHJ9+by6gZXrp1AMYHsee9WAa+S2
dgQ+DfbCXN7vHxSoH7o5BDgMdzV4LUge4CeRsKiyS4wbTgqMpJV/LvrOfofN2YFOn9WyeRAJ89mF
HTKAtS1AuLxm0wqf0dbUPE2iEcjbyWWaWwgZeBZkLqargcdBlHjyngakSsKdbNQsaNs17fJow1z8
j5jGDiRumpk7mzjPqE+Rndj3RqLIVuTqXyNt2Lif9QKQ9lbmoqpHGt+/H1Vm87WdOxJaXRBgja8H
G17YvWh/f2oJX+JaWt2gFIv1dKkrzPKP1Z+819sl8zcdaZhoa17oqjHXDDqv5xAORLVdRbDB8qF2
mzY0RKoRRUe5xrwm7TcJjsE5zJJRb3kpWCwl1iOB9heYbT5cNKteYVCcoJcq7holw71d/OirnNkJ
EM2Agm+wlAtBN9SKzrCh6ObM0E5aG4SPhS3XvlgYOoFib+FcrgX25k+a8cqcGargqq0KHZabyO8n
VTRAu8lNScfBQJvTYavZmLBjawUEz9CanG9l/ka8a+rYCGWlZQLSX5qe3VxRx6oydVJNdjysxem7
NixY8c/Jlbsbu6/9v/yiUdAoZC6X9zuVU0C/Cb2HTttX0DwKTFg0wWQQwTNcWKsD/+WOc43zRDME
d9LbO8BQ3H/3H+PYaaUUSttKW6wpGZGlGmv89lEFEfOrfj2UImaMP+I97u6Z/5GVRjubI3wEi8Zv
Sf3VXSM6WFl9Q6YPePFDW651viJgCPjcqwomh956qKkVcZq19XefQcT0YbRFVAeZsxhCbzrA9Pv6
02Q195Z9+4bxcD2u6SHGrpXdVhT+zivWzVDS9WTafjwwFIyZRf+0Trz/ji1ZaCvrFIE77I4S1pnm
3w/iV4E6xPmEJ9rWxzCD4hxwfeAu9hRaXQJYO2MhC526aI/RzYW3h1UlzTd3QruKoLi8LrvvvqQ/
owJmeDH3fx4Csyzw4Sv9LOle4+tl+AWechqj26DGDXNUmU7xMcpCbpxHC4Ncue+ggqZwZS4+Mn24
ljc+yyA2mnnfElQ7tYNQyuqU7EvZqQMun3FbmR8QuHspj6pwuOukGyEmh277kiZiQpc2CZyVvO7t
wOd+V36+f4ZFkzjds1YkrRoZ7DZs7sdtv07evOSqB2b+jF4sXH7P/MfLG7qukParakVVVD24/Q4+
EnnA5WFTglj3XfxHZJ2WG08p1g3ZvxuR+t9CD4L565h4yiwHxcXUSNUpiva4Ugr2RALal6OBQMBq
Y+CJkYrxgECreS5Bl6eQR/tFjNfRsk3g2SnduCOsk9MZhRDpSrjn1PxEEIyMjsLkNmNF9PpRMZxV
BozcedL7E20xZ+ayou7XJi9ZO8ssOzZWtQ1+0s15jiVl+s/HvBadaIKZfZz2QhTOOvMxfaC5N9hM
iazjFelqmhOQ3dmgSXoWa7grl8NWK0Yha/FTDkK/QmBEwjsLJ//wU2/l/6KPw52i5aSVhPxtRmDf
EY+gkrqYyp1HUcuS+PkvwTndPb3qJAbEVNotmdH4vvHUwH1ZEH1HbXymnrJChqzsasgfMdKctQpj
YmnKEnnieYq5B4Rq0EL5//5YWjd5JezNQGzsU7iM2xoFbR/sP8wP2GxtJ28JzYlPGWAnkrZS2ZR6
VIv1tbbKnPdMIZPWUkSe31ak5xRk5vZR/Jdj59Hn8BE7QjwybBD4XuT7voVrAr/Km898pIiYtrZ5
hnxXNV9l2Ue91Uc7AJn+7e3uAIkY/EomkOvq5GSaWjBn0bYD1b2DX8VSSACYnMqF4WUDnCINnSP2
3AeJGlFLPx/aHazeerFArY+aT99vcbTj0MbGxFD9U1Rf7Qr44yNg7xT4isPOLbLZT2MTee1mnhFl
ZeAZHiVfmCBpzUyw7zZSrkdE2dfw8OQMLr/5oUnNQc7LS+Ftzmb7rr//EAOMeeqFcQyJ33gOm7NF
4EBzSe9PRVB/ByF4DHGkOE9ky3e4MisYCC5TiS6UpyG7N5flZ9xoYUxB+fp0kQqT8TzPJtOHH4Ii
6AtPjCvElGnZLohWSzfrjFnYCMZ3cvzuXicxruhwLHTDF6qXR1c2HO9b4jOFo08e9TNGv3dul2HG
1sRna1f2Cyi7KTHAy6zn6ClV9dXqFY7AThQzG7kaDX9m5vtISo4dDtDv3k7XFW0OgaFnPCVwfwPW
k2AqLl490g3OQzx4k8t8UXoR8o3OWQvioozkxkhg9JPslZPwJkDFlp5Lq5Hw6k+fNdHT5iUqVcah
RawwAlb0YojAr5hWNHTH+F9cOeTqbt/vRxCrMJpbdMTi8yV2rHwhfMW75RkPa8PueytQMHD3w2DF
FTubtUWuR70hicPvfn9yAdAAM3EY3BpcVfp0JUU0qem8bm8lAaAaXHXfxO2qWEktnGO1Yr+VH8QA
kQvfky3WB/VzyApW4XNVUzaU16yNAKn04yDMSFDkUi+F8ANrw2n1TrrKh9YI21e7McyJT3Y+nCLa
3zKoxBYHu+k74GhCPlXxwPdAsugWpXDFf8eo3OxX7A2hITDF9jt6XZuyZWHI+DY89CKMtFu2N/k0
D+/KWqO9CWEbUbESwbzZ0tJUsRY2n88Ab7bideo/a1i3hos39VB1rcjuRz9xYRBpIYOcsZk5fD2Q
ciaVP3wwqSxCr5ITJyjTUSPjoynPuN6RzTx0t3C+k1U1UWAoJLVzuICc/nB2WwCaE6UKDERPziNW
AHRUBQnKZQwBXIFBajF8FGNrItWuWmWfrCqEwpWda4L4XKbKrbOceq+4EX7FOg8/q9qTL4sDTqU2
d7S49rob5kHl7tcrxrt8rOJI+rIGwjG8yNswWGSRdDxdexdNtAuix20WzBO3SkxYCnYKyR6CtNZ7
NuLNUOUR0tPoXMJuFAu7L5ELfXYWItgrnu3kZ9BgWjQlIncEjEOjSAWUIOi4A+hb0L7UyC0XuE0r
BKBiRNAYgEoB68FBcTPCj9OMnsLHxpGteSNzo3JEJdn4YRa/gODL0I7wLariNB8UaO/C7lNY4sOj
g4uyqa+4fRWAPsiiz14R56Fm4WURqNcYXj6YkrdtpgmNkwALV+yqaKxVXP6xVREV21p5cd52NBTq
gfdEDTcKy6X86y4txKBu/YQZIqwGiPLa8s6Kh4z5V7C4z+84mftpTtQQf3dt2NwC1ulwXSXUAVC/
R+h9YQ6dOSsZe6NjeYdlTdWVYRwmm+Ypx/Mik0bqyBHSy4/dS/pg9aQGRAWmlZq37VqlczyIj0og
T9F8vmAl1bQey6eMJlK1xtmw4CJyFY625sqe1p4KPTFIvoDJgNdqDN/VQ8B3JBTg0MiZiSnqz8rW
fBcc8Vh+WbWWe/sKqvCI9puxGNwTViN8iEsEM29likRK0lDwHCRG6X5t4bjOvYY3Ky4Eff3XRcZv
SmDcz6fGVhqS+xqov0oI0okA0HcdPTYjL8KfnCz1GOravocnit1530B12fGfQvCMA8TenBrdXls1
PkATGJ/Vu1ZJFyf6pyBy+KhqbwNQ5zH+tFBQSaoKIwRb138gQiYG7Lq3jrnwgm0X769qVAD7Zp6X
n+7rWDJrZ1h4i2sV3UBKQBEEhqVaIlAuCXZ223GzZmT89e/srV+FsPDnw5WA9SaczP+FXBxubeQl
Cm7RQ/4YnuYx0DbOe30Bh/aGWkZQa+UWf4RxVeplI5NNfN4+EQdSrzi1qQjlPV/JnmmH8wRZhCcS
IZ7SsxhU10QQa7JL1ob1SriyMgxWQfaKrObLjhhfRomLCUvPRIOdDeP4ZxZwF2p9+MDn8KVKSdN9
1ewPYdytR3sJf9JeZgH45Bk/TLYqHVveBSAJ54urYhFhyv/+ARWmRp6MzkXCedFuCogxZRVaPIVa
xmZ6NXq40VD0Q7hi77pP+CjajZ3dalutLBTRxTDTFSv2hSed3BAFiiVqwNCEsf8A3LV2RVxZtdv/
7CZrNskARx0PccAvi2Ld1dlCiDsk/mhNnvTsrlov2R7qkraF1a6MYvafmhwQKfahAWKGUJcC2Yo0
xUugUna8cVdUwaun6075hXP8nqv4+hv575siDTUuP6J11lZe/CT18WFj3PrkL/PRSyL5NAxT7KyN
APIiku0eKkENfhhqIEDMGTVSjaMDY0pY+9ubmhrEj2rWhodr26RKpFB9Jm1YE0pDwT8K5HirrYX1
oiRRr/yoOSsYX1Djpv8ucGpGuKujedUFEE82Vgw5FkcYx1SkUaCYJ4JiHMPUI6p2qr4ozh91We9o
zNNhn9jMeOUO2bPg1Pq1NMD5D5Qmn4RUT/eEf4fWaGOkchG8Hl4hpp6r4sWviyirHLWnMFQlzTEH
Z0E31VRpwy8fUzYFVz+p1UPzN8wA4oGieBmbJdKw4G96zOytsexys/Ip8iQDLQZrs5Q3+YZQPPGU
uc3MAV03j9IYm+2exkYJLzCR7cpWfU7IcsUI3R42zRiW70WsILwZMLB2qGQ+dso1NjWLlv0hp+gJ
fQC6BRu/jdzGCL853f1HuzmzG+Og42SIp5nVGk2B6ASm4zl57VQ1KAaQvnZEH5Ngx836BQmkk3tP
U09D6yaSLDCiQMig8SUaPinaHu4eUYwofF1vFxzZIFaLAXjPK5Mnno3Jpc+7lzgb+tsVdb1HCteS
ebWoDuW/MVtKjnyyM/l9bdP9mJmYwUHWBJ+wJbByiT25TFehXgkakPrGnPvO+Ldetd1+TKQF3tfx
2H8kDK6daQ7SszidN2rnptNxk7g0cNjbNC9TeCvCj57JZGiKFTY3U1dB7jzIpR/rSKvSZ2jCRRiZ
Wu4tnbr8IG6u+Tww5iomAHtwAI0o6ziFXHFxTk+/gQziJTgU+sSeGxMFB9IdOQbXZCaND7RPMpHa
n4TLFiK2pSzNzmFvqk8XeNEtSWz9Oi3KVGTsHNaSJgcfjl7tlif0XrPMKp5nHVinBe9kunelY+X5
KbhYwaRUzWrbAO2Qebi/bh/vwPlSoYf20hwaF+np/MsVpax97Mm2nenxWIpJUViVkNJKD4qd0eYO
mKA68FYzM8RjLeZL7Qh048mqufQGpT8DnVEZsk7d2T3KhmbMM0h78JB6psIoNMp7/LJMpnuOXfC2
UfPOR/B03++dGTW4JTQL5jppjG0BIJmh3ofWWI0SkrTpeGIhnjshMU97fkBX1pB2HN6/AcnWC42e
6dun/vRiTp3MBUpsFb1wQ0XrR8czp8UShcGncpKjjt0B48MNsAp3BXylp3iEu5z0hWAhqLoQwHDx
JJ6D9HTRIABs21DDWN72GCG+sRpkBPlJed31NAHJiZbGGH7vEx952tamFEjVMMS4evXNyzzIp2r2
XYvaXAetdtKFM3jOg8rQyh1n2zdKNZCBVbpUiN0KaIvKxWjp/OWnbrCsq6Wl7AAHnZ9q6X2I4BHN
8boZ6UNDoi8ybkvzMOG1VLCJx5hui/nOR1+/ayPoL4u0tmAroLTLWROpFDFp6+e6otbTcmgOVBAn
DKLuVUqvwmn4lpNKy2siHlv6RIzJuqtYSlHsfOR8V6MO1bF/XtYlHNr3sJY7ymAJP/bPqnRjgpFO
0zc6pMiiKjgNPEbUA55vrhXt1lQq4CBcJS37sbsF/HplwZWKcMff6XRJ2EZsyBcMZzVwkm3T4F3r
laEvO2wV4eWJDy5d4GVJf99CGqzlt+r0PwJDleP3LsL8XS7TsU8+D1y+K828Gj6t9Q2uWGDI7BFq
tQZ1/rIiLg99qryEj5+sQH8jMGhPhCjpM2zWQshcii7Nv8IWD0jfdJZQJGLe8fVJcw7ll2GMmNOa
vNPbydcyQtpg01wO+0A/JN8JRjmBDZwL0+dhxDrY1m32szteBUqhyH/eygknxp+oLEjxyP53gGzf
8BJGs0m5A2J3/b/od8erb8oVzq+AOd0MENIaAwGhffABjrpw/aZ8U/eFy3DodIF1feIBxh3K/Ej8
AjErcEeVd6kbs3evQ68zPBkYd+iwlBgW53S00Vde1V7G+ApcxkZO6ZIY/GZ4dY4w2nfKgWqcK3uH
6EHgqv1tYlcYgl3+T3GEkwTscWIK3XrLLgykW9oSLJgwsebs/qd/R5emXmxkUORmL3t8pJnI7qwT
aYa/UoaFbmyAZMo1S4PDaV97zKdr0RIG0+qFqdhEIt8lcWdEPxGMChG9R3639tPGqzXyegG7VHb8
bz9bZYIy/XEbjsMaXSjXs4DnobfsOkx2vVfbMZZ3KvFd/tgSAI0mkxoITqAzx64l1oSXwNe+BqTw
7L6LZJ0XDWlO8yjcQqArszpExcfhGheJik8U5lAzS4go1gcDXh7MR319i3EjgXs74uijEss+OboU
hLmAnNmMkz6M/REOpIvbWye44LzXjnsyl2nDFfhJIgYh65y4EWPGgE2FnIGgemk3mp0fZ+/oVWRV
+rUN+eTqyOVEQJ9DySSilyToB8Tn0shzPf37jV6Vj305aNNp+CCZssuBzytY7WaN2jZcOjAJ+y0N
GLQC0hDcPU2RK132f5F90N61gHx8ETC86KTdn1ZNVmkDoa4cRWHB5zlLyMZXAMlYhJMnn41k1+Uv
LzuLZ/YykKV/Od8XmpQktEIjopSii6LujHscsKDvOcu8qK+MQzkXabvby3KCOaX57YUhHayHMYp3
NNc6YSlYpzBgacdijXF3ruJrrZgCfoNyXonlnUPZKWLxoydV98NLd6/rC29UX4MzCY1UOTotd1p/
bVyA7BTHGWFN6blC7cfN/r4zrDdfkcvIiFSU0mo5XW3s1zKTRCpebwafITbSIhKC4rMHbuBnlepq
OUK8/iy1u8AiL4D0Y0JhOTgywYFu4Ur+SpglAk33QOk2Pythy/QgEdG+pa2jH7RUNt+tO60qnub+
IG20k0fSEIeOnM9kL1krHWOCfOTvucERU3XBq25bSYK4jX8TM+OWpK4TZxjE6Q7FfTMYSzZs8P/3
xpwfmktMsG6UQKg5mrbAWcPO4N33zcUvy1wQjpyjK24kiYVxKzkrUe2nNdj/YnKw9e4wlkVf/R91
+iLmTLboW7T2r0OrCBbP/LkLSxwMxELnOMfY9CKEYgFJLaqhsLFklaQDE2XdbJsh+47LCggsNMox
rNu3M7Xcn1/SJ0aWSmOrxF1a/bPU8I8y7SnOmpzKrbEL01ZsMVJn9xY+eaJBc8gvIPu0WdPDyX5o
B3cndJ7NyqnIQgYJbsksDEIyjHbCe2vcwzS0NrruI4JUe8KRnESxXULPbxu7g0qBTlfzxCn8mrav
DAUWWO4hhsshyny2GfpAj74mivpQ7kRHNUvds/nruU4eudY9/qSu2FMJ4fHESMPSVleiIYVohAGj
3bd+oOQIEhZEDLRtniDLcRs+fcfbzmGZDi5u55FfTIv3JgXqKNiSngLbGUnhTbkZAGwfRxPn7mkH
lof2qyf7gIris3T41epn29fFJ/xnMiWZZCz0k9hL7AFP6oGDDeiaG84Cm8chrCuOxICjqkCyfqwn
qQyufPfSIIeFKDDprkZZytX1ryMr3DA4KmCWGA7d/QWzMkEEBTNJ5Y9TspbxUMjUO+WZe4mLWpnN
EjNvmVkBQLDGzzMyNBzNuPRHH6qJMhqI0NqJuWjGjBywgrpAS4P5gKzuKbAwL7deobdT0jyKyxMU
lf+lUTKEqOSfbBIvcu0vUIVuPN63ReRblT3gTs+M+9gij97C/1q++7jeETu4kzwKx+Qrr+HNtHM2
1DdeVxfAaohnHQ3Vv9UkHt5NiBQO+Jj/j4kAM8g3YX4Z/LNvyBJxfeh9z054r/Y0mV/u7VO4Y6Y/
WwNKx9PQw7VQ19K00D9ytAVl5iCLx5wBrSrd0YUulxa6hG1GpWA4FklPcOkVaR5oe2m5uUMFMked
8kwRA7Wxti7Z9r6TmBoE0FfLk9DtjXjlB0L+j8EJWKXHasNBYmwi39hXNClAX0GRj8OIYsm7OmZS
IgcgTxsMj9rRRzrxu+S72IN6+v1PiXixhtDsx0rN3J2Bz0GuEPWFwSaCTGd+htHWGhjZxWVmTCNY
gtv9ZDnN85OLNSNGC+XkSqbAPph/5qvw5SBKljIxfuvtKgM1mxvLqyrs316ss45MyVqObfx0mFYI
9kOneRI0gUFDYrUWUucnalxbfcrXwtV6lGLJdR25hPOHgLLJlnyejiJAkJDvpU5yEr5TdNsL+roY
xKBw8HueC9vSzbqL8tXsFOMXFzK6IrfSLTVHrKdt3jm+frEA0xM9ShtL2A98U7mkT7Rw+i0hbd1L
aMuayW/jg9u//8XWareANKo8Vuldi/7qnlBPOvJdYOCItUecYfAHbwQj4uYx+uNW2rExEuVVUukP
TRWI7+dyAF51Oyy6S7FhTnncBybl/uWwi1LekEcBDtXn1vLduL0UOQQvb91NmXcK6mAoXj+ltwQ6
74C5ykdh/brUI+CPgClEzHpFGew5xzFcGmrdX25U11yDyI7PTpcFahvhM9ErzwuvzxLsVHXC/QIZ
DhXXYhKYwhZiTrK29K/MEcwQk3L5u4q4lRvZYsCD6+2VkaNT3ljNJaRbK8rqrDFlGHTxEjNg6LZ3
e7zWNltammdwTHuJDMvknt/WWVA9UFxOSrLfWxtzqTfc1woQlZq/we7SlGntyvkkY3aP7kwzrfX6
m3f90UkNVyQ4kNJAqEW6CqFuriniVf3NJa25RMgnRdxCEIELQ/AStei1/w1rJR+I4lhp8/DsZZpx
kH7HqZdKELnTS9wNUS1WKHcIDcsOEn1l63Gpe2/zT2zfHbbgGh9Lf7kDGld+tsUREIZX9NrEaFqQ
cFd3k2L5jyb+upDsi7xM/uw/mzT9TpIpBHEtf/U7R7rnxb1xZu5XX/Nq1iADy2LsMVO2nyGs126B
qzxPzlFb3lZ2QZ8NdR8Nhrv28/Pv1/vyQmr6ulwIvhJWADJ1XUxAfVZJnf7iGQq8gfz6M06qbk7r
GNaJ9b/0IgYs9Ds+KXRRdtTzfbgRr3WrHvJOb9vULAmmUw6d1aryQegzXxMp28OJUCN/z0NrpPnm
irhNIkaDWH0TcUBoyCc4Bi6FgfrmhL8rF2rGZWmK1QEWNZqx2NRv6D6RdlqSMKoWCbC1/loxnaZk
vAz6oxNmjS8j83XxqconfWOdlJpp+GzAJ1ah4GPi0p+nP790IDddCNPv3UrkYD9fO5+2kBOS5t4M
aKDn9hkNi/VSnmod7aOi0hOrYjaHj6n5OpXyx5LD15WzvR+A6mP1yR3VrCo0CY3vhiQRCf78MEtx
dJmIiz4QNY+HKkIp0s37PudOrgkBOcdk+nEtsMmA4/kMF5ClZn22XTYz+5c1owIu0PmK+Vh9BzgT
AyTlEWmPliEQQ7S73sdbcTo1CyD6PdJuJ5u/61nqkHz3YMXXhYlE6dqTSKw7y56QsLQTiw8OB2+N
T/UGJngO59HNBrc6Gd0ZstJ4ltFd4bwILbDeGFpRpXAzbWzFlcfMFF2fjNy30DQvxTGKywOnYw4Z
P/j8uUp91TCHKbPi8YpaJZA4L1gkI0081fmvyhH3Klv0J5K7l6Py+KP4XtEnSIj3FcPqxTRLY1V8
2QNbViLk+j0k+6Or61MWAEnkUVXq7N4Le/oMtCrQtiIdp9xXLVcCQahvS0T9CD7VmYu27C+oAUKZ
YY19cozHPjz3yHtIskPkJRplmt6iNpdNE0ORjR4lxXgJxDHyF4RtvK4iGvom+vR1wU60883mqWo3
6ENcsZMjO/GyrpmRVpY6R53Yz5J8d9CX6o3RyA5b0fLeWdQFf+6LBte0pRtPbVxQUUfMdyRTMc4n
7eKPxNrFOsPYMfj5PsfMdGpyexktEyqYpeJub3h/h6V58+7kdpANOwO6YX8ljnbwfXzuBpb2y5cr
VHtfQB/YWD9wYE/ar2qLC4rkp9EZ/F9+mQ4P7BlqN3YgmzCBr3OSVpTT9AZmnbWfFEbUhJ51ts6N
BNcpmoxB1Vywcb/nxKxtGJOT7ZMb4+jBaQH2yZqAYVVwT1gVAVz0VLLhGudZNnZUivSaH+7ioqYG
bByXwRkxZYR2ziRpcWeLjcNp+JAHEehibng+jM2D2qA/iAgoElnu5ZVPtw1E19133+hhxJh6SR9f
jaO1s5GvPFcsWOjpBHxDo67a5SEz6Qs+VVpsEzFohQqnH7koEMUesq1ajQF+VIUWec8Wk0pRMCoV
uxM7D342rB28EMfmQE8d4Ga06WGN80wSpVa6lf7HliSJlkA8G9J1vib6TetY6aC8k84n2MyVHjGc
WlSTG4I8XcAFQnsYZat5pCp893xKt8VzT20IgSOG5VY3O0meRrhoLYfU22Hi9B9wjt7mWAQMBZ1y
gKFfXnJeP7/GZO/QEb5yKUvv/d4Enw96ugJ+H+hUJAjQGbtAbYwx3/w+IHjnU0v1J9qRimvA5lsw
H2vf5vTiPuErkkP7kwhd001FLbbd8LXPHBHlE4Ap0KUSu5p5rsCU+xIQfSuycl397eClSHO99VpV
DpBbxcNdBWXKr9r5eEr+/gletatD01oQ+wRkVU/9wCQ3pfKcH2rflZMOBxUh98i1eiqspBE5Yapm
cMNzg+OhmGcsWDc205Kce7pfgfWUun6ECYRjgzLaXb81FP0ecKeYmQ58+fehLDEw6HOSwvAKBz9d
J71tEgDjE6bFglnYUmbnqCkBjakFcXYt1r3CtKPGLrynQSn3KaTnSpqeNGWpEfs=
`protect end_protected
