-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zpkPwzO3vrNN21IazqgeZQ/6mZdDBdKiS0yRbQf7ULXvuLskK9pSnLuVAejrk64rj5o+3cYTfhxV
EUD46xkSYE8IWKGemEUhjjMGw1ekiqSoTMWH+V16xYVp1Dia9leiUJaO5tL1U1AYuGGPKGzGX6j2
D843PwGc7oL2WOj+nA1WSBOpcsTkrCqzpp/j+yewfaTYmSBvKRCtOwFPCzEoIj4s4tM5KSfaMF+T
P9+6GTE4Cr9rUM8XCHThoA0L1DOwbJACoRVWY4U9GH2zqhxPXmVh7Yp7xit7hokJ2D+XoXkmeAZB
sXbMeTfnmcFNhk49qXZtYB1F68DrC/X5NVsiQw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114400)
`protect data_block
2C2w594QTslo7FQUNVtDA2hXj5OXq5YrEUa6bFeeBiyl6TV/JM3RKI2FhtucYjVqJDY/2z5iXKDf
MKuUBwlpy1yocuHFYNkkkfmrv1z+85XFTJWKkVcAycLo/qs/htV/Zgqlag/jMlN6NJcdPqCdyp2v
chc8k7OjfHjsuYFuaRhjv4pCV0f+0bbw08NGhlNH6RLy/2bnJS9ysCzu6ottdVhLUTd+BfgTAZwJ
FbddbTVNlAgqV9GajhQKMT0bqbgzD3TNnqjCwobyxgh+CrIB7DTDjR3f91/Filhi255QET+d4q5J
bKYyWF8sPjzMsN5FeeJTSEkk2msWE+WE0ON8yxd4ZtRi7u1npBoYM2j32NrSxyMW+klPE9B3zWzP
ycNTJfYuBlj5tX48vq5wUdX5zzvN92+iCOF4jLyVCS8GqjbKYKn9XbMLxk3H16VNNJE9B5PMIeJN
5rCM8mF6anS9vVeEDwbr5FT3fZgRNvDl3zuj6BqcbdEXtdG+H8PAStnGe2mFpRdFWw85JCIOSIoS
xbAlUc8apgm1830xTvLALtCIRmVSa09i8n7sbpYSjDU3NoQHG9FryG0iWP+yL+dX7HDVMJ+cnK4f
nznY0ML+f0OhmkOBDSsz1o1A8FamolHVjLM+cQKp7a+r6XMGl26pzDkkGKMXuMZeJgF7gU0GOmMJ
iljAX/rAv7A8mJ2/T59BeoWja/yu7z5ZusCISKg0pOtJ1qjnyuYGyzVdjAxdnH7DDU6hguzDlv74
M51ISQQT0A2psO0spnDgU/u9qtGpGbUVNtFJA0unnItbUmmuvWiF+shasN6nwud0v21Y3QehFcEi
SV3TQXnWzsEh1uC33IH0xK9+AknpLsCOaZZxGKUnYnAGonYlw9vngpBKxXYeOdts3+7ycut0l4TZ
faaUAMlrM12gJ8qpPoFcciO6FEHyMIw0BMr6PAW8PKNRfKP845cEYzogd+GQCwsTF7A1azCOkmJj
BiAtnY2HZO2UQEL7IjcL0EKKC2DrKUP8H3h4I+Po/iTbXprLicPzrBP4bUmAo8xkCgYB9JbdmLld
8CPnLdTQDBTqNMhFHXrCCmEoHgzxl2HRPsRoMyGpoxXS2j7MfSiyFqlsmD91uHYmUutzVFnx0PbL
wcl7xsfeyXi+samFIw4eAlLMYVVlU4UtQi5vlby8bbAfHPeh1pU2P9B1RODrVwT+TFLMDUPmSe4Y
IWZdXu6V78Zkg1OGPIx2cw3fpfOZ9TTn663xmswezhlDmtX8Eji2Px0TKuvkigjd6TSy/+ZACokK
3xProNrSuLOs8hhjxMDtGLr+Xin7dluJURYuut7zz1alY0gWXmaAQjqJ9H1lDIE4k7tcDAi+GWhp
NXCcdr8SzMmIubdBPEer6tfG++uGGSsdk/1vQE0ecsXxivsJYNiBRwjptaOjmuK+uivf/TgRvL6A
YM3AO6IdIFIRBf5ZjfWogJYRchK9dhhbKzbGRZOIdOKY0ndKjqf6boRYvNK7ueAK2JfEK2SOoUjj
U40zZ5HXRcCrIdmE7AnN+p2iim+sekUQrt1sfzTg0GyDGB2ISmYBLSAxCEOxVzWdak1/evdHCKap
AOoWrJBMrKU1wTd2sBa3D5dmbLYCPemrrRrnILK1SWjKXsTnEKBJ14nhUmeIDxnFuhELp7aC1EYI
Jc1mmmAgoNSRUjMdR9NaXntRJ4nwlujCwEissNWGZ0JvyKha6To50DbmujWbfZs520k3I8Wj+o77
RpPNhbVDitIfvIPdIVGCNYP+dSVdo1/QzcD8G09YFJOAEkRKHejknoPmtFt1qgjzcsErqKp949CG
MA+oJTnRq6/hOd4jhgP9jOiblk5xa4hoc0h5r3ZLzEXq3DR2tg7nMSi1WxiATfh/bvTs5PHzelfT
ZtnjEGUYNwCfjRkxjWW4tFNYq7/E3CNQmQkhKXSXMAhAmnQFjtKTx4Abt7dzdZTq1pwIFWREiKnC
fjb4BX+WHOtuVXEl7T+weuUtVLZmV2EXmblbGc1wTlkbRsMpdzx9fq2ImyGyy8Iw3/wMH8bx4YAX
KF7s0H70njUAkedw7MEjaMwX4y5ygWYMiHZEeDC5QJ9zuoHjZ9iYPAs7F4EhF0x50EohYdYPMMf4
elNCfA5iZZSeD1ZBQKy02dud1rqq9+//8AUbEifKBaoB4kYMjvNik3Kjtw4LkDeTP1ArMCJ62yQf
eFkm/u0IH4IyZlfgRHyErFBlXAvphwO5ul3+XF7KLxFwnICYreFX3sRfd9w0MXPg52ReuiXUSNx1
lREkA53SCcBXaba0rSwewW3SoO6Njmuzh9IFvgcISqCndUp9rvKMnsKR/9RGBl7SAErgFiWtF2ea
qTaI8gxYCIuDXGSBbewWBS+AqKLW0FGDVTBWmiqmroS0MqkhbXIOw7HJpn1mQjTOuh4TKt7pLdur
J/2Qj624bYUCos/ffrJkp5ELTX0K9XbAEZ2ppCPvwdD1lm3qlBKF4C8eOem1fg7G/xwd6/WZaUTn
bXfqkH3/sltOu2BQbUaIke8UjVvdB3EoffXu23juUOwmSQUFcLI3klS2DmyOyK8od2l7uOU1tyaK
YoMJyXEVs/Az+zRG3CxFj/8hHDQ+93wwmnZmYiBDu+ViwPMquKMxHBBk2cE6HosfwlQBLrYFWBlr
/PtM9AcPZcFpYLD/Fl8enE0uBULwtN0agwIcGkiNWXuWY3MZNcc7JgmAXo2IsE2Cl3fVA2k+1H2p
ff9d3ByE/HGWzH03UI0uNI5k39jrWSije3SdNjDkME2vhb5f17/+aZtEwfQ1MSbLW03hRjK2xpFZ
r+a3tjfmbC5xC+YMHcJ5nLoMYShUemrsqUUnMB+fLmIstlR1g+HgZeNJE6x4w3ELNudTM/DA4/pM
ri710PZYQlOdM38pJEhbwoFjjlZp+TlIytt9C8Z85wPGU7eI+ThTEDze5atPAKrSAB0+L2qQk6A/
Mlk+LgbL/bYUMA2gewy278zfdpVCSg3SFfH/DdtOiCjAML28zo7TkUgf/XhCZFTRP/5EZfLSvkRw
O/vVjdxU/JfbK4wkg0RsXPW8Mn/voaVyFZnGxEp5Jo89pKcIDtBr5EOe1NawRvc1x0crZhPG5DZc
//1YHjy9rOVCUUmLlad5Xp7+y/t66sSMy1Ea4yE2L+cXYZU/Q2iZepHmgvkUraz9g1e1jJ0d04EN
d4ikSjScFE5V/pYIkgRmzMdKpLCG3qKRoHGyfuEjf0B5PTfPxMRoj8b7Nblt6ZDpYvYjujGN+Ytt
I2cRRtHplufplpnlxWFSyDKeA4H+4RcO2gvNw/HoyZQI6RSCw2okN33PzNrwV6BUZuK7RsQLAm9U
L5TR6FI/kKMo0m9KPPOhGOQWD3jP0Toh2RRUFygpuYQdEZCEFNbQkq7DL14uR7XTEwn+k3zVUuB0
AAWCtXkxIlnPbEdXOcr0v5fMcLr7aVqZAywEQIv/ozygH24rMNoduNgqwIF4vpSuaL/RJ2rXL6YF
w2G6WHZBa8DorLg6qEnaMGT6QPn/KldUgQMPq3Ke8yk6ytwiZEBJkgq9gGavqcYwPIihE+uqzm7f
iQO2c7YRzByzcgTYcUj6tz5YshDiMl0RVbgb09UnHeOb0UcqiqRCOclIWLYtFgCG28I59IvJRons
Hirirhe1p7W9wVurb3n6gfzmjR82V05Zo3bGI4y8kg+1vlC6ADq6ltumG+e91SnrmonZP7ZtbDrF
ZYMpWkLLeVeza/tozXo5rtbcGzcZcfzbbP4PtCmWHgsJ4QRgY4oZRidrHx0U0Dcvp8D8lnJU61JE
bKvRoL55gftRPs7bG1JZ0jfmesbfsc3VXFaER5He+Nsv32eW7rFofH9SsIJPOTv79rKkt7jkVWjV
RlAmGyb7hVY6rPd9zAL+vGNZpy4zQsbWs6I6gRad0AUWoN2wIOGdB390XMxMyCACb5tyjsWNjxbF
inoG/7nLRyZRGqgPQOS6C+8k1tChXBjwwznmaoYCjfhZHD/H30ibvHuuY1smRDeUDwkd3GeU2unI
+FNpal59ZP8NebCZ/yDjX3FxI4xsGl4rxeGI0Q9BFg6ddK96RLm3/1A6JUz5ZaqTl2XHwtdfqhKf
cYDWQhrYc/yaYELodNHhBX+FVYQLNByCeUNihKyzRz87R4xPJYUaT44Q8BcdL4lJOYiUbxHmLAh7
k09/hu02T3FzWGw/hSCp4mwCmFTuUeMmJtKvSbENebGu4GMAN1szdlO0I09b7oUmadGr6gauRWAc
k4JCk1PZvgyq3NoCraimMYCsTsrDD+KicaFDsBbW786eylVHGuoqDJcwGuO8jemLVN0kSSPRbkxn
rAN6lh5zE+ipCxSNx5mNBTwiyTjcU6f9LtJ6bj8ClfSR2PNuTmiskATYG0ej7to3mkAckwodSGwQ
oNTLXuzKErG4upmPe70H4K0TT0eCmQF16v8noq1sHW6mY3g8AkH6HvjN1N0lrHJbeCM7YVJVvdm+
JHSQZdbpPB8bYwfsC5DxkWwawXywDsgOOV47RI9DTqn4OfT4sXG1+yjz1R34gnOzFxVlac9EJFXe
tLls4+akRmn8qbmCTVkww1FNSFKslpO8UGQ0z3x32xWpUFnj1KM4000ouSOMTc9CrXINhB3lLC0I
dScYq9ZoJMdrEE2U+/+y0wh8PLCtEpTUJusU33Kl+BBUh2F0FAUqKLi2kfVfMjR8al0yqaZwNvMe
8efPTRQTRodMppPKB7TaV6tyagjIA/+ppTQZObpi2G5PSty8/2txPd29QB54x2whg2b8ImcjVmS9
V0VbWQcD5YhSHa2FX8/ZB3LiXV/c592q/NF+2MWTO8HBPLM1eqHar0BTg0aCCSQU8bDN9D6tnYH5
F4XYnEt9rcDUFTQTfxch9CvN3m9EJSCij0ZFZIf2QqEU7KrNqEaVbuKXuH+WEJTF60AT3QFk+rfO
Oin7rP5u7H02rVIkIt3m8x9pkrphBeZIn63pAxUsojlucJ+ppn68zKahbesKuHFOaDe89gn+E/PX
OutW/rKC6Kk4THSe+/DkqIQX9vT+ApiLIw+SLP30Wx29dRU3DvxzH/mMmo/NCGSKeLpjG82Zk2/a
U9gioUk/Fkkes3AQoGEJhyhgD4hOLGfwyrMj6fYj6/WQkpP0drVCKjvJdhh9RHWszhCUGqdD3ztM
zXIY/fiM9iWUIDxkmFCU8+5A6o9LhmFmhMVssELp7f+yX0KWOy9vXov0RfTgKSrjxwyIgrBG+EtU
koLu7zdRqb4E0fd+oVlq6nnx7PMV/821yeFsMKz7V5dhLtTcOEQd4o9VvqC5+CxTJ+whjcnUxRXm
RnLimvBn3HreFPnF1V/aJ5+jbtV89udhq5lnrMxlUYlTkHSeCwbC9jyiYV4rOjpXqCjotZYqwwip
I/ujMc1qnZI7hEFQxKR3lVMK6EGLLJPwEitNZ8CtFsbrrURDDPWeuUReS2z0qMsHRcnBZkFurcgj
88bamIM/s8IBj24rqLGFXi8+TRV1XhHSF67orK/iOq3q95ZEqiXHwu0r4Nmwl51/y0fNRWXLpt/A
C/BMtiOYOz1YoG3dCD9XG347jkXKWw3VUcpibD++4yQvsvapGkTrdo6DSfaTe6R22cswhhZ2VYpk
BCfwVRAcwJfA2pXIj29IINO6wyUul9b3CmXBsEmBfuP6T7eCv2eRzf9IIYuBhW4LnPoHun1hvyP4
2Yn3AC4JHHxZR6G2LSjado3TWXdjA4+ly+xIh9eXs2Pxeq9iN5fa5cOsIjP2Ko4fXx8an6/OxNdW
jks+V8t1J5lZvvDDw7h3wAABte7hz+f6y66QR63eYXP6rH43dLOfITIvur2lY8ydXTMTcq7VuVpU
pTueJHwwIunDvzz1T5wQ1/fTFjXIRhtvhgJ/LbRsSJ56AjXqzgwbXVswip6N0Qn2lUUsIaeuYxPV
KdDG5QMRFS/xwWza7Z+I4qZV4g16IQvDrA61cwS0bifvetYCLu9oG6fAYfuI4+AOoYHgayfFdFpV
41u3ZJvsOVrOQGhU+99fBDBVF9KJsUB2aaEbmIJLNWB3Vs8wSGAgveC4MTnYCgZ/dze51JpZSXCQ
3sm1iNytGL6H94ttKZ1LAWCVe4DMcjw7hmg3UIIJc/sW15qNozIDLqkyNKEnYMi7qP9RU/wXS38y
q++dd+dxX3EEP456ki5npGEQ4I6V9dt5Lrq21WqW0YaLCIblePQzD3n+U2DSQsi1Ow7AK26NX6gw
zvUFUAurYpz9Y4PbN+i6zpkPxczhqNSOQvwHbs/UdSpJMqIpLR2SWtZK4YgFAk2wrLO/++jkIGYy
Nh2ZpZa1BzZYwczfiHUCJJW5K87W5amkGVpydvV34XDsyPhnyptUJOFtEW6MxVBXc4bGtNEPf4qM
1+Ha+qSoFf2pLV4TVvE/z/pxZo6Ao+c6B2mZDanyuR2qVwTyFpu71MYGLAGU2hjKUxYL12yWLQ+D
dtnhrnKFmFsO1fLfZnFyq3Vm3hUwCV207vQCntikxv2CXtRTFuGIIuij8PG4cZ9Pndjo+8bjL5E9
YWXC7ZB1oMqJiCQvh6k1YjMuMRAU7FSDd6YV8V8ij3cHCke5CkS99PpbHN5hDPEdqvsvC/RwrikF
L0oEWSx7qoEghUp5QglM0QCzG5cm0Smb89kyYs+rgPUvoejLdPU+NzjzKYXD8jnwp+nsPcHd1VrB
4JGH9hWCAtq62sE2en8iYU1AudnBemNchX8tAKelyd6pM2LZvFIP6qTxx9Muknb4grJglBtr3P4N
7UTKzzLaq8C/B3HE4l3e2inhcfk2zsB5tzxtkdLXEcmiVkBz0Gb0FdLPOD701LfOEnVd0GdMpqS3
ZKIMLfEHUgX/tc6YbfP/HTotPlC6yiFLlPyj4IK0w/f7Btn8F+sHdeIFVm4RurLk2BqOLWM9NRxg
1BjL4EuRlECYLyJe0P2oumuP1zXDFLhEU2IoK5MMqYWpi+SyVRkR2ZEfjBuA3gpanvhxl+e14g2t
onZW0K1xTHjVG+Mzt+32no2JQS0s7/h9LrO6ZrdCZogjI2Wy6gwIZuO1BsliRBa3Tpy3TYGHDPNP
RwBUWsUpyVJo8ECOqRueBKvJqK5Pj/lIWXsoLGGmgKZrpRhlplVIMmy8snnIjVRXLGvWhVBcl73v
6FZ5RftdGUFbtjncPCmDAFLogX0Ut1u/xdkEgBLu+thmdWwrH9eTWgcKxk6GADdEEGuQQ5vy4vq+
MQNG0yqdCjUwEU9jE5m8gUofoqJyWtOM40PaFtk41ymZZTrwaJ2nxmG/v19NgfdW6qLUAMvHEglE
F7jyExPzGgBAKGWIXjSpRPo4m2CN56yqopupPJN/wTrvCJp8Aw+pYAB6wF83z2R3RDVNee1i8DOd
d2EFKy4jQ9uqRIEy06q6MyE4N6aMZtvqfc6DSUj0qV4n/s1LHWEF+ZjjCzK/39UNnGjH3sIPNYrT
N3T0eWDXLUDJl98cGS/Hwr1wbBFRiv3tIDQmbwirmIuDANzJlU3RtQaGPy6HQvKXn/kkbkiikffy
6AaL67n3j7uwt5tPWAIz6z1v6nsxX1sJGLFjHyq9jVyhmx5z+RUa6kBPRfpMfbFR3srjoAwe3sbO
JxTh8j7R01H20TEr1OqLlfpiTJ4V/+VdKtgVutB5zVt1zJRwgHUirx8Uiv3p72G/P+rW6mgi2x2N
cLfaVkmJYDqqhQe9+IUuGIqctSqqaKciRWdv73ddTroBc7QrwCK0bo3fs66CVGxwTR1pcQOj6o/o
JnBBCIlWTzB4j6in+lV1LZxB/u7YbjUWERYPE8D+NRNch9SGsGVmV4AD+J/JKzXNCQVVwuGUlSlr
uTDGHvQLhfUr6haoSgW1nIJgVe9LAEGlB5NHT3RMKJ5INcgBe2QqZfkHlm/r3kNUcfJt5F1fZnnP
ht9CdkNlWhAG8XV3lB1CuRMry6QFFhZ332UYpN9URQISXgw51tl4XU5v4FrUxs8K0yoH50jBuVLB
iILiy2zqabZ8gWjArJPYrw+lc0AQSHXJ9u5tcxT2MQXBO14AOxyy4XV+/f5zZGAMJMZNSoHQt3Hh
ti/GQe1FXL1D/eWsqWINdpNS/nCdA0wxDyWhu2kMRtpV/mNN/7Do6dXCtQuxpedK85OsLoTWwBcM
aTkU+sjAO/XASZzU8/c5tOEjc6rCT+DNAoyf+28w65H0S91udig4P7mI+mYLogmnb0z/Q67/2m38
dPqNMwrUS2PUfdy/JK642n48W9PPDi6G2XHY7TEOa7FfV1h9xSIzgENPtYMzCymb6Jr9txXsJxHE
Xpwe+4hZncH+JnWk3KW4GhgvOBqOZ/TZ84VWEQ+kRNxfFFk4U62yh+/vAkAqpPJy8lER0KzoUF9+
0fftds7kkJVJCbpatPNOuuHyBmVispjcTl1GRcLTc/6Ga/w0zPmYXcm2mBT6gIRu2OerqT21QAeI
axY1iTB/DZ2PHcykyVKHoxjwbkAJ2CGbvdeD132VHuK4uTyEOQ/hcSD4ppiy/hsIba4lPRcx5QrE
33hk/HjAHcuu1sMEUGJqdNQZ5D1yIAXecBVV5OdLNmT1l0Vg58tF4Sw21gazwUU9Jk1cM+du6W4R
tzkS4Buz/eKHgLsgXMVYujXKgI7u+eB/OPSXP8j75tyedn4DvLP4Uqv2yNTKcEC6acU1abfrebry
Ov+HCCLGR533s4NzGeG5Dlv8s+nDqYu2loOTpyuH9d7644xqFu0nKG09x/cb4ZVJMgHWf1Z3l2uw
Wh+lflYaeVeSx0T+ezyCkLJNWs3/FiCEwL/yl1R/VIqamJXRY1/xHpQn2OOd0Rm0vTeHgFWQujCi
jhhgLLn7tg7TdKte8F75C5x9eQ6nEXRuBP0pHpmrXhyBMfNu/ho7KgnWljzw6hMcNJGw19JziCng
4kkxwat/BapwI12z16dha86+gbj6lJJnnmMWTrhZW2jxPGLKjffoTrQGi3TO77VpX1J+2qUyPUis
awbaWdQHFA8mPxgteOuPADfcsZuw8l5fY4IpFUTXOYCQ+Bv9Wf93/AmYYVTdt/JVDYJ5WMz4U/ym
Lo1L6qzBcX4HvB2y3EvHn5wrw/D1rLiLAcWEic5dS+X8lpbxg+cQw+3O9YwBmpZaMxX4je8tVmFb
d0BO9veTHNNvZbclaxjrnY+TL50dLKETUim+omwNOTDsObZU8O4f/Hff9S9wh2fCZwQlCLI37NSx
JA3O126XTbrmtWk03kiqrT0JWzHqjrT6gdLRMVCAgWzF1AH8ZubgtGAg9DIK7SmoULH6l1sE26ER
RDVMHLWKs5C4SCePkRYP+iAUkTFFmhH/Z4BRmMxwUhYSsQTGHwsTirOPkQOD3yk8A7Od09uibBvX
YTf1i2zK/lRWWCPla+d1LwT3rR5APyzQ+/03e1fPXPEfil6pVMKORNqpGyGbBGm6oFwox9lLrvKc
lJH6Dv0zSApJL+uEBhAvoyrR/cX2iAB6hZgW1h81jREr1+6X/665WReLWtUVuJnLwL457VwRPdMl
MqXEGPB/E4r2eRmG5nZP+syRRGyebKCQmRCgsJGHpMqtouk/yrIlGz89lRMMDjX46iXJObuASo0W
bJuxqyoksX0+yEX2PrVJ0CNMP5abXRfQdHCU8swIEp1aAnez/BrYym9kcUseHqtB+fsrbmVx293+
ZAGUdE+IkRoW0A+tekky+CP+brifS88o5y4NImx9ABxUtm8s8eDFWbjcsCpJDHJ/PmoycKKno5J3
1tCta79pcRkSiTR+nk2ruziyhWHn7VN8RbPs+0ZctJ5SW+fcoj2QHPQxwY3tz/Z0b3V3ZhIJRcja
1qbNhH63zP/hgO8QRKBonPa7iE4fb25ouR2L93UnLwMHSqTtDuTXHgTQDM4yb9lMsDuuSFzHiGXl
7DyZh3Mox1KdR4wxhDWGWaRQAv6gBjUdq3etSXaoEklO5dK4aFeHGHNcFNR9hAuRu2c6ehV4a3D0
Xu9+jSNkXUFmOPZqTaGvw9rcVP4Nq1tG7/oCBNhtxLMSZRchmWvaQxGDdAVXo0Q2J+uccvhzgi1l
6XnjLAft6pTgj0MKMWmzkGJVF0i84C/t3U0PbNPtKQ+3wadZWxEEQfN2yZkRwTXyLcz6ZdVzc1SA
mfGOZ4Wijyh/FCqcj6QDUw+GSJDOTbU5GfuRowzdjoNOQ3k4ha054VrwWFiaC5Ghn6umJfwcA1j6
SEYO7+HOEKJEakvdbhpqBwah9GmAY4Ba1eOFU5D6o4blKHKPnJMf4e4yhTd2btEheFXwFv6WqMA5
DDSRr+h0X9sLACnsNlRF4Vb8p0d6Z9aZloy7NJjHiMKtEeEl2PNbk5fkRVY+K3v7GaZk7BTKutAn
k2BjpdsQ40q8Z4x2MgS1ksoqUhFuIdg8mS9ZdY16LKrd30SOsp9ZTlxlZ3ze20n1wlAIEGFNV5n7
qOvThppKAaOT3nV6eR7Ya50rw/cutAJkoB46awx+ZGqo79N9FYDOWay450z9mjIneuCPrBeiFQ2l
SsjbOG0zFp3WtgnXCC+jsekC6K+59wPGkQvOSZnecvsg8lq/EjK/iBak8L1o78TxC5fiytLqnth3
BqPElCMdsENhR/9hpWMGJBfeVrP+rpb/eJlPIgexNWaX2NebPXUcq26+3m3TN9tmZ7Ks/cOMAVcB
9UQUx4nnvDzQnnsufJSEM/ypgq7tC7XVZWj2O12Rp+blsx+/Nr0+yXOqWo5DI8T+tNAPJ5F6heb9
dBXU/Pi0WjyKBMSOgwE3wTEt1rAyFSD/SdLZK+AXmQNEbAZDMbYazDjG9jjKACzzjJv6/rcCMNna
ciNMmZvbXvW3eV9Ii+cYte6Y9Yzy0gfPRLeTfB9vkoRc3lT+lT597E93N+eEq3XJDXq7OmJwCyWI
JYuwRM6gKOUWA8vSxrF8ZL1zk8bp2isK9PUP2KyuO9FSqUpZUIae9A+ulevnhDlicHggMip9QeOt
LzdCLwK87xFZR2WQ6MHrJKrT7fcZqE0XoxeUo8qCA8nqJQH4kAZn9lZDVNoEpD39YDSD3mbwBafr
x3mJF0QU6vpMT2va6/uFJ7FylGqaQW0RLFGxAEtU7Cx/0S6Il4wwRURGRjJqejsYXG2ybopTb2cd
wX++ZO/ieRbMTuq8Pzdf0VTYWtX1c/oP4TBqT/vHBMcozzQr0TCmPE0m4SghtoBx8n4lLjRmhptu
W6ygajR4U8EFhhNJne0KXZK/3YD6geNEaPMEt1LZWMeIYoHjctzT1+tQ9gyKI7LGOcRhwNi90kXM
6bTxCr9SmvlEEULf+Syx2dWy9ZFog/9Xcf3mtTVr4my27OH7UplohJUOIZ/v+unFD2rHSzbCjjpz
G5bt+LlFI0HFMwXQzq6ORD5R9C4EBWl+DsT+Ug2Dwcfzn/8x5PVOvi3fzcmMfWj8j2f5/MekKX7Q
iX/EccZPQw8zMZso/mNncWHYpj9lcH7kl3ZvU1EgDr3iobnWmp/s/PkDfEUQl3PfuabpN5sWaHQS
7qLrgd4cWrjLfS78EOG2Qk0+DLcq6S7b1cpy0guwa8dQy7SrLa6uUui2wKXfmlodmxNwQc7jYAh2
RKSwZa4oBNcGEHo/tiv9tSpf+GdB5YvL/ZVA70nh9p7VrLWZNCcw/KtkhqE3WY2D3QbqEDNKJfeN
XHi2SnAulis01npXhJEJEVBCXwVLZSHuqNyulvcu71ZaOaYkpideLFrLbCRdFLE2KU/IvIbECvT9
kPHsSGHAn3Ti0QGzJg8GGiFzS5uR+q/u4IqcEFgt3danU120oX7/yIqXMpOVi596Wixw7P/hn2YD
kzVlu7z0dny8trtorfCl3gulDxjZJxIAP5dnA8VSaAe/y2vS2mwnsLk4z39StYqC8rT38rwDqFFf
CFORCWx4hXPNPo7sWQlOcAXIF5QSBtNeqPM4C+Wjx0kB2omv6VB+CVo0sbg5vIU4w2T/n25NJ6vZ
Jl93pQVQan27lgOQuqmroVOiQ6MHElUgPVOy62QiTdHHWd4xSXQ1rM2aGfKoI5rC2qmADzZSBjHd
zdYfHs7WWp7eJtGt/Oxps5iuboA2W0yce1SUBwiO78EAdjV//CMRx+E0jyvah9r32RbzORy1qfsQ
Q1O5ZsZHkYmqPeGriRn71zC+XOnmpHN7kOHFVCYFKtADUMyrCQAyP7DJeYYS6Mi5HHvowP1n7ry0
4JwXEOxYd1HjnbZk4EPrODK/qA9PUzszSr0z45OflOka8Y7WKlu7kgUv/QDr5f+9rQ0NogTQfOxU
Q6GC7LBosOTVDNHiIpKP8loTNhWpMyzGSJCzod1XTrrtcITz64NKCgY62+X5aRNg4o6iqPiPjXAb
yElQfX2YSJchIgoUyCtXN/alqBRepMmyEFmBCStohgX1OPi8yXuKKuG4WlWyqqHR4WfUNUv4I9qX
kZZy/iaxWuEy13KMMgzmI/qy7OMfprreyoMTt/R7J9mWLRrAcUCosMJteb8xDGUFdE09VFFZU3hI
wycA8yVFWH+rqHEsEbT0hOFJw8MS7uMpGEPl6piaZyNh4rNINx/r5hLX7RcN5a9UmnVHkXU5Di9f
OloE1X7JAOiziSrUvp7RR6peUCPQb18R3FzRfoaCjIqMXy3IhF+EynHeL71gWDLhP+fic+d/oZLT
D+m9lc32pu83PpupGObsqHD51lWgUVx05Jlba5oS9mnAZH9i7CM5Q1YT7Min0UUNB5MdR+tOcDTH
El35cHX2wo6yRRoB59JO9nmuzpWW/BrEtIVxi22HP4zQB/Zc92zneQmDhJ4my1lVot8NqtDlFgn0
m0vQ+UPBli8xU+UgIzO6e5pG6W8JRN2TD1JxcBAhcqKGoI+1al5stPYGYPP1oED3D4bqTKcmF5fY
JPow/6b5cecfnUasNudLlcgX1HgYvqnZeCnAgHnbyLHPl2+A93P56d6HSKJxcqUS0SqAGtxmXJAb
QXHB0HYaJlXHxHXRWB+1cyqBa5+ERuNIGDFUsfLypJJVirVYjB/5pPUbKSp4pBUDL4hwVOBA6WyG
qtlRsQDH4NnhhpUMPn1BcTRufJPuEQzQqlHTOtzz8THJnGUUZjjtaA6UdIB0X36bQIKBjyH+DENW
jMj5cmTb9QCIvNKrYZ8JjRqYEsDk2SK7TwPoCdxJ6Ay8OWbdrLLGCrq+qdmkcVJvruG840ioGa9I
5ACT8/Au/9jUjOu34I0x+yiE7q4B+ggs3umrOFIPqwrDihvbzNVk0ZqR9LM8BjF4G1uS2VrrihZR
9dltmuFthXjRNVvWu2gVmEvoI/cLX/BnE2MjvhRjDMCmFapS7sXnhk3KKR2Ey3Iioxms7InrtCAj
Ulw7nYpNn8HLQRDw6X35rcXW6NquYam3jyRdOBhHr5QrmLtW/eb9MYL60Xzr//jXshNPVFmdCEWG
oNU8PC1rubv0VW0AOihC0q8m+AIAacsBYGne50uXdcI8nJiO7qNQ9SZA8YMk8mT/KirsU8FD1+qp
fzHhJjC0KzO1nLy1IzLZjQ99NOSI2EOj+9i8A7vcCcjR1yI5YvkbdevS2ys5XlF4U6rdei/tOQD2
FH7MndehszrzueKYX1g+0MFu7yoSSfG8MnJPXiSxyL83sVf4ortkqT2WcPY9gSc+IRk5T6Prane6
b9nL80WDdKbGDeDOMrtFb3DpBLo3PzXN6KDxzKNdFZxz1o2XpHtFDzk7e6YRAe6dUVJaCQ0yOz4v
G92g9bCP/vuSVflPE/sNBtpAt2gMzqcKTuFaOnQz8XZDk14HUUac7mlPayQfT+PCR+Olg0806miV
J0FhlCxF1K7XtEqZmaXABY3O8AMgWZCxre9/t0Mgn82jaXx0JKx9H2vLj5hJCRGmBeoV2S0Cbi/o
SQjEiBk5DNtmIiJbz+6Ij6wB2oKBiJeSRoKnyMGDT/NrYlb5jlPZxdo2SpoKDum8tJmIdT7LGwVy
msb+ZCQJTLZBkGIq0fWDNDFdTReI2b6DykWD3rmw/BUsPbgLpGAJjmVsFY3gGdLWIwFAdE2fXOkc
dy56NrPntmQ7cwQSXrd+aSaAMYrRiqi+VcYKhr1GnvzIrPv/UMG1OCRoxJF55Mm8TicZGILfGGQl
26ksy6L2jWuz73XC/4uKLpet41vDjUxR+1DBPOHIl6OzQ+LihnrogMl2fTYjwq5YmRAvYLnqvTVL
vrVHFuL0/v7qoDXUsdiFClKFrv8otKQ3bzaLSCImVDwOSSMZpg7BiQRdEOSz3DRffeQ/Ah01D8R6
uSGarR/QZHTQEe1wiuXiz0fGTbDjUMlrbp2WkDngTwS3m2pOxZPmhnW2lP2ReTwJEqEsEGhJoDhl
dnXfCyuZpmDykTkDCMV4yc76WQWEOn/h7P3DY2RjULj8Xyy90VJ2SOIl5i/UoFU3WISQZABVKqd9
P0oTmNl+1rxg90/Bw34Yond/7gZPTYF0nF+jParaoAQ6qomoVgygFMpiFGckmwfAzYiMPkONCXvf
UPxGAdMKcdHLjLbbQ+fiGU3XcZ1/dIOs1dNhgEKdSIT5a1lNroyU4m/JVxoPk1yhJfWy+2a4P24l
iLIY+mQ8EPV9mhV9lZxcd8E+a24H9hH4D8uzG/8UX3YnjgS6bwXHJ+LbeRUa7ouN4eEtxHrUEIuT
4CnTegNEUEDHeLeJqP9XpizIeRrabnDCmIJs/hi1ajt3yKAciJNckwDs7l0XgEYfD/aJRiOxHkQz
1ORQp0i447cRYVmnnq/4ynjw1wr4c5e3Q7RyYp74H6f9Nc72sFcYhklftGJZygMBPP4TRIsUU4rw
MddWRsdk6QmPBxM3L5a5p/EZOG7iyPcvGHnVIBDkf7Q9pGQXYR65YU3/qpETwHCV8Ql6QeDgVlCa
GHjp5JS4McWEk0T+tlonrVm+RfvHiDLtYEJ8AbTVxuVQYAVDYBXiaY7O3+TbvMYd9InXJUp3N6aZ
Lri2iNhKzURtP/14tyjrsSQ4nZX5gTkgL+XyU2eoIy7jfQeV3Nj1pzzTc2Po6f9hTXwI4Ek2NAbI
0hpD5nKTvthL410rnNiyCd35FsAbYplR70CHIRjTvHICXemCWkQujibKt4J3vPy1Us06Od2V8KVe
PX/GOzPMyaTFTKZxX+7XCGH91ZooR/jy11kqUMm3LA9w8k5hwAyFHUIUGMA8z231WiVXX4w6sGtJ
u7BUp/Feqr6lm5YuwSMJAiU1NY3CLumOnuEtvuXHG4Ra9PrD4gO4KHF79+SVb/06iRjLRTKIuLdA
4RHjgSIDvWBCHHMpvgtpD2ah7dwXJUScFkmItREWbbGrN1fZw3uqSaBnWdZZGzQ6bB/o4D2DtePh
YzrAK0XQcQ01weo8e+1oBEbeOJHuvHzJMNCkk8+WgKFOxyi6GXQ4pKulhcXch8asqB0vYKDrwcOU
h9ZIXwx+4lSm375Iup4D7m5Qw/8GasDHVhDaqmKhHfC/netV+30kRLG/LWqYl/LXIX5+BFQY7wQb
qeqY6sCbNblnC3/yiVfdZ91aOJ/AeDlHyeJXLutAetr+d1+gxgeNsV1XNDNFPBFa+rEICjMM5f3U
FBLThZhRi0N8DjlNKl39LXwbDh8VfsUmTnCXHQajxk2has3slQupRu1IA8TxhNwCpOlF/4f2UlAH
IDfSrqrN99FM7ulR3ymQkRwCkqJxbioZEPx2NUpb7oFxFBwVC//03TW+B6z33eqcokg7NLuRLUZW
Foc8WtrjcnvsAfywFQTMmp734Wfl1D5+gdq1qTLc3I7ZRlIGxbO7rN99oFYLu6fWxXrAT5/V8xR7
lOQkN6d9YSD7dH0so6WRljqzykEZJYX1uXLD8jcp8iUcTldC0bQ/ippHzlnARmzNtEJHAsENLUFs
BtD5lXPWxKTxO4NB8rReS23fyp+reL1dSW5LBVm3PBnZXV4e+EnekX/9aKS0PR58qreCcKkD3FIU
dpAj7MhTgcsSxG9hTWfLOiWDXTDKpbNBDzqu4XHVL0PdlA4duzD4Ct0VcGGNQ08JXupL3YBNZ6xd
/7BtDuaigwrkpsb1iDKnYmroOtxqZEYpEod6T5kvR45JiVeRH8WME9f5PQETLKv9y8YNuJ7W40Yy
40ZSe/YX/gEWN3LNMONL7PD0FNlXrwqenSV+1a5Zfz7R/IhUJeCpC+OmD7fS6dxATygsZf0P6Apl
8UfL7eB8tMmSC17jA+MvwOYtaOjzybx2IY1wPazLsKr+on+5Ml94I+Axcj4l3g3Er9TAuIELfVFW
32e8hwEvmwUgpAge9mg0hzbHoPa18ypYhFJ4sHpTvcKgSFYpiKhkomPnRBVItzzR0o0wUFJvUUoU
ZKjNjU+mbfN32qZb2ngQYsbLkeTB6pG5L2ll7f4zZyRjnrIMFmoy6LfSY2s2+yp8IH0/aGBGGBQ3
yg+GWNjqC1KIeqiNi3GZ0K6u+ID3ZyAHt3x4dU7EBOmUooKlIgthhEFeGNOxzFSHkxHNNE18q0+O
5BZspKIDlI53AF8VfuXvcxu6LJMg88mOyCHQgV7N3C3oLZBk3HIkP3jL4qxlEyRyZFe3a9AOgIWf
JJhpyoSehqEUBKjTeCLz4WOD/55dZI3+s2bwlgOw320UGo/kkCTwUGIcNder36AQlp8F2BwOCcuB
bc/5UqWCisJkRyoIhNEX8F1gGi86Kd6YesiNvvckL5WrpYpKfpKgYcNWKRK3zJtDUMdoIbo046Q1
HykIi86fQ8M1fPog31sOYwizKVmzeAu0m6Pqj8A52gb5uw9gdXw7N8IKmt9RL467feUQaXahIntI
jpu8A9ouvPAIkTxze6BlzEiBklnIfWYKPkAMrI3miv+Tpppt+zUjWIj7kRj1JwA0TSKQCgVXUy9T
v/07al2AxcPCQ8VJs+8KDpq9iwoVdXJ5K7PoAyZwSFE/G0Q2tIKmWiTVIAcrZ8GlEaRMrpAqHxae
5ohxfFMq9aHfdgZ4rz6Uh8XQufSrbnH6X6pCsWbKsQCKSMCTkhjrVPe12VB3xhgE+ZbHZSbf8d29
2TizFuUNMRNYVtnCYG1h1JQc2dmEaHC2GXdgBRTqOnkAOFOSmspdEJTp0S6nQVVTHCFVyvicYW3n
tdYncO46A7co0183QXQ4svO/XWlMAHLiJZkcDv8rl9HUMeaoWpM1qvUx+x4hK5DwrZVZytsHo6SW
2OJokdXmUGv1vkzP5eshWTdoiGJR+Z3itUiR3OjAYtbQxbuEtYBHXNOxqG0k+z8a9BufAsEUBw33
uYe7NEasejMydbit95Ge5+LMbg6MJM2bUcFg+BIazORCwoyfud32+Op9Ild13HZFZENylp+I/7lz
ST/j2wPWcsSaJOdpCbo2PsCCkVzxdyGNjSBU33K65k115AKivK7q314+GcRqR3Bi/9+VAhvflVhI
DBhGfCBd4LfSqomuAZLrF/47yjaQaALcLNgmbWX7gNyEOMVjWgJNP1OVQRv6ekgXJYuSf0V/v5tU
MfSj/HzUFqU2U7QhHz+OWPtrIqTEybpCOeSQQi2ooW+J5sgExiw4IEuU3FhucUenbWSCklw6mMxd
qIQZVdsFjMacX2FYkD6a+EUv60/mG2OJ4bwJHVaojYoEu4saunx6GQx79jD2ciRbvQ/dq8ug5dwn
QUxUIb5B3eCYUzWdSWPQnR7sduTM7SnasX5/WjBJxSY0L3HHZTdTVw4i8g/SRn0BDx2n3CdDXL5k
WLFSApllCrBHnTbEpHHFsOMqmAjfaH6jp5VDL9il8jKwCnjFZZqWF9soGCy1GUT4X1Rylt7pW1Hl
MV6ar6HtPsFNKcaUhFHVBfXYCwzF3dKgikEkIUTOHLB+8Ukvwro7LGXw91OFy7+zKV91tj+aWCwZ
sAfhJ9Gk5NJDPIoyeI8dIFX3uiHKMgdugFOgWp/2GFspEPtmwVzg68PWg4PlnB3+91EqHRBq21va
di7MO17bDyfjp0f+JoX/7NxwP9GUx2ClRyvU+cC2ywJSuKQW75BM0Y+1/Vo4CyFRh5QhAE3+pLom
zNwint9GR9mPcaKWPSdPj8bUeZ5AdrlY/00x9C+MRLm93DdbJHYD32gXSQ1YliV4eei+r95B260V
ct//zaLDq/hTq95Cry3urNseCen8j07e+p+XsInRo7To1ViqUYZCrc2npvt47stiFebxDOCmC23V
pcJ2J+EMJf96u8gd93LT5+BCexUvIkdgrN1RpibLSb3YV3YsYDEHvwMw47ZDQP7Z9TG61KufH/yq
e094IgsBzTnhL7NvtLubW62pZuHPXK79DfZeMqboYxsM1WWnQ3a6NfNvuQZamQN1JKbul/nsYrrL
ALMYuvZ7InFYbHHolAe2fUCDNhXLj/XPAvFws6pbY5KbXEDM4jNa1GUgnxl79cVnuzCjH7SQcSxo
PPMakWktnFZxXVaW3ONTJFPObx/DCGofhNtZ/Yx0a1Y5pfFi9G8JFh0PeobLACNdcCR607BOEfzD
2/sv+IGVG4jeVH9uBy0bQxWc6kGpVrGj+zActapLDyjY4ZscJWhRoo05hHAxTqpVw6YBSA14/xSY
mxdrxk+PkfyKMtR5PqbyJFl2NyXbwOZej0v6M4e6OcUadrX+m3xz4Qzjsjz45cPhf/pyt97Tek3I
R5vVB2OA2Co29dTmnGr/0jcL5tPzCtjBfTyne30sf/VIVFlIqabaCK/XTieplLtPohV8xQvuGXBp
cd+Lnnk9oPJIY60uBZgUTD7PL8JseXQKxV7jnhphHNPpIGrAYmkDnK2fx6mfUXUqNzWSEgX+nzTY
gY+SxzzVOwOVq93ICHnDmaJGeyyHxXuSSYsc8EVYoJ6UpKMx0AtXENa0s+ZNwxS2aWWyrrllI4Fh
iXOCby6NC8mUd3DK9CtW5gukUs8epHt6psb26FOriBJCfNqJ07agE7SxObPS2MKhd+6SZrQBA9+y
WpMQ3Wb1J/KcGgHOsFCvkcYyh8AFN02VTe12vHCGR1k79kRvLGoNE+fzLwe9qpQHU8KXnbF3kRLc
sz2abKo+jKC1vLuo/Tq26f8YACKOSdhwqPlnVMHPhMckyPmLHFU4XYFjCN3Ye0Zvtq/5bHz3//39
2b/V+uN9trYGojFE64JWP61WckyQAKo7WZGKxsr+qojlAL8VtRYNQQcOI1GFVw4fl2ccS/l5xL5Y
/9nLMlAPvzNjAy9A+eoiqEUxO5tkEakMq36zfcXWLXknCBLxmDeARXTXfcOn8kMLN4hH8QQmc+iZ
r3ywRDgxd1FlGbgs0NeX6IX7rCAxueYjx9Hm0B771tI2Axg9C2V1L9useuO+7iWf4iXCiO69hI7e
VC35hi6xK+UisniMXtZuMqJhINdCJaMzO68QsJsvxaOssmRoEUaur4IEumIqpxhuxryNzgmLvTQd
P8h7SWqs2F5Yx83ab2LbwDguDSPJoNUpbRvayXx3msBDGwS4ygtUM26J0EexIk0CMlR0IQBGEgjy
aF4R9XSAwSKApA4bHO+WVlAnPEc4Tly6HVT85au577fLIuFSo9fANIMWL8VZEqjHg9Ka6lQjZ4G0
Sj7pIO8EWfSSZ+ZHRTrgLlAm578Brn7v4ywyLgeKoZ1iFAHLnVkdUblmDO4uw6vFlU27kd2rl2Gg
/gV4oG2u2jZEs6+htMNrl0ofeBJVkvq++5ICCSlP6LjVBx3sle+nQ5FhlqVx+IPSmfYa408g1NAh
S9qbe1PobR6imkgVwjXk5NRoTzcIUie59qn8vbGmLzwbiSfEX2pw8IkfxsMf0GV6HjUjKsFyFE0z
P0YoYE6YZ8yl1gYv6X1ANwH5vyAhTXNtRQU+RccDn65NQKXmfv6XgpWv+xbooCJieci/G7E5cpkV
J6ZEN7UxgmP/zp2Aw/eOjVQvk17bLYJclyB7nVy3tFTMPkvKgKYVh2YGbIHP/QPAUu9hvHdtrKXx
c8DN11MC7C4VqMV2xFhzs4W6Mq4/lV0vu+ARc28/JrAjJvT+YwKJB7fL2RuZ1dMBXuO+I0irL24n
1ErlmP+nZ2f7tnS+Re7T7aX01P3eiWe1BseUc3a9OPF3uwZ0zTty95VImalN0+wZColpC32RKX9j
YlDyYZW3UkrUc5Nm84Kq4H3RdHBU5Hf8Tc0BoLWyDKje7KhsGoEc6oDG0xUqUTPSmQ2dlI3Yss+u
MC7R/r7zJXLL+4gXY/IfcIipk1iU92CwlqUoGR47peYLc24VoqgPtNY7ur5yTz+ewJnUUOUg8N6v
NZdNMckLDoDPjhPVV8FKQ3JWuwHaVQrxu9i+lEj9mZkVhicAPjeNubqAjZdCKpGSIZ3TSwe5qFB0
tJp1SMTbLt9KwUkivfPtm0wuvj8EV7rKamE4qXlaV8I1+/ej6Vf+fJlst2soBLrX5ONo5IVtUdeE
o/Pi6lQU/t0q9/6H/l7pu6CRbpVXQxlGPa/bLK5aJ70b8TXmpwKBxysQl9MEJuFFX2/EG2DIbwKL
bY51B/QwNPcXQ9kToA/d6f0STU30B/DNL7goPEGp7OawQTMNuoNHfWJRSfOCiE0bbnKCzMSlNL1Y
Cr0SlajzzfVSQJCBFXW2ryZhyv2+f1DjPhc/aH/BCibLP+OMGkd4OAy9WnvTEGeoVmfGvqBdvSGN
8idMW3MyE+6Ua1gI1c2HRs1OmSQdtGcF+q5TbPnoKRllR5byS5pxhc+JP1eNX774A468/Nm0NkYk
d1VWzrGjzI4eFMS/gmLbYMBvgJR7zNUW8iOmHSIa3L6+gqsjTXnQ8UxoHCfK6scl6zbRsoMa1moP
Fell49xdLBiHQIBGQNDetR45FqCNtFBUs9UPkHRNqIzkb5uyz06FrPJrOh+ks34h/zwjEu2fDVcZ
Fo2UOO7aS46REMPnazcUg2QYWf6ZvFs2mrg43iI46yCT1YtxN+w+bizVvHg8jQ8WYSwKtqGRkf6a
+pNOwwmX4D8drA7RnOsJwfXKZAd9bV3QKdzMyVO3aDimViDHZhsgBaJWwuJYw1apTrqMiVw3n1Xd
zwgWWpQR1Uqt6Ak0esDYaQIPtpl9ZvfBz+Wj9+oTkyqFj0F6eJRqJCvUsJtasjmxBDt4VRyI52UA
hC8N3oW9lePxKqyNNdZ9f2jEZDCM8n4WuldG1cPqv6+J20zcPKrUdfL+jydEIes8qK6ex5aPRAsM
3gh3mn/r3uJRAHDM9dbW4Dtl7PxTxkBSBjpDKEDDMSvIrZ8ovVFvnxukzImt8nU3g/bgBNFyTM4+
rcn6JJJRDMka4bXfVVnDJA46sJ8xVn5G2KdvOWXqnwlGA+RlToLl+tD06HGClhdyO5HM1L2w7Iew
4gm7vV0u+A8mF8lUb/Kp3TMKzgiYhj79ySLMg0+NMjKC7rX2jWhcAAIyY7uSHLtw505Uih4EB1cS
/iRA6G3ReCLVc3n3cMyTIoyyBW+J/9JV59+hmRlUm74yUWBvzRJOj+Sne/38doxLp3LtIXJho+Nh
jh4oMNObg8VBzMH1mpw79vaAIV/P+f6Ij1J3vsPfg77QBMEBR7/PXcEmgWy8d2zNSJwzYckZ4ej1
DITknazEAf5grf4yD4O5h6NlZylur5z2BhXQNaWvXKbPBtH1e6HOHtUQDVEbbzKivBT4MBjjReQo
JnQLEhwiskZFXwosqBXG/fhAOJ4IfdTVtYPcY/7YXNhzjBs2E5BjBV/nQnprz5jAb3ZK6/GnC1a6
f7y8owOLUFOrg6LW56eq/XqYR1HoU2Z6UTUHnFbaDedfDhIIe3QuA9zDK9KzxBtVKCB8lyolf3+w
9V5Hu5rv/fOu71lffaFIhxqH03/LRdThLlXpZQtHXYzrTVLrF7WVJGKc/N5aj4xiiSsD92jVYzHO
qkHqMkJZrDNEx8RYGjOLsQj52twSfrutnPMHnioTMTHLL4riYqfwTlCa9LKt3rh5HnsMva3kJvpB
AyUWnF/ikPfghF9WyvqqtUT8EdW7z6/Qq6KIsYaZ/6BDtvzpcVK33dXXefxnsuixyoaAUUteI8Ff
M3FKJD2F7/UDomENAQLQxAPfgei73ziTnCioHvO//xMCWDR8BoIPf89LDazf3vDUvovKX1NVA9V4
H9eaxvlUMj+fnl6ACSCuIfy7vbyk5hwciOe0k6u7X4HplDmoiGL35fd6oHAiHmZ6uQD9vaye4DC/
hdPvJavdCzft0wl92aj9LEdx87y6P/voSDMICJXh3vlU17IncIGxaxuRJlRNBBoKnGZvBCk6Gwha
f0AI7rUB9BFlGPPxWx4iME4GMrMa5o6XkroWuOWywdj+C0FKxiRmgM+RwJqspAW0vF7vPlaCZRcD
eAcTtr3XzlbvEFuz+kk+22kvrLrWwZJzhUbk7TTKF8knkhwgFX6spNEYmhiiwsnBd6BWvzHA2HFu
wz9nnd7H/7Kf1dvfGU1yYKrcjRCOOio0TMaLIokPdFlx/QMhCbW5YCIq+DU0Q4kgpavgjjNeSOMX
7SmNA+D+WsDlNaW/f41H1XD1MAvqXoGE/XSUEVVbfYa4OeuNwDnfoSFdVwH54zBXNJUJxPgQVMWQ
cfG69MTAG04cLFfwnQ+BVG/7kFDU+eQ4mPe3UpOf8qwyQ9zIC0cgnvf6otIroCsvqIzbrr5TCzQg
jSfi2iGJk4gXQ5CQbBSMACccZUHFesxF68Zk1VloghN/6S1hjq+dZHZJsvUQSULjZ37fyYOTlov4
BU2ZN31xyAIDNGWNVu0wl86vEpuxauNwLItEEUUIqKh8f7S1uaSGvYKTjgCT/w8VNMhB1MtQko7Z
tt0V15BKunBUeAJjKgVcOSE2IQ2UDxAf6cjnNc16CpjAHGrJcx5OWc0WfsroYc8ZDSmbjVzoszAO
iv2DAVL+hX4qmt+r888d7l3JFJLUAW0PD+h+dmsLKeU2JzrDsSYH65ICcknrCIVeDOH+pOiNZ8nQ
O/PIGP9IlQ39L6+btdocVncmwyL2oi4YXthl+o94sX1aWsowHafDI36KK7RuJbBanOYQvPfGZ+at
qep9DMzE+rw+xRiJ/YGBfrROa8lvAsnv/mhlph1zK8iTGI/Safp5PQTRIrJThHwKWxYljg/uM4sI
1X0nr+34aJ4T1q1B4/BecprdjXc7OZUdyMgAypKJI9GlvQTQGe2LDJwv2i1JzAeooWL6DTHED3HN
fu7QsfbOCDZNgTaNoSRK4CYL5pNbovXoRqQdQdXZ8m6ONB+QvHrJY6RJKnkNMIh098LHVmOuozFM
CC/eZdn13zh8i1EOnkUicie1ERYTM8YEGCaJZi6T9CiFW7bohyogt47M1w7XEtQBT5cI2YeGD0/E
vz0/9HVGDrVLcIXsUskh4lPnQ8R23O0LIaxVkA8pSN2UfOUbcVrZNNGCVq0wAIDX6oOZiXsBjplE
mu+CMWtZugv/UN7yJMZCV7MIK8DF9pcnn95s6o2GRNpI5H5kb3Oltwi3I0VtxApxaSVFPLUUCyhC
6aBmMGYaHD7YpmZ1833G4H0Gpcgg8aJgRSuMoleIOe5TzuDChPwQ/KsYP4ozbQ4jkfg35SXwBx++
f7U++1kMtheJkMUhXfQhIbpU060bLUqQVOiFcCLMpny4JVdnHnEMTcjJ+YIpDF7S5sO+8+WJ6ybE
SLtVihmlMFRc+Byd9/urfsJwXRpjHU1lPJi92xiVM69BD2W3eDlgVUGG8T8mmsb6L/mlLBlLOazq
56AQU9N64M1JXic6nXafNCOJVMavIsIoTqAV7P6/6xnFlObHp+2GLyAVgm4Rtt/P5XNx8vXodigF
k6CGD13qAaX0Uo9fIuGnS2aCeAfL6CNY8iE8I+t2+G9Oqu2DaPEXurTn+wKd7Lon6yMZixSVgTtL
rD8G0KTSDZY1ocUs5TjUYpu4QsDeqFKuNdwYMGQuPhoQPrEeZ8zFOmv72r6enRZMZu/OvNQwURU2
ZuIwDUh1fOoXdRbgSzzqdGpV1xjB7HW3YvVWh1Dyn61DQ7lTZmqHuYZ2AJ1Vx/Bb4hvEMmii2rsg
g65BYw4QP/5e03DHI8oMi8/Lio8/YKEDVrUu3prWU3+ISnjLOfEGnIqv9YbPymqBz8zdJEVrdth0
FVS8d4+icdxDE+xG9vQ+2WMOdlwSTNScETtTwh2FmJeyj6zxdR3oZgX4mzARVrco2ZaegVNRBTMm
wXVY1Pp83s4xaOSweevJw6AdAizc5p7tO7ZEcyi63+Ob/V2ZvjdlWh68R66a4kAtK+Q8EJCa18La
ORVC0WV7fBLCExRD3092Sz3VTW5n8e9oCIqjbqliJ/GPfAuI7L8VkfqmdjClPu19WwI35+6qh0hy
ro9CSGzXPHkG8QzFkCFwJdrQaYnh56vxnbJCZ/UARHhrVtIaws13qoPg79Oq4wwT2l4427NOLzqn
t4jxbyJ3joUdn0EpC1GOK1+fd1kYiTdwFw+fpvQ29frQEo82mfVyzTQV2KzFemH307JJwz5cyO8N
LaoLHR5b53l79RVSe40tbdIPqrlhoWXnNbX/HHhejIqy7d7iImoA8fusAjlVeW7Utt1P/F7+ZQpv
bKf4lb6xB4YnV5FaAWylNAl8JiDeyE7e20Jv2LtRHNu7ZLzfqFMGUxa7TJj16uKGNxaWlM/5Q3Iw
jQ/KZL7Oezr8bFWP/XAAsCZThqfHKSNRxOEUb6DtnGbA+PROth9mKNHa5O/p6BHBlGnkawx5xMXN
sz1FuqzZQTNe57POnQKcUQjWWlcVDrstaw2rXPqcSFS+Z159x85pT8VAiUTz1XjYh74xwaZG1yRn
wfLqoq8di3VR4n8xWqz58x2ik0XRBVn0yfHeHwtrIiFMQU905aY91FHmPJ+xkuimcdyVF78VZjnt
jmiJ8IJUD2IbRPbDzf3ro/V2tqlFqGtvLBpQcZWY78xRESVfikn2UpeCZAK8kE0Vrff6+VBDG0fI
vzgWot2GiNJhRquE7J8MlV1vwQn9IgKedGdAAT6gnmwggdVfwGZZg5DZTseovrCE97g+5Ov7lFib
D6XH+KLhXlNomKPzdxHYP0PGw5ink3OCsVcG6UOtOWNsJ95mFSrS62RKt/qLGBKV76da+h5XBvBT
8/1c7d4w5niSuOWZbK/RYHI/Kjvcny/Sj64kpRmnvJXYmM8KsdHnSNeAWjjgS23pBCYT3ey/jvTD
zzwGg1JeSIWbhuNbTYULtpy0fcQ0rs/WVSzCA98rQifmELWp+pzk8AUjW9UcWqXh8t/NPFLKDk1E
sTsk4KXKTrMVEqkb1G45rc/xsbNMo9r04IhBCnXAdscz6p1gPd8D7IGhB1dYur1SUnSwqggQjhKV
C9Ql/8TOBK1ay3PW85hg4NKjsb1wjAVQ36eHvbucBFDu0WM8crau0h5nUogHtVi5OVWiuPAdJg+V
ELEJxgbMQhzYUWq9I26n2SNHKDiLpiOeCmmLxNUGbhB6gfSovukais7BDT92fqkgjmwPRKJrMu/D
Qz85JcrCH5kBMew8uhKqH136DdXhuOuWjJGKwcYCldG6HPzGIUT/37ztAl/qDIxru0IxsIA9xkQS
6Fp32zhrrrRJhL/dHwz3YEz5cs+aNJjow4cPvvDjZWPaCxpmzAZZ0VhTXYxsuV17ZjorOI8saroG
lMjddAFChWgk7dTC5ydBkv7ULWuaQtGkP5e87X8aJfHmOrIwytKVUias/selNWit/tOYhSByNB3y
kbOKBmbP4XRj3y9sW4eoGIaadboDqR+3J0KqVV5eOBP7qaYOqbSaUokOlcK3rJxUARUYaXeDdwsZ
+5TGZ69bWDzZdSZ0nEibAsKHxUUnAcsixrXhzI0bpPpa1lX7EjEMo0ELPFOkinJdPyl0evcCM8aX
lLEm6kiW/Gf3bcCmGbC1LPBnxO1vYA9JbYPeE/U++wTWNWS78VehM6EueGjvqxP3nErqAiANatve
XpeLXVf5fN3ITLpPGU0FhjQ+gEScadkpHyi1VXyoYH9CMF6Cj9SBR1nKC2Flagqz+szcKQatFgyG
JrD17CMzswNt+nawSOjll34LWhEFc7vzEojoQTogaBGdjLzx2nR8BMrmXt1wc9to12yOFEzR3MKz
CjRRUmoUIpsjqHRwrYSR+jiAwV1lrLD38PXsr+ofcw7SxSpIp/mFXuhD9GDF2uvTvnC8NfNxUwNl
9CgvsJQzQ+hlj4jb2o/yzVG6H3fqCqfcRbGOP70ptitJDTVoVpStXHVE2tF9/TAwFXx3uqXtwEuN
IHAM5lkpW2339VvqAzR+WMDTh7KAZJPEcYPdRa+I9xI3vtcURJf649SVZxCpCIAiGtmPiSI9gw4v
TxY8GYmbgG85jVu8gwKJ3ZB861Yj67yk6RPaC7REQJGPBlRShAP0jUHtm76XLFrTEsg+oUyG9y/m
XOkLgn19VeVqWjiZxsKIFE7lwZ3rfLwov92XDxgWYyWy3A9hClGUTqSuGGI9wEAsDVxOU2h92Abp
PIf4zJ1wf9eOHB3hvaCQiTu5Pp1cfJ61aSkz75tR+Rw+ATQ+mui52Dpsjo63AGSdYMJrcPDfb7l7
ILxZrD0kkdBSmWhcHKgLh0YU+HDx4VaLae4cUJj1P6au55JiACx0/p9nvuvvR+4hNoDt8j5tnAfG
sPt85FOZfOhulYBIj6tHuffxg3yiEz1KYL0+GnqVLF1ke32Vwu42U9tgQLFXbapak0HVEvp2sEr4
Obqs9/CsDt6URfhpQ0Vaiy4o1b+/oHIUzd7FDGFxpipBFByTfT7HS3cXfOwrkxcKwjQS3vXE1hk3
9oGG1SNb7SksSfeCuDOnqk4j88AzpvD9z30DShXxrnCdr6OmObtg85kzjzZwTk4ihPuU22GT6Tku
DHf1HKjzSk67a2otC4Lb3bAY11FuwW9F+CRyIUecInyY3WF814tUA+vejvnCfysZcbrvC+552tqN
+Bro6NueQ9TJ+9d8OJ03caLD/5osg+D3CLWKiFcjVHX53xJANV2b8I1omPrcX6TJbtQT6EcF3v2+
gJZTtvENqLF2OnXXmrsC0dA+dAosEmzrkP5Yt2StMoDKAIQXMLR1u86pda2Ok3WdXjNM/1xo7iTL
HliiLM4vX2ybbJhsFpcwMkg/xtUSHMfhKn3uGR6PMIY+D/ZRV3gG8dy88P+YUnbrOal39h0XafuH
U3uq0UtF0U14PVbG0q4sIrlPFlKR4MAEutD9N7ltCoH8rAzKvVc3Q32g1+c8oCjik2hdbJtyHKid
9UF7IJ3FPMTGlAFzMDlhspGQewcLDuVuKCuB5LPywkGt195lKAcZL+ceo0QYxn6x8a3X4VapKfYL
POJvqo1PgjBHu1UYp7LdBT4lhLVBDL1ublQ2SFROTwDiZJ2tbsAmGA9HJWE3H+FHE6v37zgqs6qn
PuS0N8jRqDG/eHSUjZXAiKXXF63p9X9JFm24GcWLVxN+aDxMzqhiN085a3xLImWejfk0P5w5BUfW
4rvcgh+WM5XLuXIwEfbxkMR7l2OE9F0if0zPG6NVbQqa4LreCUqMhiNbYW58uB2RnrbTdeVCwDT7
ONoJJTVRUmGQxI+xkrnjjwrwyJsyzcy1oLbGCn2OyCB0KWdIIuVagqh8PV78xSJ4gVEjDdaz5z0n
SeEr8jVwcNWungEeHOuzSdif0MjFTYFIdPRER//iBZdoLD7bL02DwntwOh2YMumosWgZuD8cLfzU
eNZNiCrGhgpawRoYQs6pZWEMWAAWJQJ1L+3SWELitm6KCbzj7UoyPixx3whbsQEkHDWW7islxciw
JyLfqu7HjnJEHO64qZ8sbcMtdbmW36GN0JhqK7RqeQUiPDphDGnpmk25WhPyj/ut3HWujFTXJcP3
YrYMsWTAEr8j+KpbgHnPFqfal0oUEdEgaCuFfIuFmwfEwosKZMb6mxCdyXuNbq6aUemyxwf63zQ3
kWiiHK79Bu1V5uNCs4KAm/eZEBMsRLWCkjBvwPDftHfRns6cHoBg5jA4f8nWjwRkFecZm+Q7ZwtM
usLQqsrD3W1kiOYhxF+/1plpq9RjWP95ZwiuRjKKStQXjfUs+putpkxihDdJgHh4L/qOdkOmqFHS
3eeacGrtfj6zfSjfV8wxyAv2J9OnpbwLfDeiL9GA5LDlh+8IUvSo2HO0a3g/+QSVGr7HIIN+VVWP
AUO5WEl/1QGOxxdbimPA0J7TyuRMOubtetX1q2qHxTlVmjkSAVgIZ+KC4cut8vWk505Qn8MXxCMp
hlqKOEPkr/Vo6EkLQOXDoSC72KkBxRM1/XXdiaA0QDW0VcQdiVQMjDeLrQflzwMqR9C9lYBG88Ac
+Yxkz/ttnJXSYXJGJ+aUPp9QusSpCiEgSJFINeqHQA0r2AeJx3EKX/Ft29bPK7zrSR2bv9yHG6gU
n5ncEaD64A1vBlTRdK9h4jsSIOF8Rhpc6dcwqjI4McozW6np6JDhlUsmuynBcIEgKru0sx1l9mv+
I7wtbbzNXTg9jAazbhw+990t2qtfpK7QxKuReJb5P5KT7AazweIFnwtoMKQs2FeycNeSjdnXDSUw
zd/kYrTtJH1xUO3J7rbABE1ZNxGFBugpeQjkwRSHc4CySZQl2O3as1OJzbqq2iADBczt2o0HwRhw
3a1nEPoCOEgNebtSAl7MNFSHmhmM5/XZDV4XKLTiN/BPcgnw2Yyb720iYuPRMEbpdzMckDnlkHPD
Zcf+0WWxE7dkIVTXZKkVE0Tlodr0/m9pw3nSNVJz1bW/IQN02lhbL9LxNtijj/sTMYiiuJ/Ilcvn
55mevCyN01P1vVWo65uEO1aVn2wd7N8CDS6oe0y0mLtiHkoWmhWVkuCSRhbTpweegCxD5hhW9Nfu
WetqKBsTTX9ycvWmR+eTgg9knkqIcX3l/6TcUFwTO7lUKDQU68t9Pe1zvW7qsmtk43JdeAkOmR+o
h1qXWNTCLpiBUBEOSpQ/CDG3DyC7P45WhXQrJIw7u3jENp0oDoZjRKUByw5/kmTPnpH90ZM73Aay
UksrHxEdYt4G5aQmBf5lgpTydhX9sBpTrnz8kAoqIInldSN9nH0NEfVz+aSRd4rGPT02einA/1aD
dDtXwRy5JcltvQTOQq7C1lo8abhmDFatVfVn4wVyan653e5IdlD1xMkZcGpabWZLB6yGnaAruiOw
xovIMa4wniAksKyk68JW0YEjtY8DRnjrgHdGQXn5yKomCJbQGe3C2NV15Fg9ZFJZh7jTJJHDRaXt
XIDpaWbIYfy9uM57HMJGw3GlNxE9UmmUEBfiGWDYYV/VL2vOGVcRs/w0/QYpJF+8FpWYWF3xl113
QRgKkm1AjSe+7XkWvHG42NQ7o9ALhED4aSFUHDDhxWbcfEHwnxCipk105mkS4QtwbWkDDF35+tOp
XhFx0dDAB8AqzvajsY3wNvEy43QdvaKWrASglMpvoMeAlVgRUu+iBm3Wn9zbaLAFUmgsnEGdKah2
PitLCah/6TGzUcjwpBmeYTK+/R5hOE4+nW9BawOTCM0jdUQWvqr0Cx3A5zR+M6SzRbbpVQtqzYB3
NO+AT0abr8aghxup9+WZA0HX9/qhB3wdX2JxoflUUgr4v83qUAU/RLuyaPSu6m4Zp95VKcEfRznJ
5owrDi+wA13pWmRRV9rYjuR73vUvzC3aJnr/RcychVQLYUvZyCiuBSpI0OAYgFCGtDx/6jZj3wU1
5ub4D8pSaAru3nWOMeFsYu0xS4hqQLYsqriAKZuz+KlJZg8oi79DLz14xOJvohWNPlPLEwHvfKDt
lSunlrCPH9BZHTJp57wEWdcFEjppQ9yi0iWM7xH40/ucCG2HfT6drFtAcTRfKXtlAjinHDxqrGkt
+ouf4CqVRND3zJfpZhFAWsJFmDMQrjD/fgeZjFRNK1ZwUXaRzcRHZ93ndVtUcgcnO3LMUkwOVVLZ
AMywZL1YA3nHS+0VhKKEVO09xuLwhFM4IwMFlOkJpe7bJHGy37HQpB7m4hAYdqeHw4D8Ftf1gLh6
pSJEBWT/qM1hNoJrkXhUnhhA9PRtG4r85XA4RKmjoUvZE8XT6wAvUXzod0WW4ac0Cxd9j92kpBTb
d1kgKDq/XM+3XehYos4lzoXNmCfn264e3/Mn6BtAVM0tFsi4Quc/YSnC4Lvb94fbbKzWmOcR+mmr
si108/LVyayNG2voz7hSvYq6XfZlmtHkslpKNI2PHnTYEkGsSKP6TG5s6Bg1QHwzjmE52IhZdSNy
RfartdODRdXON8Tsy/WbfPiopgNwV1rBath9zX9LocU6AgGrfGXwKamu7RTr4O8XJIIZMInvdkrc
MgxNPQ19VUkLM8ysM9xtAWjvmA0pdH7DThuF55UZ9I4msTQCWAsbaFEMzoHodrL9XZ3djCLMna1B
7j9WAlWxYe/ZReVzxydA2OoE19HYLibVYOMO5LCgRt9XO+7p/HyeEUE60cPM459hjKsq/d6Y/5yh
8P7pnzscF9QsBU8VdT2hU1qM3u6KUlH9uhe907FXSQ210Jj1iKRXDnNNod7VI4jjWStu3eHEZwB/
Qtc2ILn6EKTG+mqTSH7jkxGDiHiX0HN/oLi4DEvH1Jwu4ReBB1v4kWfVO0T/mZGJ44CONYFwu3XI
qjPJMgwYSaR9SmaZS9jKba89wl5SQ0QaXwJVOnvkyJQ8Wl4pJoGO9dwI8HfANa/DW3JCEN9vgCH4
57dWk01oqxtld8fk4fPaMVmE/aK3WoRiC6kWFQHSqWAaRQ6XldnAZlLboMbkcyywk1FdlbBMyKcf
qv4MCgeMUq3eFTd62pmwfMf/wjmo5uMiTGvIqUUqevY1nADZDfNYh9qhKGJEwjnPK7FyvN5tYNq7
UsivL91h3xsZqJNdM32zetv4B6sUrgEkmu2h93fA3YyUqWQtrrf/Yqun01dVq0cNWRpPzRCqvpiq
qweR9Cv9SlsF00vrKoAOOQ+C4YO9MH+p4NoxQzIZizANWGViru1DhjVK+eUc9usTM31uAN7rr6zc
1tschNdGfhcvPI1+HhJGS7JjRNMtRv7SwCYdzRPLfF743DF7e/9yH4P57DngqM2rCDJPG+H/4zHA
Sac5wJrqeIMHObBA9gFtEV77l17xnU+q6zvtASMBZh0Yxbp6Dz10odaO5Pr/vVFSglPorqHYWsJJ
KrapjCph5+k2xHDtYqdRghkKo84y4S2inHEiIQZjpotNPcPMydHQmW26tKiFo5rjLSUrhEwWt/3P
GA6dN71MjhuuJnWz3PVUwR1IkuLGHNpwsBgUGADQWYGL9Yh8O6w7GLG54rjzNXisMKsU8wplcEzv
i523+o1Yhe5uE6nUNqYHpOxCRVPh/ZVQdn0ZvPJrNy6HvOnTr3YBikIVA9mwMUjarrvDoJPyzRz/
l/L3hGBRToK0klvm8Aubk8K4NmHdPFJuv5eBJy4S8tRJ2ivUb1IUTAX+0QembVFuA5ebDISnxXgC
GuDihcixBLVpObBYZtfiYEJ1HZOVQ+8wpEy3S1TOT3DUKEFjOjb2XFOFoeIXazc9V2QEy278tgF9
CgKqk2TswXyU5oXk0woJLXGz48t5F9sGD1VijWYv6lx+zdg1xcywk44/7q+KNPyhLOeEiWInzqZu
OMn6I2EBMYqzzjbUAxu3GpClcD1FTzJp6f9Tc/DGm59Ur/hr2kLziaYsIAA2Zt5i+piMPRHObgs0
ZQyxt19BBNdnJ3WD8TKxnZR0XYrz1u1JqIcOPe4QTvLaGJjzkVthcPDC6eJyBOLpx6Xzu93u/ijZ
mHnR8lsSENNxRbRE/YvktlK69BHGHs0aZVO+7w9DhW62auXyxCaloMJl4Eer0leM1zgkGksUxLhB
Ztnd/gOriN/1E40CNGUryPPQUGp8tUmJ/E9B14IyOMdtRb6HUtIHPVG0WlQhXpXcLDky9DMESRz/
c+pxGz09Gc+4r0yVZSZKcSXDhzTHHCyaKLLVoJydkfkeJRnlybIa34+X38gxrv9OvtHWsjKAxnYA
avI+SDNMLfflR5M4d009F7JT5wExRzM/YqfCPmckBeGtLoGBkPXb1eqJj/48+quHo8R3+8my7VsX
NjWCyNOqgPL/Ea4swFOlfpKMN82brMTm1o9yeij5gW5GIz2lvU86b/NrTt7A1RO8bS2zRmNmZn8G
4LVQMenAXzCwD6KXCf+7+Hq/21i63wPU5Ro2rN4ZWNJBllofPw4m0fdOAhmfOpUUnIUHz42pa0p5
tSHAtbMQbH/87hgyxc6SXLOua3DYiaZnlAGhuIMAwZ6mGz5qdZMWo6BCQjmshPet8x78X5TnGMt2
7aIjeuv0BUF8yIFiP1GUSml8Qr15c6kp/GiIJEn7vNee/c+J7TDyeAqVZsdvWMlV3Djv495qRKVC
YbteXNGyKVKvpYLP1T2CxUPtRD8Gt9oPuIxQa4n9V26/G1MW9cXTbPa5lz3FKyhGU6I1vfX2ny+D
jdVGEqRFckq90/HRQ1fnnFaW7JS5YO3B6VW17b2tQXJNThVRz8MuT46Kl9O0HyKBvL5OH3a032hh
MAU0QPvoBhyLa0hIsiO4fZMHdQIvhkk2RIuRamXAB6c39OB5Vspr00zlk3EmbBm5gi6K5cYo9fbs
2rHgaUzuy19eBmDtytCdvkNuudXr1dfLz3BIPzSLAR2dwtdPxuSxMlV3ZDgqrLNs0i16XHSwvdQ/
pTMBIp83M2tlnjNMwXt4HgaZS44VR5QiembDJTl2NgyQ/t4lodihPECkFgc2yvVJOWKXB9S++eZr
IzAzxVfrbev5nPk9oqQmKh2Pfq7TiNVIEI5GEaIcLPeBav179D/M+smZnCWNXdY5AshJztXQSSfx
jEQYFQ6JV3If73BlrjcgtApAXnNbKgIvqcsViBPWLOel9I8J1bd3U4QzQe9vUoduo1xSZk9HIyo5
qRZfDkp0AYjVtL7YrRsVYR7tx47/EpL+9PuFV4hYje2GOPJjoVuPiHhdAfoDxEgG3daKFZGgB8Ax
Y/zws5ht3ES2IY1MRuNP5hVaysipO0nd+WmfNiW/DnHdi1CUYM7cRVmHUs4la9BBc3f5xxZzeGsD
nw/1bFyKibYtjkpIN2W7We2on0FWe+RP6PoAcbim+oghTtaIuJsLJSRuvTSPzl0Ehlnn6L9ed+tw
6Qw5WpilVOba/S2EIKw5j/B049ONL13y6Bd3pAZxr5dogh4QD3yEgIF8ST4Ao/rJZ68rsta62JmL
YzgkW1G54zTCa9kqVl2QghZjh6d0fFWIDN6hZ64vOTGFR85YZ/Jth1SU3HAXLSm9MBGXEX2aKgnk
yseAqSTr6Yi4SAPi65Ev0XVx7Sw55l+CrzHjexZFXfS/GA6XQo8VxS0OS3KsO8DobKYWXDLD7nZj
zgzG5vU1NDgdDm8YyL9g6MzXpQ70Vgca5Kovc4GCG8jAcQoG4jRSDA+VNzny5ucMbLq8ov5ZicnO
xmTQqM20CRc5P/CoH70rQYBUEYGJriZ42yb6HjrGaWkPYKfVPXEepNtqmaa3aRYf73J3vq7IpXwX
09uuWZpDbAt9uDC6WvbZpZnQuUsG8JeqS0oARFihbU8EqmL5eb0tJeTjM5Wxtn6iq7YWIo0ADM4f
YnEO2DVbEnu6nQF3MRI0Xplw4kBpLrMKUF1FlUdARmX5VrnPlScJq6GKLzc9e+bofPBGWFGXWhxp
r8VgqmknBZ4sUfW2Fpc3dunpmY0EBochbVbgzaazGZZ7hfVvtUnJpCAH+Eck1DquXI50nt7PNTmV
lsMrSxcBwCVU7qgZaKe2KeMSdjb9jNwdmlDgSijnZxZTl9rbNiZbZrlEpMRwqitjH0p/QJzI/6cY
YV85a4VJMi9rsVy1D4ebqOqal/0f4/tQ/k+BBz20h8kJyUZubANo8D/ant1cSBe+GTDTxNn4Uf1P
WsV7UqB3Uhse9Z327AUo++RGArJ42rsAR0kpimB34gMwICAflnX5fhWP0WZh/SRjqsnhLwtDRZgR
mzLNaGMsqeTiiO8W0ltXYGYX5yGRQJYFhFGGLkuefga8GufikYHhdgBjaRccqlFgMOX5GwiGcJ+m
CzolXuoTtS/1prLem+3LEKoU1+73m+2Kzek1+AVIPGyQ6xgGdMgwm+4FAC2ieMz4QkPND0UdxVXL
g0VT48xBJegYwnVaE34JeMGHGuijcIRgY/1yTWpW4BFGGVkmifEXlw32DuqcSHg5p2cus3sqUvlT
cEhAfRT3Tf7fUj1z3EPk4DcDWijX9MiiGA8RM1R/A0szL8vz+I0zcscLngS7WFCAQIS8sxElVB+Z
EIfHIprVG0oqrAsEWolm0RRfyFQ7heqOe51XY4jhtRNY4836PiSmr8LAUCFh5B02Yc2QLCX5anye
sfmh+SPL80RYqyZegrC8wJrqz/uZuMrL0dV4csUF42xqZQGFQ7D1sE0R3kyHcB/H29/l9JLNt7Vh
dHlbWzD6Td6gUTve8Hza0OaKWkW/A+BYKHFnyhk9QbyF4oJvfPxkx8uVet+2Suu7PsdryvCMwu83
+L0scSrpm7diZFnRjhWJBi6rWabtokc6+E8ka2CKc6aie/VfRNzinQnp7gA9MWo3EEXCIItV8pQr
II9R9K6FstgSNLIsZ2pdTet7JWvOmOmPOSN+VL8zWTNNt23cJqEHOHMvAU2tmsE/607+G9JkbM3z
wkJXvYhIpmFY0RHTqS0EABEywJPP0ATJ8FY3UWD4K4E+iW1wQS3Touh8qS/ftiMkruDofhB06lf7
bVKmPGH57YGaPRX5N+r4QgUL8o+0O33daCWnaaZzyIsm9YtxZUtH/ck0YvwGjYPyYjOz8R5KcChp
aPzPKyuzvRuRI89vgOfpKo7PEHMch10cg44M7WCseW8I1H6ChWDpWQwQDa2xs0IAeeQcmWtMn590
kRCLGzPKvnXlir7MTsnLLlbI3FuQtjOHFyv1knUxV08DwoXOcKdS1kU0Pf1FwiXZJwQlfeyvMGbR
7YdHF8IPSWF6qRBUsM++RhccEyr3vH4wOKqh5wOxr7esQYGC4WkXSwv18JMrAGcDJnDKObc9mJzb
WYvA4awDBWPGA9ckM/K2BT3gN9Rt3zMTlgXioHrAqyZaxf4NWVpfO+kXX3rNR8ZpkNHCyLprWAPl
uwmxsiix82NR5x6Tu4rXAoFBFsXonB5w594uWTxWi3NGRc93W3tsurvFS60a06ZZ2ADjY3y3ldcp
c3vVBIEpFSvJMiyEdaNW7Nayj0B/42Lg/5UXUSBCDqcBfozJXMgLRNyJ/xYjovYn6cDi8wYXBxIa
t6kDyJYNam7Li+l+Hwf/QwSvgIZ3yd7+G52mOKrjnWcWAthd23WyeZ5MuygFZY08YORcAXRik2FG
0MHHh+T4M7A20yqZZKiUsEnpnzRAvwmEnWAKiJjR9qRw6qJ020GxNtuqagfG2pMkWt6IJfS3z/zd
bKUOb+bCrmxnqq0bEvG57ykYm1ND8A00a01XTp9asSMqygUTKP/NrQ+tpCmTlApy2oOL9Tnrit2v
oaFa978djww7Ubkn+4XRoDcmsHwXb38dTgL3JdLVkbvmOBgcU2Z1IxyQoP5rRHBegBBje1HmItbd
iTsrKMzIU/yazOzCatWPFjV/y4Rb8noTBv2VpjRGBMlZ3+ECm+G34axm8b2TDJckid3MtPlWeqCH
cteiU9J9Y4LAkNc+e6mdPswPam8+BcNbYwLURjojnjWuTB6ts7gZ8p/d9hj3vAh/m1AUjJpeV/gZ
DUHj/z7v2REaJ1+mGTTwPHV/TfX4tnrLNob05KRuwnIxGhS6th9JmVnRbXfgYL3yv/EAq3EpQKrI
rjQlr95WQLk7Fmm75mMFVr4xlNuMHa9g0gpf6zq1KB9mLAIcKVDfKy9YnEg829Im30i94RGK71GE
1GNhGy9T6/rShHQyZ9noqG6zEULv5hpxlcNw7AWBtQ2NCkkIoxRA8Bb9Gk6oBiYcjsbsDGNnMuaD
p7Qn7SaKLkaaU3rjMv1n5Xa/QVHYymBV+z0Rk7FwCmW+VXrC7jggcNfJJHh4HSChIKVsKr7f4/JI
B2WFftohQBFw9B71PW/al0ZXbXfFhtH6gToJ4DaRZw5rbPfBCe9twHsfPAJRh+7NgUmZ+0M7dLtD
aG3HrP2kdsBOvdcstsNMDTYJd1WwCMCkf08irZSgp2Fre/Op2rH3McDxorfhs8yz98k51B93RTNQ
RjU7U7NHQiGvI3y9RQhb+7wXVds7epm+ruEueTdKj5Nr24ryFYZ+dQrQ2ekally8MuHtO1xToWo1
raawNUIqGjIYl87+h5xzHhqhkkwwxVqb1HqfuFztmnW+ZMI4gCRzR0da/mXqWRpk2dLtT/uuhg3i
1rrzXUvtUWuaIQ4QMp1ssGukXWmAhqAB2rM5XNAk0yRKyEjjiBiUxNPzJjYzdK15LXP9pb+okoS2
j0JKtMoARxBpGVPzFqwdcEVm5NtzMDb4zPelEyW9L2AmIsZn4CAHKCbvljdk76sM7XkAYP14Dfay
U7XREFBLsHXYumiPPJN6T+Yn/5mRpyydonYVOuBL5voNFIqWdkDk0pKvJhFZFluhAmgF8SyfT1He
1d4MPrMIDp8ebriZYnRTR4jV2NXVWiXmk3JwGxR0LF9yojHDlTncIGxTpUBvyems0CcD1gDe2dYO
RB8y+nUdJOGOXE1+VROlaR1ilt6sU+0VZYXV2//3jCYmb9L4cmqcvb4FERrWQa0mS3G/4CpQGjtO
LcRk2zG39T6ASXkHQ6PRsrNwU8UtPsZmc5Evcvf1CSikmAWLDlxpFqyjk7JyqZ5KlsodmtgddTYE
isSSe4SGeBwjoHot9gHbpC9CMitA5vZUS/150zLUiBiOMBWuAn270kTrBARdW9t8WDu/vsOgI/8A
/kzaAOA2e1OfWqp2vANvGUtfRgIFZQkCNBBF4HXS7ClvZZYg1vIipAy4oCiaJaCTKPN8AvaLn4zC
OevOVzcfG09mdt13EsLt791JNB72auNlH4jDzQ7ZduB+5W9e+LN63SfilEqQVxXt2zWaEjeGOjZj
YHKK5xtl7CXgMvjHPC8rMoozBEgvkAVo2u6Z8sS45ePjVyC9iQcYjh5CjDD6V4UEvwlXwQ/kqKCV
a6h2c7NrJjz/WB4/yfqJwJ/C4YaFTswM3A3DwDJ14Cd3tfle7lk+ID+EH3PuF3a2yr3KZf7berhv
FD0H8iBo8PPLCTXJHxhSz2W9lCFsPhyJrOQrFiXobgBTgfmpKKWpBU56D4bwcBrO3EJFU9wkrgPq
1Cc0g6dsmKU/h+PF9Cj0HuLyvpahALB1qg8kCnI3AZKtzhSBXjaxMyRwyT/K43WE6I1ByIl0GCjp
pi0rPEoqdQ8kkfp5waLaYx76lqIxjccTeB1Igrs6xSfyD1ehm8CXKCWn+N/JUlUISa4fcjnwuD1e
lo0o/Z1drN2MYxxMJdtIy+Mhn2dERdft8ihMHu5+ZPDVaoVwJsfJxcDqf9/u9KGjlhtHAuQGx4lT
ThWsQYPlZ2xl7c1fuKZ20kI1CJv0E0XhVh0qGZJyCUHZhxiOfVt5r1VO4429R3KLBqvODzwJIjh3
cZFzQXYWfsoLd4FOJUdqKCY5D7olnkGtfmoDfeQfgRT9T70KOlEJ6Rnlm5+GzmX8J8cWllwhsN7O
Bj/gHfFnr0u2ONX1uMkGYtQy2k1OjOI7LGkp1p0CoLE4odRs+nwLUsHeuVMq4DWyR2eKzwT4iKx6
34wfWrr7ZXCRYLomvLJhq7h8OMJC/CAADRU98w0tdTxhlYn0bS8jzpMT51k/gak0IFpLjpvhpAqw
ymJRpkITuUVEvosmsEs2UR7WCJLrEf7sQyRFH3Lf3vKGW5s519DLLb7cTEjEKDkizImj2ZrWjdYT
L8ZPWvp0ThW36Z40bxLIEaYECsmbwzeruguizXtbPZ/KvuhPAJWoJWoSsGf+DeYNDFuOJsGpm5L7
rd/J0P8b1qDZzEhbB52+ru+UmrpM3yZveVMjuEIO6p/svhq80G6IjbRiIhBVNiChBVM1pMi4eSpA
KkABfDI2ZKUk5TseVDPiRjxMd04CQFV13W9NtzF1usn3+cCihKpysjNbNgi1FdtMeVjUuXwvTtjT
02h9E0il1Y/kTTK6RLSmmvCzpnt6M7b3lyWXmjEhLudYw89H3FsJvhuXY39+wKZuFsV8bVRK2Lzc
GcspUwOgvTv9Wx3zbhNIgOhZYE7hIMRGzaDbXli98xtPDx+D3dlg1D7Ve69DScGFmjSzVdrhKCNx
L3nyOJk0eT0o5yv0HQKZ8ihvfX/x9TXy/DGoG2+YcZCauSY0Inqh7hgezSLrrZoSNHGmL3lufGOi
b3/wxg51QL5jAZXX824L9UbRTyR7ZLyzzzXN0X0U/0R1WtXXEP0mBxj1ZWzw9k4EXw0tMtv8hafN
ewIIswd28u5LqQPxzgJ/jL/KPmaY0A5eTPSWTLZxxbvg6moPjtPXALsU8eJf5LlKRY93jXaJYBVC
C1SlLbpgVlHkuzglthjMHH/g5+7PeEH55UWG5vavX2EAKx2MFf7wHmIEbwVNspFdVZ19Gbf55Kay
EV4Bk+PXbSL9gGrWh521M5wxJLtMIkWWCfB9iRzqQr5h2SWFIWhCB0Ei2lCDsSl1fiSn14GqFW+T
PDKA9p9+LSf8TxsC/kXjTDBGUEaqPNLZ3UacT2hX88ILnP5uHEzXpvzLl7F61Qub0X9KWO2+R+zv
KMnPlXniNVo7BDtzU1qwwvB8d/o1SlJyJaZdARfA4nbWtfGLqLsmoXilk4T3GlOyqk4hgvN6Qi+J
EAvpLK2w7Z26BIJODyGCZwvMkiXJHn2p4mCbbzHGV2PIo0aJCtK8SK26p6d87ElBfBEEWQzo45y+
D9zluP16/hOmOo2xwrVB0+bKghPUMBciFTS+TDo/AJnDDAdX9nf+VXK3Q61RqCAFqhlH3RKBrpHq
/utCUUvyHVqf6Lb0i49/bZlMtGVWZhXcVjFxWaSx30mNPKIGHYAuPA8M5uzPv+Fn6Od/hynj3a2O
zJVw+fdugFid55GDstIY98XGit0KzYIFS0NK4wsqDHSkgFBApg3KyBAgFWlGNSse8NO0h/CavB6G
sCXvgamCN0QkNru3LMB6cmkIBC+BxpCLQDBiHm90GS9mYOcsiDa/Yckif0ib6c5vO4iooXuwr3Jj
e0LLgCA04H38pJyEaZac7pPAwoDYcxfj5VsDdFdotSNSYsKXX9odvrrlVV7Y9jMJINCgqNk3wY5n
Fqf7DqST6flQp9+CN9ZtxUnrk67qx/Df9SdlCbROCFHGNTX1ZXGnrKfvfCDiMBC6kVPIhdtCOSxY
XVdpEmX1MMyyXtPpxz1XS1uh6lgXfY/DdlyOzUi3TOXiOJegDuCYdTlrFkaQ7zq0rdc8j1d/uzbB
lVZ9KRVedc49EIGhuO+VU1bC/vDclJsUAUrVD9AAad6ULlwpTYu/z/F1OO2BPpVx+ILY8YCD7a3D
2uhNIzoNK7k6wGkb2Kww3gs9T4rYM4+exdzPK4hX8HOXMj8jc+oinpiS1EdT23Xvn//Kh6zfcZwe
RoVlbdk8OKd3S5LN6XSyR/DAP2ZK9FtLNJa3EN3nFJQyO6tJH0LPsw9WlUV02qjOkNsq3juR5rTW
ohELFBz0Zy7TeAKpNLEer3Wdm+XI+lkjgRx3QLCi8GNBoFUWTYkipj6Lyt8VVs5Y6YgY0/PJ5Q5t
9sEgRLirkGHtGAOex2/doZwZLb9ncOePfe44dPh20xJaYksKpMR771TkpGHRNX78ceNQKbMKyPMZ
P/0EWjI7wGZ1fwUSDFyF68s0/WmyS9/ZhV8plBK5qUeGeMUq03dzbgVYCb6RqgqYCTGvjdpTmUeT
8jajBzVDvnhRMKSB9bAiusmtWaFve97R/3IZnaoA7glhDw6FM65A2ZJYEoI6M06vgc5h79n71L6o
RW08t63KrFk1KqUtjSONNy+0SEdnOl35z00KK7Y9GXtk3Rd70gq72LtlAwGlV6N5OzWGOeuDC3ir
pbQGOPRhEYzIF6GPi35EKYsSMUnE+pIeMIA9JWNZCAj118I5YiWuhBnr8PF6kW8NLmBDWiWRB4BW
lzZ678/w2TrqB3XYXMl1kTTuSe3IUqkGrk09tXgEaAw3jikIo14riuiH69bb4y+YZWfq7gNM0ydy
bsZqkzh7IhLv7nOULRD0wHm8K6N0jVF7MSjPRcoGmz7WztMOswNEih/2wlcm5byymOSFChPw3NPC
+0mUWazHv8agxqSugjOKNMAIq2umH6CeYBBvU0MklZMHhJX6Kh3ZIiyjbVL4ExRy6cisspQY4kAs
RhJkpeG4ow7z9KdAPD1qxrn9iaoh2w5EfRYxjGdGqsr+TD3ZGHJPkJlLG27uSnAZkiK92osn0Es/
IBEozh5A6vfmJ1Hwgd8hsyJxWfHr1jNDsQe0lotilfnvQuf0KTcYTdRQc8bCv+y2181I8TW+Fio+
CxMYGJg3ySo+N953cGN89TzmKnxgiPXVnWWUiuV5hSc50sIHruvdBz5PDpcaorvXDKknyfCuy0tJ
elEcM0DHkPLXm9WSscvPS7Hhjx8Hbz3LfBS+G9s+5qVfPopYcwacOwy3fHGjCdoaTEQY9Uz4j87t
W1gtDhJgeL+JZ2z6mMxwbhPgPEPUkcPA69ifaflyd4EY6b2kCuQKQtV2FOb/ACEOe3VYXLWEoHsA
9f5YFPPqxuet0p7tfbRJSmyboMERsIHmecBj9TRNHCoZ09s+7st+juvT/LITjBXGzQfjHRod3rgb
f3mwR6C3pe/2jaZGqBkcIjfcZQvx0p7SSWchiTzlih0tFc3WVoyzKNQq4xoR4SQa2A7w3NoBtw6P
1+mV7df2sj3Fd3PeRIyMK8LXMgiXMCEKxX3CCsBokN5fUasq8IfxnnMJva0uo4T9uLwEF8URhs8X
hRWdqcZ+M7q44ZfyMZuHz2hXuWYC71WBE4GKNFea1o0hgIM6gqpRRdwmnOYMkKXm8/p6rlOX5Pof
3abz9wO/w8lw18fp5ZU1VG6uiDmj8Cd23jnOvMlB47ciqKICK4Pv6UAh4HF9Fr94fIIaZBZavXvW
POReQB/uwihPl/XJzWHN8FYn+kJVprV05P+8Oc19KLqSGPQK9lmcVw1LUc04aVoxM3Quc3YCkQ0H
RC92zbV3KDXXGPwjKSx9KfdMGlvFGOZEzT5+F0JY6fOMLi7Fuws9afVlHWxmTxsnRMoCxh8hfjmC
SyWmFwAMpgEbVes3KhR6GRxyAbGliWcnowP32n8cMBg/SEAAAwltqeB+Y8QibqAFT09wHyGwh68r
ZXsx+U5kIk05QMeatmp9jMRn1hJm+tiwciBPDiEnX89YWoNvSBczGuOAAAm8O7gfOc8JOIJZ2d/K
R8C6MuO6Mbo3zErW03kPxH/6XJLvYyEXZ6vttBMOL7ffjbJNdMvQDmWxa9QQl/OGpaA/iXp/roIN
dVawuEzNcsYTLDDezrhius8/E6d6pNF9XnXh8Lkibrj5Ski6fvtrcEd97Dxe7PR4Z5VgRNj0RBkZ
+S8CLzGxhCix3US8TBJmM9N6sYwaCkn8gxoNpfsWA5PPYNCF/LEZo4MYcdGbITSQ3iR3Kuz4eVIE
1wBbUI1g7FC512rKDZRqunmWaEXoqTtps+pjWtQ99VT2m89X3lqKYLVkxHD+nWFkTy6FpCwbH7N6
10j8dTrkERvAPZJKsk3D01wD7+altLbbAgvEMO8t/9D60NKUZTLiF6q3s+isl4cMUje93mNVKE/P
TxqR5VpHOFlNjSbOOVutcuCbQb+uPYDWnVdPass7+cmgEqXjN4CJ8mr9WNtsWb7UCluJx6hfj2+h
ugv6IOjlvdE1kIwHlJoSbAvNP5FUDY4gh3EdVDLSf6fmhZHOhPrZPXZ7zm6N4sv284LJcMR2bp7B
vTKZWm7GAbmYV42PLj0Afnpb7O2/F7xvn0UXxFQxdNMEVXdBSE16g4eSsmYZUulQ+gGV5BgH2OwD
AP9THIp4r3CAzP/XYM1rswJugImt9izQQKx3ANXPLiiXqkl24n5kWIZWugMpmy1SLXGlkiCHbsUI
Mb8yH+SlGU0CPgSaWjWykAQUUwayqtgDmMgOUWRuh4o58fc3fNQWVene+XqhP1xXRUgbeaUT+4Lr
rkOx8BYNLPFxcQmaX00Cs9buokl0oEG512I19Ra95f7uhYdFjbFgWWvGXKE/skT+MemyAK+rCdGV
StDpQGXVIGX6AHhTIsozpEiPHA+IKiotRnaF1gQ4WJmOKw4wIlowdyzXbqSv5kZR0eMAvKx/ZRHw
fp6MB3Gg7a42wekKyE4BRH0VnkiRJRwW+4XSRIgQrUJ87N3d7/OPoWwXflkvKd+L2D/bKNwXcwzW
YjR7ve38zmKZCIcvxtpxMU9IHnkrzAnrd060a1nDty5Bh1993qU/ErStp8cdM1DTqqlvwujAnda9
XFOOTc02e6OtaXjsvZ+MYz/m8M8U+8Y/ezJOPfs1vTb30kOY8D9sYuJJx61nopKcrFLRW2daQ1Nc
wn3ZbVb3lqlWgUX8AQIjw6JoIMt+W7w2etA1/ghAtqf5Q03/bvdv4PVA6q+20HIiPUthIDZ6Wwlz
MnDgWw6qNGCuPfL4Wt9uuMvHc2PkNMz30jYpEl2I1L2/7ghkl9FATI0tIa4RRKcHbfl/X46bWPtn
NkY8Bt5gSE4tyO6Xnt/lVZK6crGbudIq4oynfpv/W4AW8yaS+4LudYnuXIucXaH1w/Gnh6KMV3t7
wGh29rbYPlVucAt0JGbzKPQDBKoWqn7f+9vth2bYlVVMjpJ55LEJWg9DTxGnORJDedeGixqbjuu9
qz3kvMtGme5S6mzolP8Xx2xK8+pERAg7t75KmdM60v6Hbxtnu/F3sfjqpxg8GCb2Pd94WYaH1Cl8
IAem7WUcJ7hSIXaYiyTSTSsPubx6weBfK2npgMt1di/5nwC05nLaqTrUYSCGunFUcyaIivgoQihs
j3arA+xWHuvVMwrgJV1kkljQTet/QZtRGJ2AMgMPxy2dIw2kyW2M2LeJlFUq6LOuryTmfvaciKOJ
a1grk8Ckc4zqIGvTlflBWjRn64Pb+oSjdXpXqEUJS9YlMacJ3AXbD4ofxGSXp+CAVbKf2hxJo8Us
jDpdeOYcQ8g3D86nLnJRBQsTZEFNOo2o66Yub6GjM4+jgQQ4B4AO5IB5vGLqq0Nl53AFiNbVTxwn
BIAcCKtwTPyTVcH9hwl0Zhyd8SIzd/iY8ylcyN4p/+AWUDezd/ProwVpoP7IEKtKn36ueBcRznVT
3KYwiFjhikg5A/AKEzaHfOoh3X/MOzVoywksw9O0BnUV4NmMdVj7JkjP1lDO8YrMeixIukH9RIJ4
OkPZ+0nZZeiYfNC9KewwOq20IykQ9uRZLZK/Cq3jKus4ehudKFcjWtWtPOXZPesWtZpSkTNWKvbN
KJ/KofqOxvT7j1bO7y4PKZn3O92E7uFlk8FxsofLjtBvM3ojDfJVW0hNZPO7s+192YdtLZatxnQh
MughW+1Kz7zuLV74mv6iFXZBvhwEA3t4YyV7PZIcIZ9k4wxCJFkMPXolxm+IdDmXZKRLxhZ26sVf
uSjuCJZjMTNerCHKIQ1ye0vLydpmq9tk2d+bjdq04x6E1CAZByrohwoZFEq0o0qZVNhAsT74S3FM
Dp0jXn4VX1N58eqgOGd5xNX22IB14xE6n7tiHZ0bWmOZX/48hFuxkpowjQT8eG5S8zOGwjvpkixF
rfOIcqbszzAV5TzWLnGt7Fxvy7T4bs44cXn9V0NbogbQadfwhDoJNnUZfhwaWYYRF3FmF1eKV8FT
0wZ/w5XwwpHdujKlVBsKtxO7vWFOzTMHxBK/c4Mlh7//oMfaENpaQ4syr/cblsrulQtQZSqS3udl
HuhqFv/13pvTtg7aeJfxuXGxldmIFasS2sLKfyq6aaHHEXkG4wWNwxpX/3jbQG66CDXidCtdOIsG
Uf3S4mkXH8fu/jMqo/bwB/trJ+VkLNnoW2+4LarAjAjpf0a4AJ1ZeBQ2PfAueYpx2mqXHQwR+bv5
Gz1BcZjooR2dawuxTqr77FQjwJhqKTUVDfrZVAvRqa12mYT0crarLuUl/Rv9x/IeCC4dAOfYeulN
o+sB8KHUnjPzxOQMvRiqRNc9oG25Ix8tzoWQ2kqX5yVy3NfhiVIssjbdovTID0DjWNUeh/nPoa6F
sA7PHqb9CtEXDjTFHNvyZEFU1tJHuHxSElvS5UeAshrY4EvdjQskb5pWdx1xw6KiYy9Tj5e/ui9m
hfcyDT+i5KW9KUbI4p9k/tg6Ej4w5eZ/ZrjAe6AtN+9fCTWCraWtwXl4xRv/aWAlEpIjgsT9Zkzl
yb+W1ekIRhSxrLAd8BoUHOS3uuBb4RlnOAJGprDTVti0W6P44OcjD9H5gqi+uLKaQ7rg3eGNzdtj
eaos3vwOAjZSPPFJz38KCWSM7kZeng5uCwXEUK1TLempjxqvF3LC4eN/Mr+T142/iw3oG6dmZ60m
2hSiKuUbn0NjYHk/M9Us8saMO3tdoN+Z31O1Y7x23lj6s9464dfxW8WGxSqWa7I/Anp9caOZRHB/
m8amKr0jUiVWDxB+CUgBZ/4kv4uOBwYzakWdSZmAr6Db1xEhPqJNixz6y52CJrRjDYRXlMwDjg0t
LzeXzyctfeRUChGJJrTxN0CgIAkJYrQUDybSSYMqQfBHzLqOngoFy1cZ3K5JOyEcrZkBswPdx/Dt
jTYEJWIMepAk0C4rmp8ZBev2G1AgfUwHFFx0N0cN6GA+zmhuMeCJnYXGATKlvKjW62gARNnOe+BI
8K68HsDzTpFqf0Z+pZzuN7xAdWdVgN7WiAhnQGIT5xxhGycnpeg1pbc9cL3P9Az1kabC/SmF3sE0
zMibjvKiwnZJdk1jkpUSuPzo/rdrj4E08Hf8xUNucTgT66eJeoHs6NRlbXM59SvbISX+RMDFNO2i
cHAh2CwVhNKVqC7yFbcA4Ta8bpIOYy8Wb38YfmjD+zYOH8+/BOKdA+38y7Vq5jRfVSn88RYbiVtj
lRM2Al2BAOxUj9N53JTReMpjsMlaV0bHjkzk1yScdA0+jZRBbaigtT3pMKeRMIy1A6okJVSf/p0u
T388qIwj001q2NWb8FO8m7WFEtSestFdJnqms8HKBcVGZez2/RHhU/W51FA7GpHmQ4ZgrMmIiSHO
zszMKjawBnnvAZTcDoLli1kXd1Ia55GnboKs8D4m4iFrmT+baRvuNdt4ijVxfuXL8ZZNJUf+tYOw
o2vU2tnD68uIDURERkQzlJ6bbfcJEX9M+9Z31jrpxY5ug2xrEdI2fgO3wsxBmZgpJ88Jl/Khi+9n
yXyJir+fG+EggSq+/sMFsNMbulFytpQUPILQT58Auy97JZALCiUFGsE683meV74IDIZwfxGVymFz
4OVe2SJPGY+vc4xjRk4TvwsqpNsIYGJzX5ZVdACYmd7gSNlI5NZNmppYJcV/AQii1guGPMY0NzNy
u9U8TytNj0ZsKBgyscFoVQGpbR4Q9sY1+22j6dRBm3cIh/xkC4aAlzpEf1bu8I17MV1EbSSkt3p5
/lm1Csw1KwOiRHRsqNOpYdMm4arCc94wVbA/q0ylTPXpKqr++pZo4M0ziyRb+Cr9hLQC+4p81j7c
OdD7py4NICa32XiXF4o6oR+xMw7TwPNLB9UL3EQ8ADqr2O4ptS5rG96HllZJYp4LsNyL9KPdU7F5
Lx0ynmtZUwj2h7lE03pRX734gozkoNYeXCcGkIszIn+PwEpPvrzicRVRuJj3vtoHXVHZTYg/OH3M
74fvSt+GxRhpx4Md7MwHEv0UV8OVXzI6HIkPLge447VngSOcSuOxxPqPpUw2YiEZTl92Bpvyy8kD
2J3YIXaMFQS1vpd50QTYSiWEePRij9FQR2evXl08iB0l8zSdOlt35Q2yn+aTuX6boKV0tRap+kM/
N7qUYdV2w0CCDME+G+tw/lE6gxvSpUPVy4jsoqbdOyEJ3gw4YXOWjvmJ2xS44MV3xc2swTff8UyV
P1LI6fxj79ek9GN4oUdtatHg3sXU9kTXn+DfFSkFm99cZLTglpKutGd27Itcb5OnNvldGh+/uF42
h9rmMcsv4a3HujQOacy9/MU8+rYRb75TseXY9PS8gIlpCHiZpAOAo/1nJ2lnjYHErr0Xn2leYkqC
reU8NipNwRHUuhAiN9RnPayoi2RQ8lZ6MPmgLEBr4+XfoLznNWrE58Zt3bGLiBHlvhK88Rx2Cnrp
I8rcF+WTUKuyHvCfLphxRLXvr/3U8cnQdI1iuR9drGTglEf2ub1Q/yTrd2vAVtn5DG2Z91YSS8UF
TgD3ixrGTScdXNBcwT4u6RHPqFGOg3gCxQFEoRcFMTJMJBtkJtT0Ve29aA3W7WE3T+nLZHRBe3re
UwNSIVC5W6pazdt3l1jqWafUk40vAK/14/sO6Ul6LJFnLZS+7NTGqKeWwnToW/dreCy3gx2DN7dn
Eniqpf1xWRpQT8FcFhJ2ZPTgVN2sSGaRF+IkbE4P0nze5aoEHxRZ9LnFL8iSCwsyh/CKX2JVvs0e
N/fbtjxsPU3Q3pqCit99Mx2FQtVcOAHN76JiGDNjC4AnFPslm/8mOcwttl7gEx0WU9zUWJdi3xa7
SaD1kEm2XDBXzpn409hl1Z8Pf2v4YoEc0xvfPQOeNN4Nv5KwXiB1JbnfjLYIN10+hDzZoaGkzo8c
fX1wlEjV31bPzUA//sgMzEDj6kv8Z3UIxvN1ntRJGItYAZXzsTJGEsXYuFccoCK02mrNoyg/a5si
pCffQ98wkIilMBAczVIOwjRJB2M8TtprOxn6ZwGCxxREZAnW0RtjzWG8tp9dvpS1gpWui3Oyrb96
RbAJozAfdisVNlN31M3eh/frFBliJPL2wDBZnGKu31Y5WWkitkt/0fXVEIYZ/lECGjs6V7llZDLG
Li5+fYZFUiZm/Y9zpGMhIAhRslNTImxMZB9c+qf1MTLDJNM5kQHtbuBWjZavF0IVFHAb4VWLUXvx
/BEjV+2zpD0K9lzyih3zPyMdyyS4l3lbp/D96ujX70fIn72+fQkeXrcu4wbnwivJdIHXxMkoASS4
oFgh8T5Vz/5s4RD89QZSS1TJDT93ERL+dpM+0s05Cg+RWexws0mgZLsBvoxnLcZqqxcTsi/+LgrW
7paSgLhbnQ7qwCp8zwpZ6TZv797tZhndjMqs4ouHpINM0171nfdmPnqWUrUFfyGv/N95+EBfHzzX
GaNv00NdmsspHFe+loc6ptAlSDCe+Usy6NJoutCEvgPHQWbeNDRPOCQIsKMmKi6eIuJfpPBTVJww
aVXhD4G9jPQqbDy06DZIwHlO2kZk00uiYtS35IA5HH0w8JHFoC7OfsQS+DmQOHA9FgBdGv6mDSw4
bOE9WjLc2b2Ht9rX+javkKYGaMmBPyYR6CmO9bXsDA9WbXSBoBwdo4PxuX+eAVRx0l+SSmAlxT1c
okMNi3aEAj4NXTuRgiWtW81fW6QyDIU3R4a5/8mXDbnkPlMrHkf1QTFH9RIFmMhcrIEFLNWOHpsH
3GBGnzWerAcIcbA57zKM3xGKk5NBYQel13vpPg7z5+Z7hJigEB5m3T0/I9NI6M6zRFO6LtmJ/z7F
/MXnSpGJvvnLavkt4kcYQvc2xncz/RiWnKvKmaX4VDzZkx/3yjrGM+irR+3HSYBdt+79T0fNR+zx
IDCd7qk+tSNfpejJoposAq5Ag74zTiOntWYK/dpcQQgRpWycLyMInwXTaQUg1BILHf8Ao0T1pq4r
Fsj3Ngaj0RWtMdL7L/PBoRJVyAuXvSH/oQj/Q+xfFnY6k4/Thizzz7mx1z73gQjO9c4rcS5WgKZP
3z3Y33KP6ofgaFmxnDCPCwdBFIo0Neh5sgszyIRW4Uqqvc/y67UgZz6n3eW5b5d0tLY2/Jq0arYW
/uI7oDvmhkmeoCiJ2RxibBW8iuQ6kfMXqpjGlt7NgZonzSlxpee8Xyjq+G2fBUnYLusWCrFG9wwR
6sMdlaea80Xg9oZ0A3K0Y3CDFfQP0b+CE8YC45wwUdJ7Gm59suuhZTzjWfv02mJLkvJKEF7zZBmP
XqpNXnH3XBHUbUziTBt7IjyjabdbMm/i/HqujjyMqQG47YzHconp0P/KeBlqwSub4dHK/3ehia5l
5kdh7HfzG1jF4LGcptMFfQx7ErPXT+th6meINgwuaKGWW9cErORYf1nVb21Q7okZmg/aiVnk17lE
FD1LTrbXH6uYeAHRoJ8O7RNT5bSRJH4cZNNjkfaaPYUYSR2P3Uc9bHyPU97b1CAzdgLh409jPJsu
VPovERzggXgYeY28N8b5GO9jlJyGegcd6apEp6l9iztzZVghznxFiL4U85YtYXvyhCdSrL+jLkfX
4NUbcd0Ed813s0MVAITP3fTNb7DoxtnUzHUlBegMjo7lw0yPfoOVxtScaJVcJgdSWD5mn0IV85FU
ALGEv7aiiULtlPFjHELpVjaNL4xpzH2BLmGi9oI11Aer8gEMCVQTqwHjD2mbT41GsyN5Y/INVg6Z
PYxN6vE5NKxsh+gswfvbkNh1ewdWK+UiZ213ylSNNGdxS0CwTYDw8sjqTsp7Oxhu/895WyOUvA/h
eXzLkIMElElxmIFm3cZA/x5vLW4uEK4qdZLHAH+9HXN7t2bsmFQR0lnBTWOhdudVW/RamvstRytU
vQuXOTIG9vawrhtVuIIF+HU/FgwC56dxRVcyECI2ZhTNLEYDzYGCg87G9+h1Nmf6tbKAdT5duweM
QKRbE1UF2phKapONc8xsIMcEcH+5XdGayHZ2kvHU5S6qkE3o63TxXyATeqe/eZjTZiLUgh0r3tm2
+37lsXuB8Y1v7OLW7h3CgvGSDRMpuBRQikHuuKOqLx1eASRkazcpfbgGUQ9kR1hLPLkwCxxR7jFz
IYOdwcpfVd37qpADranivFSbfQcUTntgZoBC6Xdrtq7EHry9MamqRp6/GPtXy4gGD8r3aYVxkSfy
/2PL9SEmxM3QnkZOgU8+RP3qBaBjVIOSSCzhFZ44XQUjq5oFzjvVbRKMUx/bwG2Fn9JtjQgk/LTF
fb5QzvDaQuT6TYQJE5utZjFAWOJeRL5MpgTvQJCdFeBMzSkMkB7/NKE3ttMxH7pAxDn8mudKjVtF
NT1ElqRNyKvBcwR71NOEOZWwnhVWIyMOEcVth6/lk6yajAWq0SJDvBgU7GcX8hGOUIO2sb1YXo4l
TS0WsTFuiWhEc04+BDkceEoCfpulRvBc93RSjtUkfwuhR9oWqTQmVJU4hhADISLkGKSIohPrgcrx
LBRM2CLlRmR1zg/xfMtHgSboeu8/yfchOOs8nojLZ5V/7yVJ9vP9iXeYL8T82SqoCfYxDG+msS/P
TjfE85SvXxCSEMO9mi4u5/io/ESlIYXe1LkXVENU0wkjShoE+p5i1MGB/B1GdTn3Gey5IQSMilr9
yfQyUYI+oB8j9tUeEQSsuN1WRBXN2P/YycXZRPOBHLmRehungF5DA74pcWXD/DfOcHUlRHsEwcMN
QKze3NfELRDhzAZ4VlE9+BBtNGkm1BijI0x8NKGtpuvpW5/ZP0wrGJljRjNokE6qB41BMigX10zP
ZB107Viqe/UIF9UJeXIkOMFQv1EPFAcne0C9cL0kuBctOsYKJoV+uqFIFXJYREhWw4WtRrX1FIBo
j/Snhp03jIXD1fKCvBi9nphXlKFcoIdI2fnc9qg50Hw6Ob3mLBo8ugni+CoL9rdlfzpNHQIXrBF+
4C3lVZCGN4FF9amfl+tgyICVETIW6IZdmOjb3ERK3pY+VcZ34836kZ91Dvc8vrwp5IUujuvwl4Tq
XotTRX9nAT3bCHIlm2Lyh1Lp5qijxij7VC3AaPrY44y/j0zqXvzmh8/kjSqRKBPibgDcQl7wcASu
mnDSA8Iv8WjEsnUE8m07Ee1ZkEMRKk/+iXdsvfvZY61sy4xryCQDgeQhe23jn3gEfwlc0zXYXLUH
VTIXVCPvqzuuAtU9DeZZdh17Fs9CiudlbGJikt88sz00LChrncg/qN6/btDl4Le3DmEA6ZudosLQ
olZMqTJTfuv9Qkk0/uAr3+Kxi5s0m7d2SCl4Ou7ifGMTfBblb2vqU21XsKWEJUpmMneJE1hV+wds
d1Ci1II/M7+IDo1xa8EGi7QnvUoK2kqip1pjpZDi9f8GNdZClBvy7SdIGaVcgsThvh7tHmlxLOwE
yJj1sL7Yl7DhPiaMPU0jQSyc0k2GPHdDc4cckktzLDvt+Z57L+3ztVwp1gzUyJRTqykCxFgDb47G
gF01t1tmUW48r4z1u1upMLrCAFkLKHCCkeqMWnKMd47oBpEhUJNzDuJ5rGRWLns3E6in6pvMAQ1K
/N7sIuPFSLMxWXZQU3AA1ZVyM+60NfTmUhvLnkgrfDe62UlWHcj5r3fvda12gqyhyQH4kFte7YRd
hX+bGUUtc+h5igm+fgrjk74p98ZoOr6bggxcX0wFn5iZyDoq7uhKUrKSTmC8O/N3Cd/9CoD3DzZQ
xxaV39QgnqElmah269fxnsin3pazMyAY64TwF1sILPJVxZ6qNvyx19OvqqVdkF3PtOkY8XcCXk0o
SSQidVX5kWIE2fTHFlolM0j+8Ig0G5piVuLbg6RI1oKxYP2OO2UDVWyC4uRRmIA7kisdCsS3aeys
KHgw3PNn8S/Bc8zc00gcsgRdrVrjXUGmKgsm5HZv8w8aVHuA787AhjrTlk93kUzC5WQfo7BVCoHL
xP7yD/c0EcKM3cdDo9oyFJYx78t016d5o8x1vnJHIOtWc2GOtoq76dDe9obuCoL69dXlQQScnRBE
996VV1tKUDRlFpbz6SscVJ/toRPbjLM60hi3H2qmpQKmxy4mZka5bLyX1woOrnYGR7PzQ4dBdvbH
u+ANRD2OWERVtdviCbGkME+zFktTfFOSP69zcy56DpviHwHkqjqtunLN8Xsl72Gg1Ioc+p85wABI
yv66QrIqcYhgaWScM92TmFA5KtiYEIUNSJk634CK9Rnzi/oZ0rCq/VfFgCJu2nO03Zv89NX1DW0k
PC0rvMJzf1K5EXT7O4vki1rLPd98DPvOvAeQ8ZYn8V6fqO8fvosgvkUTMCmJXY4gVKys3EZlqFCw
IB/Wa5Mgd4zxyC2BSVi7e2JwHc7xztpvMQmedPMAj9Oqt0/6aIIMif3FV+8MItqa/WLo6rsaNG0i
J1ap0m98QsjzQEXFyhskhtHffKII444hz0cx4GkfzqlkzeuJX0HYlsMc4UeTkcSfOrM/WQKjpOW6
5bX7ZNRX3gOdBaUHPPV9knVQMSzHuGkfKANA3hrAPSycgw4nCFXtbJlWE8K4yZtyqJnipfXQx8f2
9MvfLSBbRR8mEyR9y+wqwuQHBymq5J7W9DtT/93xtlLbO+HF/AUH5RxFXfnKfqlWydzP5k8u45lj
y435SBjZXVYYDJUC/04UeKDivz1EAG8nK3vGsCZfc3aS9StdzINdWuUKU8/1BpYZvNNoRtjsQXW6
4E5S5DXmWhl9CnCCdnd37ZSMC0KHDJCwAAPaG5UwuYneY19nRQwJQDpePGcrvxwpmE2M0L3ys+t/
5SEajm80b2HFKiVaxJzl0W4n6GqKqTv1rQWe1ghZcxW60Yzd6hc7MzRdtAk0eUHQH4sV6Ven9gQb
cLj6mjtofCh5urD63U0tkC5xmXQtB03jPhn9iIHwwBdUwkFn3WlH2F13J44AStsc9a7plY73b0x7
ORDWNU+EflPZhvQqSPt6NkmOvCCT24ljD9MSToWz25DSiZfm0xc5JfxwX4E9Lu8p48YvGohRPJGD
CRLIK8ZtAsGy0LROJeBsOsDfySC9dFnubs/wH/EQ/zH7E84MpXr0UONJWIpuTOUpleCxApp7b5Bj
c7uccJ6rlNmT/mJADypWa21vjrtblRamxW9svfb5+imFP8BV0VKK3QHt5SoobeY9Vls0PM5wrt7q
S6o9oSTgKBBRaKa4bcoXKbxzrgsn+/pH6YkeQN0IShIS5rmuFVC7eXMk2b5GqBjzhDrpocg4xD1X
mqgPvJaXVqTb2J2GAceGqhHfFOoSLdtn2E2Rn9GW3oocTPdiCVGLeIegMKAAXmFGk7StS/wl8NsQ
zSxCzEbr5fjdTrqfeMnirCJHWsUeIvnwsM0yNduGc/airKi5GqizCXGau7A6qhuSJNQas7UMLZsm
cbqb2uBONxh73CR6pGCkKhLL2l4d0+Wx1S17vvInjTpcCo9uuWMS5RmByxTB9enLqTP+vxhFijPV
mxaQDoYDCZbiDZl8JK7NhFH1/4U+2JJNXMeB8bOg1c2cojR+MqGne86xF3x7LFdGuJOvb0pR/Goe
vDDFBx5mcfIQa9srF68Fn7vBwduY1IIOCjNuVBwtd0X79qYDCru3DkgsVPrzLw5qeqSY2NMaczRv
NLxW/SJYZUj6PKg+TGT8B33g9C2u6gERvP+qqM+nedKzq0K30q9j+w7THFcWHhTLKiHLvwGpSz3k
/dGDQPsx9itbOieG8EWteR9sXEKbKo2hIIFhfzGyIu2/3McvR7eZeW79HtK9UFPzrkm/Asu6xoyj
kYJK347wxw9rYH4T+gtD5B3g1VgRxDkD6zj7ZTN6Y0y0iL1qZksVMQgIVoWg0kF4y7yoDwoOyd4V
uzq8OUv2cVM0eIBsHhi42WLT11jbzuwlMfE6jDMViflJ9bty3zygYZ+WmW4pl3BaqxeTwmdpg1iH
5BjktrqWVi8BvvVZHCNB198hPbFVPYRkZMGlFQni4sywAcSn3MOmczPfHyH83rfA++YfowYU2Nmf
kEt9vWHTVQQktTTwBiq9zWVWaBuuv2WmUPmCbHJhre2zED+6RpXYE07wosZJ4Kz/vG4jQWn+szvx
TyLGolP0zortl1chzS2dssPtdh2e+Pr6crElJ7WyANHa6uHFjjqch3iaXO4XQEgqOh6JY3AleX2E
RCK4/ShdlgeQsLQIy6wQY7rH7NZJzNjwE+hJVvfdOev4CC8urZ7rPS22+tyVFD+CvOV2Tv4/NbB7
bSkovS/FTrOI/GX6jNhjjGOi/11f8kMHkfS985neQpMr7ZTc7PrrEeLSKiyRS0/LuTEpN65yUTy3
2Bk/gXndLQp2yhIZHoeiDM4NP76s7ZFcJdNK8R4W2Bh376HzEurD1jG9QM8bqDFfrQIVEw/i0tIC
Qbef19OmD7W5/9kSyFWF7Hyy7E/Lo1+Q1OdXLjgeHO4s1S8rVkPU5mhmxF4oDoRd6ihesf+4aVKO
c7yfVdAbf1+FuQVk6j/1qFKSU3caedykkelwbPynmYmg2fdYv8j6xZ9H+idn1FHEM8scD7sgbwgy
VrVKKbIYfpHWw8Te4NAW9+I9mB/5sUHaj4Y6HRkPeQmw2T5W4ALppqChoo09NGIudXbANuhE1j5e
iecbIv8RBzrip4pGwVyImd5UH4ik7TMzlHkrOOLjN0JWsotbzlYEB1mGKsyg7/r7+/eFqRCjbxUH
E4lohudR9lbaVHFoazAvuFCt4Mb0ORr/LiGAowjoTBz/Cs/2RFazSP/sBITnWJR64uOe/WP7ZG1Q
0lLKWhOGQXoNi3QXM1pAJQUG4jIC+JBi/BAWxg6zasWF73TI+HrPw+MLgMkZ4ZNK/gtgTN8EPDpy
qzFNfGvsdZiLqiveWDMr20FqaCsgKF7oOnKjSnMHaNRWf03lh7BM6cvOZrRInJTS8wkKbK66nQwU
q+Q4f7s2F45U6clY1lULAEC4bwTbQ56GkeqLIyDqhOX3BnjFpokbdt7d9uvDO4ilZ0j3JN4TGVNw
DJi9Gp1d+2FPlRmdG12c4R8Nc3hxHm5TxXHQ63+Yy+2e2VNhgbiVf2y4j8IOY4fle8XIczaI8/XG
0IMU029BpeQpEHJM7r0MDvOJBWCR/ac4AlynauaBikGHHtmZ8VjhCLBDidjUjHUzkYKTH83R1eVW
QO6YboxRWAYAJuyvyj5qfq6TaxNJftU//Xk/5clM99fvx/Yrvy8+ozAwFZkd1sYM5eivZNSkuhqw
WRXQiz+l5t5S//RMkCDwHZvfsjFlvN6vxLsH17UJr6daeFdlWkQ94nuh6bOn1hWVN0WUWHpsxc+a
uM8XhL4BG/Bfvy3FIUtfzHP4RaUjaIF88G6J2Y9XkETIlU9Vrgs/o99PdO9tUbb9fc5NPE1YqrWH
gm+oNftO8JCUqlOMGYBcQpRhPsTno9tc/H0CeUDmFq0En8jtfxvEPnfYddmD0yKnBMBN26Q4TNIA
mnF0VN0huCt6WwD1CjPYbf1nfZ3OHBa8fXXFQCrAmYOWPtCyQfqH64Azb8pWi1FWqCgvY/8CMt7m
oNV0Ydr3ZCG0Sx4N2NJ463EVlR/b3XO0oqsIAuNsPzfd+tDXLGmYPojxO3wkLgjWUri2jDISKECj
JCG3OdoD72u2mYMRDHw68IjE83bBdcYBU2mnvcsJWDlA8+m52/9tiPJbbbPQjaQOBZXcazi7+Mec
AGjkE0qXanzyYe0ZT98PNalHsETrnBjuD6YxmfFcPJGWY4whfyAOKCVTmkpr8cdfGfl5l8m63kB8
RKLidUgmeqRQPa8JFnuNjK6CInAXgDdAyeQwzmg8lnTVmzHXZQOHu+umWj3Afr3/V4vR7J5NZrRJ
ItfrKclHYtaMpgOm+HFl0TqqJOdWDW54DPogBszhMw55FHKJMgb6mGJzJyP3Aq6gXe4OpwVT2a2G
YE1B0/BWgmraeg8335tl2wZTGOwVJCdGdL8mww6ocFn/Ybkb92GBIQNGNi4PGZfYMrvW9KCedVkS
98mQqo/uj3sRZ6BGKmcxtpNES+wAwpDju0gSMAKIi2JYJEzVpNcVDuG85X4gRyw8eM0i2uV9CthZ
VeN2cgvjkMNSFmrgn2duscbx4wwAOFAskL/QDXUaKJSgQL2/nvdCVyZZODvY5SE7BMgethg6k5c8
jIYWOqvNlrylDfHTN88yVVJKWVEwqY2KTLXOQ6WTXlM6yM+uVpVRsO+cY9vED9nqoEW51quB6tX7
tZRryuiZH8wnslnfFMu10uL7WnvCpiH1grq98q9IlYQbIiM/6YAn+EduaJyM1/6zT94QY0i7XbB3
ZxuT1Vk/G8zMjygVz3kRRSEf2RYhuNbYnYiHS/ypBYNwVm9sjZLGSZgLCbZMitANEv4WaTJj43I/
UwUoxy3VlC++3mL9+LzhITeC3D+UwA5Js+Prlj66p1O8vSRbXvazS2Bx3NmELhh1/+jDN6OzWEuu
Bs/eGnM+WIE77Yt2+xqglKstafrdZtG5GSI1qyF828jCDtcF27M9KoG+Eax0z7FnHHXD9dNOCyMo
ZL3FiyYlexL1X7wwq9vHgZRt7znPUmxKjqphed1G2wl+PwiUoWB0VkFdD9n14OAE2FNXYdvYhv5j
qro0rw7lNr8ZUVeSo9lyvF5J5/dr24tR+G1cNj9fYuOKP/aFD0+ln6rFXyunS5YxJtbMFXyJbA3B
c+LbejDA60DYC9JSRaG/TlZzFodKSfAtE77V2fs8ozQg5kmvvnqhVE0S87doYyRcof82MLvdNpwN
rIHytbD0cBqQppm/pXXOiv6L1DUm3KxFGXCFxUcOIkcGqTHXv3P5lBRlcrAjRDxS83sNXn6P46OD
bVxv5tSieKLIRit4hSIsGms4+UUh7Vhx51xFWGF5zAWu1YxfhMBr67vjw73kk/g5Zwtf22F+/s7x
4WUzG0ob/FTi/oNeRBz/xpDXmQloD+n9ABFeSoc6HNf7WBnleff0PzGLvqXJ2CSH0LR8jRB/UNKZ
HU/vf9aZ3/cyCvLa3eySi2zh3dE76Y0hNSgSSzaNxNyX14q7++C0x13Q/ZFGIoGU0e7lWuZ8P/Ot
j/HfvKuN+t1LC9u3egiqJTZVPo3up9ykar1IYRRWFk7fZmAI+QPh8QtqoN1vrsT2FhuZ2n8dquqj
pdOrSMJ4IX2xLS8PRj88T0SC3CdJ/hgR4kMMnwhMCnEAJ9n8J95xpvOPNho+T/0ZPHneo7y1mtgg
9HoQTRaJVGUGXN4fwIgICQp0JZLU9e5KLy4t1ScIPrVGTcM++ml6Ub7ZTRGlb9TkgD+cOhHAN2rU
uFnJEtI5Vyp0bBW3tmaWRRqYj2e/khKc19tToKK53SPBmGC1DjnXDwl/HRpNXCb0doa10K6EG49e
tI4kBF6hkSkEao8hpf1+wj5KhXpLbaPoVMCPtg9RkeIDSl8f4OVTwq/Lf1necN3/fyfdcGOhDkVQ
IaS9EuV+zbytfBpdo0QxCESamMYnVxHLlEQO3iYTlw+79jQW6K8i3nJqQdIto9gyaHToZrWZRuT3
Rr5SQnI0PlU4ZJFAJg2sQG2NaP1PEbJ6mu+59ur3qCRF47ny576owxOLI7uMprvO5y8rVCn7rq6+
lTuQxNxR5FEeCovJ11l2bEa4gAL5EJTxWSe/wcTPxRVxHamomJZ8Jd83IR0+7Lwf03yDpEjgSXbH
TTXDIB5v4iqk7oDt1byEJAL2TvQ7/hStImv+1Cu5XpMCjLwf7k93qdllpLg2uLe4LIM+FhiuVAol
dQA8oJPupH7GE+00dzhwTU3/7eEiQ8uX16RUhSauqjuwrYvHy8jNAkDrl9XI4M1W6BlPpmKiNaM7
G8FIBvMeFARXM+eZRjHfWsBeYDrBfGPUcsZN2Pp+VfriMe1BGfAefohjel94PbczH7ad1wk2myLH
1HZAU/3KqxlDL8x2vufL6GViVK//Ye+NI7uGJrAzZQyiwup/Z/TzC1TZSQubBBuqUjNn9st6qEiF
p/JZoAeQ/2YfgERCmbyKO5Cfgyv0C3dgSFsHVnR+gMxrVe4q0ZJ5lt5cp+1dv2adZY9Jx9FqHvCb
ZxMXHW6omXcxoVNTB0mDc3Vh0kW1IY3xlj5q6KimWgVf1AcnJ4svL9v5+7oF1RQg03RTfN/UWFDO
554Q50rGV7TRj0t679lgqiobaYAKc7dDr9yI/c06z18Cpk3U8T2zVpgIQn0l8zG+GI34pBAfdm1O
rRIwVmEV0b87rPleeIuJYiQk9Qgj9CJk4UrajZLaCDzmKJN+8AqL3BSkKT/w/BnN9q+hNw2SRydI
PK61MFk3SoXqmOZbfS5EPsmuy4/nNAFNwUSEppjpXays6Dkaec/4n5y27VzULpshcTin0Sx4LMkt
Bh4YxjGCi+g2DjOryL048aaMAmmMFITfNn2Lu76gzq64tnOGJW/VZSTQWKcxMTJONxYSI/PUw5Ke
V4LKTiq1fsKNFcWi+9gLzt0qBl1c4OgKhYkSiQK67yoKshRrtZ5S1qOVBT7jx/9Z4NRGgY0m7msj
kWwMZEL1YtvtWbGKCGVIn+NBa8X0cenEMVOtWP0sI59Gnz9KdHIlBCnxM+OjsxeC9NRm76z8VrOD
7IdxU/a7CPvSWCAbeUB9fJ9VvuMnVUITNmbURTLGJy9TltkXnxVlIsgtXWxi4UO0QZVhsOcY3X1U
XiXRn2EISqAq4RU2jFyljO47XRP5kHPPo/sKSgfyvS5Dskv8wjpq4CjB9G5mpLJiYKvqCmJKM08/
uCtcDAEF9762MJmhSnQ/tGVgl8aIySYQgYnVqboMtTuj03FdUT4LCvJN8CZHn4rTPv37x0h4bAsS
tD5idEY7mst1tYJsxqbR5nzGy7l//c8RcqV6v9+gRwwKxE+1dq5XniP2MeH4ayNsRa+kuGKNRUYI
DkE4ZEqRVRA8z1WyjPJKPcdcBnDZZoGGYb3S6eVpNBBtKXQ6kHV55xXjVsPPGhCMXhZ/dRcY/+ew
4dh2nZymLvMuMMGS9VPc5KtY+uWJ4SE+VNGTrehhZehuGDmmOGyxBTfAGR0AkDtxK2JWpcZKRmA4
ZcN3e+e9MCuylUA8+qAsISXsskMLj5CF8nusptGjYv3/lpuMo3cpB/gdZL1U2OsTBNIVCfG5+r5V
w3wd1eqWDZEq9bs36xL4Q+pFnBj6+3+mLjLxOyDHrvUx5mJ4d8uSzDMzY+lMTk+abIeY3YAZp53O
gfYuIEhAGZWSJCUKpGG8nvirkkrS5BZVZQb7Olev0+TDfbdaUiUnSXY7/vtKnVj/kcxsMSJxFnO3
SmAYqLsX/5X+nFXJxxiMCu9QioI3QCRWohec/gYISMdmttMN0VfGvv/6OHvwDcJ4lzT2zLSsSCTO
0d/pO6KuL9d6UguA96Bpkwkma6qg+zbHlnHsSDWmitGBueoux962EC3USnwXtOQbA+T0KtT17DxW
S+082X0as5x+AA3r6xQXXVaqKljl6jXaFHCGONiy8YG/oV4cYbIOyCyThRC40hPm+lEzY35chQH/
vebIOM2zbg8gdCa3PzIjp/yQLXLY8UIa08BmyeEh/xznsKlDOqaKtbC5Q8A0IuUcC5KBmYgN9Gd7
xSoafa3JM8pG6ZbWHXH23z19DLoy82s9NHbYvDa09isw87FDnw+ZjJz/G4qvrEBkqupeIa3sQuxO
utXFXZVJDmDOMCfdx4a6tfiZI4HXajjkDprtdbzYvGPQn+tyJ+Fcj94WNoDYRO5b0hv8fkvaBYHO
PLy+r1nQvRNgbfMiRc9vZ7wwfMJcG4TSsp5fQUc+TTbxrshe/VTS1iIjRTd2nFXkJwxU56+VtAS4
7+nyModgzcCqu4cv/IieDqnbkM+lXD/aNc3aLCt+kZ0zbXLhpe9/T1qECbXMZBA08bWGLSZI0TSd
ljl6F9stin2OJyv3UUwQOLtPllPBmrSsSCgj2pK5mED+A84LdUzMXOxK8tKMScSmRqBZuEVwArn1
6MyX7R976RFtPIn12LlhPVfAnm6A3c9xsqskuzQyRd6KcJPDDZB49Ztc+4Kewe3b3xTasIBA/yhm
fW92uDiWm/L20EMmLMcTARRqN/umNJug2RO6ZEzNtJ7funJbvJ4IiJG4iAFg/B81b8X0uhCLBrYM
p57icmG4zOZCsPXZkVoy53TuTK95ZwWAEmNTKL9mrBFAqVm4LsARK9ImiEkAk7QrWNCx0zhwbZUf
8pfaLLZMoMam6fOFVoLX9aMNNP5kGHKNx811UY8SaixAoLyWahcFXrj5JhenUEDTW66ChiaZqNlM
xTxLd+lflt0HfhU219mptQAL/yNkhM9LdarjaM28yzZBXGDiu4ZwDjdb1zLoHMrRXuT5bUcl4Fud
nzP6OBY+0BZOpmXqVS82ag0FzPSklXwYoyvX0UJrOBOiaz2swhVAm8CH3+7kTUZQfqt7xOUanp0J
ZLY2G6IidoukqKS+xUjMKatNROgKKeSjwAWqZIjAEhm//luKxo6MolFps5L7Z2q8EPYu4bN9T+ZP
CV1whpT45Tvht4SQigBn+9dZl0807RGAbF8SvnXLdWQrL0LV4cNHAuKXeXbvT4vLNDQwzKjYPT++
FIpD9Z06Ylv8tJDQpFrcKtmAe08TD6kteqJ6dAQkngjUjpzq8g6ysUVI/mPunM2nl0xw4pY09YbG
V2OA4s/HFFBXe9pjNgqNTYXWjfktXlO7eHSrmcRAIr8Kru3EJUyC7FCNq/NH3eU9FCkFFXirceRC
eZZcJvPLcs9cxPKSiZro0Zb6Z7HD3FUoYLNE9mTI9EmuPotUC2Q3rqcKDnIkMUuURJ98ZAB9fqwJ
DskUgFy26NPrVKpYhlqsTSMXN7m8Oww/E08grrDyJ9XvdCNe+WAQFBLldAQN/t8xd1eCSwtbdML1
KmL3jY0YYg0zR7OCZMpOX41/zsTv4kz8IQ8eVSqBt0aPTK6VpL8ONSLO7ABDsPXY2F5BEdkptiA3
hSBC08BrKXdHaXWBidVU0QXyUzQDaSEKt25irBRN1oSN3EJgTxOIf7sTzZvhtR8l7lVQ/jsGBrc/
Gyu+yynKND0TSwa1GXu4rPPuhtksloMFwS8tYlpwyVGM9XlxN7a24l+AeDVE2ZljLxlJHts/8+Wf
9EuIN8XGN260fTyWeZ0pADWBgxXdxqD7MlEFV9qSi+1BMrAf34eVgfAUGXCs3JJ3pzWTcY0GqzIT
+fuwY7qDeZek+X8GU8maOAVtlJOEcDu+MaTiV/QNOhVrGqr2ofjTekejp5xGWdfAiYZd6JNj0m5Z
dQWbqQ87UXsJ5Tn9vEnSqGFTPE86sctVjobBPzaEFbxXeyibqvk64k648bI328PtI7+UnOHw+9AY
ZnVza/SfjnW3QF/5JrGF0P89SX134ggitgWCA+fmwPd50oAsJKuu98oUxq6ExizTrOIoV0Mq7eUP
3prYbVslE/v0zs0av9jX4rcqKeq8/A+Gc5kwLxo+ETiLo6cw4+kV5KIaUEXeGvuHbisGAwhWMY4V
7GR/+y2a7cN1r1TQabUrgVY5Ejup/U98ogTx/cF0dotmcaSv3aSY687g9F6RyUXH0HTX7HKyUwSN
bwDn5x7TpyFFDqZ27A4oeh7LWxpLiED6KCrlG1R7hzF68mlkcHzdhXEkKh2d3X5YAxTZPg8HMfWx
vSs3K0TeOCwWYFnEPj2ZlIaWJJWUJLddO4gbbvp84r/D1Fxu8yk3pDG8hgDTvaOgYYbsWUAnUskd
gZ3EKqbE/A+Pn+rwtHIZFHZNBGpUH7/hG/0FDWNBd55QearBAon6rdmNrdQ9F8TTjhAHrbkROv+b
QG3ug9iNN0SbkKgxqHy1gmooQNNSD2a4t8DUG/jaqspg5tAsW9ePTn9pV0hova5JBncXvzacWRxL
LZeO3qPGBbg6Zp66jDqIOCDW8VYyZcVILB+7ht571S7rp37iNi+Q32T/CArbEUNeru27y/gMYKSO
MiTmcFowYtM/KqzM/31OO8TZXSsWblr00CzCrUb7WqbmYL6GukFl9WXlj3d5MTjIcfyLtQjRReue
Wnge2d6r/MYc6ovHOrMPXlsGGKnGTCArUwSRnDhKQ1UXztEo4C9VOOveT54QDD5WpLdUChr8ywWu
fY3nyYUCgWN9ATAnQQm0z4LE6p72D7iayrxjnTJjOWTKia3o32oQ5pPva5JOuyDeZNPmdKqmDvaZ
/JXQpF9Si9F3zffRs9SvO7kYF5fF7sXmBh//YbGcuFXL+hA+63uwy8E4UML23w9tjadI4mxeSrhf
qE13QAZiJlznUdNXFUYurOQU4u2IS4TYFzugBogtxoDkzfI3Yerrfw9kwe+ngte2kbINsl2LDRel
/yzjV6SgmHQMskJfdYwvK1O4DV2RJNnlwXitS6+yBjeuEr0E6vFnliDl2IM4dwbWUKzrzoMnaw2K
I1jl8RT01JpF7mMIc+6J4hFc6CZ6FLLRhp4+YBnUxAK1/i3Ww/7XxS9IvJ5PwhwVWdxNGvzK0xe0
SJXybOb0oKWcdMnR0QykV7o5Tg31lp2PcSFVKxpALBU1RvEAjJdwffqILT1uybA/PWLSWA/A36sV
qgMAGFyJbgJrXGHm7Vryjlu9r73VCfQmp+hy+OgIodQamiu7EeEUPciuAevxRsspMZVOtObb6tkr
BTYIRIwclyvK6us+UxLRAUmhw5W9s8/F3xAjEQ8MB1d9ilvxXrNm8BkFdNZJlamoKtMMfHcV5fUW
Ik65INm2Vj31NdT+lf534H2txVx2ICajn0MbRgDg7f1es1c/6balS5bcxd7KxLF/n0M5nh/puAjl
NW8kAuxPShYd/NYFwXPZmOZ4Kwc2Ho//4bP3XF/hFUgY20fu1hzxWaCNU/DI/mO9BxkcfmTZ3jP1
B+yJPT0hqu5J2FkSX4ybT6kCDQh9wYxCzP+13lZ2n3vUDJPhuqYFfr/WIPaeeT8BfnwwFGThHtI9
QiDN92eVjdvjqPjarALqs0ETD6FsFcZX7OnWpLk7JTL/dDNpgHaTi7Pp6mUCBrp6RWRA/o6LngbG
WiOVRggIn1LnJaBKJQvSKsw7VcVmpiy7VVjDVKlH2dvWjQH8xmhnB4iz4/8fCletJ1AekJZn+Xjg
1bJJk4kABrEWc7gbR5WUKZF+ZZYIqa4VAM5ndh/CFINmtvQIp6STlptluhlj3IM8lxLN1Rhcq34u
gz6WslrjMNh4GDHBOXleK9joqP30GQCowmVMDX8fhWtaQu0vLmKJ8cxtjw1kIrBwAv0fCnXlYkwe
bWFvsMv72Zig/Beeru3Bi3ISDcHohsIskalMGNwxckf4XpasNYHu29VbflCh1ipBZUiPIW9vsx1W
/pkor29dfUx2aLMhBQqZ6ZUnrRZ85ad+1Y0QA0+wFieD4o21IBcJ3elU8OfDHb3eRBw2wDdaOSps
ASMhEnvFeWDkOZdhACT6AlOPDi6YEa7vqrUuIf+vR5oP9S8gu38ZxFOOsfhYEPmTzaAOguPYJqq/
vCCAtkCUYVbzR8f5D+vaeiaVsFI5dndzAF/1a1/AY1wOPz3lkkctlhH55BCBtGOb9eApmUbCWvMR
d3vRrtuG1oXdu+zY0iE6rR+waUmtPogNnRJZQgKkuTzrq1E80d452Vc8LgUxdKnSW8EUlgRFf9XR
0eJZiQWfxc576z3ZYrV71036aduROiQzn+PT2nPgeTgFx0VGAhpysxcEQr9h1BrC3rWO9N3voA2U
msuyVDfC/3yF7h04hi8y5yuY3M/N60MO+tCeQOEXsFbZy9d4LvvppiRpMOZ3c0lw48jhrAXIBRSF
pxvSNE6cNH7NzJ45nf1CXU5w+5gVuE8DTsDKFSc8+pfG0TP0i4ia309mWzy1mPAY8NdMZLGyTtTP
S4AjcbBRoXHzP/VvFSpCN0x8DKbVkIxqPCQmJ2+jSwYbQpXEc296I4avd/0yn8FtqP6ett/nQ3lk
bWwj8OIdAv1apAPEqDd2WM9kGR7x5YD83jJEP62AjC5f43vKFXn++N8vbueAG93KKxoFT9AY6QDE
ktJlKmhtzhPEKuCLoHS5igWkDCuBeRrYO3kjePkPvZ/dQ4X61YnF4OmOXMnadwjp7lGJBsYL46iW
TYi7GwTk2SQs7/ybXJhoxqJP1XUg+Y1ImgUpxae+0ArEas65szZcYq7EEsl/U91dLAq/cVnRtEpg
QsbztnED3tJDlPnMQHs4Oykn4ijBhedLWh1u/VKWG0oxKH0pOYdz7cIGjxedQvQ/1Jc9uQdTH0Ae
6/M4zD/wJQdO+bhidtE9FQUsknKhNDFrtJGUkwB3LlyHM/Yxr0mtO6QfCNST5bXFl2PuhnlKE/xH
YM1atjcdIOGcZc+9anft5zXOg8xTWwAkWIDDAKqho8eLCA+Z/5eC2O2hXdkkZbcwVULAeBAqQNsN
DxdfxAA3+XdPrTtxwcmDxnR/aS4W0mm7vzpK9haXY8lKAhicbeJjZ3akCu9p/Car0psfv3k+y/yN
O579/znaAyZpt5qvQZsXpt5VGDvH/yhnyJDW0Ak03XBML1PV7t5xIBpBgBS5UfHa5MrkEh+hXdHE
rdDdbHgbUxfkDNq90APOmSdoZCoha+Qxmme3W2aIIFigk+stUyUYzKAB0jy4oNN6HSkDgV5QkSXS
oQnQP4vlR7qo5xx0oS8VqlVySJKBG5t3Ku0nGa7XAqI5WNEPzdyNJ/AW78UmCpb5FSxofo/Qrutt
pwwzdaHCv/a5RQ18cR0t8aog/rxxmLS1W0L6VZnw1VI4Yc4tPpS/brIK82Kvna0+pDojKNglV5u4
05WisCj0DyhX6Q9J1AeYX17BoQlPEy2xhcz2sJVDlxzOQZKBMvIp5lBTPZbk/LRyUEQIO+CN+emt
HyZ5p/10EGJs7gyshJ+PEl5WU0SEHj7B3AYVAA6cHm7ngW827gTaAAQqu7wN5qszsDa9uG8QThD2
glLBovTpyHMIaErFlJm+MZ67BW8LynG6rmVbDyhfi3x2IpQdjkne5WrMKSvQT4nIwwSZ8Tr+UspG
T9lUsXJ43EtzREVw+fKS6v5srMKaDRVoM/RpBX0ozDTc6W95Kj/jsPyvyoBZnU69jVK/FLviRNWb
wOeixLHytGDw+/2qpdqgOU0zRFlI0BSh3ZW4BpBq5FzutJdDU3pCC/R78IcgH0hVgNCuSjad/Ml4
FXv0c5o7k5PbRYZFxuQ3crqDqyePYGUXuOeHzpVqBhHyqw6vwBPurcJJqQKSILhfSiVg896k9nxm
FbLfokJ6sC/xDrtEPm38HxxTfy+yXMpcTjF0tvmay1xgY4EmjoR6VTPp6/fBl1lX2KVRiZCX9ZVl
5Lp4H4fqpyxlRtDMmr5jpF1g46C9labo6y5kod+CukuI2704PkgEDUX6XSwexALxWPCUjK2ou0lS
IaC6Dg0uofVLLBh6XizybPxrnxbS6ZIA8BKDjsJrLRhc6d/cEOmntB4Qp3v2IoNcXKZgX1m7MNbw
nZfSw8opmwUiHXKUEIP3my6BGM9pKhMO1TOn45GHqNz10POtFb8xDkMxvhb8WFkY8bSz0iHkXPfC
I7PIljks+/uEEU+n10NBOaefJfc2jIlwf9X0kJfux7bavXfnr/jEU2J68y1/SptFFdf2wp8uSfnw
8nNXtncKRh+0S2Cs/2RiXcRgiVNwoyn0RuFpuy8SVdHQKTIoRAxrFah6k42knbLuvA5GX68Ck8Op
VxVhkijhvREJ8QYsDI3mY5HN5ZA14MwfLAwvfI2PDHhISgLHcylqkRr5ClBi534xusAyslIMfQQg
Rs8haVZz2NT6ZIr+jYdEFdQ5o86V6YUldT105//JpMktlkyaJWJB3AIU5Ovt3CRRfnnP3BjOSre+
FRqUDrtSSgz5VRJ0iOgWutSgQEyn0WgU8MYGYy+hCfazIgly9h6TgOBZOnizrHySqRr7LHZtj8jj
N+McLRZxjH4iTj22RzwAVno/MSKWtZJy5cssHmTt0FwW+m0jzGRwSIJT0FTlFqn9Cg1UdgmN7aSn
vNWIXBT6cmsof/rLnCrq1DZ9/z/5bo1IHL2sQGZ87uzM19EUBVjBjbzoU+VwpOB6/DnaBdAKrCAZ
iHGHkxJSQOU2/Nrf8n1byOD6oEzPNe/z3wnfxl6vbHfqC/nGTQzjsagrdqxeYz1Dn9Xekf8u845R
ED5XnmNVhO/T25utMbRbAjI4At9GdaBiRuTRBGy1ISyCvHrKxDK7KQikbHvuuzpWAQfxGN8FKVzu
tZXXht+TTfGFCJ7dsXpXg46LtKH6Pv5PAPaTzZ0xWfVgrh+Dbnbct4tefHk6igS1+FmIi3M2xcJz
ND8s0JQc1TspWxkhVd6dX3D8kanwVk9zb/ZHCUiz5YPTWWKoJ3cAG8f3BNrj+QJbpHJDeB97T0Z3
24xqR+q6R2NgH2qINcPTyzIUXYlO5AmYta1NzbqR6IEJ/0133ExqO9XCwISst6xfU6iOh6ffznUQ
FmTNIXUs/62G6b3MAiYm4729YeW9DsDMsmSD5fgQGA0wjvFFLeivE36VqTvN6wCtKC/CX6wQWRSm
WQ5jdCsUGU2dDNA14j2a203307TmSjzpKE46obfsPQRs52f5VmyAE0JcBHvmuXfTbLdtxSnxwINz
l3ixnFalQR0k5n4P91GxQdwITebPOB/2KAhvidS51Yt4osC2M6BJs8T4aglFCjgkvq0p1F2uAknT
UO55Mw5N1Wh70AqkUzX0IMoQ/ITtXtye5MxqywM9WKHkfFqnvKLeEgpWxSuReh7hkOYPyNjScs5t
TQbQWcqKno/z/UUQuelOUJLnCM9vZi7Er1WphVc7d4KztQ2k1AyJBr438s4fyohV39ZlUbtXmLAd
89fTeG2oec3Eu89POAAZLAxgm9k6LCnaQHSPiJeSta4KbMbVUVA9gxybyd7Q9xSc07rYfWysKUgW
8t2X/Ei2wr0JZKV7v6tfFSd+5TUrMlVcKQ/4kR2b4OJWR01fsdMH5vbL9BQOjMpcrB3r9w5Vsog5
xJRyHrBBXSUmE+wSz74bm3NHRIskXnuiDclEkHy2kX7eYtxgvpACrACCaDlC4tFm+XOE9DIWHlWA
VNRkEnQR+huzEl1XGOAjDuZnNSwk8JNYo+5xyfgSwZE6i08wNA0eiliysps/95CQi5XwHYHiWfrB
4Ay1M1I/uxI5I7L9qw3dzySF9IBkN3dOgW5mz9NuuV+yKEJbpz/vd5CMA+lUaUBi72Q+k4SppPW4
fkk2aJD45bC8jPX/MqivFp6hkRXF5XTZ9dSCcMjgs6eJl9Z5JEvsIv8TYyevl5q73gtI9tXJKboW
tzTiYZ/gVaaRp6J+AWm95CZcd9nLV76Ljza3z1by8kHbZnLjZ3ahTcNGaJVpekj6sZE3QFiBUUTV
A4F7X+6cR8RuYVlPRrO6MfqD4mgjpypWbFBKdSAuVWQamt7qmAkn/VPraG+b4m7jnV9rXmmvJTVq
ZtaFuiPuF+apkRQ7ZwcoD/D/XgpcBzlaDau2vtQFJXIbtTViURTiPzvhP3jXAtCwSt+qpgkmYU9X
N+3TuhK3az/Ss7JmOCAUC3xyzUaSfRftQom3WIu7Ufh7nQZ/3OmUovd1bgtGdCqG8qkjZ9qeLVep
u71mN7q79fMVkLmtaNbEZilo9zz3TG7Zqvm5lnizdgBGIM2kCNB+R8lkXF+Q7fWgPtgZMSUlP8se
nhQdkxDscCMfAuJCebU0HwTtHtAOCjyzGzBA2B3EQ6ZCPOAxARUxsLlUAbpyn1apzkg9+H1+SiB4
dlaFHpujpa+RyV46pVQwmJ6xMQfr7df2XvmmVyc+VJomauvU+3CXOW6Nw/uTEo3F5etnaIMrPJpM
vYlSEYg7k8x5Cf0KEs6k+9qRlVkt5kwjftu7ooUMzqr3kjuOYSABAvSPy9+sk/11lSC6nByN2wpq
K3tqr5S6qY21YRdcP6ahgnitBuKAhCgARMnBUg0SJRPlhv8zIpp7cIU3WQ5IgS98SRACZ5+3CPrS
1ZqX8NWjaQ5GzQCZKVjG+1nHhxmtRbq4/XyqgiBp3TBwq73Ga9Sb+McCEYvmTtnZ0cY7OzwvM+Dm
Pa9PlXum2OYqIRIUztAsDSUtUdJuat4/DtArwdcHCO+7q6FrAAi0YU/VLxSxCYe8yCFDUbNUkVAs
jSMZVxw9BY6yxqk+RElSYkw16WkCAehPvQcAFByQhr9ecivSDAUUI5dKJodzCwR+7MaEh0blCxBc
2YsFnRfl/631LJoc8OG8wE8+e/1u7s6cB0nDkgkh5cuVKGLT/r/xoqJ9h+IsSpankICTs8jkZ20P
29XtOiMA4+UL24vNPqdBO/DGMWdtSFQsbDSXS0VRqVaWud3jTgQch5U+yn5hhwEP+j6KyiV77HgA
BP9b+XP5b7cFlgb7vf20okQgxw/0qDsxviJOIAytG0+dE6lLGDRNv0eg/3KiuDdZdqJHi3MHSaNW
v89UaJ50GqtkcjV5rau1SCrFSIS+6Ugm6Q4i819KfgtTzoGEFn3pRUUD1umyRcSBEe7ox97IpnrQ
JomRfr4MKG71nOYSF/xuHGuPvkiRIfNV5eBHEwfzMkDQ20b1e7k02EOFKLcPJWKiv7UsgWwh26IU
Qhd/oBB/qwoa4+Ntow7ZGjTOtVCGNTSG/RfZ9qkDhzA9q+hZRj3HXYfScl8xAi6gTxnYUgtg3hqs
7v+dWC4KKvyuSQIXv+6tSctFnrnCQs/fu2OV7Hr7AkT5ALKetHxyx72HSSwv9/4bW7Cl7kkvHu3h
rTW6jBAgqw+DwSIFYbgTh36qVuOFKHUYL++R2nWwJoUB9dZIkiAGvgOydt40Yf9aCSLCLg7U5T8r
OAbGoAptvesEP3pYeOKge5qXM7kFmkrZjV3ufdij2em6TVb8/rtlWlVrcfvFi5Yt3U43oAnnBjGV
xVVA+XiAFEnuG5kM+I5ki9pF/IrABwUVbrsLkxAoxndIqJL0eC6WWGIv9Cs4vgZeid9eomY0PeaY
K2ZBuwBlNXWGJ2R7SgWWfOGljx76Hn9XmiRGkFTdb2jxi7fpgR3Tc4aegAU8j3xS2TVx+aGslyuu
136XtK5WbwPzmeGVYXQVSjfU4N1wf9RtlOYGVS6m1CVgbjjuXMHH1neB6hyfo9mjRWgHIJ4GtRVV
Q0kNfQPnHpns5ZKLFm5PTPFRqw6YHeCBagXOAm182imflJsPvfDry3zT+lmCwbCmHB0y6Ryh6AGh
aPZJgQgiwe25CZzvWanghDkTBhk35lt9LHdx9HQhlO2e3t7c3syd0OV4DkElKtJWm+uy27N6no5e
lmTR64O+Pov13DQQgxSEoY/1KcK7ZnOlw1hVRUkGyCtK5bpOzgmkXSPBLWBFDUkKaizFiEXYKJ11
kMYauhoLZNw/doP6VVAQvgQfWAnn3bR3w4xVkqaQV01mUFnohwEnwtI/mKAAZLUJGK/rJ5NjvB00
62qYkYA0AQchIxKgi+rEgMYVrrBH4IuXXuYi5mVCCmr935WXBPyffuQL6u99iH4zCuSKwDuMSUAW
DGT0FS9mYHiU256VRIi9UnUx+1Xy7zmM0M5vs6SI/u/S3ZXdP9CGjmP5Dvh64frQ+0pH9HFmrZn9
agTCd7hMuFNgjBLJnMGlHJzb2rT6xVOIXSRQazx5q5xNXzVRJYkMyKGuxlC02IIuuFr4sZJCPlcL
IG3eBrhDncIxLTuiZnLY6nd9lS2x2F4JCh815+Q3VdOtEysvsyfMtOH+LjOBoSl7w3gcSEwlofoO
KrbyADTteW2Cni+X/PI2ljooG5Y7QdPHdFJ/hsXLpVdaCmvpqhCOANF9b8XEX4ZlB/DYfm7jSdyr
ZjwePAVyYj1I4wcfiVm7ia31ESrDbfQ1dpBZygd/4sBsANeu/wpugRHJdR9dB3EicD547x6aiSju
RhKQZFZOR4/2LxmXnlU7QkIQeMof0AgkZ1u0ISSbNlLpY82ACgnAcblxjAwU2dmZEN+ddwMUhV4M
v4yV74LJpTl0Mpb+KbGtOjwQR7Rg/WIFp0Na9D9psgBj1oydRtFk2MXVUGLRA3CMxUbsR63gm+K+
Obu2rd4C3GKypH5vfFcdjAwhjWzs0vddAHRvUIglJFxFw1+RvRV48TBtAWref1QJKzWnjTpKdRkH
7kpgYaLsQmbzlCKUuAOhxa7xWq7rfY4I2wjc1d+jqcOS6b053zPVschE/DMocDsWq0VuTALtOaNt
Roj4MDEF+rIYAgLMfhGs0Tx1489eTYtMwKKJrtMyQv9ovj/6j7sE9O01OWxh27DDX4O94xIdXpxJ
LFEnvxlXzQJNB5Nyczf4GainDM68hzcrAL5sqvDWRJH5QfjhSAqOZ7Kk4Uw2NkzwtymHKSkko6Bs
fOKv9VIfVFPpFdEN6aIJ1K3eNF8gL+pTFS7qlFgREJDu9vG0XE2gBF3rjv46ZE1eJfTVgBh+dM9H
PDMLSgTmceBavScKYPZjw9cPNFAhx0vrFCJ8ky8zi5uJ5V4ZS05HqZNO8PD/qCdT8MEXq63Cz4ho
yGJpA0lNUlhtC7zwoaunXtz8bHQ/wT6Iaa5GSV5cG+2mQB0Q8u3CYY4bx5d4sDD0Qhm+2wYrsvme
MKU2/qMkbfXEBuypTSkouUjTHdfjyCG3Z3zspUMhLKJQeF0Wic+cCvi+SCSCuk01vv4L9kvE+kRi
7sWJIocBAV4DkI2n7lp4sCSCun2R/ICrKaTY1fhRhTfAFKcHdelJMo7dngFyBliYtOzGgotiMJsV
Km6mEsRYgSe422j8vcaMfN6So2XYI8gNQYWOvu6MH8c3efMfAPg7msnCqNd4ZVfuIkiABea4sNZE
boiB3NX35DTgvTgMwNOLlCxUPB2esH6yBAu4NGgQyi2ljP+o7nQ2QyjhsLTd2rGDB8cgtlodRF3E
ulJedFb44NR1LoaLf4XyPpwPq2r6roKp7JZsFyavJZHdkZSEkcuV6gaWegh9dDCBzeKghiHSG5R7
b0PrhLvvX9D6VJBTu9JpuWsFVIQ1cuWDHEARWFxoTJN/mnq7BSCrpP9ioxPisSDYxq4fG/Sv03o+
SYQSTyOAGALJ6NT28FDbca/e+J60JgeFExoSOuzAHBJNftvnix82kG/oeHJzkXfHWGIyuTnBVIO4
QL4PtJiC5SgD0SBVXMF7RcK/QTQhePzSi78OGGs8YCJVjQ7KVfWI5U18SqnyUufxo1WCCswr7gt+
m3uvfzV86qw6yr3fdqDjaJdZOUbfhyO/5CYp23MT91f6qR+sUZqKYkuEdc0fw2VoOGBYq4Y/oxYZ
IO4hqs++hm0UgWyuDj8mj63HrTFJVS3R9XDptioTeUxhrfQP8rDLu0XWptdJ7EDlHf654fi745uN
ZLbUpPBeAnD86ma+h13mkIGD+1UvPOscTsOU1IZu9WHkRDC7MPzZb2GI333PnNbw5408m1aZ1nxL
rHlYLMe0niLi42S5+OU1DLEc6Lo4Dhih3vSe5RXIBi0xuS5D0UPKTP+J7FvkAAvn2Dav4K1XbwqZ
ky2RIe9jY7LOmP3xekE9Xbq5Jlkf/BfvRHypBi+pIAnqwjbfaIX1Zka0iqDhPEzYPp/IPDLoaYbD
Mbna6DKCuzlVAhuEqR582FYz57Yj2yy4vKJg8bW3HBp9WUoGXlKozXwJR1C3WVvm0bFfKdBw//is
RLSAnQea+KGIaXWFEwZrQBhqHmJEF+DBCtZnPUL9BwnkpBa9GJMqvV0PXsZmMUvKR38Sk+496atR
du7h897txqwmvu18D4pgTyzEeW+3UcIK7pI7iryN26kt1Ag9iDWnMyIsLJXUvNfAXlk70uf6hsZE
m8zKabPQbzfv7CJ72uirajsND73BB2aZPNY8vTRc7Aj12NOOlWV5br7mbTmckcaUDMnr40bviwPz
71bi2WxmkO3oKYVRZocuWB4FacFjUK04giE/PgIntDQSrXfF7uC2Op+N8ScwsLLVfhzHihkvN2C3
iYC0KWpmTiVfE3fLFlj911CD9SPZeE52yK7akl+/P5Y5bFO+Bgn+LGBAWCT3jAq7IYl7jXBuYuxg
A0SHaA2gY+AVBBD7FZZ81dHRsfmK6WQyordLGgT0XV3bXRglhsXXgaYj962/ayXyatEI0htjwKk9
qyMlSeN6Ozeh21KbSK6l0c0gPnG4PuddkZsjhC6JW3kK1wbVjnejSzo51ka9V3Wa3TolzMVdcv9F
3FjAt3VlgAdVtP/tUkF2DCv1FQPjX37+P0tQ0xNnnJg9yES8aSwmCqAcWc6LUqt5zJJuNALetyJ7
99N4JI0KIK91Q0WC6mToZgec/96aLCcBKswvt8pB2Vf38uxgFVJhRIA2rgMYQhIVuGYZYD6BozWz
zFKbfWJZoRvsYxpcFJKSiSP+YyY3kuXXvF+bQOBDhZrsvqm8BEPnOxVO2TZRfQAKf1ix/yrhS6U9
M+Si8KoVMORAk89hyCepP9FldigjNDgiAcJvWXtO970Tx0EPqcAN3TIiSemBNwV6CpqE+SIKsTA7
uc3Vc0XOGGZG7MQbqCdNuxRsVkXBWGwoElik0V3sDiVKG5x6/tqZUeLGrGBM9YmIP0PiWxYvYk4e
lJrVrNb3zCRzUR6OAh3ESrOaTxQKD7u7XGmufOK1bQiAN092CEJknIQd1ZWIsvH4NKILXag5lDvW
9I4LjwfOXyS/WV5hdH6isMagSADmlLDB3n4w2drq5ZPRbCdqoGwo68O5fgiBrT/aUeKlySnqhLQ9
37ft03lWDm3QYhW4d+eOl0ab1OOHZ/YCxqL94VsnKeYtYfoTtjzIjuiGfBBw7+rg49AnRZsznkC9
K672c7iyr31q6fgQlmZviWBQHGBJ6jOAuyY2JT/UG1t8NsAA1x9XQUfL9JxvJwpz1CXqdPcGZ9nr
DCAxD63HISQ7lTN9JsL47kQ2vSzUNH358eTf/+I0NFbyTV1xSBrUlhbFJj83d5rRUwfeNpqy4znd
7OUXetkBW21hx+p3+A94O0vg7d3uVPCCwf0km+1q9T4M6Bk/FPFOgi5/jMV5zyegy9+iOZlePP+W
r5b9VYZ4gxvpwp5Vn6fg1+rIfwi9pVRudSWoK3PvxRcDXmTFjCVyOTjkKvxjD5xWpaDVpq3cdiTL
iVoxOlD4qexUT2jgPd8p/8oTgCmWfoV2U1f0nkh5038ZVKDBV8YJpjZJH9JogNiqbqo3Arts81QP
qEhBzv9Ew9tNaybsoYGz5eBfv3n3FKtE8UQpku0jfX518k/c3N12NZPmhbIt1XbdMiKMAxwtBIfV
A/9j14xn+zkiSfGrDA36ugypb0B8joJ9kipe9MR0+2df6zVdRAM7Y1BrT73QLnAEWDT4kd7U0/Pu
0kaHKCRNxlTs0AQZ7zQgVF4O1PMwKcaq/pMj9/rO0y/RUg55Tm3lyWCle9LjbXUOIE1IrphXPrth
Nn8SX8YeDadhdLI+TjTASh44hi5k91+lraaV6MU/7BDK+6aJCDFYjDi93KZCuSzUInx1mHe+Omse
iSF4a7CiAXlG/6ptu4aaCah3VD+pCfHtBbWkzFD91njBsQeYPV4jtCdV3RSAR5TRP+gTnnjp5b2X
BoCBDPBCmHRX5JdNvdrNPOnWcJRFOVWaT8+r5KI4rKWp4SngcIMv6RX4CV7Ix8+kHkKiyPKvy4Ru
WMxrXCwsyEDLU0EkhCBbNiY5wFjIMG8zdgLXxthJaJeE58/M/n4Dj0ewG8oaya/YLnzIHWycpj8x
ra12mXf0GI9OZQzw+B35FeQ077ZVY/bMMUQPxiC4y/rMqpDQ2QjFeyq41pV88s6uN7HLQaoobVSb
LcB7/MFLbgpX7k9kmjRsLSK00ls6eOuMuLVtE6iDHL4Xqd1aWoVVm5zzUTUI2iNBFRs8OrezuwLQ
S6hANJuvO6A9XQ6SGU6zU/IQSbFDuHB5bIfPLFWmIOO8WZk61cV18XPXODEeI8Is2cuwNmbBGdbL
FSg2Hkjpai1mLt25NNV2Tmh8CwTVaJFPGwzLf71os7ldvhSp4eqhKBtwohNZKWm9lNe7YAvDtWkC
nla1Qv1gg34ee5Yp/3R72OU/mERnoNl65qc3QrAaQ3Sm+bqDfK9OfxytkflcUOq74rJvKJX4Apuc
FGF3uvlrdScPSftqbR+FdbF+bvWYEPeZxt4h1Cr2ylwZhA4NI1jNKf17DNO/ukMZ626Ox7AaGPFK
bzqU8uM3Is4h04Nyg6qImYPKognnPQxFxKfBss65dNbI7CkYKLJc7/II9upgydjHJsvw6dKg7Omz
jIUZv7ZumO0NnKRsgL5U++3wsoFgR4oE+O7+97ZNUHiPbtQc1sGEq8GrMcMlKlwJ+HM32jMvBILE
endi8blt+ESnR2ziHwMuoU7XZRw7S2N/Nm8kt/DWp4pExpIO9QqL/LiDO+1kgVn/5fdwFF7gAV9N
lZwC+c/KUMlPTLTAbwyJ69A2lSiRHQgvE6h7aFoZT5qOE4h1jiMfO8GpdyeFTkYd5Bgy/jsGDx4f
+IDwzLOmC8Opjk5GGIhMpxNFUXDlScr3w2q+UNda4BRRxbZbNKNTAuHzUpLimUkLRY94XnUus80m
sK5khGIL7I9nY7lhPt8uGC2BQ7n2OuadmmaNHfd6NI4U1gXDvBpfBzm08dVZAxQT6kvm77dhcSt2
BQpO1AHE1sn438FGdBLWXny6f4BGOnecebtBN0Piqb+PcN0E6gSwBeCpqtTSscroy/ysAlZYnyA4
7PAJBo6g/+hxkdPtBgVNlMDVuOewCGY8NP5acso9luxWoU+ePJmWVWd06l8/z+bspiuifUuLK8HL
FGp829amX7m+J0P+CBWvzzvtTiyUk+BeqK70oSsgJcWi0Lwa8B3ceBaX0/eTOeWPCXcvo0NIu2dW
76n/emJBSHRBsJ0TfBpiIEC7an+k3Q6vOuhMA0iHC3sIbljRKXtTGscQBpBKZCBupwFX9fU/WQ3J
xAHHQ/DRkk8NmaRFAlzeGlZ8jXlAv+5xTXd8kX1U0He4y79kTaSC5XuQtK4v4+26l8EXzLpiSyRp
RbjzSbq6Od9NnqEauQJWldT/4GuJJ3zHiZBuiSGcwPgi2cl0WdySUKnL1Aqx+uVUsU4aEL3WSU6l
dcmOccglpHvnGS/vsgnhG+SC5cByip/UTJdbudWvjPFiN+svt0WRoWEB+J+hCzcISnrQ03maaJLB
aYOgAFO8VpPvXFyAhWCoXuXJcIJdkNjjRz9jhVe4GnAMwZFvXmSC06EmUC7P6DtBfeDXWr6WxxAD
GoikACF0mFLQNV9O/IaYrmeRR1wiIT6lvNTehy+dm4kFPSrvZC2YqPPHnQU1FX7FjlNtwAsNWBb7
z+lkBCOnjAvwtFEWKBx47XhozMRMeiwmcOhnSuUJraU+8VaGvs3e3m5oeS5K/RKei1WWxkxXNoWt
txbwc5pMAw4SwLy3O9yfRNYb3R30lryE0nbeO7UqoUlYxoZHYkDQd4u08uzzl+VAUCx3AzkIlafu
nyPAzcOxNRPrGkWr/mnycPj8/QrCJ6WxBXnAT6RYoJ/eaNDvdWTKnplNj+gfp7qpDie8I4SAvM4V
L2rGak1bQs1BTfJg+68uOoTZc75tUxOy6rxYyeMjys1IcSM9CNE+o0ZDKjWeQVH3/ROcGrGBwdCV
8x1IHj8FssAFvoRGeJ93/IEDJ9ZU8lpwjGpp0ISLiWPRLnanCaDCGAgH4m5R1prlP/fpQyoaaj7S
Eyn83mXbe0JWzk8kzZg5I/Ho9MhTvS3PVu6oG4XGZti7rJjwStJm/WPrD5yXuMh+Dat+HXPDULxa
FDs5y9j7a8okCGikhaW4ek2J7Y0VeH/tA1aIwflVsOJ52v2w/WjU9/RMEzKY+5EYld2RL12HphIk
y/i2wgsykNWFzpbEvqq0e0r+z2UZgU1GCgLKSIZBUhoomH+6jRSBgPqo2VpubWDJYBRGfjXHpeM0
Yj/XVKGSQwancqvvpexJsIrLJ/9YtY9rEkbpamhjv3QO6agxgHysn1yJbgFBMAUh5xOAEji/p6HP
l0IEERdk+pcf/TX3lF/0mh96n51MD6OM2VL5FevPT4J9ZiL6SHCFOGZCiPXPN0BdnZHrMsHmBgdM
9mevR9duBLLqZCbiBRKZlPFz/BubwAdUOzt7pBEmMXXTTlbNk9z6l1SrbbW9fMeG1zZdA5Iibgxu
UcMJfuzpw0ItwUqSjIfBH5Ofx/uxhyCNA7ZkUq7i9/6Cy/IuVG2bqqrE5cZSxo3EmhZZJeG4nw/K
VySwdwkOftFgPu8KO73nXQZjlm61vCN1cRoRvM6onrgMZWaJVq9MdG9Te+tDL2l1pzLA6rXoGHLO
486fFiJrEcTO3ma00iee5aYXG+g9Q+ooFfVTp2zN5Bc/hSA2DsOoZ2THeR4P02ndbUgoNo+SYSjU
KKI/8Djb0O2AE9GafNmZHbZO22pHkT7DBKZHfWeqreeWtV8hRtYCz6QcoTW7633smGGMK6/XSK4c
1BaKwqLpWcyu3cnuRAa74zbxaL+wDwnFP1S0H+s3XNl7/t7fdJRAmg2myb9a+CFPbTzkBvNZaHBg
9a1G+3+z6hfUYtU2IMR1KbX+IbpRx7rEDGRG9qULBFnjRycIaWCtJzzHIfyiSKR2yWi4PCI5y52k
9cOt7+9eLjhVIFHPACILq31x5xYaM90ygfwqrbukWxw7DQnygcpHab1QIVb86TcZ+g5nWpyTFGQN
zBYthd36TnxcjfO9i+BxYvS0RtefcQ/D+xgx8u/tCzrbjiS/RRxmUcuqf0YB+KfH8L+u1OgWXQSu
l/tpm/QLHpiDj2yBLder28/KYjGrJbRe2hSy7EM8fy77ncgIPp5xIyc6KluwtSSXujeUOwhD7Lon
qVVafj2S5SqKT1rvEco4fTbbXrEMsf4SGdA0PSBG01BtX4LR8gaz1+F6UVviDNWheVT+p/HsxXDS
EhbtW4rZRq5yzwUjuHUjFC2dpXGWvAIqwmfqb2Hjhiklx8p20ZznJRl1tv0WQZQ/z0qbGsTgEKCr
l4E29yy3/Sn5YoL3PHKkXnpMLMHZgIERDtMxIJzIvD/bdRXPWx7aTM+KaLV3b+vngJrXPUEJIXkx
g921tR7G/G4J5a8hn06Cyn16StHjpX1xlJfIfCrprvKl33VFcmOLWfZt6/siEn1Ls48XHZ4fviWB
N4t0PeAcZ0Qh33qowKvul9hakYEIFxK3pqIatbHoA2et28XFvJGtba5bVCq7RBVRhj4Sb7GzArZ3
Vn8YSqstkjvmgxU4M/MISzhHxsP3MaH6bfjDrYRjBsjNMiofJVhtRqXm4ClIiJBHHLLhTL2vpXHu
eyzSERUicKUYkavJhf5AU7La9zZQKtviBSqyRPCZWt2JQvYQ/aY5XfFOvmU2hk/hs5nUysIgPHe4
2wN0KBOfCyEc9dE6HGE5ItydT55S2GmsvxE1qLMcBgYk+grPS4ur3nG5oNBrh2BTMj7jIrUUHTZG
pRkHaQYpd8vqNt73d8ABsbkTdoBEZvfPir94law0Jc7aKbQCItGQ1tUBYebHXQDDhgeG+wFTfK7m
A6bncIKBn/sL301vtoe52VOusGAU3GQjhnekkgMGy9K4TT+AaPJCE0IE3zKCqwVmLzMWwVz+QfWH
YP1pQqCWNesRibl+befJKEZtD8pHPIfcmge/U+8jvGp1q+yakuptKPG5IKp47QZzSK6I4mcWNDBh
YJh6jn4OP64QRLYvUxjoENfNPUPq3DwL2fXjkLMOyGkhINzZRZUQHBKdMxeWz7BvTzda/epvnIwQ
gCsDzYRUdHOHIagEXexxP+eUfSKRbg6nQYo9xWfZEkqoSgNxDCrDWBu17T/Pm3hL2PshWigBLEeD
Kp4r1wlAw42HQXk8eV2OFF+aHdUrokISkYVfT+8kBLnAqRWBNl6AZdZN78DCYP7QZd7akDbA54IA
C8392qRKkV7wSSh2D8h7JIBj7Q4kXjtsyIeBmKbdzVboSyb29eg6bwdqvNs2f6VauRsLbnu+PX/o
eVL3Yj4r//HQB1PHbWJ8h0a+dcqI4SEVFWy7wa7yvk/Lf8WCSUg4MHmE4dZ/bdS6dmElIGMupkH2
MQtMeHes/fnX1f25nZctyDZtIu6gn6DxF6MOHMtyNoUj/bzhjzlpXsCZMEnDW7VHlgjl5qY0TIg7
3v2epry85/rtISBB1N4IZ3XuCKDixgnOzeUU4BsLamfEpMtfj4P18ZtfZaYr2sUabCp+UYsgt2B9
upgutRHV73TKVZp8P8Q4pW0IcS61SqXQvnoK40lqTSnBRTtbvc9JdhInXie+hmiS3b/bsxGkY1YA
Ck1cbJmZf1rPOKLrJBf7mn9BpOLsdr0QRPnlpkgtjCSP5GU2LqoTPBnJ1GZk2aYEzd38GCXi5ytC
hR1yI9w8o0Nr291wwIDxY9Rt3Bw8wX+LXg06u8/MVtijehpJ5QwRq55mX6LtKraNf4r186fwqTn4
nnhaqwkWa+PGi/8h/e9FyjZyk67+Rz2RI1kPfBFRq4gtJOVTzdhsOoIgAxJkaMc5ulk0pNudBveH
GZmA6VStyIypu1TJX5kH2+5iRm1j/ZrqtuxGOCQMD1fOmB17jFIfpxiMidUCbKHCALB0PQZXYGyB
s8PGZs+h31IGjc0CesZNYPEm2Pwcq7sCYNVScsBIwQKdG2MMmjS2Cbj9USEvPso8o/tz+yQMxmHN
WWwl5/MT5oJ53y2cxWhE4u+yOZiPHZdhQ1yH8FUNGrgFCTo/3GFJFmesBHYi1FplOxn/XOI2FYoI
xcH64ranwO6hCq6DIkiQK3n7zEcy/YWQeDJ+dHmwxknGvjZZoXB6Z2RKTsuuye1N4/+lgNSr45M8
TAd/V1IxABFEX32Gk7H7JReGZgFCvyxvWgbgMBhjzqJ5p0n5VVs23qDOMLOKNRjHIjfGuWhhcfz6
1ViWs3bF7ujhQz8t/Gx3jtP2gXVcl/QRqh+TiTpM/rxUuN+nLO67J52XSjloQYOSRJVwhWs5LAUy
sD66MttBqYkU9czGhBRvu/Ha+C207F8hr/4B1hV7/YrlYCSIZwZOMONHj53h5HX6AMWYZuOss0Im
LMR0vRJ82iOLfrc2ANymFFJw1R/PR5TUc5FchdOp1tQwvBZ0DvstUECuIw1D6ww48x8T1c8agfYD
i6yBQlWdBYcUHWxGyVGaxb0g+WLedt9BfyiftvAk/BCVC+MdFOznn9l27rVmZFQjD0+N5TDUyP/i
tb+3VLzCnSrFuWYG1VocCM6ESJIuojVT2JuD/20wiDXQrdkKUL4HpxuD6ZrjsPPnHOFFMdT+W0y+
uwEq/fhK+x+Q+MpcT1Oky09ZxmpA6ok1Gh2D81EDEhwNMmoyFEUoVlMnmenCqUB5BaE/sIrd32Z3
anwvnnpcRngkgkE7zLEZWOHBAGAtsINuI4ilpJjYRiWD+Neh19/DQOUet079WMK0YvbzFe9SQ1fR
yuZTMvzsY7im5nrWONa1uys39ubAzP21ofzTTM4FbY4LRYtY4jmkqdDlFDE6PJALja+1Vh9Or2Tp
pbUKnmk6AhgQXmGDdNUf/LMx3/AozBMitOdG15eNNHqZnfnKsvIB93BED/9N23s4K0RgTAbuuxXl
nVfswAK1nB8iLw8OYcqA17fHIwW0aKD86WpdD6TNGGjRHKKsrtPveqqWeKUyPgEoxeKWnDuI7KoN
OwzDlFgRaNxl3TM22Ul/WKAws4eeuB8VV9hitp+S35rQ27trdxxIEKWbY/dWHejTS7v6e2Zh9s6J
0D5oJ9lz2JL1w6hI4U3bTNz5iPzQsUSI5Y580/V0zHCr5p7HXb25uzh514oL2IKkZgLe8/Ggvzdj
cXJ5KzE9YwttIjU51Cl3dFDGm1jL5Xw2sje7fA7SzSNWdx2Qhhw9vC0g5kZUEltcekxNYj/iRkZp
o/WyN+Nw1JW/Bspv1Qt+DgrgesSBdH0+dIrkuvI1JWgXdpMgyMJdHe5nmcjmMINGWcwRQvBsbEFB
p+inRkHMuOBbh1a7DKlpHl5hbV7TJdbyAHKtLGUP++9k1fNXwgiqS+ihdIuE55teLNdc0MIOFvVK
omwgQVi/yCKOGXgR9fXED6HEyW7p3KVYICotCPmZ8iPkGTKAYV4aP0fJO7nL1N4ThwGmY7c4Nvr7
xVO8nMDxTrDnZ7OnnCuC0+qLQ8kYY2vQqhaw5nmRSK4+tLK/QCillRo/zVhVaN4U00lKZ59h9xzF
26OQsMxio6tQ7DP+jKXtMRIylTqJaFSBzYJRI5d6hJb2P10ltkQjhKrax+bhjwKu3cl+mXxZZ/Y/
blUhMh5pbmzwzGw6lFMGYMZ4wYXMjqJkyZ0FDXrS7jnxWQQm7Q6i6KA2JTJylWFpenCQVByihADa
yPQkNKCx8zvh3jSD2eOYRr/ex1rRb1Kp71SzYoazm4TanOmy/KvGvdftgEIabwjzCs2DgRNyBjun
6rO2MIdzkS4wCXueFNoEx4Ijz3ysXTD4u8NRFQMcS+LhLb8HIHp14BoPHdk7IsNhMJOXUXgsAThM
nJwpa0zotTGOFCHeosPJboa+9X606QmE9vqBd7UtU0lKSC2pqBHDX/wrK8bj/kpTW+znz5sw0ASq
CgeCL13Bc9LnVCbnlShsNfWaPvkye/FMF4niFkTcKnwMz51V//lIXxkX/jFsrDs4snc5vRwDALQ2
3ZWOkbQTlhrYkQGGbat1ubeZ5X3hSLsZQStCO8obDcYYDYdo9iKs2XjAXFBqLYLIKkRDBUGM614b
FllE4W/rHMHVeRw7e5SRjSUXXvmgZESFrbTQZvBVYNNPa6ZZ4qwOI/sKyqifZNbfo8gH6OiDXgLw
7W0cxsPTwy3/tGin/9fQduUE+unL1EqyMadGTQdBvISpkJFk4T67lvCOn42iv1MZgzHtQDg/3X5e
J2U84PS5ihXK69/oAHwKmubUPmjrHgdT1IS3i0nq6p0l/+SbbXxbinyiyby6PO/px9bPrXW6DTJa
3bUyvoC/0twK8u4WlccLQKNXVhpI0c0RHXFLxiVa1kaN8MPQqC5Pa96GbCTtIBxucJjO7AC/yTCy
VVC+rAgT+8pvHSbbFyC6YXl5lhLAVEM91r6e6eganBvDAg8vjrZK+35+3MdqArTBz095+x6K5/6y
3tJPLFBGBwIs3LysFdaIsIe1NqhQYPAxSkscehLvTsHeIm2h3WdC3JsWkjuplX/SCgPOiHhG1LjK
F0DXGSeXoa6pY/D7Oqa3C/W42rAoRAn97fmfkzKKVaVW9uLwpVSkhrcSFRV0jNtIWV1Ig6FRw5bS
GUbkUfQ4VGSj6zWGa7YDmEOKROZS0vgBLoLNtemIaAJbOuxUeUks7OtjnGiIuQBYulbBQX8N7KYW
j8lt+Y7dtF8xprUC0waDqWLVhUIoiRl/8PUXDVC5MK/fmhWeee5vqHUlhzKq79oUsYemuSY9jVYY
NTsnAFiA5zfTxSl36C5koI0eFVZralOvpwSM1zuZjQXyamVyT4CPlOI5nfc6TrvSN8AtP9tWjaiw
gQtX68otv4DZntRZth4RX71DIEXrX8o9P45E27V6UgPbV1oppzo4+csEpodoGMEzHt2pySsZRgPo
LNMCA+yCj7TAMeXMLHIvI7ZwE8otC2mwH+3A1pqxt8gFGJwiJkfwHTDC8ujPhTR4YGjxHNHf99MP
GijLc1yra4uU71hqHx2Roul/SPWUkLGweEZ9svgjDBJopUAG+nPQAaaTyPZcPgXYK22KMwsr40kC
PR13mts7UTcr0Hnd3skMwIOC0TPr+DR/nKBaS+uhSiVbsq4C6OifVAdp2EJL+WHUPI12PfdgCqrE
d5jccHYM07AHDcp/qBR+CoZLPaPw23unX0Ojb50q7dt1hqdqXD7XIyE8Af26WvO14Mwe/O2JXm0j
5zcEvoHBjZp/C/5SDysOT0TSl/Jao20J7Wi30Qkggf25zUg9F603ikRe5L4JGfzEu56Sw9pFPLFy
FCzuef9RDxHWc6FHXhrVyhHVDfwylGrCyondbC62TgLl5TR3gk5XpwJR5u8om784ZqZ5vvNMr3v7
HveWSeiIKAsggCQ9aLvQI/TfO5lPBiNIGPPYah+A0NApwfrTT/MM05lHLYGPtiF9VbWsyPLCd7gl
rhA4dXn1Xi2T6l7K1/g9TxEMqfsl3r9dLum0ZqGR+zuHNHQgq1K6QvtXcipr2dAANGJzTEURUvHJ
yh21Y5Bblyl0glaqSCePfBqomuDTRSvWhdJWB7TpPS4+r9B7nHjpYhwg/bbdrwZf/uZzywNy8lBt
C1eMej7awjevXd2BVsGQFdpbYQ6RMLqTKFYAD25Y+V80AyM8ZMPow1b/ezPC63h3+1CJZcshtnkQ
2nqCoDYEittGmpnrZhC5gwc8AcMdivZU8dBaJtd54T+FCAn4wOfqGA5p3p1yA6wPfZWLSuGKtxp9
gezGkt5MRa1qyqHfM68Oup1gz9eaXTK8/BGQWpeOq9Uo6UzZafns4KvZOuD4EASJyztgynklUlJc
mNDM3IvkjUAEjnzWLPtspnjHbkCCzEhSG5yVyEMYbcVaehc/xTNq32dXR+aNSfMjSeiXLL5j8obl
vGxwGnUAMdz/msCzM46odaO6ncKy2gis1q0oRBCY4gn4v/YYV/Ev721DhphjdjtPdEFlBcn7sZky
rx/XOHTgPbadpi1DV/9C9HOLIErKhODjXLjEu26+bkBcIxbuusfi+e3SD82zIEqFA0UlA0IMsV/0
KRt/EBrF/BBr3XmrZ9P4xoEzv8TyPZMAmwM83+wwKWf1+BweTS4QLTX9QvLkm2tEprtRLncglIUl
sqUyl+iBsDpuQcaykyOdEHN9t41E1CxCeTfi8fg595YSyOFllmU/Wmwjynxlt5sC+qXV747he+vI
vSwz9HVxQ3iccxuwGVRSBMdo3bbkUSZhRIzOnQ3cL8CxmunSrDLLfFTRa9s5GZGI7t958F87VWil
r7+rpucxn7T4T13fcN5LtnLcsPn7Ab8jwgjz2vnaAddmmJPGDXHyUdCeXr9NyskrtGL78V5io3Yz
UCKtpdZTB5kX+BZ8a5k5DvXmX9kyGeztsfoafg588Nr0LNoAOrrppJ4EPpiezT5rSThOcoxf1fiL
XOckCeho+L5yFI6AJZYvspWVLu9yviTedUiQpCSiljJQ4kt4+XNb4nNainEJYzB66Tg1jnfkXFr5
Ut34mLa21p+prOOltDmRNFmdHqyJfuyd5hekK9T0r9gR7f81VorakiMIiS+rVHPeZIXvFnVgZ5ea
DOZr1n4/3LZ/cxLUhOFHAuwFzce0HejWJYuUBtcD8fq/H0DpObIWDSLfrIMRlyUucfYLY/8QfsJi
cRj0Qjiv6/nVwTEKNYvtUPh0qa87/dXNvdIfEQziZDzLIjdwpa8h+HPimFfaVDzJrK+ya/iWzztw
+Ve9s1ZmsGSPaCKYL1npd22qIeupaza8n6z244hKjuV8JELNyH8RRnySDoi8ux592QOzqcAMvVNE
hCRDfbF8i38lk7M/dQKTWDyzlS9h2KisObEf/x9hhtaSiWvY9LYnLBcqOFifPIOLp5xy3YPx3Fnj
NSxgAsSXGo4UUf18GMCq7Zl1fBrkm6KR+DHdhzErirp5ziXytKm64bvKQDKlSoew8V4mfz8l+V3B
aMFyZCftOJC3ydelhmRpg0Y+9vmtbTFHZ9E88Wk2U1k15nMFJpbNQKbxRPTnYoMr0hLdppMuajdf
nhqJB6gVploq/7dix+g1xL+pQiqFGOVLzhXO7TG8r+hy1kNeAMIAIM7dfREdwzpf8NqWr7lgY5DN
GNyWsvIJWEGpKSnurTh8ACm9Vnbt4PFnmEyrDSh+1XuDQxfUANdhfIEjtacum1O5AWE3Y0+sajFS
GVib3nMBHA7aaXRi1LV/SoRk96sA4wshCpjRcdvUpBplmHqPvF5UmFBQvjakbYmeIg/3FgY6nAOf
wxwsDOEMXcpae5pQm36MjNdYnTbVUnPuxnFaQfoFmwKRPU9zN+mWgBBQ+iApatUgFR1CuKKgMRd9
VbGxEbDW7xWBub0X8IOvmkWnnLmTBuV6dCqanKr09eDPrdwQVmTbCl0h2xBUu9S2p6AbhSVfE9q9
ceZdEYzXXYlttRyOU3Padsf6Fik/DnYpJWJ1BHW69PpwbS3H5BMZ99e8sw6xJ+FNham8DUZY05Ar
24zgjqPCkTGp/OYZHJas1KPH83YCxde+gDiXmAXPnZXc0+1gW4Ehi9BUWLJIuZX53/85JNCfuwR/
p9uGjv4XHEZVmF0cYPPuJL3f9VtDPd7ncDEcNbyEHcdL+SBy/lRbweG2db80k4ZbvoG41Sn0VuYT
e74MAJBcK6hZ5H4ypCzDCqfQPOVckmXObf6oAcubuLw7sGL6iW1e4uIAniUAnZxvd7JK1TgeVdMS
gtKEA4hMndz3cPdZnQfjd+86HwL2+IUG23SsEBXRd8gbrifqwh2GMpEqYOodMcJAni1AiVmPKoR9
4yTKAoFGjRswbCpW1IWSLKWD3MXbS2O506nTMj+fMQ7QN/L+Ur7OuyyvEDCsDz3WaN7rwoA4qpQe
YhKMv9ymxuJInsox3Vah20UwejRzmoA0F57/TlUGTbKAzepEt5jOxQ+QQy1U9M6ZE3kFGy/Zw49m
+0jVileXUul5SoXSDNxTijmZElev5NalcWDDGhIopUZY7ujYQB6OEIxw/ny20778AHb6YjbTRRdM
i30Ms5HZarddFdzR67nd4/onNeasz+mi8HlY54eFOgHiq0Lgu1IfAUoM8DQsjMsJBx7KKXhaiGaf
3wUIATMHgsJ04gtYTQtCG0d95GDIfCTeY/VisbOFFL19TiAsBaLZYbwmLQXHnQzdxezdkjAE422r
rUHSXqG//iRK7rWlVVaV9P6oMU0SJ3TIXC2hL7Y6rIvERKVvVN9t5+rlDSI8TgqnuZYHFgpt+7C6
aIjziOgmMDnbdTm7rqkSW+7OtvextapLlWfrEza3nxUTqygAJ7hnMYhVZtSoe61NqlMeZxur4QlE
nWxJzCrABoxUJC/x2wMnnM8zvgPjYvI+DDPoe3FvDRaMIPrTmR/rb2wn3sCq7ooAqy8WwNf91MYM
5X1GS4dHTfBc3kq1kM0XAwQ6oxpw921tEL8pSoLDHRghTGD35AVMfCGUpeP4ve80SrJCivJ1Naau
lJgwz6cI4qRKEJ+URkkiogElWXKcRDy8lArBpfSeDWIyzXi4EK5Q7rMg/5Uv3zN7Oyq7hFvHjX6J
Fzb1u5g9THENAQRhiuPLq+P329iECLwxd6eBj1AeosNNU/CA20P0vpkzRLhry53w42SSgVpdkGvh
cQg5ri+lPJ0vj3wxQyKXjwCt+LvPfNYeT5XpOHUwauU2vhebIwdKPUAAPMjMJi2qT6pkHn9p5yL/
5DosKgLy4am90FbjoJeOcbyc/C6easfdJ6hs0Jw3qwGK7A2GKjbq2SWDTciTXMf9Ptw0NLdaRhLb
fdYIn0xuYlui2lrr5Tu0cERIY//1vwzHgb0LlzjkY9rcj5NL6lZfPqVNMmATENZ+kbQONE23ZpHy
dTiwCHGwH/pJMd89wJJlsc1ZG0QtSnb91ZehMc/YVdfB1fDumM7MB618bff2Jn0IZWn+WTpqT0sY
e48OwoaeHIUuDgM7sRK9nFgVuBtYnqleYxjeK92So1GKiE+SucMI55nVSS9IPWAuO9K7amyNDS2A
GJehVXh/1WlE91L/ufGFchnt5ySuxWu7UWeHC+iYRHi9U4e6OcCztGrdj06kiJBPgEZTzWLZKx0n
JIQ62Aaj6XgX0/QfnioOA0DLNRM2T9RWsefHrDfznfTw2yC0+LhaOBRLCpOvIJNfGLOKAlJx2cpc
3k0Z1UnUCDLA8AF6kgDfhHD9IKLrSmQSi9aRLlcqCJmuHanTiiBrUhY4miitZ1sjvOweh6AEw5Jp
rClksz7TVZCtW3uUrwUypOtTAuwRLPBgHoIL25q1uuypp1dHRZrIcDjePS1Qdc2Wknm14lFpwN6P
4mARuyKpYVrPv6MVrMj200OALL8cRQZnEv1y4QcRiKZnJz75+7k7FQl4KytacQLqBubGauvpzXrg
jDdZz8A1qvpKsbeMGAlgGBWRV3yCPPvtV3zG97jjiNsZh8Sikq0oyh7WoVtTtl4xMkdAqgd3mwjd
PnNmxYuHtgGpE7HacpZIY8Xz9BLXjjTPKV6qZrSWJ0y9yL+mpOxozBskATcRiYZQ1/3b/IgZ1/fI
vPJt0VsCOzbE2I42KHuVqlaV1aRuEpPSvY3nmo1zylZfVO2aZZXlFRD7QlzT8/vvq10eYnGg1p08
fq2jfbcUbpTFurECi3MUejxlsYJMXQS9P29/93Xw6lgMuQfR3X749lzdTcpBPS1vu/25GX/WQgDr
3O7Mk/3kYuVtP0MnOoz1sT/ff1gfP14wNET+5CSiWIlwHwNO1R/mLAopaf1LYPB5P2g89Mk+KUE5
OUVQfLh542R7KFlZzfwDlQ31rVpUtCqbbP6nIdzIyYt+Mgqr4ixarEeNaBnKV0A/fKi76tkFmASY
FCi9n/g1aMvpaqGFvd6UU6WwbfCX8PpPabiUaZsDYLrqQaEP30dqEbVwgtxtx3uf7cepqK5AZSrQ
/LdX/8cZWeDoaiOJkNUv7Ml19R34wh3AgUMKPg1HLxTKXyzA145qgXyLVl2deuf2rB4KCubZ3zk3
EbPwEnRdLL4SFVNu49to3RPYfttR3ZaYt78zY83BMiG1lR3WM4ZSUYUO1m3v35lTCDZwnGbRzqTj
sqJnIs3D3WnPgeUSaIaFnGg8vK/opnmW9uMSTpPc9xNyf1a9yoR2ZeSrS2zjM7nzhiGPBSfWvMRF
i4ALt6WZqVp/7NRrDFBqjlwH0LtXEr1DM4wNLevI3gvkGwcrmmPNW4u5SSMNZ7DRQjVLnB7a/QMJ
VUANIq5fhY/VQCcRvRyH2s8NfZGZa1rDxdIPIz7m8TvLl041nQY6A33IBU5O2isO6q3iH3AM7chX
nL/Jcrrngq2EOnwlmQybXk9f4rE5Ra65hvULxE4kmk3UzRy/oNjHogHVTi9Km5vfSN26t028ZVSY
eG524V0+qOhDUAJrGyfUpbv9NohTL0h6te2txh9wZg98OV5pjLluDZhlIl2AeLn0pVXaiV/HCR/y
C9MQ0DdVx5uFVsPR4qXwHfRmvM5uAOaSk+4ak6FKxmig5caoPpBOuCoOi9XIvQAiSywfDAn1AkHh
AzPJRvovjrm6C0O5lFQQcD+EJmSvR22OCSVc6Znwh0rzhka/bNhx5C5KZ6dX2H3S/QIwkC/+rwkU
YX1McWEdv1FVrYVdLNlI3ZD+lUP9nGzJI5I7Ofv1c2c1YrFpYKzox8pIyxgRdjgYlUy6lUBCqYMk
7YhKuQj4TftuINnRdxc2IydFlY7upG2AUhcbPVM3gFd/FxyeuipNRcu03sAHjBOkMLshnDZjpOi7
D7OT2SXCKJdVTF8fCpJ9negFYNlHnTmFP+y741DADuhRC53nu5dcBji1saudSDckoV2TPHEY5KSn
/wwhB6LsgVjgx+b50gD96iOOanz3bX1pKtgymMqVgIpyCJ041tNp1KTdZHGHIzDrlqoH2I80e/IF
8jx6rQ5ppmUaWVUxqb8yRbTGxMzF+gGkpky8KrTsOSWuOTcsqscgGpBSOhTuRgcZuKBUs/1YfOEC
w9dijzeBJgEwElft6beDd8grQseJxOj0nLMzShUIb+8j+JwtbFwMSG9bzkuqQgOD+6skDLwW1X6F
SwyvW1p//RRVqcFLfqa51BjUx6PfsErHDT/AnELlqhaqCS9Oo79zhqbUj4BOPMYf/B/1lmP1TYXb
RLA7U6nB1m0o3myJ2I+JaMVIU0JJI0V/6AmHED87XxwUg4DzZN9GkYHVb8eZbAPUgv8maWz+D6WJ
GBY8FoOC7jaLyTAGnNIjjoOi2DeBbYihMB2q8tM/vbLds2d/dvgXVZk0FbPP4UIQTshv9ABsqJnU
aHnFHRidP9/98chy0IAp5+OBJyU+52mG73MZ2ylU/4fQHNBBiOZQUmmJpRWRtHnPdIYb/YZYjmru
/TN8mFo0BqxeBse8CikJLSMtIj0t8lwJvkyjeYJ0pcLX9tCKrnPwKzZ/OtxUZgFIRgQvvwoIKrRp
diGSJazt5uCS5f3ZH9Q2GA5PNM6meNMMQSMLZtcF5kfeWE7TiCRsLddLfXqnVAkZ5TKIN6lmcmkt
N6TZTk4NVYDZSqKPT85PNv4OANh6f6IsjIRrFLoC4SjFyiwn57HfHxOahQBTqnzHPtiMzvqQtSri
jkSjcx3dZ8l+8YGD6ub5MoWHDrFFse4L+fcKv47o/n4EK0eegq7hKps3WoZ1qdaGvvi0MI33sgpo
Zkt0jJRVRfc9rsLiPTi1u9sgMYpEzxXG99BgkzGevH2lyqye5FnemJy2G8MbNd+cZOaecb5EomDT
5ST/bZP8j4HBIg85RXxx9jkW6qzLveWy58PjPHZVCG7xBqrg4qH82SbjIygzSBz4PX13dFWWm2MU
9M+hXmsnkijd3Q9398PtpFHpnIuljUdg6CLJL9JOMnTVhE791+GB8YkYzKBPbXIylqQySWKmkTuw
eHZOphz1duT6pzJnWDkzgScuPl2Ziva/mYWAYGlBcv2vuVWFaHstDJdG3DsAhTwM3CKSPFuGyjmi
NO4jdH7ktfp3eYVh2td1LZnHgp3XQ2+egoXXlT1bu8olB58C5vnOOVrYDDMSurvCGk6CMiAY3kdy
7xzhVBOCkt0AiWArVwD3Q9LyJn80GLUieiOsbB5R5B89a8BaMZju4FdXsP9l8dsndLsuuoAbLYCA
tztLtmFqJzznQR2Fu+ckhgBKw8DLgh7+Zxr32sLc2bBWerROWdqsIgoA6P58NY+xCvquFJ4yvpLd
YBLwgbg1l3ODTqO1i7sheOrZarYmmUFgB5mwFxrO9cqnPiqSqtn7p+weyzD/avTCfSQZGRsj7rAd
lI0KPigy25dJ5SF/IaxpjRSOp7dvRPG+yHlc4yImyzM3DfjW2ZUvcsc2CGfBQ8zuGwDU+tJGedVC
5AQow54k3zT7c7cIniEZLUahTgXWoQOO3GOt1D02Jf6OaQjp0edgGdhQAFjZVSRaMveQN+CeZTgI
0/+8VylXV5P6bgOxDxzY0ghjbKwvTgitK7juTV/nrcyKhu4tZTDK1ONAx+WblCPS3Y8Ehuu14SVV
zJfSJpuwTWrXlRIKQJzCuyrxtyMfpIlR4jNKB/hgoJheeCLRUckDpr+zHBst4rI7K4NIHLpi/Ldb
OQu4+iH41t0fDgYuNGYm0Z0AmjoZdjE5dxQ6+GtxkNGJ20uDaU3i5YhdAeKWxCUnVxFEuAUKmn0c
J9OY3DTFIO5GY1iKNp11hfEuWR+5DfbirE8lZPTIoXcyPFRZRX5q07IngqoP2imEIF7Tsrf7qP2I
qJ2bOXEK9wzZmAfaivFunnz978alEBeqz233tVQ+95zmx35LqHQt1QQLQdzFox3LbHrOSk0MyJ47
lQZOZxaAb84d0LAcrTCdAF7gMOc0uXsbDp/9/wPakRUgFHRfBaFRGORz1RUD6jHhe7QPS5+AjBSo
IKG+z/6QcPRIYK98/oVAjSMAmS7dp6MvXfUq0mxqwXl7IJk1tAg/cTcDKCN60yhF6zsl5oOoPwrl
vK6lt3aRhpaXYP0ZsH8HiHQQyfgDPN/N/lpR35Wk4kBua58Dz0zLhN4mdTyQ82yelx0CCxX+IHjQ
/oYXRZ0OwSZ1s8+A4mR0tyVRCbdVl9L+GXMX2UiYYkmPY+WBnAPqLGVwNTkQ/yY0IzUj9LZ9jbXQ
Yex3JbMmJ54JRfMC/iZkzqr//dWwU/7cfhDu5jVFdj1wB4NbTRGoWfR5bFv2p8kOpOGhRi63LHc3
L8OJW0D7wwMIEezZicXefZTowLxgLGi2kpz8MmuOTfxbKxg45fRvo2a+GKo4ao+vOrdgjZZ9yfLC
PBbV168KQGBsFLb7G7CAdz8C07CdcLdA0PxfFSgGhCY8bmxg0RibnwPLorzCD2OC29F2g5ky5Ay0
yQUrJ8lnSEOnedvSXJ/x5nlh6TR7drbY/7r51xFlwy56QvkITuvhKHM6QX9fgwv6xFL+IecZ8Gpd
g2U/Xpz8trn8Ng8nLXM8wOX5Ceae7GzVWNyRluz8WJR9wyvRUU10KOb4uKYSaitBtFiVZpoDSVnY
F44F9/aXsoUeKJlLyETJUFDINydEwxMsOxamaU2MORXW5louTx06pubfZv65fa8grtQlMN40r9UP
9oODfwm1fyXnYdOqJ0WDMwexGQqOWh7JAun4CYSd4YcrofVo/4TyWyz5ImAel+rSudxp2FA50QzM
ZD2A0vXowxoIHFLJ/Jr1MIaqQXS4wO+UDV9ySCe1d4PUssSvhmWCdhJc1P8iyf4DB49cl9FuodRH
WkMU1hL+Ya9ywRnn76NYqrYqVgr+zXq3T+dIJSBeoaTwshrPF7dwKlsPLEnAJI6h06Z8lozuy6YY
EGPl54lmolvhjTFwaFyOLywoG/6m82pdmL0zRzI20SjQ6pwIHXfLiz0r4+ra/5espvYrPAuIYZIz
6gRa0xfhkZlpJrUJaTkkwd5qyUcxH/5APgDBB3buGetM2SQlZRr6s3jRuV+GJRawAl6vWYXpZxoU
iVIU57Bd5Mv25s+kGKX5XTfaBz/hScJs2da7JmEFJym8CmSuEYHVOYJqE93T4ClWe9WIJWwpF+3A
2mFa0Ri5t2L8OouepMo9/6F66iNiUvdDEQnIZUNKDZSHveieds/Sbcfb6XeWNM7fAQCGL4TMLn7t
98iVdw0zNfBfdW8cAKfNf0k+1gPL9PrsYOmXmqu/sP0pEs2yHLQo5la7aISzKqNgrHvQfvW7daku
SGgiWz6TfZjAWd0KrdFRFdcVdu7UnclaNSOxVY8/6q5OMjCJr7O5AkrpKYxCfHXprGwom+N1GDuu
e7UgCelcROfBmbfbivyHiv1hgyX6hwr14GjiXH2bhD8znIazQvz35zL+hPQoqjYQjgrY1tN/7zp7
p3e6eHwk//bDoktoBStQc1uXNZSE0MqsCRH/O5Ou3SuDq0dwrEkX2W5G7TQ6p6AppLIF/QwwXhK4
xvpj+o9QLOtLoJ6jRxO1FkhvJ4qry72OjlDL+DSUO29sVfT8sABkFzTV4eR3Ugxx9J1P4p2EM9Pr
k6sYl1VNxljdREsStCFWQDxxfqChkUVoXIECJqvwH/T9Ngx1mnB1qUpfCvrE05lxgEt+VEdI2g6V
r60eYFTS8rnABVtwzIQvCxuXSWZBenrHW1LnpkC65yrnBKdLnjDH9PJkz8sorcsfSPzqUx19Zia5
q6FIMNjWEQ3OZ4VetlnBSz/1ep5tGoHrhzM10W6E5i2/7cVe4BCGwX9uEE2JWAexOJ6iyvwPzhpe
EFCO+RVmJR62gugZ9qN8W9/Zum+jle8Ytff/3bshR6rXZhoOWzQ8QIzutInpBl0Exde1x5Rnw3Y7
as3Th6fughrpUCacx826BjXJEZVxI5wHt4bA7kwnahG+9TrNW/nHyX/0Tc7NACmOumeo03+dGPw2
jlXHj1YGGzjqD8epzLw8S97F9RBXV/kAk+UwkPIxWF6d+qH26jhcCueV3DcCIlTRUYyaUVOSHZ/d
L05A+Dk7zDjPCMDZBbffswdo+U31EdZXqWq1Ff53451cBWYPfMhOJq5y5OX21i9+x7WnMQlgjjhl
9RI6Z3ciu8vaIhdUXwVpiLBrqJmT0Q7RBzZ+/Kiqpw1RplUnxGymaCq2vzCzI6a4trcXEaMiff5c
AsG7pux6+qAZHiY2L2x1lc7OkAWy74O+lOpVJ//VrA3PyzTRVMYVU/mNH7H/fEE0E9K+wWiGxNGK
osO0QDeC9UzI1bhYQFRe/vg4e3FrLYl173nOi4vikn6bbzjK5emkr0pvuL3E0svTvQ00yruXSTCT
q9HZU+OPmdqa7Sb44EQp24HBISvcb2tuuCUoF5mrhOIuZEwB+IRwwFDOI9vzrfJOztQSYQdWo8f+
49SfxDLAs4b0EK0i8uoockDExGosWWmqhKjs0Da6LX30399NUznLBGBQzhACDW8YYqaacSy5UwRX
ItgkPD0qjXIN452S/YWa0v2PfKEnJceRXkQrWER1OWSsPvQCXrhJd2rKO3fNuLjiPEkJbPVlZD3+
TTs5XcFcfXZiwdz2CyDOmE1s3r5PznBuEaWKwT66VHpE03SPen9ifhQhTiJSoYWCT+82bacGxOxl
u6jB020Dn/Y0h3ZbfQs7VT3nY/mbwV2G4rc9w8KVzpWpBUHL4sImY/ATJ4Q40b6movT5oH9VkpSz
zGeU4H7A/Cy2EsBk0tEOpMouWuU6iZDgpPGn7o0l6aVcvnBlvM9K0dng6CXFNeMsGu5vMuCiQyN/
3QaEfct6KU9R0y4Qnft92VAdj6+euTfyBVixR/c0lhBz1HkcsNjK6D2hV3iRb7yUdn5sXXBzJVEX
F41zRF+A5S82ZY/SIisVSrCD1I1hWauDCKAAQq3KERC0YWincWUoVeZUXexxsH+GyT6/IPqS1E0g
+LLCYuR3uvz/an/sarBU3VRsNZ2g/mmfPYKsXInGcdRvuMOW2+LOFsO9VVMcgVXRDSaR1BinMHMj
TFEVcjc2JvI421Br8fLRgvXkcn7POZEx4xiu7aS9wpf3DS6tVwyS4M4CxcRvbXqz/hrI4y3Xc6Sy
VLZkgTwwOSd06IDVUnIzUTf3ZFD6VhTRvbkXF//VY8hQjAXSCrHf8D5+Vz5a/o/v/H0252zFJk1K
CHADM719h7dEGsDjvNHaznkn004YxBREA5XM0kZdRlGUBPcMuBhRXMmXCrTDQ0XO6BTtcVggjS3p
9M4iMkGD7nlBXyVcFtrnl+HT3D0FfXACkdza4TCOMzH8P/RJtq4I7HT4iYARRHMU4LmIu2WLxVok
atdXAPsrCJ8yvwiSYDERVYM5ityOHtJRBIxGGbuTw/Dp5um113eKFpnz3jPaRKB923OWOBFOmYof
+wADwy5J2FTa2JSsPbRXnMpnHKvcEL6dz+4sj2OSPhq+t/pIpzCgM+rMxaVD7F/xi63JtrXLay/v
xm9ZV2VPm4uOG8F8zk6MJmsznyTLcDIelbxZTvTZ3XM6GkUpS4GhRArfKCfv4SSxzqEfIg625W1z
eQnp2O7193ZIbNUuKtijVoDHnkeU8vAu2s0EhR0e4Ga4puhJYHgA4xYnBiaa/YZOWIihGRCHSqLu
kuMtgBT8X8aCWxufTL92b+wxPgztTzGMmooFjSs9k8YqjSaBb+gjpafxYM2kdsimIgyimXnqxl8V
ao8hAGXmAhL4Lyah7giV/xCwocVyvypYPjJFm+dhpC57D18YszNDqZ2oHqDalVylE4jUs/XwvGDo
STOnoo7Za6peeLZVfH3MFGSjKend2C0k4CWTS/m/hxXrYZdCyFgpywtfdM3fI2iRmk8kxFbHLYAy
jA56ZbqlEg3rW0kmkkmlf9phzTn7W/YvxyPZrzk2rkPpItSTCwiSfH9x1vLzDokT6fwzky5mO8w0
VGvuc7noHaCWF/vbb5Wt97z5VG6Uz1Z2KDaFTswlHuSDkcHqGq4DLTd3Ffzdv8N2798Z+X7qfN9P
Jse0F5dlv+affO5NFOXo8AO2kVwA2I9xrH02hNMyHhBSVF5yfhjO37JyXwqmgMy75VxPnm+jdVkA
hkwx+2SFzlm31DC/yvLGyMuVfuAgVpLk2McJPnBcLRe8DxdlEuxS648/Aum5N7kdg8LhkwhV70KR
Qskkilx6KAs5VNDgn+87g7Wdhq0D2bU47nOhFnY6POs1xWrSgkFtaD6mqR7jYpu+Fmg3gPktegID
LiGK/zlXwa+3Cov5XfIrzuErI25AiHUU5kKdm/CY7AKdYi+EltS0BHGSg947A5EsuC41qFxzuV16
/Np7VNCRU84Go9PaAIlaCB6gnFpE7rMVAPDt946bK1Qok11UZzML6JsCN0PMHrb6kcme6IjsNkjo
AtFGj6B+Y9QigoqgEhRKTj45RrrP8lCqdoyXrkdq6ODa0WGOU1hVO1lJK8myWvy1y5jThO5xv2Jt
HjHn3mXR3KANqNvR2P2yEqVrSJZ3C15xmAfnFQgXK3UDaalMuJZ0Y4OZvVZ2ErtyKzTZpPkvMG0R
7CEojJzIOEkIxcAUZ5kFO/dlWqmiH4LgncxSWYyC4KKzZyHZUK5IGed/ylKlyl0sUc94hYF2bCWJ
Tjt/sziQNd/OirlaSatE2t+uLvn37O6ZP623svu1nx7NS+3utjkIcAB9i0TVmzhRKi04MLhwZupA
H9PDfEI3yPIJJNmHwzoneBmwJdR6WarM05eq9/ea16nQRRrl9luLoqmqlnVenF6C9pgrfmBkzSR2
6Y6vF7oRznFly3r8tsAOMMnyYUfAk7pmFjEdOmQTh9cevSDFLpfIUX/RooldDtGbYjkEwt+ne5Ec
8UzNmk5dcXlSLIHMdFhmMFZU4Q0bStVeyqUFKV98tZIouLyf7BI0Nwu6zJAvOmstl92d8QKY+xir
QnUlK55eNzrI4qIpDM0CDcUQ3pHBp3VybRSecb3MZzzIOce4Z9e2zWoC9KoeEnim9JNfkil/ctrh
CYsk8qcpIBUr5OipwEc+tan+JAVZ0d0nN7uOAm1r1rooVljiCoagMlgeC2dxWNfWEpOncXXhurLA
YRnmv6NqNXXH0AnQePpJNO/gaeeZSciaS1szricb3rV9PYvvy3jRFBsqoNtqlCEoFXHzgK/7EFj6
zzUxMe14e26+anTGQ+U7f30F6OBHIvnqUHofCxQAnpsvpxtpoiKeQp9EYbP5NXqMYiOTgUYbusX1
MME0VznV9PCSDOWhNHDGNBIR8eFNSHVp+LRc3hNoBDC0wJeSGJeb3ZOo5gg/Vb+7OAf64/jPcZ0N
QnDav/Wf8/xLg9gfjLByxfMvGuQdVfgB5k37ci1keG+4dl5fUygb2XGOU9ZcEhzLVbVuYwu28MXd
8UHLj21iucY2g9qEyAtsU/nbfhL+pmU0e0cejveQWa8ZxklryeoCpd66TNxbUHdhLBxeGgkeAfg+
1WXdtVyomlueombus2h338GRmP/x7/E78soJoVDuWstQ5h40cYnlAlBoUaFw1LxZToALK+qnF5BO
joLxiHDMXcLTIdMcANs5koCAUrlz2bLOdPCRnWHiUvdvG+kHKbnVonX67Jwr0BYdZyVPbo6/8UFU
znBAxgFkm3L+WIpEtb44NkJSI8F+viN/6w6F/jfeBa49TnHcyXRrltetf5sbRDGRgqTghk34MgQs
TvXcJWAsmwEdGZ3j8GsS3tnWdhejR457CrR+FjfBKPcwwCcpMEG7rImJ2bEwa1t2hjo8XwpGvgtv
sBWr0S1w3hnTtrA92QtHM192JLcVZcxJPo1EBTYN8q+D/17Tc5NMJbIRUYP1xz0OuImaUzD1Hxfg
h8JSud3nxlRtQRzPZ/Yai0l4rTdA+5Vkyom+LO0gRGwpIyfmnro3wmWaCbzw9VzcHDw6qrRJOlVU
AabJ9fVKeOmYqhVwF83fU0Y3fZ0ta5wwW02YldrSU4ITcrneCiNEL5cwTWDck0At1f0qtYKlRAdJ
4GV/1w6CT7jSIzNBBSAYwLsEicyt1ZC/1TkG7X9hDP6r1hiQN+5RaqUwEPKvJnfrW/Kd9wz86cNB
ihCBULz+B71dKJLdhdO+vQ76lBnweTvP3+rzpgx781NIybd5ftK6WRYcMfTfZQeYQtmEq0YXC/Zm
WQQwhj6/YOWadHGUg1QFjczMlq2g0+yE2wHc5B/NSigo7qLzrn53mJridXjNWKimJPaizKfpGncw
doYedERN18oyfJk0fSC+/kpBO9fQjc6ft4JuryE6jb4cgfO81SvhAP2KuQ67e52RlhW4oa6W3qyQ
Suq8lobGcIYjkcbiZb9zKAoK2S04H7jH2Ca0kP6Ns1565AhIk1BJ/X3rpWgeEKvN6oJnX0r/nTzL
TpQIodEIzf53O3zQ8/HMRGs8RjZUqI9W21T5yB1G8SVq35LP/63BoYxmruA4xUdFAHHyo8GEQIPH
QNZA425tf1IhlaiahjSeBJhbAVdKBlNddr//9U3AFUEjOjDGo7comO5uExDG7+fC/uParMXY1BZ7
jZ8aqOF4Ui4JueRZMQeL5ZDAckQQY7MQ2PnvqiEfPDnjfJMt/jH0yA7V1a6hmmgoCRkZFGP2LdjR
B+pjXXN/jMV3jW3hX+sQvlXmcjTh1E4wV4WqG+NNrExK8B8ueAuiaAk39N1c97KMACQBCHjpEzZF
Fyxnk1Ap6Ip1Hpqdya7avjSyYnw3NKm9JkPq0ZXp8SJ5weZt/GrRIhcZnhian4zEbgr8y9yyr/Ea
jtSlWWohNmkbdDH426EusiO75BtdxjGLyF5M7yIOAvPzcCM+E54ugDUwYWDrzSNwC6qqKU8qrbWO
yrNhQOvUkWN9V5GaIFjKqTc3+0D6Ot4yySMKkyKEGCARD3fbfuVGtr5aOZAd4J5wT2VZ3Im0P2yt
TdCdLYR3kOgF7sDF/Mu4UcfEOzzvS5xKHTIJnG80gxKYs3S3lQDZEq4/4t7949A/VPahpK0DxcpR
Er0H+jPAUEShlx7c3jjV9jKAZIqd2ys5b/6q6kLVaSE2GbIA4oZPeL3kAHi7ZqhCjdqdf1Ju358G
x5ZMrGSmyRd/9BH+ELuhHjz8JerGH1a+u7lRVey1wLlWIA+LxaLrMvgS/8JPm+Ugjd5Gc74pCZ4R
OV3uRQcFMhkAgwoF+sNIy/lIqptxebaJMyK1hAf/3WbraI+eMQRcaPLpS4tr7WTW2V5wuprLA52B
IYisRI16H49G4Vc4VGrIpG13JLYYtKkb40DuTvgR6wvFT7yxBoqbebqYMPPclGfsErOXMulm/8Dt
jtMOV1UvAm5ve56cCTkWtNU44p7tnTT5pLOFHngceqWuAO9JhUeBFQRbpBx+Z7lEzjs33khgg92n
/wcIE3sipieSU7do1iUR/neDFUaZT2pFtltQru4dFYtHrXfQkFElPxuankrBLE/MwDG0iXV7E9lQ
fvJ+jFx1GztKvJ7u+MF8qlFheP5AWoBUn+bsSAsDOA91fLSBBR77LXqZ01YVfSvqtWbXkbKU5hN1
+8GXm+0ZPIBGglJwrbMtrW1mbwWX962sUmGmPBlo08nvigqp6SmhSEnegpwG3cO+PfvJuQPe9Ds1
b6xUGA+5PYSZ6iE885juh4qAcw2BPYu8xdrTVuVXviGZGSU9yL36kqmnoDQ7bIZXn70nXGlRXx7H
Ox+chOs16zkXcDQjmtoXd1cKCpp2NkKDorNYzKEf3WnYVg+yAevIjY520mcpK0IqSCBaYW2oweTf
3A3e65cjF8cSY1x4gt2XLp/KV8QxDo/GSQ6c0PCN6mOF4fdslOAdYCVi67G2EGtUeqiX+ZRXDk97
KU4j3EWJ23yBrxCj80Jkg1slFPUvNCGv/bMKfSLcIxZZ3cMkxokymSUSq2rGd+fDS+ZmDp76Z3U7
CYirfrcIiNfR39XZfFs3PbbFmHy7w1Sh5O253GuAemuiqwVyo3JyB7LXyiKKFV3TflNjnrBwEpWw
kVaV7gxIlS06D86FyRYRgShsBbobn0no59IkUtP71gV6G+Dhzbj2jbIA9gvON8Fk8s8kxhBW8HLL
wp5rB+j0PbjTCzannRrUhSCaD/ee/PxEOBCeWM14OlHWbGQBhLFsWv5F+4dB673Sw8eJGkIAZhC4
uPWfOg2wvI/oNXtksbgPx605gofA/jpkgH0Sst6Pp0Xu+AuxKrCNCSOxBwp/TIcyLyrE+iICqb1K
khrs3Y2q4AB+ibkLelhvxN6P/jIjfM3kC7x0R5r7E/HNwDcIZRIGsTxCHcQp1DeJDPkvkodzOrMd
aYbLh4hyyBvKJ3ZtwRAO+d9tG+WNTs+n229S6V/j/w4yCFQ0E3xMdxIfU77wapT3FJZq1ZUSBDSu
7pwaO1fPrK7XtNvrtmqCPS3XDxao/UUt9OtgmPFC4vHv00AvYNkVW1g/kdpF7kSESR/j98BC0G69
rJ/oiFLNwBJExej9gueKx8BNzZFZwQeOXbfMZnMf0BTipnWy/FsRHx6E9LKNRN3j+Xg5ioMNhfQZ
iHTa4UcT6zVvgBJk0lygysew7hV4bBmarbPKk3N/gx0y6Jqh4nOCBsLrdHX75B8pKXX7q6oKdsEv
4TV28dkVPFeTviQRouJkltsiEzdH1Kq97bjOCTFhd1NE+r/rqsHgnIlDsFD1S3ygyxBUxHIqURO1
kh8QTMFOck+IB/o59P4ucEEHBHcGtkt/hynMsl+e8QKXVdRoICUqJcnhIOj+MAaT43rTv8kPDQt5
L+m/lvDKllb+BFpy6rbrQSD+4l3Uzggw3BfMm7SfetTHXPtVnb8rRGcGrUxKxnqatW/RMO8nBXHZ
A4UfNQB/OxCVodu5wSmnUWKXIqpvkNK5b4LBcaxUKMbpjclYe3CTtZaELEhbK9zh+hMtx+W0xlXq
qHgdHk2DxM6TXagbPjxtJF4BoMKkbrX0BwQJC+FvL3ngrRpXaF2H+oflH8woTrDuhwJLcm5S5V4b
tybnsJuGWhblh9ZrKEzEWZJ1vs2deo15reBtxmN1YW+HG8WT6oWeRJ3Ng28Qjh8IqJmPoOGSXY8T
S5OtazqDqKrq97YfdNTmzVfNgCpGzqOvgNtiNh0rI1AOvr05fb8H3Ko7hPMJpHuk2/C0jE1wja/v
tJLCWvbMGikuyYuSCpqYjt6NN5b/hZlonhKcuHamUrwxJTRGtnHP+Ms5YBG5IgxVEzizBwQJqrw6
1YKvBYyEQUK8P8wuWCRogtPIg4cPrZaIJqkfzU1T+qY6Zom+l0KJYyOVwaTHEDthC+RgmLxPrtrq
ls5EUSRIPLXqGBfyCPmqyhuR+2ei6mUR0DwLqYZvfrHCCRhBgAc140exky0h+QyJPyNf3qdxiQk/
1MYBKX4R32mlArqm9KK/RRxdLUrwkcVEG9GDGADHBEFH2niyWjlyFjwKGlvfEyoSCsV+SiYdIXVg
fwj0iKU8BzGP2274sCXxh4Ue/sDQPQfIAfO98nwCjKWde1dxv8cZc69rh2P7mn2FYPMhIHq1Pbd3
CpZSJOo+m/R0Zn0cdeS/jZkxh2W01taQs9U49sgxXvosGNGNKkh+4GQ8oHNAQZN6pyGvLtE0g3Yl
Rpn5yonCNt60yQbVwyjsISJrDFHdhsvUxaAi/bNmfqxwgkLEf3lqZb+Kp9A3OdT89QkUj30F4Zr2
Zsc0rEJiw9Pxn+qgXCrOdUKcq6hmC2T9U0hbZwdDYRgLINxMJ0DxSFOQ/LrGv1SVYGrp5lQ+16Cw
H7SXS6ZisrD4BahF/wpJTpeLfsl4RouOQ7usLCgwyKzTXLJQX/asddRL+mFqmFxqZKLaZZki7pc5
ea3O77RwrIOttda8XPHLLMFjASMWAOUYhhmeU/xraNdIXLa9OWkHJkNq5903UiBMTtaSDug7aQIS
0RWjnNCP4T0JRnmZ9mVi/v72RKS3t499cz84tuxKPKsQQljnl29ARqAZe87PvEouKwK6/ry6o/iw
tz1U6odrTrH/qguZEe6rvFXyQLYt+ETywQBZXNV/jyhzyGK2Uf8mlRSz2cCWpOS2J7O1zcyhlGZM
lQB028DJLkgFczeAgf6lzlOeW8Cjl3TtxC6PmKSbP61QvxrQHqc6p+EG2pbzdRYYZKAA06N8EIX9
m0IEAI/oelfJeEH73sO2FMk70r9rVq/63v5J0R5salB7qmevpVvSosfPIO8oJV4JjOFZ3g9W6doQ
hQv8dduG9HSEMsTx4uJdpecN1nGSJmDBatLEVUvWxbcWT9qmlvdhS8gKHpZXKEaer4jcTZ9OQl4m
6FCuEaLH6aKHZw/dVCLW1FD2r0o2jZFTxqLP9wEU3XhgXzPuVNCo8416wDAViPYqPEQzA5L0cUGI
fMWnyB2WSwh6aaapn5Iybh0yZwcpOLqkpHTuNr6hulowU9livcVTY+up2sCa+XgKQx2rvqXUPdaD
75CRV5jO/qWd35fyt24MD0VjBmvCgyvraUNoK/94D/LG30CnnDzr2VHIc1+8j55CXIvcsBSZNTMZ
LCd5Cet7sZrHQibiBq5DGmGV1DRWupT61b4UQZtyY2kCIgbngOsx6wP/SzpC3rohlNLLuDxtOUcW
AtjBMW6E7qoij5WTfl/qPE2m9Czb1kMHnHMVu9UFnGpyMORm0a46Hs44v7u1F/hgtYU6FC9hrgKJ
muP2Fc7a6TzoqRXuoLbA+EhGHWQh/WFkEzbWj+i0M5qtt4D1O4LHY5U26YlnpFZwX5+Vje1n6rwa
6uu7nnLTAT3tNwHejOzXfJAVX0RPYaPAWZDFfcNx3Dfr6PKYM3A3oaK4gp6MYOHCSUjtG7bZKHUS
u+u9+R+3taSUGtc8izPLqm2FDZotVSRQHElNGlx8BxHNxFVbs+IDuRnrBGOEPaGyrsunA40/hvxr
tf/1UrqSWXQklyriCbIdQQcEuwk4pcA5cvRgqP+SL1qMAy5Zk06+OQDig358d2q3PlLJs6XVqcPu
8abjkUK1XkeeBC0Eq03idezSXOywQuTORwkbX+9mWBWiB/Pz10bkgpb58R41dYQO7DeLYGyD0O4f
AzLZxE+7rhc4sjuDfssFcqmgs2ufbm96SfGtCcY6FYUxwY/k4NRSCcA1n3hrIldIZOYMp1PDjz6H
ij4ckRVgKzOc45k7mayQE547bmd5b5pKe/NAgHuEmI8wPHfwlfInGiTmPuEIsfAnCwZ5fVh1JkAp
SBa7RhR0eP88OFQFTNNct3SK2mmqVpy9xnLrogvqdB5l6l5i1zaIpKWLMOnIWVqt3LGHoh4J6CdS
HCxhAdYLViGEXbQtX/7gStO8s4Oels6BjB6pGLnAX7xb8NXgLSUygPf1qEczkkR0ZM1IZbPgydOB
qP+wxi8VzLao4Iy9ksGQimm2JFZc5HSjrFIwUwfyOCqOBmyVEZDU8dNqFsTVTDEdWwv1CUTsd/Ta
dfdqzUpCcZQ5BP1pW8w35WHZnT8nqC4YmEIya85bwi1VBX66v2KcwwWrL+FmkvO84ce+/moHTt4B
6xBEVu3RjxNXUQsEH3jdAz50QK6BqJsVmhhAo+oYgSCDcDoQEaEnwq6fpNyzVr8TPKCfPLi9w44Z
DM8NKBNDrGFBh9bC0DaW3uM3CutHczZvAOygXfmGbRn1hxK9kAPvniFsHQb8tfmQEviFYn6pLeb/
s5vILMfYfTTzJKz5gFDLRQQ0p4uBZO1hrqg5hRUCLNKA1LoFbNR2D8TSCPYIOEFbckIie0+QELAC
JDwTbRy3WtkCmdZ9DcPDvC75DmdcJdrDHYBRUm3QYwUE/oMRiRiCI2TZKjt3P/cmHvwQ7tfqF1Op
pF159NR5onz22eEC4vfe8Jgs6TmdnmpaUZaXkZcPcCDskX2/XYJ/HxhC7YpXE3sewFSEFDYXOdNk
qclvLd/mA3rNOnCFOowXFVGwK2O/sWh6PlLeflxY9dpgDnXWG6LrqRdVdIefBd4xFdtrvGDgNMQ2
BeA5+UmA6kgRLjXOytxhxueXz9m1THWAMCoMb/zszKfJEq1aMjjZZuP1g/3KpoY/gYtpEyaNM6NF
nYz9fHtqRPevMWYR4oii2LqeW2b3vTIM5k2Ubf8S9/pfrU8kdkaaz2Gjf/BLgM9nPvuugDMFjjkD
IPty8lPW56EGgu4QRpZh1p2I+QjfBcgnB+XpKAPX0QGyT2jGWKGvmxbtUMXWJ0nBFJButA679pVs
x4NXangCEcX2h0Tq2BluWDiC3n0REjhp7NCDRdNh79Vc0OQhWTyp3Q0qTn6KmPkuBH05vjKwm9Yp
YOWd1WlQQ+1cbFCC9T73FNBHWrCnb5cq5NPnWMcPOlaPiA94kfJI7wOlcQeqV9II5zaQ+qYi2/L6
ih8QBd2PScY/1eoD2scSPKjDh/c/+n5fm8/uchCdzl5YOwLCgo1lVPnCos60WFYx965I1uu+bdOZ
pEtyZYvDxBFsi3x/cfvgOi799z0IRhIMXFkoMP62mYloFicYgwePehML25CXbwC46cEYuDuNrKcZ
0Xtjzfnp0vYvb3TUVu0hHunj8KwkzQgXyugsFYHBBJ9iifUVYj93TwfEltxa7B2hRSB39x37voxm
qvLHA0JyoCy+afKwT06MYK+CWaXkgkn4AensKPDOMMJPkXE6Wgpmpbz+MOWhkgycAoGfdxg6/pfR
cw3BXXzjxlBAukUVza5ehHu/GsCSuN62FVql756j4r2geGnGA2OShLt6jNQucdJ26Ty5mkM6Z9dl
ctGb+J13UIaEckSrWDtPbhPTWjnqT4hpSC2HcPxOHhTUixXHkyZVsX3lTnltAskqEsn1oBxYU341
R3O7RyO9W619sT5Fie7yPtTkp2yfI4iG87VHqDBxaGfQToD88QIczSlsSJroFJwkJZ3Z4D078XQE
w5DP4EwKr4BcYUIdE+w/GEVKz+pSlndUuNsGMqheMxDUNEI/JYN5yMUYBGHAmhrX7QGA0VUFbU+A
E7EU2wpg3/NN/I4YSvoaSs/4nGbocvbSgHOKE0Cvd1vJVIrUPATWW4rv2q1CAWmMnO49wY1zpDMP
BCwnLCJLKonnORtRA8zkfwm0MuUGYvLKauVlejKgT+fbG4YIcSRCCp8CpqvFIiA0kytYt5DXvXw3
TseoT26Xg2n/TwzIpT8WqMJ3QpHTl7PblTTzx85jXYW4qczonKcmqiNenenx2xwSyPK4qBE+WyZ9
oFNVIv9aUmrfkyvg3qD5BRjk7nuZ/UE7H9nzVY6HIPYGdNT/eCPBvoGwRIoAoVQsVgA+pO1vlf3v
CEXspKL7iEHlOVxyReHucfkcBY3y+imu4UADLSLBroHqH9mSUYaB9xscc9eT+hB5uz6lEutqak1Z
DAaVMRMqoVryR7DI49I1RkrUDgVqdA7Rqsv3GGteWVYwWEtlGEhMtvUvwnDFYeztI2tQXgj1wgnJ
scotB3Q/BKs43I/pfwS/X4/Q/HEIG1bD+jOnyLxQomQiAtHsy/yXZ9a90Vh9gnv6XW14rj+HDQHO
k/L1N3S0TUMlZ/NasudzjsHUy7Fkk/W7lIJ0kr3+aRyLtMhtYU/dWF2j2++NQT19tSEWsiRg7P1m
p8qdXwsNw8mVwiIyDablPgC5ZpoCj5zHiY7jK72XM4IP+tVkRx0CR6l+uFtieAyPkJWFCa5g5cEO
pTU33jK8aD0nd/HaO4KvjZ993CHqxMD3bMvgO3Lk6F4WvkJgAbjqorReMb4CZWI0+AVhc6U765hS
7UlCoub7k1pUQoUaI5GU3noY+J7R7Po/9/AXuVYrH3yBt604q9H4MGQm/6NBTtp1AJ0bcKTQ5xqX
aD1vKft6xsYbUgZatJYFqdJuENdaYcJ34eod0DJ2C5GzGQdeoHQqoyDQS2jdNatZd7jahGuULqQ7
xitygCXsU/eQ12VFBzRRNQ/RrqnCJiQX7cLcoOdurcNwwsj5a/9/HhVlNUHoGWMOp3yeKhSxXVPW
WPSvX2TRfDyA+8y5KdV5RqTTHZqfSPkuCvS7iDaRxrSMc5ssX2h144W/F3bO/jh4g8rJGPwPvLuO
+gpbTo+ygLVcYik9QQaJOblXuLMT12KD9QxKnqR1qtOm5jifFWDL1OLR8/egQNPSmcT8+/KwmwVo
7TPxnSmXVBDLNVmQf9+Zt07XQoKFtAbB72ISnRtVTiwbcFd4G6zPSu279Hud4rC3OTOt5Gf88T54
34czvpskU52t+MDd2qX3c6RDz1QdjNZIiAnaSJvAVyUI15RNZUnnHgD+3KuX42K4kuPfvwWx+QRo
i2cQqaiaFt9ArxvUtVwbUTCIk2bHX/OPblmTNSOkcPZ+Ci+c4WdllCPQZ9uP7sPYe0l/gLyFh2T9
yVDDAJCdmZFujPrLmPXoz8mkW0tPf688Dh49/y0iklTEqCS915MIIPGev43hMscY8oH7dMbcqzjG
QKcztRyc0LCtGK9QsGBpKetr0kBASOemrg1aOdcIpaSWgkvIG80rNtiXD3U0NBEeYKz40FGMI7Pb
lcKXHkUUlpH5PNPnG4oOVWksBSpJuMnOOB40Zh+swarxa5XnLqqS3KXvqOiD4lWjGowFqshBM0rI
NSVMmjqru/rpAGl/EHrI0OogDbkflOXGhT4I5GltfPjIbwLfp0Ub0N7jZQJNyE4/0y/y/a2q6v5v
PFLIpaHhMUw4OLnsPwj38NbWtlNHhyH3sQd8ZIU7vmc1LaYWKBXZOd/sC7U1hvyh0khyyqr4quTE
7nQkT9DZwEGv+mWrbOSileK9wiVG6wfQo2wyjgWAhWEgnW78fRiF5Ep0KkH33gfZyHcs4K9kvYbR
U8lmOIRcgVyfX9LSYGQ4icfD+563LlyUX6sE4QRBP7foUuikNthgmqUFwLOxjesfti2akYdQsvaY
S/chSOQDWuwlOGMAeZJj6FkbUwX4OjjZmK+XolLg8m3qr/7XCO//Q2taKCWzMJ0xbI7t5+sjRfuT
sOXoi0wprIk5s7vEu3Fmt7uQsksgs8Pcm4tNcFe7nfMZcUvPcf9h8FF309wvx67BcbDMgdWZJ7p0
IYyYF6/xdP5eeu5W4Nd0N/+Kc/BqbUOWJyFqwtwlJ2X7H7H0jYfrr6iSK7u0jzN85aaCjuC0s716
Cq6fg8tETThKBXhWckMGDcv81ORKr30Ny/n6sMmgiVyPRiLX8tDU4x6cRKla9isWi7/SXV0cq+Tm
/lNor6Mr3WW7tlmLUAZ4+PcLKzQ/WfsWohqITieSRsLA0g4TN9iqvZdGXGui3NSFThOG48xJuWLr
TQ13/bkXkPrS+r1MnpeZhuID6ZarbvPPByqEvwLy0uGodiDnvE7k/oztYfiTWJEhi3mDrQyMNX5S
rvvuuCioX+StRhHRXBN/9J3ESsP47JyXDrbUXbRT5QZZ98Gcc/iuT9WhNNS65gqbZpogfwDw+bmX
DWBWgimMECq0Y1Js3GRQz7mqVkLIXVAoWUtCIc/DWokLHo0WDDwQL4YrKGg8oWTt4pGJZwGPQmpN
bVjNaq5tNJMkGoWzKX2YsVkZy+JUW/jjaS3XijW5KUDfifPIjqkhslZ4YlyGMGWvi1UhaCJB5/ST
Aqlfl3SvUxCeAj+i0jCGDilSc7NWcbI4FwoNWVOvo4/RERYyElWQEnnsuloB+6bQWwo7uAZ/Tpne
iNCL3CSfUudXHgPT2gwIHFK+A+mGNYnS1IjBzkS49h7YO1QVPaHLl6SO4J20TJVEPI6usZEiYmNE
wD8k5Nlehbl6CgtaNg7DWT2c1yGHuwm7U2eOw+cmz+1GLwXRcsyjuPaRBa2G9t0QLSARa94+/qNd
uOK4ySxP5Uc80iTlegf4FW3rQANT/Jh0MGJV5hvts3IG9+LXVPsuCIiUNuSrQVdwDGDtIHIVnDS3
SaqE/WfRV9nFZkCz4/AciED6Yar1cop7xClhIeY1OvXYZHPvzmXO+DOEhKO43fPGmaPr8aZrq5dW
FqOEOm0nTtoGS2GTKYirG1RRcJ0/L1CqIJhrgDWqCqq5ApF92HJ/0dmPEJj/rO9z77i3smkDhrqn
xBlmTzicSo7EQObGCh6OvYJei5O2bE7hAdNbRcaNSgtaimvnrBQ2DpvOIbZTZOMJ6hQVqrTLBjOj
6n6ID29XdsA7ME4XmvHseuajtUZiZVgqxmSnHBkXcaiDw6+KDYM7vc0IIay+BqufXMvMA3Su9uTr
Nm5S82P3VIQEtaD98ZbMfgCaCZl6uluY1YL5pyGfKTlLCNyazCW/FBjZsIOhmeti6ThhAo6r80o9
z/wluF54vbeZ1tR9IC1eeajzZBPZ+0ofAQuCQZlv9yERNGD1bywj9FfPoKjDqkiDqQz/GG5Jv/E3
KFgx6ixCtGZxCvTQbg9+NH6TsP0G+indLMdCqZ2sOWeYrKrl8/9p8wGF6A8B2fopfMmEDFv3MnRy
zTlwouauol+qxpO6EwJReI54QBh+MHDlgTeUA6G1YvfHcyOwsKDj5gf8tFexbsqXu3q9Fu5jFqC1
xpqCg3eEokbL/Yvs+rhNLq79yfJv2BojrI/EwA9lw2x0xv3B/MPEA90fATN+ybsrf3TXw8RtKh11
64ZABt8RbTBxCzCnMJJtiw8gMt4U2QpJzu33k5EBDiZ/XxI2D8aakBJOcP/em1uASRrEwMZq/PTB
7JxLYgsA88SK9sPclQp9xe4ZJwM/WNtLt9iQ/aob1g3rm5ReH7Y0kI6L741z1j6nxrdUA6dxcJ0A
CqLWU6y/jdIqOC3OxUnrxB1gZHmvYbNtUttGlCrBg/I11Bu9EESvtaiA7E3rzejW5Xjhk01E+NyH
yDPE1tZyKOiRtqSiPaCfWBmc3T4LYbQLorUJs4i/ESVB0WiynCsgHBvLkgaGmWyOlCN1QNn19EUf
sV53zbcN46CnjZ0w2erWakC891MZy6KWDm/V1dHFemV1OE3k/qBnOboE6OeosaBblL706PeAnoGW
j1sgo2Y3VKZjhIjG8bnj8sthcUuaAZGhJsL9MVMwWOdLsgHol445Qsz4u2Xjq3aAixFaSDsu2VtI
Uf1xnGUm005CR9YkjvM0waFA+YIm/KM5c6uDP7mcHyjVvlzUq4tfhbgvu6tcqbnKCJuEnCOeLROW
+NI/T3FJ71R71J8a/yG5oRTiXgdapazbJlutz/OHxLviqHtbYIrY32kQ+5JyJsQjM3srM9WhobAd
E5z45zl4sRI+p6cIcuPTLalIVeUdE/IJiA4amrM0Zl9yXfnW5ExDg+zG/kmp0OR4Uud3DabrPNvr
O32gAuU1g/QdXbNVqDlYkT7IwkXDjD7w487G41kDfpKPr87MqB7JmQ04Cl3ZE1d1+gGPfucUEyI0
X1vrE/M1zgqFQ0lbSLpFXS0EvunTBpsGBX85Ow7TuZQb0HK68SnMKCsLTUNxlE50FH4jlafPKdKS
Y55fgAoetteIL8eqGl3LI8yHDph0Zfai4L/NFp0bR4VtrAE7f/STac6mg+Uo6blomUZqNBw4eIOB
gJHFL0CiUqQFyQq486VgthxfJBJr48t4QA9OIJq4DFpP52UY90VZL46v0ak+Os4UHCy/WAUMnzNu
IS/b2z7UQu8Il3HL59zce1oB5+1Pu63vdUiMUPKAz6K9wtnBn/Ii+/i1j6FptYoRMU1401baVKjE
ClPQIt3EuwvOtP5Bq80fAPi1jUBqkwQAP1p9k/uUJfEoDO1LYbnyFwDqbVwIzoYuEPrUlhyEkd/n
zwj8RJB4oE7EHt+LIuPGumxvqFBhU6Cp6Zech8Pdqubc/TkRfCdqulTPtrwnqaXfYYBsmzI5ummr
ReGF8GhTqvBw/bd7XdRD94EAsyQtu3ND12eLT+0FfC8p+h5aP+rj7EamEBSX0fVT7IJ9xVLraxPp
z0ipyd5a9nUSNEoq3/uw7pGZtRb57phj//9UJdZSYSJS9u9884pe1VAlYYqSLpIQZRfbWUdHQgGz
CIkExo1vUTNda9VKWp0jLIwDvFEB4emAvD5uqXo6CdipReGNZlP3ngWdvFmaLdRAfLcia1t2I9ve
+zZ0knLubGQAusdyJFRi+x3RFlOB8jDwTjPjh8s6Sl4gKpKCZiP+698NgN5FgCaOVoaWyLTL9GPP
7uEq84HoLN2OfDho7xNMbV7R/nGVFvnhzDZ3PFnISoH1cERGK0o7W0xtOk6cowGwHC+mkqk/GsW+
7daQ2zRBpYug2F3JkgCv0P45FaMR+vLonueDdTny/bG86nz68/Rvs+MfGDEelWBooePtuzi7QstA
J+EyzqYYvsfDkLUp7isJi2yVkW0dn/6j0Hfgk+HEgawOJ0Cl+y9DvhdaeYn/Wv0tQMwNF+gHCbQP
Y8gSX95Vk10YeolwPAsYZhxaAZ+2PuuU861vnWSFuKUZ5+TImQj0sRZ6nG4+szp5R5+/tNLcJzoB
fHxuYHvD60svUoMsQRwgbYhFn2M9wmMDM0dzNtpjoyfwc/XxDnGOIgia1tEDryTCu/LC7Bdvr45g
Ic6zRLisCxmrfPk8hSSIllZRDXLmUIu2/kTTwqrZbfYJ7925OhOobj1GRrgWLHT4dhZ20ehs7hSM
rq5pTokSSgrzGm9gEHncotkOWZGluh+bW01Xl7ChQNrVwLeRdgXJ/TI5422vbbkgz+aPusz54g6d
PsvD+/ENYiy3sqIgYbXGw+txX2Gd8AfwmLpcVDiBQw1G37f/RInrzvBHSEQJ/mRMWCnuXfUpoWst
THIBt94AUHufL/k+G6Fq0gp2YsZHr/7B5eUXglvvwRKMjJJjCTbG4rHAhPEqfNbsUYNYq3Aiuzq0
HTZ5r8UJddnuhxaWOYARdUFhUSC6okNNiVYbnV+E/2iX4Gl144gJ1g/+efCI7tqL2meB3hxzFjuZ
jFesJ/lq36ulCGkbxBIDDes4cWZ/BChVcEvKT726bvnqF8/PaV8kRURaUVZ3ziJHLurpeZ6ufhDZ
mTaM/OV/k9UOWt2ke5vK/p25RJslOHYpfiy7E+5xBXjVeo1UFp8MeJivaJl1TREbforxhjS2l+xU
dCoSFv3lWdDikc8HCbm/TxUbw7N18LP5l0GT1uspBbc6WokWI1RD1OMSEu3xHvSjIj4SxztCTyLE
PEasc0KD3Foh9hRl2SCUKlghM1atidt/9TOsANnKyQiIKVWQurfxSH1BX8lXY54HejYmyluYvvJU
BYTTHjH+L2fpDp6dgdY6DREoRWCRAHW3/b2xEVLYp76SCrNN8bfIorZjOKzoElNPeKaJB7/WaAWr
+Jx+8BiMQsb1y7Ck8dsblTLAcnwEoJN3AsbI5IbYOkXQLIqwrskIwNj1UPU+nKO/PV2pe5ikkZqB
1ziC/ZbAcCVeHpzaF2/NzjYjojPOcC9bo3KgNuR4iM4mJGdftDy8L+/4mqDnwgmrXmpL05qgrzzX
hghTyBR8ybK6onjoRaKG4Z71lXLNSTKwmv5SDeUvJLpN7XOeXXqJm8Pfl19w96UUf4kA+MfNyDH5
3spk01R9SXfWtbIYMc4iSMyH9ni9ybb4rQNbhBR9AawFFmxbanozYYoBTdZ6mfcL4FdMYOyzuWEh
3p8DoK7B8jsyjwZOIO6tlbtfC7F7mnI5o6eHUwGmSP6wnkG9ygwV+rmnRO5nbIwaDi3XjvTwtmEA
1AeyaQF0yI9JNfs3gJvVkjxX3ipqxMvL/cfY1Mi1bHn31uKU9qENwWRNT2MfwPFHiRIcFHW7qdFC
EhVpX1c1xfAowlsqu732ABiqyc5cPXGT+yNqOMyKT2YfEIyJMBcBgfyFSNnHsJ4VFQwvAoZN63T4
arBzVg1Txh1t8zCBPn4vDcxPeVDpGSAETZ1daPLzYqK4TzSuXHAoVLzgW2f1eNVHKpRFRzSvyf2X
SpfE3YAPjWActOl2oqGe6ocj4QD/iXrwflc0miGSotwxJPmutOgHAuCz2SHQ+ISu1mHuZ5kA3vuY
EHMHZxZ3jB1aH0nCyQiXsTniwCJ7gOEhOklHnvR5zZ012zzeRGvIAQgrh4xH+s7b3Hy+2d7KLktV
+GATzfvNVzkJCH9mFQ/f0Xue+9e6ifESJh1+HaYFTBt67jyPDc8bEUinXEaEYE7GV/5GKZjCiBLB
NrcziyakDxi+pXVyE5lW1Wl29OmrjOK6YaRRh4TUiRcwbFoaO3tKtlhzOaNytxx0AmfUON7kU9mP
kz9NJc26LLnl45UlrrjzKVRhWzv8guoKphfjdXtkEHMB6XlQkr+Z97y2UQkN5HL8xBzBvPxiF4FI
o+gsi5oWHdoqq7wPJjmFnVpLXleU7l95gPvbbmc0v2R9IIXDw4VLoNmNJ3opCnt31X4a7IY9fnXO
TFFypudljtaV3yFZfIX0S/DqfWUgmZGjd99YO+WZTHJVUOajbbi7jMafay/Es+TZeIKroIHW37g2
AyI5X68TkskC7wdzmt5eFY8BKvKBPK1ufP8DUBxeOW5hltV4c6S4/bW8hrEoG5DfN5FuU2E2v7oG
9C13BEGt/Cos+DAklh5sXVJw59waVi/Xm8P8+DVCkP0dXOPV2htFC90f89toSqWnIv0W5M1fpm1I
7szeR2MSbYn5m3XlO7h+H8/hX8b0aOCrKj5fFNnQPfVABJa7KLMa1ua120SgTLAnw6jAsTAMvTpu
KWLHb4OmzEHo59iF+PCU8vVOX1OXEVkJ3HidWEav99M0A9p6BiN/Yh8geBz2lowDynl8K+DWQcCe
+HjbnCSyhe5PvyEe/CghGRc5eEkH6b9hNps+cSyeSMOkGvkzHoVCf1I4EzBN2ZR7TPNVq4VAe03H
jT6KXjiE27o5Od/UY5YgkY7jII9QVrpN4oNDBg1A6o6qDnv82xNilxN86JeAaTj3sZjxyoI0pBjr
eV7w0e5JDylSGAMcfTKnUngDkXda4uODSxOLUylXzhvoUtL6jQ88Wg086kdYccFUV1hpO4YT4+ZM
Aoo+vOMULo0yXHrJQdxVXBSddU7tcr1I+V6kKuMDLrCJ6H5pTN7ztB0lFLMduU2SqV9Ex6VVgD5a
eKpBRR2v/QlMwgPKWVg5vtqMFWnPPDHoToTpz+MHShSo1XAxlCZr/HyrDS+I6rzZEqamRMxNfgtW
ZIcF/5oyCrsYKlGUj9XxIhVW4iTwX1YJJXTgakU9RDImhjMHsr5rreKefORNaTRK5hjPlXsMkmnc
Zpffa6SW4pNAq4sBId/S7sUIO52kIQUI5XYKVpfbghEPBeQWirH4Gdfc76hpZzKYhSNf7rH+RDtD
VTkUAidPfprMvcLmi7shtcM7KqLaX2AahIUMEtaeHpc4Lft6EIHWoTpy11QnTxfDbSn4Og3kcBIt
QO1wN+N36aGDqWFG4MTBCLcjM94QNxhZQs456oMix9S8iJHxoiydcyebd/JS2DrhCRCcmUyY4ggP
6KhGIteBJiGpzTvK81E11YZhFOyAP7ZbhsJvT4Pa1mg1mKkbxi+CRopaQcrWaDl7Mu5bplCVfmfg
i7suKYkJpcxq8A/QuwEXZ8DKVTOPjFUTQSo8WcTaB8vy8o+Q/qWkMfJlKvhF+Xm7B54OyVbqkNE4
DiOPLyUoeZCalFut543MZi4ELXO+/mXce+/vdSNuhzL3r1wtTSqe05pH1qZEIyWRFt0EnK7ttjKa
MKGbNlTTmjTCaDk8GTrO+FDiXqtKZTb3GZQ0ZODcxnQWjAA/n1xjkZYdcV/nC+gN4dxDYXtP3H2L
CwIXujHLlIAdw0BqQR7DTDfTAHmOruYh9kmkaKoEp5EMjqkZJ77iyBheLbGPPt+9C44yJKxnxSDk
F1FlbXvOHsjgFewuNa6QlGzvEQ1uCLe7ff1i48g832mzI9pPNBl9ofGFwFgSGZ9pxfacOXgrP1aJ
3MoSMKtBceCylHkyCAS/sNnFH9cuzpRP8R8yzspKHcxQPjudgfZSIawGjMHo+QSn8WV3wm1xQ5VD
g4Z8Di9I46qtYGJMtJKJhi6ubK5TjevIo8kNcVssPBo9JA29ZzxBoXJaFng6phbBKgRcT4Zb/El9
EjafZz29ImkJ6S9ThBneEiWcRkX6bB5VvZkgylJla53CfxgFbdADT2k5voKmBeBQ1VNLuD64+JCS
hee6mVuDzY08ZfZ9JhCQqvLIwxc8HcXVz5K6gcg23kUI33hL5gnXpMkMa3cOH9SGoxqxmoJGiLSJ
cWBTIZD8TaxNBIIIt/9sg7JhKD8ubKLr04tMkyW0rK9gwCe8VdVbj7gHSW/48N8Hm5+fBfBjOx0s
eJpiLRVuKJJVfk4saP+qd3IdPpjp4Cb9dYRtBQnvOQoa9W+6yrOa1A7cnKOaqYLf9OeRcUyVIJvO
EKwQVreEwSHHb1gVb6+0qhONtfFjYDk+z53zPepi1fDHhFuoOlWGZOlXlUZCkuF2EUvFQ0cAqJZu
YBV4BhK+G5sIwzyjEVhuLGl4rbtLaXwP6fudWrtNcgaCmaLVFwv2lcWhATnvr6g56XXLGKFVfkmz
edXCla0rHdhFL1cFmLzfQmw/b9LQ530WRkDm/zK/VEarpgtRBzFlFlgKL9ZzrFeUA3UQnyskoYE6
l693L0jUmZOQDFlczMI2RWslSbiGHdXGKg2N7Lyi/rCjZZBsNG1i57pIl/SVvAATXw2dCu1b6h6p
a7AbPpd12m7AcmcPfxWJ63KYaYqQubIIdUqEvzgjPgtEa9b8W48bgaGweOmuKmziVWAbnSw8E00P
yPLE5CyVvEjeEca1GA5SDR2bJbId8ZCSXpZYojlTZWDL63dVjV04uef1QNnfPRn0RBlkU/U+XhGQ
VZow9ntGjPSORsnPRgZdzh9ev9It7fmyqbbSPusu1zQBi3sMJKZEjJkwOIW4jzT43l8gIe9+6RTj
jmghYNYgh9ouOCNG8egVLyb+le5qEbce3MubA8IhG/mXyMRZHuHDnSK6psYrvMAYY02/29si5rPe
L9wXpnlIEUzyRqIlOGeu7Uh/W79COhmd7becWiBnwcruyDk0AbS895SzDsJSMTDTysOTEftaDT2b
vEuXDuz8OZPOVWjR7GWCtbAmER55eZW+WB0laR3cgsJRyrn+WUbI+BsWCqF82fddKtHOkc5uG6fb
P7vOMOGQhAthjbcI3DpMQ5NqdWQMplwFxm1G5j0Xd/50isZ7ZF0ultcoqHULJRX4WRExESpVjN3J
Dzam5aHeLjyRPr+9Xk7C19w1LR0KDe2DoWkusudHB7GXaCG5oRJwrRrXAlyjXlr5hM3skZuRFGDx
XQZWeU3lXjYcVMZ3yBbMdtDwThJ5dGIXmsVnQCI6btogzoxg09TWb8Pkt3GnGt7jYCf5se/iDbTX
AEnV1qTNTdvGOAphphY/gMF3BtYRb+Y/6NBKybww6ywH22CgAYgZMJC5L9w1CxZfFCB+jTPFg2o6
WyDSXWj5Hm2QS9NxaRFSCCSd8KE4LfBR6CZLKdb6dI+/H6Aa++lNaUn+EVHo56B6jX4+v63dMPYa
VCZBTQtvDaolocUwxKsrmQmPS9N5ZrwQuerNfjoyECaZlO0dAmquwXO2ZxYytx5aA9IZa2CngXgM
BP6FY7JJ3fFxMZb0lWjwH8wR9H6hBLhZlot2c3IgAW/ZgqGEQErNXsaYxhfKAuHn4moOE6WanIZ2
6ccuCHo0gmu55UtfMn6jNJ3ZLZQKwVZ/Wcz/0KmU//QtcRMcnRzxzdrvjvQuyClWiOZemuzGt9HA
hqbwAVt9JShhmTQFHFKlxC5prxebSH2p58lLpNIUk6phDklJntDBufcXSkDtfetwdjXswkht7HHI
Lr1AXPtNLwlVLVDOFQPlUbCJk0vd8uORqhaaT7GjLV97aWDSJ1IP5AWds5Slfli+0hZZM0TM1iUq
8ZGCBxd0d34RsXSPSH9AELYTeGUGiIsLhTvKsqxGUHKxSreMWfl1HMxNgYGmvY64/1+2nayioNEm
GKYm8cVNtWKrtZ33JVakaMlHetTzdTmsTTxqP1ZCFLYpypLqBStoDI7kfy43tPvzOrENvMAHHF/l
kycMOEu3KnvpJXRH29rBHBldCY14AYAefPlgIGkydCi+onYw3KnSC11X9HSq1xSrA2bJBuab+Lmh
iyTSXVwhne8eht1dEwPpjmTjBZs6QMRTDPS4ioxC8xOTQqVYh49Pzu9HFTMTyJadvwu8bT6ApieP
/JxFiic2mzN3nyK0tjk//9V/FItdQaSQS/cKrcjqTvz2q9HrpnRGcKgUL+dkOf/nxxvcSYmuBRji
btQRiZUlZpq9GBKW8rajNXnNGoUjzI5+aneRWqdsh5tW+HDmTxvpZc5k4IdbFbmTau4P37jX4wpQ
pCi3H+wHCMuWBOSa8kKZ8DRGNPONK/5WlOiymkK2Wh+SU4DJQu4y933e9fOEZSoQUEos9KRYPsT7
1MUy+v5QnWGzryB9MvENWhNh5FeGys3yj6duT095vSASZZgAOC3lJ/T+5v40feYR0YdiYc2cdjYb
vb2BSu1TttW0LCU6tIrkqQBezFWVZ+Vm72yZP1uRzWVIFPTkOHlGUH8NZoSOJ7EfkBLao0OX/KnX
cZsNXYK//lww/wtbjGPfiHTvQb1T/Z8Yyrdj43ZzvNYCa7nZsxjPAU2TxuCj3RCIEomZaeAaE1Yu
dhjfOIENwNlzg50WPJYX2q/UYkWCafHZtNQT7AIi2s87BjEdlSBIkxMxOcLXvJ1NVELXsPT/aSj3
n0Z67Gp9Uyng405qY+iIofdIObtv77Iwxxoye5E2Jvthk3kbzAdAjBcNcKplb1HVL8k7RgB/Bpd3
EdPptS1Ql0q1R9zmw46YoRn3T5JA792PxIcx1loe5ttmW56LOw3tSFMvPjgqgJTI+QuCbMUkGqgi
qhjhQlLt41goXu2Vv+P1Am2Gf2xIznL83ZqldYtuY2t5I9uycrVKqc0jJYTFUZO4qhM8YzfBuBx5
lYhG1EYC7RbR6e29WFrj0YBZcGpEbJVDh+R+qfQ/GN0V0j5bbnjQ2JWjUEfO6Slr3fBrHKPBpcae
B03OgQDjV/8kPO9ouKpZAkwW9ZVqtx5V84s6GBj/6XZb3bQS34BrECL2zScdghbemsXdxKHGvCR/
7fPc6y83df1RtljidvZKpwYp1QVc6W7JQYohkbRtM/Ghv1DSZmZuc6peqtYxbtgd3H1moxIVuU0C
zxWq/d+0H3RcK5xZQ2MOmTj6zxZOZK9vk3swY5YSd3Bo7ixYyE0d10FvDxRdjzr2lI87WMWcTLS4
mhM/gSX5gdXvWxdHkCM2D6b4TYex5snoYDqFrdPY6y2Iy98ih+2w/vlPUUSl4A93kmCgcmg9czu5
8m4BnQ14eIams0qlDk27NHi2qhxM+2ydDL8qc1YaTcXNu2e6lReljrC0trGR5OonPx7ywruLVI8L
bVlp4b2KD1lSFQYJxkOzWY3IkmVTor8wHhcqXYQm0KXobewyNgr+1deiAZAyQspcp24c7jqKMh5f
dZFl67iCwtmk0ZpNSLgZCqahT/T940qCUHysKBmNloSDOIctOLSZH4so/nH0LYOmnHjsM8dKbh7u
otsC5M6zFpNhkmU29oSJi5LZHb3BHxTX5d6XJoLn+4aczUpzKGnhcPjZYKId3K0eMmWRjIm72PIi
w2iBeZfX5NqFUti7PJcOkmN5WM9KJDEmc8xnImbuwMY1HN0QJQbQatdrjV6rnn1CWkrilrYu7Qbh
HG94NyhiEylqCXtxny/6Fie9td2X6FppMHeeQXzf2K1EONpIt1RBiR0I+JmKMQmM3gPXSW999gn9
ZhPoY7VxuT4uKDMT9u76EoLJG8BcvK5vwwwVeVVfi5d5vfpwYL4++XYsglt3BGMMcwdum271RGBq
3kx3VIvNUht7+L3vMMmCbR6BqgNBLuaASeRjpDnUFZseGHaBmCTbkXeEkxxC9qcOQ86wRLvXIyvy
8yuPIjAqjYJfw6bhUc8ySfAB4MxTUO86Pa0tH71WD3CKRriRDxpEEFMGAFavADflFKPuiwGM4Ykh
mm3ouD6BzsbHih9zU41EItirrv6dN/gKKkXkRMiiYkJ3IW6P91xBo3U8qAUACjCENGP2V1AJP/ap
TdaMpjxaPd9b1nwmjCVHMLTkwO9wei53IdHJKmL69agHwwaPtbJQMfYkFmAsOk9OlXN6yophSrAg
hKeI8ZHispYvse+CgEawihG7Pm/ymW/MJuGp25j/wiJzi/4KCzwQGYDvT8AOp7JVoOPDzEE0zqI9
FBiAeR8d8GXmijGOKLRFPNKGpYCsEasl2c1gc7bj7D3tTl+xSwfdpLLUkj4hKgPUAO2QYeh0qG4y
WkrHczoki7UhZ7gZsbvLxRFZ+BTqXuIZE4wP2swxgiR7XqbSLjPsPr8tQfZgB8OvbEe9otSxs+Vm
E8F3y7Sj4HPp8DwtCnVgnmLa0KChuSpyxb1Le5IoZtwgEHYhp71kostF06AK4xFbIVmGE8Jxcu8c
ZY1B0N/+JuTXGh575BUUPlIe7CmhflOwW7MecXlIdqQAQ5V7563ONqNL4MUBk7/RFo/dRX/4KPTY
hEzxJmMZbqghDJFQVWLM1FLfxQxgjxfi0k9aUs9CinYECAjFmVq/tLqe0nDOE+p88VQypHJ/rL9h
RmEpfTto5d4FyCIOIyue1hRHO/+wzkNRMK822sNx/Jkr+u+4owepXaNPVaJXSHgC00jRF3pygc0m
WCmZwSVXhEUGN4zNLyf8MM8ArvsHueICHSfN50s2BX4k+HnM9KBwjUGKggGwhYqLE/4I7em04trY
JJR0ki3Lr4lL9vCq3ubq+tBqz4jAVUArniKlKEUNb77nH5EETRfl6gPWl8Yt4Z9Azpr3GLfHGPx+
SEHMMaFYNRwkcogMYN3EHdxsQJ8YPDRWdVz94eSatgRAI/92qfoA7LnXTFuz+fe46uf9BANypqqy
q+09ICIJkD3oJ8/evpljWmWGuvhrfXfufHk7RtOKq6thPo9zrz4FjetN1GD9Attw97YuuJ1baoe9
2GktNTU5KnWO9okspbelWGhHu+5hKoYaoLOUU55najDYgIFWHFQP2Tk+otY/IsuNbxID7dHD8HZ5
3CHvI+bV94WUaV10cNCso0Ue8imbr4w+qhKT6470PiCVeTS0wVyyDGl6svv+H5kS4ZfEZFrfcDYz
XMfoiK1EF4Iu59l/rAXFZiJh+O0kpjc5h6KPwmwhAbzBBVEmeDO/ZtiZ5AU8MDx2yjKzPNn1cEUz
L44J1TVxfYc1nKrnsghfBJ+lzJEcRuxuGobbaYZuAFz4rpaEMTHNGW8SgoVG4ojbSPZsu//Hd6hH
p3n4kvO1zBFznrL8CJ6QB/itaZ5WHtb/OkUigsC5blpds1LPSsrOHrH1STM2VwlvCrG+NWrFgnKj
GPeDmXz0J9gGew5JJ5PsqTO7URc/JsHzfUEeG07oVD3ezkYxEuhtrJH959NwW5YI03t/fxeiPXKO
CVBySU/jwRvKOcR3fAltFsnDLMcc/gyo0gKNXsNctWLA0+84lVSZz/eRlRc7EonJ9DHu003xOODr
CtoMEbOyP48LmWU6979ddhkH0jRrcp53G3FZkIqBlLZ0JsiTgTQ5oStDUXHi/66yTHe3N2Kq4lH/
LAHQsjxv+PxDgDJ8Y96+0QVtexydaZG1OvepjdbFU30ny5veWwc5uwojdZ93r5v4FV8zeE/kd3bE
dONQJQHxAxU58X+126Po3pS3I17XprpgK8Rrr1evzI38NkJjYWVIWKXBHMgS2PIsP/eTIW0JzS52
bi/ThtWrOTjZE4ApCd921JPcEkvBm+Uy5gqGcOVoLf/u1KNf6eUbOy3uLArGUCILcgYZjS80sxv/
mtqjCWjlUX/1F5XJGhPpPoKFkQ0sw33TYxFLv9lNOK9coguz1tl0ZlpoKwKW1mAh7cf4MZuFMUyK
RxGDcLj+N49CQ/KHRjIc+zQcJyCWFdfJm15QXSsdMFZrVIpOHxIKQftV6MZ9p5JMesmrGMLwjDeq
FDYdt9k60jw3c1ww3zHjg+UM6dX55O+vmxIIZ8e3K5oBZ1CnQiHOaQmE21Q4sahOiZAGT+9OBJeR
Qe5++vY2Xiekmz2sgPOsLcPsL2NKEsyQc2oHXqLm+svpUB20TDYbgWqnwlYDWawg9ZoPeig3woik
/yUdDcXD5ZHva9OAgAKnV7uoWv5DXlAP0Zb0I5Ixuba6bA/NESwQxkhynGWwfK6YpSZEETwgSaDg
F5qP/yCkgPvMgavhfZuM4lL5jVh3K2d4UU9H0PFjFnQ4/LqZNhsT2fo0MaoN8mjOZ3AtDNAuV9q+
l3WEfnGUyJ3eI0KBiqNfaSo0/y7UmigDybRxh+fWWnVkVIPLv8gdE5zz1ntR8ReFrb5CQME4Ej6q
TbjFIKxctPglCDuHu5GBwlKk2tBHOFnqAzNO9psOeGaFziymuWAkM1z4s0oJ7tCU/X6vZuHXXKuP
3F3M91deWAye8uOUUoVaK58S6EcUDTCOpf75vDKDmzH7Qmnb1NPkyYHtBojizS9Tf77f+uCfg0hb
xPJZC9EunOCnQqIT3u/ogyWWHDP3DoocXLViCGjssa1zaJAROoLhBD68vVU+zKu6WC2JJA/I2YHi
m5kty6d5aK8qU43uWEbB6OShHHjpaVtJrGoTose63pJhvx+wI0Owcevs7PS2TwU3Fh+XtHrTkQGQ
5xcVGKcGH5XmhU8QqkpZVLpxR7F8F//7c0UNZhxUAkmzcXmIUYZSl2tEyz7v6z1t5D+pNpQTWx6L
0xr9BfEmsnm7G65Z/qp4SL9rxsd2YErdci6slIVvorHJ+/ROTCDXBoN16eDDtKgrFBedVmRW9iMU
HCwUcsA+YaUWQlh90k3NkZ0TO3VMSEtreMPirsZkEPThvOMC0OJqr+vec9w7QJ8ADepRjPb1Zsmw
ll18fzWgB7d8TsTIkIQZ43qPMUilNh5o4L8NUTv+yTg3jbSkIgoQRhXCUaRXI5V5g4XbfeTIZQEx
8B3DGW7OB2ZDC82qj8xTxMoselPeQ17GjCPe+W1YYi8ri1/uCq7jNtA+wT0FngKdRh6j6ONFZNVV
i433Y9d4b7PluS3crzI6G+8bsksO15q5WG9P/QACcft1nd2Ei+jlROYorNo4FzMDyM9LzbsJVnht
LPug7TRN4D+xJp5KUKKFnQnikg+qfqicumW5xTKYao/tQfIoRlCHHYsuNC3ExzBuO8y4ZwguVyth
3RQUyK7yYIaCE9vpi2zEFdaSZeEZ3GitxUGXF4j6iv1Q24cid4ILRI4a8+qSclI1NPtNn8VtqpRl
yd9bKAnfhW/KL5mScfdR9rBQ50Max/LPK25axtpyTbXLfHYjkgblj3jMDSZu8THGISRQBblID4xH
BDahy1v+r1LI5aYbsRZLmS3EZGITGI40VcWW0xYMiMwf71w/8Yc+ajGkVNp5qjxWgFAFLPcq27Gf
2LhoVqFUhsHX018m/NTX6JxeiJ2ijLO0KJ+VogF5tmXgnEZEoCdxAbjM/hY/QHQCiyGvzTlJ3ZHF
qqbRRJebgtzjE/Hx/hqU9BA97zXqy1UTgGzQY9GRde59l5YuilGdCrRtCjhsICy9z1gJGECDUzVz
3NEYljhTNzOu5CTT4ESjgOoTyIQPAghTa3PNUY9CKkdrk+Szy4j67dB2uYl8ee5H0TUmpl4V1OHI
F514i02vWR4bRsS8U5KXtW9w3aAq2p+aEbHAqGm9ScttknkUY04PRVwRWROdswYWss4M+tBvUTZv
dlwPgSoA6oRQhvKTACF8fF13GgzzhfOJevA0LN4UNY3fj3NxhFfqdzmQCelFPMT9uMKmadGyqtRk
muFJWfKKR/3znSF9slT+H8apRVV4LAj3fbIJyoB0kWoh9rKK4XjXTntYV/tSq4dnJo700Za/BhY+
hBLj7O9nteHp1RALQGd29NVs7C1sKGGBaNUOq5e35WxaTi6m0ehhGnbBsTBiXZds5Ud4qhZLgk40
O7ngXak5ChYcnpUamrpX6k9e5HWVFedvyUnJCvSk+S0Ja/2x3dQMYg5yp9VlSOq5QfzfizdMh049
GGXW6g+hPyu1DCd9XNR3EUWHib2ohbg0EtfVOR+erqOxxauLQ70nFoomrux1ecgYNd32XjtAgVw8
tqTZVFD1jfFkboaWSqkJpDt4R+csoZDN5gZky7G8APOv6pbYnT8vr0aw47feLHRMkuJRmO5B0+Uj
nxdiqvPQ4aHpHp7XIYU2bfT+chI8BXv0L5Z05GAPR30e/R0fjptf55pnwlhiCakRqkw3YSNZPFh7
ix8TsP3oQseJ5xJmFIeD2bVzPmr1v4o7AKojI0T1FbDPM9MQEGA1L6nNFWByRjce5UNTO0xO3JbK
x0pC5XTom8ShBva+akZJkybdnSLEIpZIM9phoM5aqmkEus91H72IufYCFII1J/Fju3y+kHpOVAff
cRuYG/T01/BSHLZLqO9QeKvGhqyXE3KN3Ra3vkl7+p3FYFGhA0SZXbGjHtMUFFYx42L3U7USWwSK
mSM3OrassPICUKkxpy7E8VKW8pgBMtydbpxl72oYgzngr9jcDmBKmts1hE26oRPoPbrYG45UdvRR
kCEJs1u1p0ipKla9Dx4K0yhuJdgubMgAYOBH42yPFz7RJexZK4YULGz0gGAqIMoxztJTsHLvWbSV
DXFI3EtDpf0mAsyf/AS3CJ02Wt0NLER+owIdA65fJu1r3Nyy8Ztoin4nsNIizAuftKsyBZ33FrYe
KBBUzNhcNdC/mTrjP1u3+wrQKeM6dsQNKNrr5p2IVoVRc3F1bvD55FjseBC7IQUB8HJHXoViBkDE
X4/aXeKIZCcma4DZJvzI/CzLuELYwdW4uwMjxi0O1H/cnhlxqC6kkAsVjJI6c0/MHXdbRTxsKAb3
9VJZ8lGmlm6ISL48xf4Ez9shItidB9tO+Tlf9PgrvJ4ZO7e/gZTx7v8rt+HaTZibuk7pwARXJKX0
uisgb8DLSX0czN/RFnDBmVE0nyMPURzxBqBVXtCZ6y/LeXxwEKQm3jGxAFtVEHjqte33p9RDV8ni
fuWWVPk8ICVOxpd/KW8aveSNrgK385Hlddoy6AHNJZSVOPXBaI50+/fYIBApKrXRYiQ5WlXxR7PR
yy/+7ku8rQFv8J18bzmygGizYdBR1vlpVkTJwb1f2BD6MphrfuuX79TtXYpE9Uk91HnyAokGpZdV
HbE35/hUNkazqjOnhamaKB3DaDSdY/5j9wbaH3ZuO/IjoLsn4FSG2Ted29DkXIyJ2dsjoOQ+TNpt
+6ALcS9Cmwh+8cXPPK02KzoQ37rXhhmUb/pjJA2OYTMrzkwK8w+0lHuoQBIFjrFFEBl1KNu5t19A
lNohbLJHoktcoTjYihypdPzXW2GuucquOKRYMELmipR+XqzAE3JKiJHvXyHsYzv9PYXsgEc/l514
hFD+MuuenbOjMpEVViSysNiF1EN6WMm55VoRvpmpELiNMKSumYMCWIGf8BqtmmEnqCKwfEvt6dWk
0vXhh+AFy+qVuiWh66Ym8dOHA4XuLkn4nOPRD4AjLDjHEhvmWcjNar8vSAw8MIW4vNrtZ4sJiV4i
8g1A7SQ+j4gumcESH4zBymUS0g7GdQCAXdL/CDQloGseqCM9rtiK2kcIzGliFmG5pgzs31isD1Ml
jkB8dSycgnZqXyjwMQFCNeyN2SMBcBzMtN1C0Qwj9mj8jT90ZP9Q+i6jY5Qp81hGDFg7YdmDJIDb
JqpfxuGRD8ReTgfPx2IF3PMnDLRuyxjnzhMPvkIGpZUSNkmUHIL/K7Y92Ag46PvB2KDtDrQqR3kK
DbE6hdEfna5ryxKyDH9/Y2c4eCrHzTZdv6BeKVBWBrhlLUTjaf2NZHv+27HXxwYOIoOkzNmRMhHS
gjNbLkYj0MuDmRUzMHtPSTojh0HVNo4oNVbsnsw9J4j+CoIpCD1rzAUETUdSStT7ST3Lp5LNJyS9
7E0cf0VLpWF/b/xMzKAU5R9pKhqzU4Mhu3wstk2BN4hYKwuMR370Dfq7VlpZ3UgoBnjL4aiqZ9z/
uakE4WWgdzEAt92MuIDZdNu77ddxlW4EXDZWkj/OYt7ATHBxnYBcLNDBUdEP1gYAk+zbneLxjeMU
YW00gSj2vfc4er3cJrbx8oJVFbdsgaEFO+wVMiPdbyR0iDvYKLevIzJrxeqtWrOloeJCnedVXRWC
rZPmElmGZJcXVhcgV85iRG8LTQMeo8Ar26QyOEcpzOYScVSFiZgswTEKIJgoUtI3coBzVPiQprTF
6SbqlXyOkElGdGiFqI3rcvLmiCqQ1hJilmVntzXL0vJ1ufNbsudEMuv1Dp5OdvjTyRFuGV/Aqd2S
DHmSEVdUSpbNLZ77sfZDvfyFYrJlT4hLuVa6thwxQtPAffGjpbsF5bGcqE+aU9nBZQOiUVHSTnDA
GOkd8o1s6eUTv/4yhxDIyBjqQSxMJIhfgYAkOStLsL1dLa6jxOLgglVA/S5PbacwI+fhj687zVXf
qXxm1H0eIeiTbJChZNyu/TCerAioESQoT5yoTbowDub6XU3xw0T0wuKJpSAVDC17aUVnlJydCOv7
TCl6bOM94gM2nw5GkXgmoXLSNSi0WXu1nowTLYufg2osYlkJL4ib/C0C2dtfEUsXxMZ0FoUwws/O
BmKyxv6l8Id1maLvYEXU12wPvqVM8kdVMWgjyCsevWV+6hklcSvPYAnEV2xqtZ0KJqzLU5bJw+UD
mJ2KulrQh9jMsYJXIgaJQBzb/0DcmDA2Vhj5pnihlOdCbA3stZ1Ozz3dyI1jHej0yEYGsdY4YBmi
VDsmv0NQvtv/45OeSFBZU9Td8FOQ2FDxnFBvsViFQYP9KVhD/m6439Q6H+ZEepi8ce5IYe2zcT43
EtZMmsQPv6Fna8wro5Ut+zqdoAnBJVHBJ48Hp9zP88Hm0CRI4Jo06IdI14vEANWqPNjMuYYKZneW
iy/cYm3TCLL8RZ0SkL7kv7ly37ngDx682cS3Frfqzp5By+R0okbD1b7xvlh7sgHM8b3zy+aDyx0j
z/5y+R4cpa5lay3tQcfe1TmMOsQYa0X7SYiCxPGgxDOmdnxWgeKh8XFH4Cvclgdn/oH4V0/O2LJM
gUDlU4/qgj8fWH9E+c7uJFA9CHe8aU2U5AJpCfV+KHM61caSr6ba1oXguEAuWlCcZZMlo/2bDU1Q
Gzgo0LPX4iKH+urx+RA2ZrMa+lFS5P6vjmppM4CaDo79bSh2c9ZkN9dEXQOsBgqrxfE0c6FMwOvm
z+OgVnJeOxPMWaoUm38BLP7SWgIu6plPpsqXx71v8CoHWRufEIPtUlvIAK+5/qgfu0IY1CLg8cqS
eZuTcHCl0axUUquDvHasVlgJyTYoCBZ/Lr5dcHXvpL+vM9a+oIxHMo0GwjNuxSnFOgasowJEJAlV
fyxj9zAylyIMNIRqsdxx21ncj3HEZfeVqkOzjbNTZOfv+xrO+OApEEEdj2rUqHxkdNyfjrcgzCKE
Ykf7iijyYHRV34RyYWjVq7/2JlthDosDsE4ajYuiK3veTt0jMv8ZJOo7LuS35IFcjapfXLmkROwT
NLQqHFF0jYc22yKsG61zPVab1/wIAv2Qa1LUptc1V9veYNQRjCXVeo7F3qEbEqWdDMRUAUzHm9jz
eC4K1HLSK8Xg9nF3BJkfbnQmHetb001dRuK0EDyyKOtWm1xqiyR7yQvWNw6s35tyv0Zfco63+gpm
8WvIlmM/5uw4m+W3l8wfBX1Mxsa/zH3BZC3FTYK/DNcA1OZ6vebtDYgaMwzjzh0+SKT5IB0jMK3N
+w2bd5ADYG9XAekWzDUAKnx1waRuFs997etUg/6MKmv2wIH3V0N7GJbzP3ddkMU2k/6HpqDLq4zE
DBg/YKvDAbaEbCb0RV/vcTYUdEMLu66AJTcGk+PjBOmL4hBdANMk7/l53+s1rm3PasZqowzz+X4x
Tchy3D2lJQgcwV1z1pS2tWDsVDMjr/uur2GWAks23c1IqOuEcEh/ZerMKldMgpC2TRVzjnouUGIp
A/YTa1YklFB2iJVePv8N7Gd/0Nug1v6NqzbFNWQog0lL8TWEebYFJhw4S+Y745wFwaxmPl8YbMF9
gJNg7q5Oev0xPaXuAxbAP+F8OTNrLqzjae4GKhyNY9xhQd5hdMfOhcTvncBgFib/mJPI4zyFcdo7
A8BXOhrB/BprvCAR0CwT9hei7k/+8IIh/FuxaEIefmPzaA8bFQKW6yq4htSMHv3zWlspie1PeKPQ
fmcJtsFBPSwqPPMxKpIB0EShOVrOmepv9qIH3UvB8Vk7s/bzO1Jgv3kZFtFGUgkc4+oPG2YVRvp9
LipPONsnhkejqKKS5kYUKC5k63edrAfJsQEvdmZ1m+nfdlqZ3gIYMOFzOn9CUU91bHX6tLyAM3rD
A9eGRH16wJR0DAUqJQ7dB7JfXK5fsIY0/ebtHlLk/r7/awFeuSg3tCza9jeu0H2+uDAgO5qOc95a
/KiHPhXWEmKRTGjuCJ0DUd1CQksKr2xRD+9B4fXWGmTSTtH11f8cGzalWiVZrqnMhjYidS1l056Q
ZAM7ulWexA7lyHBFLRS0d7It6LejHSRssSahzbQhBpj+soZoVnHPSJoeytisjo9puWjfd0AIQ3Sp
wM1Rti3u5e5Qdmi0escjSojhKdWUvfah8hdfcSo0jyLeUzo7iyAGOhlNxwM+5FQbQUILLXnAS2rw
73/53cvu6jIFm8rGJF5sFRhKS9xmZjlC7XTG65WF7/hFUh9E4UvSCF8HYEdTvaDeUJZBHlb5m4iR
/12cydWeXz6SdkdCanGWqgGH7IoFwBnGO9ikEQZhGgt/YT8mb/C0UZCoNry5TLLLcDjL8dlPWCfY
Ygj3DlhHUb4yaEQRp7k9ikXCQQY3yydaNyBvQJoLxXnWZcjnVYCvh9La6o2jZj4dr2aAoXOSFNu+
oi2iMQS3oBX9bK3Ue/vHspmeLsnBWAoOT5pMJBVtGFGgcxiBHSU82jFN1iZKJz44u2FrtGs/RTIZ
FTWRSXTXVd7Zqn2AYSv5xEr+TlGZ7mZIiPenp+ryTl1yNfv4iGH4bQ8E3oKzHvWMzgLB/vaWvQ7V
QIlqD0XZSiVRAajZjCbY1/Bq7s8zi8nwNgyBtwALiaFGMhCZzuAVK+iflJ4291suUL0QREiSemm8
PdY1E/8mXpwyR0IQxwgI82P57+qu0s3HcxnY4sX9GIrEqBp1/uZZGPzHPAJyKWExbEAtVGjLH8Ov
Tgkfz+Ts7SKvp4LScjXKgl5OF4zgmX+YNbfEGRzdXvzD0jra48C2hn1dYIVHSZ44AUl2iyqP+sBW
bTVfBXf44Be+ajMgQuF2u460JMwamwtYZPUQ/W+fJIS1cJrROLJZI/Np+tB0j2loSZ4jyVxvBngT
KAmH3/GDsgtYWaOIJn9+Z2FVxrwuaOCJBgpkg9Kcr2OdKnSiDOj+g8v6Pnxtezrdgko1T5i2WvR8
GSBs8Z9YwtdmXtlrl81t0xSIW71vnqbykSZ2Y0VtGF1hKxIIlWCJ7zk4y5xlsblZ/Om9q48caw8x
/Gmn0RX5KWXVCcCGXxCjqZZ3DHPJ/kD6U3XpjiMxpRD+hrUaHJ7nnm2dHUoSn2XAxTzwJWhYMSh1
2Aagfyx8/1/DvCVrOk1jXvo/UFWnKOpJco4NyjLtxoTVjIvqbEnw7gMqj61qrdOjsIEUq1Jw5329
gIMs3gJJmxQr8oZAIPCCIyppia4dcNfueVpEarldO7SroqwjeABbyEAaxZ2UhwXEbe312RoDTeRo
j65lMfW4t9e1U7jj1ZR3i14ouB6r0eIGGXbVxsWbynqIcu+SA9PS8eBuDDq9lWtWzitOVO9BFxKB
McOQdYB1coZ8G3qUwHnb8w8ZbkHEjMJRlD8MEMW+YK2HNPH5GbdQFZkebhAfOh30Hl6iu2oNlsc0
2bFFNsjWKW8+qLCnwi4zJTEYNDqhoMS7PImRTHtLb2vlxUPRzw6S1nQ5huR+f5R9Z9G9VRojPGZB
ekYK8iXpSy4GtdyhVqJfkWCxqcUdA91A8oOf6pYrL9vQZ4sodEk8u9Snugy2vwApIaJiAGBe9RmQ
1sEvJSmM20/G5o6YOzHLRyz2uBDuCgKeGGK6W5PO2jKVcfHl6QpdUVqUrDXX2ED+Q9V+UhoCCKms
vwih0GPqO7M7x2+NiAfwwskN1tatNdz1Bj1If/aDeSgzfRr/AmtoPtwaINnF/KBs70jlmtqgIXzL
axKi/YV/gWYb14d01mqt0wh6ykb7jJyQpAZuIt6TjADVqk9gbEIafBK1NUxhjBBl00+bCgLTPmRQ
XViEg6aYb2iQOXCokCW5fYsuAxWy7d6uX9Nudb5/J36/z5soEYeGjvoh3b7K2EFRuXgai99/0cV5
MRiST569xyOTA3VllWHoA5DKNBAGaVwKQD1xtjuWxShKCEanRKws40JVSDuUvYX06AraMZcOPdwO
1MfQH5zmvKj106Cjw7kc59o1FR5o6lfxM3a9ZK1TfqQb7pEiZuwFm1l4UiDOjiyainrBGu44zwvH
Ki0HIyZx7bXCfvd+1wGEMt2KrIHMOs5YeKCtr008Ou+h9w0UtWIFwP+G44ZmxlslC32hv2rxO1Ez
e1wES6XhXKmS20QwK6iIsfTUZZeSArVzfNX301UVeQe8IX3lHxKxgL8HQ2KeURlwKi11AzzmMKoD
3JAzyX2QUWXSU5lt6rrIobaILvcXFA5pHHTOzDtlY3tMWIgtzJ2cjRRUJZCN43W0etRiu4feMLaS
IbOZl45U6UaDlSK1YF/Ucq2effj7x0H0Ho3a8lyatkRAdAfKcpZlRxhuYoZza6b8jHnfErWgOoX/
neVvd0RH2HcZfkGOfZMVAxQzc8flpfcoYRSnzHVeG7n5xyKDuCDKGPX2d2hQV9N1n5UQpYrZUczu
VCr9uICW+kdVVn9zJUUK5MDJo07w1G9TPGiOQ17tuaRK0+R/Sm85lyhiw0hJ+eHWj7P+Zwfc8Kze
op1d5G07557VwIs1n88SbWjC1+/GY6/EB+tcb1cQ7n9W+NV20edj37gR/z4slYdiUKjL1d53fBC7
kavHxUyNghMZIhEDxJwoUxFMtQx5+HIu/LdkG10CFuB5U98M6xJTKKNnWYmZ9GxOS1DvpNTIvlhw
+k91JwaTkqjjtfje0NEaWY9R7av9NGSqM+h4ScNwjT9yIP5oGMl3zM0ffXORrl1M7KvIlSJG9dQu
rIf/KMHmB9SAC9U74N6/k4wySWM3UfoAh9Evp4KplEKcVJvCn4u9OlEiP/+kaztSrsHaOJQ3Yddb
pqi+pxkE+qjh7JKcDOfvzK+7ZrCeMUmy0hzqvJ7JmNOpjnOKuL+2HJFxUckzFgsnrOegweFjQq85
P4ZJtijLIim+ePulGVWZ2rkmHhxgEsBIq27nL2URA4ldteV/GERvUMWq+NTCNleopgH/aVZVqgX1
spTcRk2eAtlmjD+vza1tIDgIh279py+a60rKMVDQ8Dcmp/28+Cq+L5TszPkI/gWEUAWsnyPYFpax
uQyMYmiM8Ww24eY1hQfJId9Uhm8Y9raibG6UPAsBuNm0a4cPwVCAMWwpM9l3xjohdd76TsjcQVxb
SByD7ARGQAjh3eqAqQBWsyyj95lhADaKxli1EmPaKrJTmQkl+fXFX3dmkhGoeeGea56CdHs45o7/
UTK0r6SGk8BV/XzhA6KlB7Ghhsy43jNqU8Qc5Vi3COsClMqQp652Z3jpl0aBKQggpBz8rmCtYKmp
QAIJEdzXJmbtDcv0OJhB4EGXeUOxdWguhQUiNwTgMNeNwKMjUPkiEUKffPcNCnDGk/t/lx6Q4wRd
1NMOibVmE1wnRqHoMWiun8GuVWauCCAG02XEaYm4mEREe9WhKMoIx8zdfp3x0hcZZmNeC0127tNX
oFfc38d3PLtVRISyuunnys33L2d1np8RXEi9/c4QoRkqAz3ap3nYMUayMaUovidqr95iu/nitZGF
GgqNrARsjNyiOyAifTTvoNkLGwkR3HVXm1vwTtRjyVP1yiRVdBkajsUrl6zfI4qhD7ALonQfVwLo
D7z5vaUC6GKaZUYvIAGcSgG1Ddndo2P2zFRV0Q1yH22rOvtylmCpyVjMIC2VFTkz2KRspdK82cFG
fWuJGbq51aq8xJ7t9YBFDQ6o9vNfU4iCRRAz4a9qzuKQIy/cJAezJSaDhAOPmlk4Km5tVAk5+3Ei
WHl+78VjPAOlhdlPyIo28TNYxfg+bp7YkLYkEc0H6ilMmVQt9BgXzzqScN4tB3igzF6X39ZQP3qx
4WRPq3esJLcbTLts4oO0V8sPl9W9lDjIFFbrniJ6InHlyNvQOtWoBHv+1D9xcm+dnOmQ4KER7ClE
0hp31TNBtshA5qYf+TtJbrLczRIiSoDN8MKINPLN83wdAkQsQEdJIUovKzMLhFThBUgCP4niPOEM
m5LA28+HbiKjl6qBgkpjKbjpDZ53oEeB9WlS0dojeYmH0Ctz0+38Oc7Q8y9uYUtrhb2fIS0l4wYw
ZEQWf1hOdZFPOqLjl9hdcLk3tH8klXi3MT7WFpj5B7YqFlzX1DswxmGTzJQTEoq1zFxJ+Jr32kl1
Em4etSqeRRDBc2IbKqB8+pMR5TW5wFopZ4WcFCKCp5OlBV/9/GQmKREcxBncj3ctOp25cd4adT8h
Ca0Ty5XOKh0FyuuA6VtloHEUnl8dlCs0704F7jE2908ImteaUB2wpsYcRkMCybusvs9KrGKbfhf9
IkVJ1malKv6KfoHJrb0+vt57EFx4G4kg7kvA7rqX0mRBKaVAGfUUaJZGJRG5qzgPKThbrxk1Deke
4AB4sZ5hTZfnXrQkAc4PZEUmI19sWQobtBQ2RnumDGA2qmQgvv3Hcw+DPM0GTvMW/Qrcz7FcTcsw
k9qeBbyzQfDlqN/yiMrGaL7XKzZlu5C+URZ0XnRiCRmgvXqH2v/JN8rgKHIGvcp9CgEaRMcYs2eh
x9XVCXE63VM6heGlWJeRZ7wmoaFWQ0TSi6+1L3UlT4DSYN6hogP9M0f/1elnMjh6/AznR7TPl55I
0NWAkOeYSIum511asP0GoF7xjVYqzlueHforD5dppYdKhkO079086A95E5cDiHu3nElJkRJL2leG
dAx3Qs2T15RuwOZnZU8OwuppvkBPKQ+Ew4MwP+iVtqC43WmjEpt4bHGy5MlVBfElqlJCpaP1p5LY
Ffeo9091U9I+wjZct+O9jkdGXw8utSHHqAh78//qamP181dhbooFilDuUIdzQnCrm15n7ess/Y6U
7g5nJ+kziyx+IAvNQNnt2yihN8Ilok9x4GtyE1j9napQqEzOiE3hReQS7AxtzRfils+rFrRMfu7u
CS8KcPjBQzg92spmHTt7SbFLMPuEGpnjAFTUAbr1gBDQ7DHjs1gz8enBcxmztWyOiQsXfY4WiRPL
TV9SD5euAJa9ygysXDaqtMfOQl9i5EhHx+JG0YASuap92KyrqGKfPTnB9a8S3G0EaDxFUG59v7IO
/m4Qok30A0EyVhS1/2mBnYC1r7ZAFWOBfoRivHBmerx0qXdZeI8oDMVzzjHtfufKRzsS+JEx5ilK
c7eF7R+br/m6IKUYTm0UBByUU4aOcAxvOWb8ENF1nrhd5mF5tcLTnfl2VqVPJKNBV6S1caTPsmUY
npAJUb/u6P94s0tB1fWXfIVUbIRJ/9+ivEHiM16tD+Caok8KbzkuU8exq37DED7xUlSEEsi3kBZe
K+IyPBiHR+QeNqnffceZqn2o3oxvXSpXTT+187rVFXBjQHusry4a9dacrZY7ypFiOB3xRtFIDJj3
hNUbxqa6yiwHmUd0vdUg4x4eLvlA+OhnkLbvNf0nFaimreGR4hwiWviYkNivjuiqPvActCnEcJw+
BB0FmJcroMDPdxGet1XHeOkPoVnH8yJca/lGO/HGB2Ap/wJRFnIphV86EmgSf22PgmAAeydJFnx0
TMBcUbrkBS22ObtV7vcZNG0B/GL1yVU/tQQOFyaLLRBc/GrZdiGchT6xxSkIAXPcyn9GOmJ0cvyo
SjTsoqPTGbFKLgghM+asIjhJrt5e7GwcHNOc20TAL1YEEIc7Mp9IDK3S2ht/cxKChdOXWD3lzrtO
6resoegviQdL+0RULeMnNwHJoOiqef8r+wJnZA3lTGhs8IXLsLECc/OZpp2UWXw7ZPRFDx4l7YMl
yNNpyeQ3fXgK+HwjHlDMK2MdxMzjobtKyEartHDZu0qFNITV/P4O6+q2bTXMm9j8wtfteP6LgGiB
8oqk4RlhPJgFBZwmZvWvQgKAhx/sODSUHzbFVKDgOb88k5T0Y7jMzp3skFI912bCJSxkdXXdnSfP
FqQkuS4EsRbZwGGxulkCseonHyVWMF2wqX+vzGe1xkb0uEHY/KfCZM+S2q+6WUQFVjB2LOia+Cio
hwPEXZtNswBHRixfi+KjWIrxVB5FekANM7hYJTFIRiLlth2KstOqFnK8ReoqjWNSICyLps5qODOK
J2qzr4P8MLtBR6UzFTilj73ZaiUrwfixkDejZNdnOq/oJWwchLOaFxGW0D+Hh5gB7QF+8/Gq7vsg
PmO8SxUWgF/ctOxR/FERA25R8Q/sopYqUt2ecKrX1SWlvwz0cn+507q4EVF9EI3ZrEtvfPLoddUu
6RWcBxcI3Pl1hdNJq8DD2tt4oTGy/viyek4v9d5cQQmEFsEoVdAc5jnQvifVjNCb5mu1SGLvtQHd
VGiNdypmoyKTB3xcbUJpXCUEE8ZRwozZQpjINt+AZ/N2NCMKBR4Ry5MO9GiNRd8M70SJv4dw7b+2
sexd7WZdp87nGuEBp/1dIrw55ugrGU/GAVYMfoxgctpGOsJc6CbNqGb+2BBn0QgpbUIzHPeOyNiB
6OA1yoDKQSsfg8ryZi8Ju6Z2pjWgRHKznWOyIpXbotB/Ney67zypqEyPMKHWu5jmadaaDJ3XsXOZ
xVCd9bvQ8kjfQd7K2hRO/sCRuweBJ/TOkIOwvb9W46PGw0P9gzlGTyIIoZ0Rng+3jTEV6GUp1Zl/
j1iEcEweoul46FjoKhWpQNIUfF6wBTuOLcPZvbfG2Ee7JGXdsccQzPN0c+zdkiga4oVbndEMqk5E
5bLRp8cx2ix/5pDxArQakx6R16OJqxU8NLCANku3syDPPq2pF3moUPcdkj7w8gxdFSInxZqhWIqz
/A/ROPQlZSCm+Klqo+ktQb1PH4Os3LYXk0kVotG/ZHRBwR3k8FDE4vvi0xxwEudPOXqtuXG+8102
wIy64qQDlgbXF7QhGGlD83qkf5pZpcKIvj4igUsEu3LIX5QCP1ciyTzzvttzLltiBahpBskhVyd/
49KdiSFEefE17A6STCsvtciDqEmbn18fNxD5+vgxwMMNGsZkcmr4DoAUm7q2oWx4wE2fRPea7fd/
ijslC+IXK7rf01rACj7lny/B0ValCbnG6zsX+sUoB1yDSHXg4k/mFZtX4R8CENO3rnfaiOtB4x7z
3ER6qqSAsMGNLe1/8lKUEZREcZbzmT3ZEUJKA80/J4CHbN+3ltaR/QVc3MowkUl22WeLGWvQoheQ
NEkGzj04Wa3NgwLMv4kVV25m5tnN8sgbTSYz+nWjpFxJdQBRUcpiUDNRGiqmTgVVyHPqc4PTDHWi
XchJdfhZ6i8VKPMpW4X8ovS5yl93jUWitMAagowea4BPSHhHsqRHg/M3kdfjl3KoOb3qOgNMEyY5
X+E4mTR++UvoT7IR15UtuSKkYynD8ZCNn6A2A/DxS2yILwlv2eGfamjD6wZrEQvv0s9oPcIoqpVc
9x4hhZgCzfVUZX3BIXVqEs89MZfRtu22o5OUzQLRqF9SltC3FzNjF+CGUAiPeCRns8WTFScLsK0i
gZUyHMWbfVN/jllyBwI/kXthLicCbKXTbAil6paBPzHGs2u1FN+dmYVPnumQkERIhONeQLucJl6L
nubx7OKnJeCShSgXQsd3F6ZWO9EtrzyzDZQ3PFFsIwZLN0XIInNf0wp/p1iQDqXsIns9dS8HPwcL
3pjCeAq/71pUtE/N/+rpQQ6bwVOxD/29eY1VrfddAH5SRDyQifRk9jDIcG1gIAhpoQYVl8R/lwlO
cZAmEC56JJDJlvgYiMeJqltLVuBG3Nn/XGv7oq1k1lJiJ5U5MKcllPWcsfU/XiTVgXsffrBwS0bI
fLpnfTXCT+zkud0g4eZ636zxto2d96uLnmEid7afmaXptCbrgc7dnH/r8PfqA9PVi5HN7DWiL48L
OgAEsZMtHa2ITGkwE3W0fwrs2L3mRqECrnBk66TXuaXs2qMtGYr9a4V8FdyGAwfwi3zT8eu0I2fY
qWg6XXw7LKcQ7gmFMJHg0sbpGOLaA9sprSc3FUF54LLG0KdOVyFyS16ACjyo6sTlyOevvesyDBKT
kAvbBnyPQz4TZF+DLBbRHAKmCl78rmOaoR3oTXphgGUwHfI9Ap0QsFQXFCvVD4onFCcM2w8kdFTa
noDMv7WhomfAOQmN57u+45LJga/b+hlk7/jCXM+KRN9LpqRV3N7MNSI6pz/Mfl9bIPSv7r8JM1oV
ZBGll4dqtBwUdRKxIPaDVN287/QTOTIkZ4cpKQTbHJbIlPQBtgRmpmLWgty5lGnLVlMXjJ6ZID68
PvDJMfCwR4kh7jE435knUHPaplV8FLa+e/6ExO6NiMAjKDGNT6AF8JGnRe0FCeTRi+n5DludKQCa
/qKiv44zzln9iPpbVuPsV/U/T40LdJp+E0fEyXLt4u7SylPKyQHmzlqYAeY2F5ZIL64DnaKKrnnr
oNcmaxHIzggpKKVOa7c/wfKqqwn3UuQ4TFXTfknXexRRBwQ+N63ME8mVwvgHtdetS8HJDxb+ngIB
44pcRCp3YQR+DJExa9GuhY1/o5vU8zqrhcPcPuB7efq9rNI9cxyAGJ8Kf7Rz2YIqf4I9v8nYVgyp
M/u0iiNfdfxEaSXAhZ4jhD3v59sX0eSjYE9aH+da+hMu7BpGrmtrSzZX9dbbDGl+Bmr8IrNb4KGK
C7yxUg0CYMLS9aEg7ZPIlQxJl4bvBNPs+dk72x8GPLQuTz6SbCNFifpHn45prboNTXaHPnfxx2pI
YMVskqZNtsLp0xMhiDgpew6bAOhN/f7HDLb4pxcJ3wZis507wlyuHFw21ZrcgN7PPpKxViFrEpL5
nN5PM04xYxlYUNrG3SFeRM8WEiskgykwwPK72GbFli0vsN8KptvI5TKVJi/9SdTUdpOtVG5/Ocau
dsUT9pgyKDe7NXC356clE++hgDuj9JL2YrO52upv366re+h6nHVVKsE/69DJ/KpCl0a+A8lJbW3X
JHlqscShw2YbNE5X39LrYflbU4fNeCD+xzBrE+C2lKDD2JWBV5j0Tz5pRYqyLGeecuY9v8QSkih/
c4Yuekhq0I8rBhpQJFtytuD5yvJ4ThpCQdD271EuxGUaLVWAapR1ynNQyD/RG4xkvNKSU4td4i4F
/7AmjVhwJdFzDrbQgHrkFUo509DIkUfssPyOTkMe1tVQ/AlBTTO52oRMCrCdI1OQo1Tr/u580SlV
BgullUhrTzBRMxdJgSud9Y4bCgI7TKfmg2r52FhxyoY9yxx995xnpOVcsZot4YisPMXEu2K+cHMH
bT4UUy7hrCdApD89s9IjEyG+skPZRqnx1DW/r6UMSID6D0AcGfqWmesEr33Tgo+nbx5frufr+w13
C7B8uxLjRJJGm1K4rnBnln6088ti03SpisSPVMOfIwNTCBM2TD4OGAb0OiFVr1f+iybm8MiYpSM+
da9BtiHi1cE2dZ3cVgS4vVz5xdIbbHCWWAsXU9lh3FNiJZpwFGf/FPsHPqoTSr3SF3hYK12vdHee
i69NDM3jMlWtS8fxotlNmXVMqJN8BzDOgGPGgZL+dXasEulF6itDmmQxvJDpuf5dRKriok10kRSx
tMvEPtKr7z12yZTbfEunm/rS4HDBd1ee+NAV6oNA30iGwzKK4jlm9CzoC4d6ClhASp0ULn6k4t2A
6XwZgydknysqobHemU6USe58eBTacuLCkoux6J+TvqpiVxxhQI1viZGdXLepQG0Pk9/JEMLjgmfv
H5Xwdh+Rcpn5lhePUV+Ft50KBc6+JrkjPFN9BzLhly+ZChrd3jP7J9310T/B/VWue76EEyHoGVTD
5kgjS2lh35FVWXwIHZUo0Ev66aeU9dTMFJ7FIZUBVcEbYAKSiXSYVLdO1I077jjn8MkE+v9LySq+
klAIrTDnMr22IBkqfvPXseSD9Bt2v8ZK5VmBRvI30Tm/gLhwP9GJPs9Z+Bz/I8aM1GrRCgHTfiE8
8n1YJUeJHXiInNl48SszPMQkMlPN0Bbyy3cLHy25auDWGl9KIXFLMEPWTG+rUAUoNs1hTJUtStSj
sVa/Blmql+eveqfl+4n60Z2DUPDg9dljFPcPk8c7If2hFVk7PPUoOvm+MbKYpuIKyCuj5lJ2KFp4
pWCdk1CPu123vMJ3ii0Rf4T7hASANxLAI8zhc9QHOs+bF7z/y7fb/dc3zud1ovo+cjp2D5jqeN/+
XjtF+YQhrIFWGGR3jqotld+EcVYRGJP00NPSb78dlFSql2ZqHQ+YRnfvaF9mCCglIVM+LkO4V/aS
73RILSPG46unh4DhpNLBhAlCDay1fP76epklpUgmr3xhd99i6YuxCHe4VVHQKWmZgI6ukJiPZezq
iYTmfPAKiDMxDV97QMnL2gB/c4h0m2pojTNX2m6ib/zCX5nalMX26anZFcqegiWRSSop4RTs8+EW
kfpF6cObp8LGdUOM039gjTYP9PWv+hlUyTfLCv2Ftrt3nJmcMM1z2slKqIPD70GPbtx4Cs7RCDcn
+yHmIShGAh9TjVitV36c/4l0rjxh8TBo8OZI/QTEHgnM10IEAwB5js3j6BUo1eg/fn97fsgdBjM3
ELl0nVkHOuxsCm3zip0qm5YPMeG3HxfW79eG61ibKn5UUcGuCQmj1L0QWYREX2OrO0P4r12UUVfk
KsKMMSER67kb3JeXBIBBZFYBN8DRs+JDHQplpbWhEioJd4kPHTJbqN+F8CsHssXE3uwEHQZIKP7f
efJXyCMKjGDOt9VdeQaY32ydanxA5a1LrsBpir+3FW1PRxJ3vOuD2fE3NV3SmV61F8M/Vgb/HNfM
HKLunf5hsYOi9qxoq/qg9FCf/F/sdpwsg6MvUoi7DBmI9uv3Iw+kJvkgKlq3ysI19Ak8EHbVbWCR
oUTfVLPgIAZ4GgtuTnIGmMrKibFbCXBbywcIE5z7tQwBdO/ZGIQkvzOJqpvGViAjrAoGIXyXchxz
7bA3Xnm9eNv5/RH2v+e5yl0yqL5a0BF/agu5jC62j8PtXdREb915rWMeqKPUbiBp8sPMS8lwpFLO
nPos+wP7IRwdURtPnyYghvIr8vlLjxKQBaMNKnEBKP/GBpmQaIY2fkyyulJHnqbZrtMD8BfSATRN
jd6WwvX4sOS00A9sIw6SpV1LZQ7ZYSbJ5ltE8U7eiXv03JO90At3/NYYmjt55aqOFaLHAf6Bd6G2
bEXJwcQ761rJsFCEjJyruq0oOp44bsXdnyq3cI69hUnLvum8I9SS9DGqP5qjWd+9EtBMuUlm+0BO
zr2QnP8+jAVpPQWG+KJQfOzSYeMuq1GmAgBn+69NexGZDvBxvSw1xEwc5LvpXtm790EYb/G1r5YB
bkYBvDICq8RmifWc6VE3QDO+Zy++5ZnIWwKrla2cJX2+29YG30uHmxP84AfuztsiiLB0yT1FnLEb
CwCgkCs2F411Cw3+z2BcoIkqiZIDqnRRnRCVzaXqC3VJwKgQ8mkiZkgH+ZL1i6MGzaxDpE/+TE8v
4fxgHUnMkbQaUZFTA7xERVlkrAM2Kldg4JPU2M1mcyBaXDSNnbsK23DwsDp39UhJKlOtW4vNd3bt
shHugt4wo1lMVI2hl3HZZFpWIp6RIgR4cDIJwINcjBlSuBotnDE7FTdiXhtrj9N3O+7cIk0FjiJN
JqlZKnIJEtsU233tb6wXIYduk7IDwUqUNbpVsBfe+qb/hBev8UmqZsIX38JI7nrlxuCo+M61ciS3
PCZfp3UCbEEX7v4vmjTuflkP3E8tQ6qJp9VWVL9rFPg+XuNJbB4ephJJ1ro5XOLI5jKAxDrCBM2p
qVl3wdaskJKkodqiWYb7Cy+yn3acWGKIKgfuzLMBEXTJ4TqZV9qwGUX3V9ckPbgds45LykFvfM21
5pvx9r/ErusHWdMshdM/ZbAuZizZUt2ee4V8OVRD2hKl3xJFcnmHrMGpmNZm1cmHikQ4q+jhkJXW
oVf1gxedGHFLLb5yseuvErkYQKhD6Cnd2/0ZpwerRvXP3Qa9Casrs4SOvYK/i0nN65JiUGIu6m4X
QmgW6Lu5epaJ4kjUnHn19iiF1TWceCWaujrzy4hnYXiKsKHIKZfD3vvgknM/AperYFsMHKbBUh6e
gAgwX53cTemzvlInHhVqWw++avpRexRgTomj3hrnSkcIj2G1NXJsnxVPASDkHydGyDIaCGdOYKQM
37kVexEKY+D9ZSfA219Hl7y18Gc7vfdSFHWbi3EVDAoTqju0JQ1UGIeXz7Sy6L84/9gLFQoz6NdP
+A2HtewpEzcrasHU/u6DbWDZj7J+AAow0ODj5bm3iJYEvdPxWyMVr7YgGhBW4kDJCjq8//dc7lrO
8p5TrbXWrz2/4thqgtGwBuP1VshLAhgixne4g6v9qDDZ0eLqtJnxTmbpRU+NzFystncbrpTNSUja
ioMJ4Vn6iYHi7C7ks//FtsyNjZvf7lkNQEqHMaOh6RhbTtrACvl4GFAQR1jU4lUY8nd72XkwI7jq
D7YFLmmd8EAwfM0UkKf0NBLEz9TJT0W8QzvTvzwDeRzDaPXre5KQ3hri5XbaYFsFuTY96ulSxN8h
1Pb3NEk/o3JEcBfnzbAHbiqTiSYyvu9S9/nzoP0h73tfk1QOSIvh3G06xsXx/v7XIZ/19qBoHHPE
Rn8u6EB6SXlWTdwhekNS67TZuADPDzvpYFcYhZhJg7y92qOP2AdfpMEnnXwcCQcEc8w5xnRbfuPu
wcDrXA/jBlrKogiYESnUsROTxkNOlZG6A8rG26RNRSBeJ+GTKpr40dMsHpj7SWtSSgRAgzEWJ+0d
4GDjGzHTDKGyXon/a+x5H/8pNjrb978VbB5IcvjrouV2oqn5lkFzQofBv591axE/T11IN1NBA1AI
lpzNq+3imtaO6V/PyM9pCdx9yE9Dek4gyV5aZXQoQq4QJ/dNE4G6EyUo9KqNS3XC5dZ2PcFI6xtI
rw8VvERyfC9eiXGoSB8bOWBu1DOxxWKSOQpPhGCg8/iv3bTHjamULaJw+hoTU8mbBa/2D8gyyUIG
no0HpMrY0cxXSXPCnZcSn8PBWSPIQa9CWye5FU5anOkV0P8fcIutq96Ce+jxiyj5Zwjcn9sdIqWU
E2wJsrcfGtFv3Be7Ig70hMkCZjguw5xzzZMlZVqJbY69tFQW6m6ovfyFpUmYMefZV565A4wgM0Hz
iR9djwLu8dfPcTBRZuXKT/wzQvM8zdmzHX7r9YvxeP1+LbZGEQFO76iOKl58jL1toqsn0HzsaZSd
Z8jTWiZzlLVSK7FS/P15R8C40tWB3I4JJ8l5zT/0LzvMnOJEUCsQWmaxUhKa2Qk4RmA6NVe3lVAC
qBiPTSzSdQpf7cnqUjTGoKqkcfrWa8Bpf7Dw5WhfVcSWju56g/FySfxaCS2pSOWUH2IwE1IXN2Zx
uGSCHH0E9YeADNcdRjJu1bBPrx+bkbMzdAX0daUsr+Iglbp5ewrnMVqYrrOe9Bdg+7wxWnsy32oD
68Irz05xZlDxomqmjzIupnRmtjUVLMPa2kmglg/IibEPVtUFt2KY9voF5c98Nzkgt/fpJf1FtqcN
KfwxwZ83AI7D2Zmx9hevaxmRDLBpAO/JgvoiXwe5pz/qA9lLRSmAJ3cMvVv7xehTYadEPBfyYpG/
4xiLwzfhabCAwaeEBX4p8kkg47s51wjL1RYyDFsy05ZsoH0gAd2xnjUBIbesHuK+sQc+0frpQ15n
wYeTU/sMS++UU0fkAVpUXEtatdlIvSuljF1FIkR5F34vXrEsYzFHSf7bM2t1UiMCb4lJ06B+Yqzx
6a/FKoZ/6wQrI1Vm7EG4DfK0zsChwWZKhlDy4gFh8/eBXN19GpVy/AQpwyiC0A1vyD2Sra+4aBEN
aEJ5BYpCR1x6upScsOwQZWYeix3SMZjva0PSil32XxcEM98aWUoIUX6vx82zJGqsVtmPY+yUioPk
APHMsFhq3+MLylxZXDSm4mEW/P6nq6Xd/48Ub/xBW730UGaWQxk/BRc/scybYSdw+D7bZd/8tpsI
F7HBt/G9x/G7JeqA5ii4KC319WAIDroulOu8OzVDGAntaT2T6ijxLtFMKYlJhw4/1fSVePNvBPhs
NE50e1Nbj1Lyr+LDMZ5+SNQTgBee+BoFZ9rMeH4W351QEdtNa+HeMTfpY3uhjwI9hDJkvO00QqQS
h2UE5vcKxru6RGAAGwMexnCYVxP5UOeoyJcjCasXK4YIWB7Hg2P5D/kDkp3X2LLkG+iOpvwgsEry
zn3cGbV1Bo9VlsQ19CRkmAvVYqvj9dIDhZTLasQrRj/TqcoO54h6D/ew9m2y3pmSdcLOU50J5R4k
ghjmFSZY2/H02A1XHNtf5EHj5Rc1SyUse0q3Xgg+n9ZlU5rw1tbj2cg4ct80sX1dQXl8HqruytzV
WtpUDdGN9KQQvY1jFbWauQU1OR6w9gvi6cndzOhRfgF1yedEq1mSZL6O4iG/zBBCpMqKib2/Zj5g
L0Ao10wUjIXtTV4/jwX9pqdEre6suMmLJFoTacDtdrxVkH6JPTNsFpWWBPetfXdwilRrahWxcN0N
Nb+eUZNaGgM1CiMuSyBUAlMhdTIXSHxi/2UI+Be11rd3OHWMBZv52d5OICa2YNuq8+QvrxvFu/VJ
3IYs9T2dqsyU4FX0rkoyEgxYieQsRY5HqYz4h3VXMK8I6R/kbdg7tW0K1QSGgxkorzXVC1AhxVxc
AZ6VRtu1jmO/MYVDvXqpnz5bKE01itBaDjWLMOCqyF9Gzcg+cosZdKDapAGocD+kssvjYiVNXcrq
we36/gCH8gLQ/k9csDST3R3euT4q+yLcBORg5wcdrklRphNZX+Xe3vDOm75FUhi8KEXXGKevv6pM
bF9JuLcqcJaAhPNFuQTfqfaQCHPj1dJggqDusNwgGFt4+6qrdXox2hWIIyexLwdF6dIf6lnC1TJI
tD4Lt3rDSjbqTmmA+aoU+qzNU8NBfCd5DR4siyWty4JyCzR6uMXLsGRhHCRiOXOTZHwwbvfMQjFX
wrmuInUvrwWo/nxsbi5o2dKQQlVDxricQrDBAl8KbnZBhUDs4v5nZfhBepoOeknyhfTi743JRcFL
rTam5dN65uFja072beumoc3uaEPkRtq/6n79Qh10CIfYwgnAI8AAQwpNg11N6H0mtPCQw50ICWU6
n8S1+swEJnLFvSrY2K0gpMiKQ8JgLhpHz71rYqm8OL405UUMfFcFxD4bBJAM4ui1oUpvcikylXmc
idKNjRe1dmahFEqGYBjvYMat0zkssS1DiactrV/QuQUatTcW8W97jbTumHFv9OroecvufrezXMwp
WwFBjxhtHjnVwk3V6g/zA0k+3LcsHHgoKQAeip0uGZDwbhtsr/mvLGNCtakt/d2C2B5PLbx1lRY+
uzZaRBu6vBetunXlqpVKCewmtpY7vympAHj7GGWMSSGIRaiVkOLYASJ0MnoJyb5+ztrdV8eYoU/5
m8XrdpYVp/1RQTn8yTPnzS7wwOmAh2VzLApAhgK2jkWkS+kSKL5nQeID8pwZCkGPShtQ1oUZf+pC
3+TUwbDZ7NzGAn2rIiSQ12NycRRl7eORiEIP9iHZPBopD57BN83tm7kDeqJmDgf3xuDQpBudxaY7
UEURt/U6fEQy0zcGWasIHEH5+WaunPQKeFtpwqhNVTzUcNkDCj3yE2QRPypDXw8epgKel5CRmxoa
xr2DNhzDfpYYY50v48es1kfm9SRh1ORnf+IsClxjmjAa7gS/WuedQ6Iha4+Xk/5oZGoB/Yepp4v2
i/m4A82YvJOQD5wAsMKX/t19o4GSceFo/LoIcxAQY+4lB7ltbdNkc/AuT1HF+9PeLClFBdyk/tsv
Nmt/rokRcE1NQn5YKbrx+5AUeqq+CvGK7s4RAI++U5GD+d+uGT+C+aNw6CxqpI+f7Xlvjy7PV/mp
RqmOE9Ua3NNxi0vAguQP+F45EehcF6NfA3rwntAPTNlnacY+QiVnsoz7QIda2E+qh8kLkwO85yNk
UUAFNaob1kNExUMgtanwBiw009Pe5hisBinxM10nEZ9liIymnntKEtfUxIpLvZwaVPFeiH4kZiy3
ZjnNtIiN7XFMYd8QXQWlbcNozbB8iMJOpymSoipiTm15ivMYUxZEaHKO/PSzFphRaOuvr3jPf0ot
D39C8DlxnxXBY0scz+jK3EyaVXmRVuYz2KNhNkLkIqHlu6Z/98efomHBNRenfPOfyUkUu6AGhidI
b1hih1tkfBSWsj00b31yX1qlUvhfR1jMciKBvf7/JRNATqXQRqs8mHUGCNvM2lq+vvFdkmNNI3AN
qLGrjj4A0vEPXUWV0KPa9uqKSpV5SaXn5vMwWEuEiWqZuNmTpiz2XDoPV/Dg8NanFx8xigTpXfXa
maeLMD2lL7GQ7Xggv2J7ibi7xwyOmpqGQcwpAUb9QW96OPsa1zZzzX+Lg2bcOgndJyzDQFSnzS4Y
nQQg9ytgXw9kfg98A5FcGaWRSkLyOAsB9vkKmY+RabMPYTV9wWqAyWUJSyZjnI05yhosXo53AbIv
vCLuSmzJ9FHfYdPeX9oSh8gBei7m0W55hCEDzxg2W/Pon2sQlerIW2BKWVKzwyKnRhW6lODLbMIC
b0qBPyUK8sutoJqKo19eK4FO1ttUSLsC76AzKC3GdklFvPgTqqzd52AirJ4uVdDN25MwlD8TsHVX
6N5Pxab97GUYH5Bf7dO3aPyJaFNvCNzARAbV/FkBytancSrFZeyXo+l3A6ov0+kXkV3FKeS5jNXi
w51OV04OXS9hqPetRkUkGJWAv6AKPOBupEEYA3c9IdO4Fjnnk87o57QwV+v9h6Nj0EL/fDRGHtww
yEz7MxLEQiJ9bCFWwC+XPTRtBr/B2S7o+kVFsxB2im61jekHVb/iCUFsxdsSmoXmk1Do44KDHcC6
yw4WAo0p4oJC+Mcei5epDghjzvEdSPOwY+XFxYgw7LCp0yrkzm3ORL4ys3ypyaJ4wdGPJT1urn/v
oP5NDf9xjM1YqGAB/F/mE/6wT4eQEyOOKniORmW7bFkfKqgE57nyW0OhnSNCAD/K74JxOWoZTVxY
5iK9saOLpGodUBVkrzaD0Q9RGC8Q0wesU2ucdp113G0qQSP5DglbeUY6PRogguInlE49NKK79Nd0
3ukdLtP5fECKMQ/LVoxN5A9Qx1FuKRFGCy4JKmczNgrszwN2ApU5rkl6psop/V2JBk65UOiBB/Dt
RyykJtcECoUoui36+h8faGV0I9kqrVfd+GMhRRu8azb3fOcIzh42sShPLo1A4iWOKxzw2Jea+iGp
wFOteFtQ9HPbREhTQsW2EdIQb/5XA3MQMES2dWTa6d3E/uNkOVlSEPNjbflrTEJIZGvh5m2MN/fM
0NwhQb2NvpycJg31FKkRcBK2jHd00xhyBZsYV8AaVoXS2y4UmRYAjJHpPnsuVQ6F7NxLPnBrHf1d
T4cT6g9DdsaEavjyzmhT2szGa9+rstTGDaYPF4wQ3wJ0m7/aA3TwVBcimQY9sracMNqDFQF0smh9
J/oPepTh9A6Kj1haUlI6uLJ7+HEgLSi4YFgPohT+g+EpAefzgoFZgYSo3QfR0ngkMHtTKwiQuxbs
TsPbMZP6rn6LFCMGcFlFNgH78mAknSQZdzuTCOd5IjreC8B7H1T9F9AVEvDAVpztCzzuoisLfN80
JP/t0y6ARMTwlyzXs4owOyeQD3rDDcgR2TrbIKy8uGf2wwy6z/xeKeEB9qW3jfFFqrNlhRO8OnpX
wPU1Muqnj0Xd021k8LX7GC1+oSwCoWdDuH1iK9fy9xGqIQNjeHNYSTiP6W1qA55d2rksMIJW47QK
9X1EtP4MfOq58P1/7LllMJ5ehyRiQYaHyQgsCSGH3a4rLPo4vOPKDZ5XxCKaE+YeoVLZiEum6Q4r
/hOs0K4rBMH90/fpxANb3L7vAKrK+AI9MCOrylGKWnlFobKxrYWRUP6TIuMYDwWbrlqLThvYmHKh
RrGdJqLSwHEJ+RJ8rgahK8MY9XWfkdwvgIb0pfMf6bSJXsq4t0LQJhjf4zc8lvXT5NzXiCHX5xgF
HFezVa1wGO3KKK6oJNPxOaLGs2PwOnMR/0KA/k6Pt/zyal9Nc2p5Uej6c6G6A97R2EB8NNQtOhiB
bg4RzqXnlYaNhG7QqDAlTZqoqEFWTTWWw3yAE8MWeMhCA49guZZZd95dCEUYwJMNB0tbwRNbDXvA
vAR6nyogin6nTmlFvSXmRYVeXCkWFwBDQ/znvlnCZZMi+HUq1JtsyRXZrOIJhgaWOsj+kQX4csmf
rIX4z8DkZpUP4zSHN84TF5lOktwEQdgXFlYT2VBTYFvkXOOik3ZdlvnkZUpBNedauSMCF95Qc3Qq
wQWYK0gX4qO1jONOv4zXkaW+Sri/Ti3LQKmwDMmyAy4GSajOEGqgtYfmm1fb/Bw2BoKCHun6rFxo
ubJ1Xwg1X6hk4uiw7wzyAXXNh5emWtzVt1ER1zK9U4uO5Cza8AX0a2chkBbSxFDhtbS5A0hNQ9JM
rFGBNML0+9KU/iRaepEOzVGUhlXzIBisBq8gZgoTapwT3V8LGzGL3ammPKK1X1sG5FsLPgBgTwL6
RdftS/KwFmQxdcFq7pc2QFLQf6dtauZcO8cjoyI0AoQNapzRtlbBqJMnu7pM+Vy7NH+EvINxmozE
OarEC7G9l0C4s7aAnY0CFRycVX62DPrdJbedvfzBW3QwjxbjnUs7kOx8mPWSjiDLXY7wX9fSwH0E
g5ibS8M9yLPusOgI7aYU3nVrzYsFbTqamIRkQJ2SoaeoY18YQPwnaNK0Y9cyPPwY7izKiwJByaep
J6BLgETRme+4WnQMsDFLJvgsUROvF0d6xiNQ8MCgoWyOVaPsLGu7A9lnPo1i8q72zCp0GX5553I2
WdRGf3w1waYeWa5oExrpFxJd//ytRrDWQYw8n1rpC2L6no08Da8fA6YhU8A5cahlb64mjFweO2d2
+2/62g6N/tqBCo3LjTsXEUVsRZgbO8nwOlTobShlXzjKM1uAfqey2BhWSN3uo7YF/ur1PVWcXtp4
NWa9xeCQ8yrDZENkUWisFE2vdmj7wDp7JTblMbgMmmTggQNU9KD8ZOkwHvnifPJA0p9ws1+P13E9
2GcWT0IkrWX7WlwsqZ1MI13BxrPlIuqS4nPXXks1Uxdp+Xjv4vjXjoWJ+g0/zjp0bKOa5iRFJLEn
IIXogWOJpl4awmKjuwA1Y9C0LZ0YvyzHgDM0/6Nvl4dYU0cbWI6CAdlPRxnSjCNL+i4E5A5ZNmRI
yRJ/S/ZJcBxX4OrtEBIntA+IJMlfW13h74TyBP97fPpmiSrUdHl7iP+lM4qZA1Uu+vB6oaVrnJNu
SM5i80XxOKbiT+fzU8N/pNXQOkpLIt7e7367dxBGcZf7tbf9RBxZQjhpRfecrQYUVfye88ErjU/K
OBLBf/aNoloTa+UWgrEEOvvu/BjcR5WTUvc3AlUnWTAdblE9VQmhFSuouknbsD2IF6/74wQlMNUA
zz164Xal6TMW2qNJLGaXhpTvZev7D0zbjGbugfR5sXYILbjzWqujOEALsWNrwPvNPDbpYucYOFDI
1Rk0eGZZiciRD2h6XtdpXevrvA22MPq5rxBzxsyGuZTAhPBYD3ttmYwTbh3fdnhWBEJ9w2XbBmn1
5B6uKOCGm+dS2dQHDetju55RwMieXYJrJvSDqOgkdT1YqBOdJmjDb9eig3gfFplzasCrNSJiKDSw
weOE5OlUvgchu2h++3237RTk1aZVugWBEPQpPrOUHp5WcLJI9bHgLZDf6ds9mrWpzZIYucbPAlLc
nBbVCcmC6N/nI7JaH4gxkAUEZqj70xeJgFkh488nz9wwhTrn6YTXxMMJM4luIWp4mw15hndF4I3M
Qrd4A2YdJmMWf0GDnrVZ8HCS4pDYKQpOxq7AUutwMCsTWy0HYFD+GqKeBUMmtC3qkKcu4yLDiJKU
inQik0RjVhnsKwDm+OIv+ZDGSOQlJvNIQDYWsMtmcOL+vOgPpYI9dOINFRJbLjL66xc/ZuZnlJ/j
/V7PLaBVJgC+ZZSFgRRY2Q3d/32WFiLS5gbxj/tpmn1k+66fH2UCCamD1EDZHE/ykPz5ZcjggGQE
YwXErsEOK7aZzd5A8SwEaHSaV1/BlVMf8JiO99uZoE6Dm3WOGAx02N2ktSjRlKUk75TgahQzqp2s
PoGBe+fi6QzfC8ccd8lUPGFmZZKHqjpsutzgNIX1mNKwiKzPXYQmgLzZUuEGZq6OVq52dctrT5LX
ji3UIsLmMBXYp8LyXHaV90PUiFq4yuAp5I+GP7CMKy1KlNDKPLI6fNNMmMaRUKoxvZ7GtKaMrnzk
hydijHJxZjPocbnQYAQg9AV5vRxgWgyYIQkYidDltfnSdN2855UcBQjMBPhHqZeE3jIg/egzMrR9
eDA5u531oWVdWuKa/mpr/p0aRx+SV0/AQouosAknx2Oc40q+FVsv/WrdkBZg8t1EoGS4LcGEOMif
+7rYSlcaGm143aDJTKZczwupV/qkSgftzbS02dOqbseo5mjuqkBDZTq1qjixk2423VpG5jiwpdU6
tjEL/z+XA4uEDA7+ZBfNJU/jWB7rzghddHwIqzoiqNSd4ku/kjB8SQRAaHBitKB06eb0a3S+KA2/
buhlYPSFidh/5yVIVlelnlhvdREoohPItvipn+aelVTIqSnVThKhQgliK9j7oxLxHY0XFz9Bnhxj
roEHE9sZhoHXH7H4wGiWx243tnvVWFTbTf9GYlKC7W8dOWFSZeiPJwrW/VkS+g8EyyV0m8JGXbEV
X0wRLlyQvoy9nGnl7JGpMNSd1MdTJi9AAxrLxRWrsEhrAk7D1DdCSBLQuTVQRK086uaU2OSrbTyI
rrzuGpRnTN2AkbeuiQ4FNNeIT/Pu8EroNj/uiR/A052enJWnZRYRVAE52NBjo3Bsb4jhTDP9Akn9
pwEjPVDpmRr1NMGwDfZ41wkDxTtHxxskk23XZvwYT+R5346y0U3779pczd4DdJEeyfj/88Ch5tw5
zoui2GFYHNjHEgzhMs8lmXcUxEnXcMyHea0trjU6Ard8eHAj2UXI1JYgKV5n0+C+/1qj8CHDc0xK
Hgyzwp/dRaoV4fR9hyV9kEmeW480OxMjcCue0W11TaRuONw18ncBrGwcQvTchIrRma/aA9yuOJkh
IsaNDf9Nuoo4lnoYPKAecj/0A7mBynPh9YQwHIbwXDScrw8jsViDHuk2GbkEUrG2ajw9RO7F6gq8
JWNSLPrzS1c+RcKo6/jdh4Q7i/qOMfhgMAIYSISpU3CFoJuYq5bNIEd6Oacna4bLVlOzCTW3p8hI
KuaM7x1IfzvOYpaJy8JHbni6hXI/lj6+HsW6CkQ26LhU3w4jd98cIKLQzhr5TN4FaN1XXnrjGAqh
B0pRQyxKxRLf7EbihCFC7Kjg2NbA2vSN4I/fMuI3usIKI5D/g6PLrisGBpgtnS0MIWDIKLcjhaV0
Qt8i7Ab/Aa4kIiVPv+fj81CyQce69ZhC46wf8AlNyNGmBX6+c+3A/WlrRKx07tBqciDb/gsc3fOz
/AT5ki5dHU9Q/e5elXfN+/lwQkpnzKVUll5PxskXFulIZcYgs5G/PgHY84Xjyzlp9yVKZQ1eQeUY
ogxyf8ni0V8hc5FyKlOv4rWG2DDV/wvyGxDxr9NvzzcqJA+Ue9xRJFfMqKYu6zwDvNvCFkq8CQR+
9D7SDBOFeekHJAOP192uZqTH/yDcN9FxoAYT7Snj294xKmi/Q/CwXiBpPjwMJE4K3joSKKJp/mBH
eB7nQzkq48QGOyNnTwuyzxQEZUqkX2bkQ3CqC5cT/IM5Y/vkeKJveLxsf4pjxskf1ypSMpO+9a6B
JvywKJaUAnJwbdKcurAPTWyPsbSlYPDjaWMnmCI170sFEi/lHbuJshVyE3WEzFxq0QRLnu7ETmbE
cPozWsBVwGh5YMwyPmn3czvVS0i4L7BCybEUAoeDTU3ZXxuHTWXE++Iu2ThXBhO5P/0yd7uhV75G
JbIOCAeluTLJnObneuNvaSIv7rCBBMD5oToM6oOl7z6D8RQraDRMGpD6eoNfAyTgpb5vU5LsWsXY
HOuFUm+VYKRZG8q/FXvyACl10iml+PmN8XZ/LXnEcPnCxm/AeVUh1n2NtH5hArS23pd0J7UN8a7F
ko/ep4iiGKfDiUhtp5hAifXHD8YUt8GmZ6wnc793v1inP5qjKflZXs3cCTsXEQqarpu9L5rUbFDV
9intJFd5vpxq2fe08aopx2sGBEWZcfrYTRCFQJVr84PeLIbbleLMhmZxIo19U+tH1FGiRRtwJEmW
jMZUpUHXdqMazHZiWnCjaaYJ8ZXTRD2SUu4earT6KPPCGvsxmDne/P7ekUF12EGapOdbuvKIXSse
LXsUb30Cf/8rS0MSJcZ+BBOd9yCHHTp/IbZNCFngoIgnj+VrKRxmqMZloo/cGI3yvZZd60PDnQQv
iIsefjmx4UPWqLVVBkdbpypyhtKX/6mveYTaVJxpfP8dW/wRGPLFiZcmpRMPRK4kly8O4XtNDyyp
Efpf08OmW6Czd8IPhwPhjg01Pe0vcxGFITUzaMv3WoZEEHzxG2p0z9STgKIHlE26JEQREgRgkXIW
y/YT7Q9ujfIxAGPbN0LPDM165jnApVJ+6FWnPcgq5fnyFYtXOfHGalQWvRNDPZy3Ju+8+Zbr1gKk
WlBOpCn17Cd8OqmTgJwWGBAb1NvQ+iKFSvD1PHQxuZ488EMVf93lZGKg+V0zunHP7ZyXHS7VLGlr
Ialpmi5dTsq6+AcTtY+iWwZnAGd56S/M7RFX2TOJP7TQacz+xQ/1JNgaAmEqVpFUO/7H8wjoFo3n
7CITyB9f1p4QGMW/sa5LxZxBfil7TLaEhFrgaAx4yWVQ/aFe6CJ3tBv0bD0vwwk+RXlk+MhS6dDI
TkgiV2cV1LCLt0wBt8KnBowVRx7tKZoPDD/JIe9sFtwp1PZYvdCUXIcUYwpzAeqdTCXZ5fpGk6Ba
U8IBbttsF9bxuC5sl9hAoTnJ2J+u6AWyM5a/RKLpuEb4NUKfmN3KEWO3MsMo5Fx2mcC5CUrN303Q
/rQOGmvi5gJp18lYz5dFnAswbrSK6l1PPQIq9m/Mq6azGQz/DfhI8c/gBFfgf3wUQgCNT0hMfCvO
el3iiXgnZfT5O0USHUVXxkuXWDLJg3qF8RV6RvEtaOPTkLvRS3arrskyCoavI1SfIROv8SUHwJ99
9SU4RWJzpRlJQVQfLq9GBHMxVfJeRVuZxKPjE2FYiTvocpUSQcILOQtwjjeHTVNGQqYtoINuGIHu
7aHLfzYHCnaQEqExsl9P2GAGsQG6JbH4zCdNP2mPT9+++fdU6m+isIPvX3S9/8IIiZhj6vXrMKt2
FuP86f4u467tlATdZsI9tcVnGh1ztiySjZH3JFVP3BzrSTfxqaJ2O2+EmD8S+L82nhXoMOQYgv2k
grNvIBZ+PhYaAyfX67px8AyWLh8V5OgjS8ZBtNFZ2aWgZaCJbyit8htmxcyA6baaXWXCJM4m0x/t
dw7As8g8c6t3S258N+skUkRnlUKa/nPNU/p3/DJ7fZs1euVhYn0m5fzssHRWMLok5EeSTsXdbnQV
0aWM2q3M4KuS9fh2XARxjf1hylIZdFep+S0Ww+odi/mpks8kX9vo2b4/YwTEQpb7ihlyuoQ+jysb
Q8Sm2FsgXggROpeO6vOX/L19Z0Lj2sPas7hPAwq0OTcGE1jl0nZ62VqO6AqhM3fDdhZd7J2de+Ib
w3spE1IgpGPnDeZzw71jVJBwYUFT5MkadH6uKHB863JPqp/5fhLKzHKAnjw0R7TkH90KDS5/Jo2u
zFKUs7NhO5H0xBt4f2Cdkq8blz94PWa8g1FZUCwUPpQK4hmf5D+FODJ54ysHaguPBXyj2EDwwtJ4
7KoZcmrqlbuQbt50XposZ3fscLuMHvrRdQFgQvLYcKfTjWa4wAj+8tZgmYdxok+0GzWqSaczFOt0
Udh2n/XQR8MjgZe2NJHQwgpzD3yDBAoKEtSljLDcFFIS4t8jYZ5fJt1bPfcFzJv9rhLSF1b4mTxj
iayWoFbMRDAVok/gHeL86WNhcr9LVrMSgh2FzCYccZksgSKxoR6CEEV1iv7xS/b1gZzMrlNjGXbV
qIkiyZRIondfuo7S1ffBZx/sPek0YX+S3iYZPoxMt24+Y4zEK3sL9Php/rl6oDQMdF/Nxb53VvmV
lr7UZdKAhhHYd0pZArlsZQ2FXMzxlXuza6cS1Yf28aDbb5VuQuqJWccYe973Lp1JuslAP9TGnxkm
xSBUW9DA+VFG/L2mDuJuZzgH1LDbD3GeLdXAJoUKU8Yjmy2PY559naklDvBZtZBFhoZUG/txMP05
5aEdx++foO1lm/xUpMjaTuW0c0xLVePrHWbzHFKde1OYc3oS1JDN6WYdoTQ1XWugAk3XJbQ4tmJb
HnWvDgDrcnaPrZKzBPxJqo58q5rDBGiFKwR/+LcNPMtPzhmQ64AgAw1xB2b8novjEHCRrFqa5IsF
mUp3UG6711xhneNwcMKQk5GesU9cfjCebYONvA0DwnP/T3Vs9TYCbjjQzKpoYwQr8Zc+7h9GSc6+
cmQY9L9xNNOu1JJrjLNaWtOlHV5n26Jw5u6+BalYLhM12pDbY2CrpOYirkwwBdjmJVGRscsKV6xZ
d9O3gslYsOtUqUe1MhJ52EovcYfIyoiGV92HLMmfG69t+y8h2J/5eTPNfANb5ch+IUiEYEHq6PqE
Ns1bP/7QzaKt+ZJt9Ui/UNv6S3Mo94QXy68zyeUp08QpmFvPLuCFbaO6weacEr320hvqUosdvvvQ
ohKoCz1CYSqtJN9Vw64ZpoiJfFlc8/QK46+s5+xwFGtRDsLYb8S3orXUqA1wx9IrTBIBo3QEQddj
J2UvN34j2tT5p4Um6bUqTVwT9le3fae+sA+LPY7U+vwIa2X5zqZ1hhnRAcD+A2aBB1MAh14ii5qj
7nc0IVbZo9VhAK/MVw4oHweSGLrromo5aiNmTzUluQreAhQ0CeUkaC9IR2NNLUUbtf7n/9GEhH1g
3qWSKqLP9qNu0THuVmUY/BBQ3JqjOuEHrTsY2Wvy54C0CRkl4/J7NQsoBn3X8WC+c8QuefKukFs3
npH45Wgl6DAHvtK0808MurBT5CukZdNlFs9Kp/46ctav4RfLYc8MnuQEHk+TKSgMVO8V0MVCbkMj
TGzpXSvpaE1BCpPurcuJTyIHW9S8jk4ODIrUThGN1Ms5NqhEKGs3dVUoRuiitS2BUKcF93a4JVjW
WftTindLArf9nMWourwOnhag4sxAYc3QW4mzo4RsjTcWis1LiSUwt4DAMMr9ACN9/4GSATy5MXyJ
dLovO8/odv2nKdSGWSRnef3WKEURs9CMjpu0OZIs6nNMnD4ok6p512JZ50XlTUv9KIjc1CmSU9Vh
z8rYZRvNWxz6XePMx48WWPFUhbQJWhK5oCJSl5jqgVi+vZ+0Ro4BmLl43oVzCm0i8lJT5vuevdrW
+zDY4j4zQEml8X5U+Yw9T8e74rdFptErkt2zj4epufIZQ6942q1fmqy/zPqa6HSSeKgf9lHRlNV7
xBLTu5LHZQTtFzVr/djP4gpbJm7dt9Y/7I4Ag3Shhur9dphJijscMYVbbDoByLzg0eN2aO/sh597
oTLE2hE66O4qonBHScAeKlGJq7u4z7Y077PXwXI8iw1WBqhmEsApoV/9GNQl+77U6rm2AoHcZajt
tSiK0Gak+Bx1i5V61zcFDK0Oko/zbKFYDDcROTn5SLNi3/ygexnHAbAT8dbi6xfc7iE+h3bUs3Bd
g+zJwLRzjg+CIxsu2SIIWDIs/0NsU9p0Q8sCUHsKdyHBfZGsCEl3tZjMo+ZFudPTkYIePS9AF2A5
nl0ar1r0QDDYqTNIpe6U1H+jbwgMSjZpdOPLnWQhYbTNxP6L45FmmvjcKGWpqyivN7W/Aw8XM43K
uiJOGyeNebMqmaWgQd7iDAal7P9wD7shggzc+aoGBL13PSHu1gxXe2H/cKX8sgR+6AqoCfHcRNl1
AjNQVp+tHpicUDUubJUk2a/rJNWINeOyBpgmiCbCtI3WXZLlcQZutAgCbERFDS/VekPQkzBkcPdR
Ujyh3+PwrqcH0G3R7TYQfylVig6GkWu7JtUtR9cd5kEhbLN5TPVSvGMv3W60SwGGh2XL2U2+f0ja
31K3gtJ0k6FfxjlD/rFPcOSxEnC8VHgd8kkafxMCg61cdB6w3QTr4bQLctK9tgZJa1k7isYmLke1
13yV012/LBYkMOcFEv9uQWE6umD/JrDIGxo+j7r2VDw9jD0SiwGElTkS9w/1bd63tVdtiHZTywT6
OCykjpikO9jPnrX+n+GF5XAeAvqXz/ytmv6nXatB6jW12NqkKF0Ew1p5oxVfxsGxR8dILNmfFDEj
0i1ZvdjBQ5B8CRAeqqHx1aH8BXNsaIvbuXO+ijG5/NpJHwWtRSw+BEfMqKIl/cuSDdURbsjXbSp/
zcLtjQU+Rk4bdfl+Qfh3ZBXk30frLuNaKFJKaI+pTJ7Xieq0pmhFTBz/mQJrk8OTZyghMGoDG23L
EUqCqQQ+j4pqdkqlHN3gNQz4hy2Vc3yNk8QtJ0RdeeB9/FfvwumoV0KIfIjSc2UZobfPYoFnTQCz
ns2yO53lPkUsZDH1pSw0WXb8DpwsPNzQUKuMwk2xPSPKcGKkUmeGBTpOVMuC+hWY1DRxyAjVGNWV
8Nx9DBGoDyWJ5eMqPV6uWxBPory7jdbf9TKx0fWsaHbz9AzYORzFqoiCP36kBbU1g2uSbfwA4Lpc
O8RM4plp3a/5V/cjXOZxFhFQgu0R66J88/ZFxFrh1vVy31Gz+k1X8d0uCaWopvIeJ0JRyZFIuPtO
2cLDTgQYFDzhtQeVAuiv8IfQ0mnirKMT9L9C7lsZSumMzg3QviyN0dNvyWmzl0Yhy41REfxpf3eW
F+v7Urf91E0EUaSC72QsOpePX2Nr/IEVLbTbSOxVyvFhuRD+AKNV+DulSV8i6YrQbcho0Goz75PC
M/3+iILGfAliq2p+fbLLCcqX9hSoce18R57AADQZZ4KeaiGrZnyprxeZwWmKMsT8Y1sKpwvrDCFH
V3NlCkkO2qSlfpFN8Qm9fSO7Immg9mHhM4yz5eF6skzWiJVa2Ew68xjatUykGjiVGEGDrbuGHJr4
rUFma7rtYP3qDixdtLAIiI2l5/pbpQmKc/Pw2HhWUU7BWyeuOpYVhKchy+j35A10Cf7bFoL/fcQJ
mA3cEQhPyWU4pjgqFV7onTNyEE1ZBCAcWnlWMpY5BRrwIO6sNWS40KbPgMYxTS811tfB5kEmb4n3
oT5Dcx+ISy136K4EzWXhGIKKOfXt4NVAH5fDtE+smYLpKnWee5Szeb7wgk81htyDcsU8dm2jLSPl
wfUBvuiBf3jE1HRJcJRgRRExdUorTft9O375YjBIYAZB2gCfqt4RekUAzNXtfhj2PATUSYLbp2fS
VyPVli6TGeF4kr/MiTL8clbNthem65y7DbJwWiLVwiyzRjxW4wUug9i94fFwzQLHpqw/V0egd5Fe
CIxOBNXRWnzNbVLBk9E04BH7V8F4o0+ThnQbxRAkeBlelTasYXEb7pGIlx57AGGbIDVNxYj+/4Xe
1E27WutWwNlXKzZiKb7USrwAM86FVcVFyAHZk6NeOwxKntLniMwKTF0YMC1ypmbSZfMBRdHKBmIY
Ax+9glduj6fXm9gcPSRR4oZua4tpyli8Y20kzTcYPpI9GZIPfI28nVjmh+yrtqDWOATBXzrwArFS
s8WtFbtN6lfNTkb6E44qxTZyyPSBr8TskhxETh6suQcixO+X1q5vcmg8wQnZMeMjKHzOMk5LYioH
yYAtM48QXi18ZyupajBTCWNdx0dxM8GNvr45EhYKmK59FwZE3pN52M+3MSc4rTDrOJunF1GEXxar
zH8qP+Tuv3E/eWUyVdmrivPY6itWrebu2prgMVQe+pnXqSwAXF2Z2lDlmzTxnTCvpeRqGSYjUNEU
T0YkDTeQlhMDqaqM6tTAArOeVJZWVXpsgLxljOGjvBu/oN5DSLZvBlJtNcd9LEj3vxjudz7oV2qS
9LIOfHDrYvLC+XA+Sg9W6nIQrte4t0K4GCO8RS3vZMYYuYWYbUk5MpLqcEYWnOFIEbsByFgtKLiZ
ojwE/YknSMMknoWytdqSozpPdytacq1fxYhLODEDHXu58NVNd6kILQWQYAbiFmblunuFXXQ/YYuk
tqHX9EK8RzyV/0gsEvpeR6z4/i5BOTJLVYMcyLY6bs6Tgc0ADpKRV+8B7dw3rvqrkHnwQROtZfDq
XmB/MGmkq3AshAko8rYoBRH7eyW38ial5MVP745IzwOlSsTkiBslJV81rEU5myALPuibmxGCypcQ
Aw4/MyPOVedfntD2wa3KoeqGBt3wxn80o5FoImTB7OE3JkiMwxYAtZf8GVD+4mX0dfWPQljsDSVl
GM7IVfYfUqjkM/MeYazUsS5qROaIDS63KASDja8BEsuX+jAP0HxcFxaciZJ8UkvDR0+wIzhuovId
2996FZUFq6/U4sCkeKuU/uPliF9srGIG54t7AKTDuAOVcSESTO2Equqi5DIVhQ7eWL2quf7rJ7+S
IpeCTWiNhUknoF7FSdx8LlXuehrhG0wbAeTf1Q/WP/wJJ8HktZO+1lHJRVoh+7vYC+UdW6O9r5JT
fYw3zjRDJLb19QBq326EgnJWgYlVCwI1Ts3hFwSvlUl5p/5LXZ4VJTTQ3rPkQaP1YfQ36lNasCKY
V1pY+SwfR2IIyDf0coSLM/sexpiNKnNb1X5aXKHQK4P8sDY0383lio79L2AyUnCjQ7WgTQ7uJA0u
xPe2njXZIiuj27w3hVXjwdnSCtWvYihD+1WicBbXd9ejKbTvoszgiygzwijMJ4LefCBDcKSOCG1s
zKH3ueg2Q91QbL1HZgdLbBqs8vcTmx31hiw9ZlEu8Bc9hoz0MqSKyvuIu/Q0PEl/Gwwojwm+vzA+
dmhgrF+Bpby6bNTYSj0CME1/RHChhOs3ZGCvsBmV1LQ+FK4VCv9cYiEFjk0CtaB8G5NhgDHYoCNm
1l3nff6PEhZ7PMD4SXmi1i7sQQkfE+tLBMVXUe/OXMQ0APcvhdUgxI9NMP1uhJoj+4jIKbcDY4yc
2B7R2Yev9PoUQSN3Ow3CFiBJ+acp7PHflBOQQIf7PfW312qjwS/rA0pogCh813fXh/vBSH1W83dP
r9gOfaEQbTNpTYDwMGETHsohz1+G/b4NqbBY9uKZl+q7S9Rj1f1/5czsmKdyRImpvGCkIL4NTNs/
DIWLYAbSh0lcUMwNVxHheaQC/V8tZcUiuJB3qmtDZlOmB4xgMCWUDdg5xXqAM2PhH/ccLwtBZ0N3
NPGcAEF7nChjeQenOdhRzroLpIgwwgGHOUjRbFQs0FgO7N7fd6iD+gvu9A6i7O0VABMUHaqQmrzg
zP55xJ82LX+Sbg6kU99kRCGfpxImMIKUxxp6o8Tiwrc19eDFJiK/gnNFToYpX6KqJ6JeIfRlojG8
HF43JyHOet8cFrF74bmOohB6+kG6L/IHTNqYZY4RuHSkTb2RH7tTIPSe+OcWsUVTnRnpZIjNGZ7K
+hEBOxzXB4KxuZt3SG0bu+XLV2fzA7QSjPUk+jY0Yv9OS3dSvgfoeTwX5Z/Vhg8p6SJwuodYY/E1
haI1T1kTFgL0wvefCG40jMybtiu89kmXW0STua5Y2+fX5RbdMM+xz4ccgI/slV97YDME5ynxgBw0
v/QBX2qusbNg1J98xG7WkKe303Hso2u6fUluOzHJM3Wdvhz3xUAzi9U8Y+1W/WAFdodizjVXs4lo
lBROKmOurRqOcq4ZCnYZLWRgJF6z+uMONWWjIvRs98aYktkb6xmPusX/OwZSzb0PNrrd68jUZB70
VR/An8a3fukxS7SYn4Vo2ejrG1bYeR1YCKoqTkr3d2Z/QULRnqM5Hy1qL1zYVwP9FFloyfK5E2Lf
+Nyqk0lNxWia2yrxzvk1cbRfq0Dtp9tJkShwhfr7IMhDGd1+B79R1lBZKuQKAdg4j6am2cF7j17w
mb5/kATd7gKwxaWfp6oL8qlXbI6VwD2KCZRw/t1g3K61piWt92akA/0w9hS6FlehT7vfEWE0lQgm
S0dNSGPa1+K6OVPIVX/T6NhM8eZHJDqXvz2Xh5O/YTqx266mTxT4eoQ/e1ZzkYRmd43yM0ty3aMN
xo9N+PzwJg7y+WfJ9PThD+AOki2WhALsx/cVvy4D5OSeEHsH4p/aJohwESfKHnhEB/OPmtKpeUM0
agizy+Etx22HQ4VnjUsn+/jIwSqAgWjqSq7Fd1pUVxxfKpuwJ66WUlHtSaoYweWwFPKAO+wKkJN2
a8k1PmlK/y3N5OECggPjQGAdQN3IvCggp8t3eFRyn4mzPHGZ55sUcDlJAJ1Q/R7lZgTZkyXSGODJ
F3u5tPJa3SEOMvhkI7mLIpw1j2GhN/dnncbzzt1a4zy8Ri8FkuXNzvrxoJuO9UFnEPUlO2FPKbUk
nA==
`protect end_protected
