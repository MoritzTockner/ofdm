-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pdPW5xJORtVyuQfYDVeF9DXBn4Qc1s9y9jp0QgXo0NEH4QnHZMqzb18VRg5AgOXeLgXsvdtG/F4p
nO9jNrTWbbaUsoPG38NARQfYqdomxYl112I3w9dUnA3mE7idivPwzFRRATp0k+pkT9ygrBHBiBOd
zvcdt4t82V3CyPwOtha4p1KEFYeVac6SuMU/i+LtEYU0MUSZ0LsCr3e696/zRX7lJCqiIxAZC3Rn
i7gii4TlA7QQ3ies29nOmEnihbw//3jA6EQ4Fsugbzq8O9tvOBwz6R3h49sGJ8pxNWl/WnipsQ9x
q0I2foCe6KmYKHi5RgKw7V7x13zNHLo934eUZg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
H3DIiuP5Hk3IUz4/SehSYX2l0Qjc502a9oPcF2iJtwvd/zSpjGA+P7gfRrNKFbj6Y1NfkxFBAYw8
3nfDqyIqOQ8jZ2d5V53CPu0Nto77faQWcRJlErYoZW3vcqQ4O8Ra3ZHVUeAEMQ7EuZIvW2gZk3dk
xlMyrMdxcXHQ1pfVZFLPLGJ22vm9k6WC5Id5KQutNTvPzF6SeSZug03io06RcRJrj+Yn7X0CcUoC
6Zi9lUdCTx+V9a4CqDWOoRPZtc0B4EPfiNzQAK0L3sHRSLEmGy6nbZyz+O23ONre46GNUO9pVZgU
bJ93BdKSmZ6q7+Zd4Ucc7QgqBJFrZ8YOwZHDGrUT0+gOlduQLwT99E9w1PNr9IQAxtRshU2kI1iT
meLXvRl8Fo0jOo+JJRQpiCT6tjIeb8HoGUCDjTazGUgaGmCtp2nS6FM1pbKXsR9dsxZb5VlNtEmk
7wHfUTmQstjH5N0Vfl4N3f8+oLbmjnFA1sIjZZXOLMlN+8KlAZhf0Fv/+g7FQYX++jY0xRZsCpUJ
Q1i2UHV+Wo1SNOJGLuHXAH8nsMJRGrFWTd7fllgpQL4bH0cjAU+D/UhgH8tMiHIpIn+YwlMQqczm
P8hufwp76Sz4mkCru/HYRgTQ7XAkuNt0jj76LD1SmJvQirBTj8yFEyreIvLWRIGStLVuxFCS7m2I
YIiFVD//e8KD66L++owSmcJxGnDHuBWXoqrkmyFaVdndYS6c00/z2s0dbkNXoJTA6yxF1WmvhnaI
BnOrTJolZUGHDKNtR1BvGp8q7JQ+g159snQZmN/VvRY62GzS9/3GpwmY4wV/6Pm/vLSeeVzITBWY
e66okpU3AB4orTBLxsyz1vI46/mxMJV5XlUVjwWqdEoHVUUbxMs6PNnz3LcHz7pY71dKV/U/b9pn
zT1WhPv7bVspYWRnyDNFbEqjK7m0g0po13gRj3m6Xs6mBSdo9y6YiHvuP9ex97j3mFJIjbC8D8JM
QCr1JM8JOwfu8AWJDmqoGzTmv1chWW0a3zeFxg/Ys3TvQHGWYQjSR6P/1CjvPOgfIWfbXgPjixmT
80+zFhgjNzADpll+FBx/zdn/lb5NoZjWHj0bMM/X+p6vvig5vya8qR0jlpr9Ia/HSHcGtSp/bN4L
7rfsBcbxLP8hP/9+77OnzPhZ/dU7MjE4VcHZE+ZxvIj0RpV49BGVmyVdH0plYO+hnh6eNfQBW1s2
SO4wmVNalI/fgLBcKcw9tVvclC+R0HIuqUBCMt43Z2hxkcoy0RQ9uxuP6sNJ05w5z0XLUrQV/hNx
ycxr/iyPsIbnsAQaoYoyLtA4Ji0g0sm4DhrXN6Yyuiy3zB+3pw2KGJjGj5LTJ1bP50SCdtNkQc0z
VMVqzBxgVLAOOPGe84gj29reurPtAm9lCr064kNFwDoksTIcwf6vEbjI6j0ow84yX7foZoaj8BbV
p1zzo44OV7+jhptLhTK1dFJYKwgcpIcC1IbMMmbsbCXWZVQW8rxebXDsmheoJZaQWxv4tq9uckbC
0YYOdDPXoonsVfEUxQgQaIZaeIEuLqbUbxGN9WzlKLURTiN09M+jAgzboJPsKX4Ug3ohHCCFFexS
TE36p4n4J3T7Ubgk2S9FFHIfcz2OXJB7gHjsi1s//9SOPpOmHXvlzFPDa5LaGK8DJanxKTja4CVK
Xyu8yX79DXmaObLM+16+jD8vkjOqDUM5bBR21L46MatWYQXdF23qTDGKZaRTjXPqBE31rjmau+Lv
ayWwxvoWGB887qgq1oPrK2I2sZldizwdb0ej54aw2Nk02CbTGKzLX0AiWnGthJtnES/ICsuUXdDW
Z982Fwx5fdmKoqWELtzRavEyejZIEyMXA3jpImpBkNC45wc6U2rakT49u/m5cMbhg2wQZFGuiAxf
jHhhZ0KKC0mHwy3q18PgUWIGS9+2z3IYTkOGa+w7fUdTfmg8efOHZdOwaym/ge7FALdyfP6Xb9pG
KV9TVQt/M0HeL5MgajFf9OaK+H+KOQtlfFB8cd1JmaUY8nTWUrBajwYEn41ww5QfvHrsVvtxaIX6
CZXdWbcgIApt6GiVBZgWZBtRwxakgFaj9C23LYdr+fnjRrHn6esqNEFMq3jfw/TzLmvuAvZlxh7A
T6uaoeM7wgd1Yo5zhVqSciEeOu9DrGlkTxIj1lJN+eIeKjSC93z5gnrSnBFg94VUmYmEF8CRrSVv
LcHAnajsavXtnaHo8xj0AFd+v4+FdZOFIq3zeWPTaOIKxcWPwehLASzlqdAAvM2PuiTowsujAOf0
Pny2RUOVR00rrrPLdWNGmglHxK9BRwTVz1ygErrWdq+zYy9A/yKnnF+EuE7oxtr1dss4qsYOUBzV
+vz603qu7R4myRpppGtcO3rUwVA6nJzQs+VOyUf0R9TC+tkKNG8Daf1JoRQZc3Fsku5TEYzlc1h9
4GHwo5CDJ8Po1JqKf9kVfYLDzEwv4u8Xbpe42SJl9f+H1vFLchfUABsfaVVUIEWFb3vj+csL2kGk
1aOiqAhMn3vZZSGKQ8b6QlfV/4PWKDajK1HXYGosvru2YKo3URtQLayJqYTdDSQxYlZ0o0/Bg5H0
YNMMyrdNlSidY3PuCLamLeTzHkudEdSDP9mry5N82B0J9hhs4FIGqBq1phs4PHhvFD92gfnSHGgZ
IzT3VeC2CaAytUjtQF6zEQF7LMkKsBzwThLiGPJbkf2ECLBj8ctBJaY09//YYfGYCZ2rv8kpqufG
Q+ULXzubyapYhtZJcxv9ICslYqYYu4MzM72XQZ5xssekR8kQmC+wwCyXyp9aRpWuL88X4jkOtbjf
9ZRZN8P+h5mXVmssOV7lir1JGBzrU3UJJiylmZh0Rmdv2VV5THQo00X5E9rWYYbo6Dny3mh5m3qK
78HTMwjwj3TdRb2DyCiTvoIukss0mfdUqwDTbnXSNtvOg7lTp6fpzPPaPbf1qDXi37Zs8sOhZ4aL
f3wKy1lT5Ek03eSH3/hpVFdXq7VQXIxfCU8OkRrZOu8O/k0rOL72CRlmFcfd5iN/j15ju8zb6doJ
xf+73JTeL3nYEb4fPA+YQPvRx00rmTK7v16ZOLBWYNgUHSdUYuuMLZxwLnGynYQGyH1qQEsCBP3W
UmULelKPz5rxprxkxvylFwCk5KbNdDc98NYA5UJK4Eqh9yHAQIg5fXl0LbU5+944Z25cW06STJXF
ihAhrs2oO3S4kQCBgHeOJjS5pPR/+hC5uUXAUAGGIeaJbtzVYpae4Q7pDVWcO6HY/jdYbz43Hxzy
vIDLkVpbkP+NNOkTrtnuO4jjD1i5qjVRf4YhfXz+G9EDEBTBdHphrdaNzeHzLfvXFdUscXa+z6lY
3LKADypN4Ria7G4hRByW1/Ogsrqbitd77Ha7azuW4W1arRPNJ2qbF/YtRywmI8gT0gO3bDEqYvNP
h6PtcgR83AB4qVFG9HnqD5Ea++uNZxwHYlfAd2w2ejprbMpNYOPZp4tkCGMTALD9RoMOKKTOPtu3
ND/Hcu1FPqWW2oHLs9VJXpMyifYNU0pes56l5vgSqrBFUwvPI6ubK0Xpmzc8uRBUu9uu95zTaTfE
V5Y68MCGjXNeDHac9JNwKmtuiJ5zDirFNIBv+mJ0KW5jafZFHDaHDQDQoaLHvLCmcOdn2iaR1Nn8
1pvCl99diY6FRHBXyW+A50N2mAT2xx3GA24wAkWjl/rwJOV7g+78+kRidxKMVU8spseUEHNnQusg
A7Y54DQII6M0CjeKVH/Pwo401xq8vvsJQqR8ShdC3AfxZLAZTD21BmR6f5Z+Xl+fpfRHyuy23p1k
O93bkciZlvkN1J+CXh8YLYbvNHQUsfvH28kpuQq3VoRXjlJHu0KsSAvQA0g/JAgz1oqPHn1NTq97
5RY2e7c22FLNNe6qeoMoLSy6Pz+545ToTr93c6nSw+eyEI6K8r9aeBDnPn2j7cpOK3W7wyZN6MdP
8661hCd4tdxKFfHtP58Dl66w3niNIs0ZsW6XesyYDzMvmgsio1L2bSSD8w0RF/VDVwpAdc1RcEkb
e0S7op00wvyXRZ8ud9SNWamwnJ3iSMcLPy8hxX4+GRu3AK5XK8/IxVaDHK5GtNkfnVt5alTKoUKp
RmcfEyKxY64Gxn4sQYfNv/EEmfb+F/n8gAL9qm8UFy8RWnOacfmwls+HQk6lQYK3Mn6gu1Zjdzlj
1+mHODWzR+L3nnUo4E/QhYZIvjsWvsluXZZGvXeNFGI6wJmUCOROEklf5vMTf1At1JtxwOq73pLE
1lLc7w6n7CsdZ1JG/rBfQSVXsD/uEBqWFUD1rfmkEP9Zi1997tOZL59Nut3/AnFi0ZrPy/cTLUCg
CNhrmrxFg7ca2addOXSBBc75FF22lyT0nRgBQh9LFHUfSkqKF1omS5Y9lnv+TbxnKTyYL72enMwX
+jSsP4/KW7eVXmCEFjRcdPcED1bacax1wOBYNdeVb+6cEVLA6ZmtgDM+cdvBdaN6FwqcuVJqHMAj
6fKtwrZxsDWlrQ+j8OeMkNlqjvd0p7S/LULB51kX3mZX3/BZS/0mu2v0BYZmtEqmF+c+Ww4Vj6M0
795wtDOF7gXZCb7TDhIpw7LuueD96Sw2aq4OfV84i2zFP2cHNixaeNkn7Q8Jeao0vuSIH7kBC6N2
iAMnQJ5AbrG/ugETPdWB0TiLAFUM89ORTKeAqAbeNarom1THhvjz/QaQCcl4D+8jy5eCd4j5hQGv
/pYgjqieqtGzzkZVfiPd6uvNlYoi/2W3H5ryvUJW4fZz426rY0ZSxC9m4M4vjjQbG183Y6uyUIj5
wvbn+ckPY45E+kYfrUYnilnhvNKo0W0eaAkKiOQOwJXjS8wUq0HOHbTtgyjAmvf4WceM+mm0U2ej
Bvy5xyAdt/6AesFnKpzzJ47f7G2WEWtobxoreBITQjPU8eoc+ralKN7O26mbIM4elwkg9Em2iqQS
vmrRMeuUKTsOHy5A91ZBKpPGfJIik2plYF7bQTN3ENvBRySQfWoNcXK1eC1epKj53K5X1SCfcDH+
HixR9on4h3/SOGtIz0p4GzB9lXdszb8yLB9YoMKd7TVp5Keuddf9syJDsUPwViwpHhuwhQWhZb9M
yf1EcrB+uXZOaDc2tCxhjodLwlAeNEP8bdlPaOTXf+f6eGNyvezXgEnlodSo8AdGtATaFf3W95Yy
2Sd+/TZYug2w6JcANiIh+q/CHyRb8QBX3MDJFer7yoMAsD3ArKWfdDHJ1o1/FvcgamPyO26nmGeq
oQILpfO3J3Rep9SvVT1A04h/eCPYGq32+XtEsEcN82B/q2jaGZH+jjhc5KC1he52ebu4Kzaf/MG6
fGez6QLwUHgztgwjAr4CSKd7UgRiiwdo1ZIXpP7XwQQzWdLkeYMMIciBfuDBG200aTibk+K850aN
SEVzIucfuvZJOdI/8qTFOjti/BRlbJ2PrCCFdLkkHehjmYOJP9s3BhNZfsDZAZFHoClX3uMFLtKQ
aCCpIlvF4rNlk8kJYGZ5WrtyDShK54GieUiaGO6X1xovT1IHiz/rfEWt8XHYuoZ8oFwNpdvlMFJ2
xLKkODKMXV0S9+pr6vSqTsEIjoo3BkiK/7A5/RglP9+8LHPUnSy6sSciLkx6hX26R6e0w24NbPum
PC9/Qm2/wmka33Yk7e14a7Anw2GSwsM/SiZLDJtwVmka0tnqaUZFzLekCx2HN3HQsfo+1VWvMsjf
K4kgQybj9RXZFbp/W3JGlz58EZ2iPVv8nwOKOuq3rmP8QRxO7hMOVuIJCObEFJvWKPLkkcxgeTyV
UH+ZpUdwpbxDXeSKozPgKcZb27XRUgIZgL5oBhmn/+4xoMw+LVfKNJjgNr6QN1A+OWmLtFrrJl1O
2oB6Z9xpk7iYLB25Zzwk+50dvrKbr5Vhnbdyf8IrsuEqTrCNHt/L6zkw7rUgl0SOgvY8MzL9tHn5
OrCla0vyvFlrz2/KPJF4evVYLgkNJ6b5lp/HmCpOCqzMbMh32+4d4uZ0Hz294uHS8C7FnTX9OFjN
ZwAfBwt5IWQ6AlxgXxV3mIuVE15UBvmJdsekjvFBFeKdRrzBVUbdNfAOTlrVSBAl2hZp56ZbcTTR
vsiNfXMRo8CwrRW0M/5dNkPZBJ0erUJkC9CzMaxc6qqf8EQdfBvYvXBX9vzz2iLCZX7KweXmMFQG
Luuh1Fma/7TxNaL1YppEEJZTIg54DMh8ul4oknCtxLio2RIpzcxgMKL3hX4WsiWHEnoZWV+lM2A/
38ur0zc8/nqz7RoF7Hdx/a3ViT11QlKfGtz1e85RaZ9voQfSVk4YZdfeTz9//PQdRHsSH5D/sJOd
PvbKUuqZWpJKYPwxruHd0b4KkBonDrp+WlqMp9Y5Vc8WanbPN+VVQy57m1qDP2pK+bhFRbHccTvH
aYyk/72X5SjWWb0qfmVL4lYw24MxvhJ2Bw+meRRfPKKOitip0MwmuQZ+8AhsgKTuE5xOYWsHu09E
7ZWZ65GMmpMaLeYkxSZxug3m9yvp/toe/J8F2zeyfdxLb69R/WaZo+VFyCG9/g6YJkLn8GR0vRRw
6bmIu+LFrsHWZC/CFomHyMG8WLRQ+oFnX8kPaL8XbbVEuPA86AlHNgD6nwfEAl0zBjUvZogirQuF
2Fi1HXDLI376ZzhKtFFxZAm4xpims2bsKyZItQ4n5BYuNt1D+l4EH95T6P3NwHJI7mRX+UQOwR22
sRT3TyZamYrGzqZ/04ThQ+l7P4Mi0L32t8ysfLsB0+Bp9wMHZxJY5YQFZLj2iBX3PTbOWGXZxMhq
7PpWRymFM3agPmavI6Qa4vn+pZgWv/zKVLzMDUcjIS8he+8MY+W8FBaQhxWABA57h/Ca0s7Rracs
c3IZRFRPCt4wq/FsvJoNnfqneTZjSQP1rUTTqnR6cZ9PQyBIN7qm2T/qDpTeIjqkAHew4DwLj2af
nao+npjA0Xu+l53d/RGVG1LKa0beU+ZxYYWaNgyhuWHIbvxLpp/IAAL+s8rL0yHhdxkmlJJ0latQ
lHxaeAimBoJbBcMd3HlxepVLX9JA0XuuUaXpRAr9lkSZ1+PFTKZZk1sMIW3mPJJYU2MqQwxO7Ge5
4fRTX7LCnK0vovPddAmkFf0oTXNzj2rlzcIgmtTOnAZ3Fe2L04SQw1q2QEbEBPvhVGSzBT+YOEmt
6vsJ69BWR3msu23v4zsmKczO7eUWX7zaCCPSPMvjXplMMqaLyc+BA152VnN0+FDI7Hun4UZrcUr8
llV/nt1WCpCo/QWKSMAwbpw+eqdmJxxIqZOBVrqktCdr3jCC2GLIbRfS4OBIhw7ZtbbZkaXVPUm3
vk+AEDIGy6D/k3JkRxr14h2j5rHB1I/6fMooXemrvhB5IpS53UnJjkHD/j6yEJ5K8eUXAehASd6R
5hDV4URt0FANAH/MKR9ijIZsut++PH5vJAx3lkCO8XfwtwS2pkqTn0y5YtyTF8xR3CXDi5Ba5iCu
SpJc5kNiYIWUGTdVcAG/ntKHL8ElmNRDAwpyvHMqRLAMzIx6H6/GgXICO0Kzw5QJnxjoRpTLYhVC
UDQVoV7JkFUi+jVR66aK9N3YyHIccZSnp5eArNDp+KwuEBkZXs95n+BcxjLPGHSBKj4cA35Rlho0
EYeEIwVFt4UZOAmFZoSmJ3aP6tfjGTCRiTwux9SMahZY9WYJrjDsN10mjA6a/WfnM0lBCL59Efgm
V4xWsl1M/APB0CRbJ2/vA1ouCJngocr7t8NMPmfzqzozkDjFt7GKTR76Egh4bQIvmrcdFV6zqzHX
qvhSRVcqtCiVWX/y9MK4AkWWC1nOFJZL0dH0iUyxBIEpg+xMmFVKGlvlmUCoKFUx5mOGLa07yRbs
sBXPh5qhxzX24R8hzbPE30rS5kRihR1Z2MkaWn5HCUflnnXYYAblvLxgrjIeh7kHUZPeROChba91
XIXvFEQJw7m/YYVjJ++rTKShM5bL5qqEs5SmH3FGdYSc5vn0im406655SMY7rUYUHdSdwV8lTwLN
YEJALGm/8fQArKvvypLSu21kcK7Yb2rL7Zfc8l/VhNr9ekNfvPcIokAO0+ry0Ic3FNY5QFwiGDux
HOTrKXjb5jz2z4C+prAS9gynEWhLCdnsA06WOp+CQQx+APZUCtBXv/qFBgFtwaNSuS97AzL0Gw4J
RpyDnmyw3VlL+q0CL0PvnfpQphuAVrgsuEmY3Jd/4CTv3rNE4LIX0lM1HtRv+ONbFXvZbZ5zV70Y
tJ5fXjVQfTcbW9YC94f0+LDaOoOynEU0SVbtj5L2B1eQ4G4Jxf1eVkLO+2BYND1ASR6htlmBpoRo
+4ri/Zz/qCT91HK+RU8/d2wOKiF1z/glv7vDTzqQCgvjg51d3GtrXSApIE9GeDOPjfzcWXJqR+bg
SyUTdZlPCopTaCTdzK/D2B9lV9Ct535zGd9Nflhg8qvs5CV/IhsXmviATufQDIE9u2MjtcjDHkcb
BkAG+meEq+BuoLipRthq/x66ByasSKtRDG9Yxe6ZbB4ik7AgSCuYCycVN77TCFelHi8fhRAnp6TO
P1AMo1F78hSjZ4/vR5PRUok/MGIjlNuEo+zrSmc2lUJolAQW9xL+xZAcn3dGVFfZaq3l6JTjoWCI
gWiac9dRVBD6qWzpx+nK6tkPGJ6oD3V4qI0xeFW8zOGr5SuM0rQst8BSjd9oeuVuECPUEncmnEv/
CbMfpv84gj9zKMIQ5+VwEVxy6pZ3CDOJ8/lkHG1qyBAZ2CvH0lm1Nr+nYLn1Iaq23OkmeEWDnbu3
0fdd/cYilBRnNc/+pFuBje6IcK/RS36Q9UoSfV9qH3K4uQ6i5WRZS0vFnHszPE7kfMWn8xOenuhr
GLMzptf/mDJRYphsjAq2LJ8uM5t6Js5u2BaerrtaHh0Z7mWd3r0Pt2tNHWs=
`protect end_protected
