-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x0x6DYGWkhiNJ/x7ZMAbWH9L/NropElxVCxA1NypFTiClmXOHNrofGR6nd4VCBupLbZfEBhuJerj
VJ4V5PhBusnX728829OEYyqXrsISTVXerOpNB1yUuYEARKgkZtOfGiAF5d4JEI2b7HhTBQ1DhKTa
nylwPA4bcTajWqjwqpIgIAYwuY8c8g8xY7dw67YnBLPdrXSCaII5U8cy48TTqx0bxwQFOBuhnOKU
ckEFcd+suhLcDdHQ8FQZbvRQsahGlqGWh3seULpSjw9qfvYLGWDZgrFNzeWU0wxScbrBP/INe2/P
DETSjDlUhdo0RMocK1v0pnqhnJGdrUmdKGD4Eg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
mVsSB2/YrrKXfHjUjViArJv5WczpDbc+zNs4NluZZkSQkmKM+8lKmRUUhVERwme28IW9ud14XG6g
DQcuOF1MfFWAU0lMjOfJ4F+FTW3JXsLRvTHhV2+Eic3k+KGvwWDGveTW8R54MZ9pd1qRKNT+UgO5
UUTd/LolKfrLFKDdp1vDCKWW+dGw/Ic3ugz7CXgfe9MC3mwk5EP6zqv3dluQydNWWOWk3TNuvPcp
flxvAtbssxLVaQuK1RLB1yJy90G1l6ZzvF9RyEmK9rvYX9ZVmDuNSkoq+4D4+hDC4DllBB4RhkKt
aiXk5lDbILmslKxiluQf96Hqo2NWP7yN9er7Y/DEg3SAEMA+vhS/N2P4as7EXUv0aludpBHIBo9t
ruQpE7d+FWJaljm5EyOP1Ij32sysRU/88+G78u4RGLFbhlgKceOWoaQlAi0quxy3mD9dEOLZj16Y
t6tqvqOBUbXMIvQ5RQW9VunsGbvPLcQUkP7k8Hg7tq9BQnyYt+pSbZ7RCkLXoOao0rCRY12JCpLH
QtgJ+VxGBGE/Gb4HF7t+DSOcBdMYb04HuNwuObgBVwGX9Vzl5bZ3LZPsAW5RjmnOgPIrTmgZmHNP
RrLWKQBW4/KO+SVehsDTpDMBUDkkn8PHtTPpS0gkFRekt56CahRPYbcWU2a+ZAl3mKBLXjxWRJnj
IEq54P7ri8IgLVdbzIYXE5f+RVvAV259PXup2mZ0LdhiW1Gem9QrkukaG97UcXq6OP5mxw8PMi4C
KVQ8POpLjS5EziTkqJpZ3cuHbgapMGxSINsQlDhKL/U0awZbF9diTqANKdRg/hVxzrUJId5KWFZC
ZCH6cAWuPyHjpqmv/EhRzkMAQY5l38hWSx/JgEhb53JrqB2tvhLyHPurUSMRuAP0leDglecjw3u9
dIFDiuuWfL7CYkB5c/c2hlmcFd5RmWNqWDmuFbvHRaCjdaV+U3Ck5DONg3g62bZhIY+geRK2T/FQ
2xtc9uegaoJbOUYz+Wn2XVCr0gKF/q2gkZ0tCRe6DCXWBdchv8DNvxztQfMs4PAAoa4gIPxPi8lE
tCrlGgqwJ5Er7D/4W1VHQ3xSRUn3N67cXR8og8vJJwgAWuSxst13+eshMUaWu8zxsd0Ipiq5DpyD
7UpsbgUCMrPYLAQ1P1yB29OhQFA5dtX9ZOpC+UgQlQMuggwIVMYpEw7mqLbxO6S91UFkZ6uQNlTn
ZTPzkRVahcLz/9TgVPWs4vPzs5kGh49H6Zv2pVA8SouvX4DEC6hNswRaxoM7QjrFtLtF0LeUwE/0
UfBuCfEDXyHaOrUodpjtfWgrBFGQ3LO9NqMJ/8guUjgdZHFLBiL8gWxrtVhJBZdE0kJboc+Ffa63
luG2KcA2Towma7bYhe/I+QPC8IDCzNIrctJKzkqh/PaBjks+Dnh+mDfie6fVHi9mwBL5poIbCq36
mCLClWNVdhuGhdS/N7aX/Kg9a3m9Dr8yYSzckXF6fqj6vgK1rxcx/NlZBG3MROeam9qzUsiCm3tT
XpRGVFmnbXmqbOQlewad+n6UmL6ZTvY9UpyGSiMgq+L10xRqn+khpelZqA2d8Iv4rzxbPQAmJWIx
+RDY75L2cXh8J4i7w8U5216EN7550QUAyDa0qU5a+Nwnv6pfx632rH7XKVH6Id0gFxlX+bVWPmzV
TqDNM2pxVKGxDXQCtJ/C+hbOzOsxSDV1av17/K76zgAP5wAZgqJqEJwDoKQa5VvsfOuRjTguPsW8
mhAdloRFhYt6PXD+UTgPVPqER+A/FZhkNtoqwi0Wn/dhoqLniK45ObjfxqgM0lSfD3PJZJGzOqtn
EbzaJ5L9670kVeBNY9ikLtv1WHic/tpG0L4z1/JEPaZfv09EkBd+6Ssremw8uprKCqATzWI+OhbA
1xtL4Rc7xYIVVKqBw/hyQiYDWZPOEWYez7lCDbY+gub2x1U9Wp6lijVk51ujvNreg3nAABX8GlbX
nI8+JzfixzBcw2l3+B5cGzLmBX/FMxbjY43yxLtnv014chvBhrHPgsboRzhHSO4IKBb+WM3g51j5
MzcskmvW2WqOF2CyT7JSDHlWSPz8cwVxLPp74ziC6sTef/0cxX58IAURJncIGMVuWAxHDuo/iCoZ
vrsxCQQhgCsKqtB6m9b/UYLCRRCKPPtJzomwLut6zG1/L5+10s4hE3RFG4emlR8dKmWbEYxBP/b7
9mQ58CCBJ24ANBncfJl+T511UmTv+GTv9G7zXJrSS59nrATHT8OmWVQtXfm1rSEqNhp2VdufUap8
83KjhNK2xxXXFUubeAtJCGZMfEGjCalIVNIBVyGlT2TmlwAN7Oib6lPX4DBsZCVjAd5bRe3TOLe7
6TdrrlcJDg76elj7qNnGy8R4EoevuTWGYDAEdeI0eb/ShPW898IU5cpNHt504MqZ3+dB0Kip+hOU
YbTkbPXl0afrF/wvouIWyRCfhW7vizDgug5VogEktD0MYJA3eLKP/DUt1rdDyyMmZsE3YmgmL8mA
VEx+fLS/rEXiJSZxpc7xWELe58hysw+CTDAKt3UF+f6caRIZZfTPOFjnC8Ei3dsYkTeMAsyiZQTh
rY+mvUaEbvYs4wQ42v0XaTIauGSzWda4Wh66A7wtYoMdZNtxnzMVfGXPkctPdCaKx1nT/HUe9lEl
4n8+qNqRCyP1HkQwgj4ip4WCD1tYKDuVdayV0os+CLpbxzp0O3ObqaP0NQ1J7i5JMW1GUTn//UEi
W5fUupjWkozLSvmqRtQ8DnapqPLSFaRnBAW6LjlESgufo5db4oFWPplso1P4C5MqgNEDBWbNuyF9
/YKbhPzs9j+FoZ7Lq5mhgODyIBOllfjbqe3kS4T8RSeqDJj9WU1U3g90kbIV+n0UlPqPdLT5edGF
ZTnhNJp1nuSjgpb4wrejCI6ieINeMPaTu9Q/z1m1HIj7Mp6AFekLPLC+JgKywEGZqbyqueXrCOys
hbJ1X/Ne3Io6SPClyIC5v6pVQfHovn5g9+QBJg0u2SzQR2dViWqWvzOkdGSgw6L+EN/DKSgFoQze
sVTtRCp8QpSNxM1ro4Ux+UmKKpbGBMpO5xEhc3M8hSLoPD00FcqjjxoYX5uR0QsnhPQLsFlqhj16
2yOtScX9881r+d63XBNRVJLhxfzH5QezyGr47KP3RnQGbY3g+OJALmHKlnoKRSDFLIwKHhiPWE6r
vPhRoa5kTrFo2YmRkr4EqYZYvaOK2nl3Zj6t6LID+JlSoQd0w7QC1tNxzZyqSDqMrBHr5B+Q2N6w
WJQQnsMqBUESt+6cNXcmXK6y6gNl88AgF6SQSgCrlieqoBob3/AY0KgezkfNgaZs5ntpZhBnaRLV
GChemmlFqoXdamuXlmSmnErpdarbBpP6216pcKybVOX2sV1VPwO6QalITCu4IKRcqtn48jDHSGSV
TOj5xSkWo/dRzqbaSwObMqvYQZhHo3qulb9vlk2dF6sG+KUZTZwvj685mY/VU53vU6e3WcF+fqCg
RtNUb8x3m2BZLRMOG0WnqT7gxKniRqQE6QWhO9M+e2eF/TIuSFWBlXVzEumJrw9t1Wc2sG815MFh
WgXksOri3GKpZP+8K4vdeGEBjWDXV9srdN9ua8wwcai5l8N8HTIPepZZw6Wt/+YwIHJ2e9zfiMMt
2yI+HSzeEOvMSPNfqZ6u7bUI+6y2WzcxsE8ejPoH83RJTsiCwcVPSd2e+7wQOfMwYZCmqDMY3aHv
Afqk1ZHJg39jABwSv095woK66GN+UtETuF/PDLgcUaaXnf+tE2Az1NDsEfOQKNAH2fqAKrC0nzHI
LSkAqk48ZVIAEqyokUj1dhOPOumXC+FEsbVKKOSHh8aahMLX4lRLiK35n/ptUN0bqDn2uP2BPnfN
AgflUyJ7pnCxf0ECB8xPc7+u9bJeW2N4ktTvMNUIF/eG1hphfGrJXiRG9zO68Qu0HVsB3WDTsTk0
GF4c3vCfGrjemGisL49WMujxco6MUamNGoDZGL6hR+s+Ycj8zSsS09XSggEqDgQcqvzFGkdsm28D
g5XA7hG3S/CGyAbK9MUqt/HOXf6hlkmiDrRucDgXWnpD9u+KwF5xPVbkIkg0fHhVMJq9rHmdtyh5
aWUOHhh/33G/e7ar4FUJz81FMglVlT2uVZmjDHhDpzJpcGjkNKFcoshqJ8w1cKn/2+o+IBZ+csgD
fdGKjIj9gJpYCcpKs3H2wMyScol5/X4hQBp682NWl+FopUyjGISGkCAHCza4/Q13CRixww/PhT2W
2bBs8Y50NFWdupE9ejjQvLnDMCQRck9k4GFzH0eD226fipax9A+xFetGOG/lT9LMDQ8eA5XIesWO
G1uyLCLXDmv+ElcN2+wAeO3PxJ9mzIHbzf5GIhZjdGQ9Xaspd30MPI4XN6eNshIbBwFapaOE1TPP
kWHE3jgScNHFzRn6Kir0uvR5xdvmOL1m2H0gS1OF8XS6d4he7jrbsDZpfggRjo4oWgTDgO8WPAe9
Ck1N+pbKe/dauKxcyBnw0Gz0+taQwOH9eXvCN2lQ6wZWyNZP8fjexxn0dWQ3+KUkY0LQjnOOcn+C
orqA3E5elpf2GXrW7vgUmCS3N5slI0gwg3gVnF2bheAzjCgC368G0FtaHRsYZ34Tmsxyr7g0BOc8
TBi78ZAM7wCtIT0yuOe5h4ihHyoADecrqe4YYzEvbVS9f0d4b9kwk6lZmdVjMVOZBKK7Jh4eIQie
mpu803rHWGXYg51QZK7neoBSCY4fdH+kXN1glO//jCnU9gHLAgdCWOWebUWjAzkqFB7+1609/g1f
A1yOnoNj8K8PPh48bGc9H6ydgoeMksyPlfxbQjss/YnpmTDizzfU0quH2appJrq453N4dWVvY2Go
4kSorya2jUgzVnSyR5RqDUF2GRoYk6ZE/4SvmzzgHWh2eiNq4ANgGWqXdAAEiP3hRAebtN60QXSn
VOEoRbME1LDwQ8P9ii36M9CAwoyf7XRz0ELx8DVUKEAKPzoL1lmylYZ8isaY95GH6SVy/MLB7dkS
EoP29G2cP+Wv4HZY0zBBghyTWq+voONFM75aU2wa855EAQeCdpCgbMKMk5ww6cZXk1PpbeGCzC1N
eJMh66ds4HMuy9Fz3o6IenPGcrpvsRejYwJcquvzwWNPd8YM9z/mNrAAEN+ay2tgsKgcQN2+ci0R
rPwbzMKZ2+iGq2FpsO7/ZOh9qCIwLHqYsIq0q+Yp32v1mGpoH16o7YoRJQFAzQgZMkk6u50F0jUg
ZgXHBuvXyJQWjA67nb7lThWLomKYQlG5pqZPjp/G5nqwoYbeHFAgFSyJbOp5lSQW6CyPogRRgoVX
pcx8lDDO2z6olPhtMTH4aXKEpCPIUty0ZEuewUV82SZczWp1lkazarXoYRE69P693+pQ93DH5NyZ
5OYxvrqGUuTsr4XyRdilIIyK7FFm1+ZrOO7lilFEFu09CMSdSPJ4tcc81p/y8OuVzKNfKSLwwL/M
j5Za63w90P0l8qskuyP0bJg1Ym+aCwWGyo26rDLntrIldXUopjTirJqzhjnBnE56MZpLwxDhOKJ6
h7dsDy4CwcpMTUEPts+BbNWY561DRN9KQgMCx9AKsi3wFMec46u6n2JqJ3YamaaDBaDuoH8hU++V
9KVRu8aDjTrTHEs9CJkXN7g7Gn0LN9XrOS5PQYgD2Kq3XIWa3IB9u1CFZcEPAGGVFtdEAmReLe6g
Sy3Z2AeZhDOD5R6rooKOn/YIh0iYMqrSYB+z39EOdleTZNMrJgn9wavBJ9/FqzbgFLZ7a2A6aBgV
2DpOz3ky3ByZCKSSZTt9K/LVpBY2zlUKV8eCGP2KCqOESFsSZokzvATUiMr8xDTsYH7PXbgf/wXo
mTr1w9she5+TnwQfeyh9n7ntw87efhLbBHvkyz5ZkADN5nXk9sQaFzKBLYNjfLinTYg9uStm2Rpx
IHxrt1NDKMIhvHvPz4cz7nLzqy3R+6z1VFZQ05Ta/Pjgby7AdwaiNKQIqegUn9gJgDEAiEzewv/5
ODAKimoyRWWCuK6BT2fP5KphVu7WDbNd2PwPdxo0FJelndfDJJ1YxkW//h6e0q/aKVNCN+8ItVJD
Fd/OHXPnaqWQ+o/hRJLEFzjB3fkh3vYU6yuvo7yPw+kF07aM4omZLd/7784a/bjRfj0vQ1geRhK8
QIxeQNGAQHff/9JX2hfxgFDvCwKwY9ayuORbtQrt+VUNZ4RS/K6oKxBEA4d98D7lYog3qLlO5BEo
fD4rBYnSj6HHO1gDoxY9WEDnV7Y2cdsWOqSQgvkf9/mQ24tabrJupW4Q62Q/niqHWijsQV1tYQ6L
BOdNbzqR4J9kRbcbV+kBXCHWRwr5gr7vHf6Z5MLA9g0cHxVMDT+uA/MfHFXm6P2EYYrIx3+wmBjw
N0ftvSHaufnEgb/r13Go/NYqlceFfSXp7n7Yvjohl4XQAbGsKJ7wiU7u5EIGu+LyP4QfvaCqbcLF
JOsl5mj5zKusIOG5k67fW2EME6I/RKQv7iNJrSXZGeNIbeuxM0spUCfZfmDRpvXiJcrIwnt6ykpg
dTMRVm0jPYAJgwx2gt/sqFa4KiteaEVpvn4GYo7rSY/LhyqU5DD9vrD0+AaXEjm+peTww09SYR/Q
zRiYNCvazckReLRcnYFEMIuj9V33U9j+qUSOPJGa7ox1Ug2JPrC4NzoIyILpAWXDneA668mRzRz4
YpajFQf3kePUOV9Xr7qMCtg3LVhI4iyFnZJSba55ch8zare8tS9BHVkZodixX/fNCiuNUQ5WZjRt
x+9FY4x8Q+RNA22NwnaX9J8r/L6qYM+G36EjQO0fPK9cGObb0rqHbMyGrOhb5iV9kY6dlFIXr/Tu
h9xd8QUKlfPA5Nxtn/RneNM0ue+QINzGRM+OSCwSHFrsGAjp9TBjar8WAMfr3NZV2lxlcvWrCwPu
aLa//las0cmJJ20XIZJf5Xy5uqK16xzV3JJCVHKCWayJ9RrL+7ICBRg0GVO6yk3HgGLC+KU3oAJv
ReU6COIBgEZBCAfs84lD9ow+ylktI2D/I27mhCuVBwVtHjxp1VNb5rHLG3pk/4/nmOhvl3s6uN4C
jOtQT7cvbmluLNfJl5eC/JM9PuKxOfETdGLNzHHS6s8L4WZ/VIEnFFT6MYw+OlwAnkbRsg/A+36r
w7qQbxZsqaAX5HGfAwkuGbtBLHs2lyz/nSdu11th1a6XLOPBWHigkoLrAeXwgni++oxwJjZe6NJ1
eioe+zkPezhNPIBFmPhe55WeOnMdnsF7N7TjzO2FFFnb6Jo7QH4jIj63aNTlkfUyQxjReY2jqV2F
Vq2LulpbKnpSU3df8BnC5wvBPvAk0QAiCJv5+AlYy1is3Ubkblai/7QytfLf9XSPpShgmuq6sx9j
a7btKWvLwOM34BTvoLmKVwqyVBNH9stw6rSigp1HOWhf+jzFSmKXcR6AL86eHnf2dF1aThiSPQ7C
OUSQIisyFRYK+7FJbfqtXl3h0u4fCknTP9FP01/+0XZDejN5uV+yoFKgg+t8gKpYSz2+oddNr68t
mhMCRb5ti7mn3pAL4vCBCLIGC/G25p+dJ2c255KBjfYGsSt9if72nL5mk2rpzIBqUMjweboIWyd4
PtLKXLCwL4lK235OsLOC0zALovSSKydsjlQ+71TiO0QpyCRByb058b0hvNUwy3kM08FKu3AxCRwV
mZySdF8UQGAqpjESgiuGqekvD/pX38kF5RaUN5gRTvmULSSmyFhuZHjvnHLTTnrBEYzuKNDQvPgY
x9BZVUF8HmuXiUeah0gaj1MSE7Myg/v6UAtrYTx/WsOCBPd0IS+AWyxMiPqqRdt7tv6jLQg/xYEN
H2nnVhF2a5QawwBEDMtbTLcnDzN94/1LgLrY1iMfz9GrIHCZ+r6zk/Oxn13TGx0MK6fkY4u4yvXi
pYxuVqY3E4l2fPQVH37W9MvWyGXmClj1ilrD7mvDwsxcvB8fSXCbztvGTPOwlvQs4uAaQvU6xyo0
caD38a0Slx4htAXWOWEKedrhFHfK3gbrflkl37K2tU0r/LqqvB+JGKwRR5WkPKcGrgDMjgAMwSoq
dhBDi1U+WBHmv9QyfC746tfbcblGB+5lVnNINf140/XoI1cX6Obe2n050uHpLFQlBwU9dQbChxkP
L90RgJjtm5SOdReQ7hacLJ/J6Fo8uVvbhT1B/4FL7zv06EU0ytRtHgxW9LpzQ306BfKOqY4gfbJr
/ReQgCja1IkpaQuYIpFIb/XjM9ZhY8tLNiuVMnrV6GD67IHbN+nRcfu37wsp3Jq0Gc8hRkhHLKrh
XAansqZfMbyNNwohhtkrvnigkErH0LQVnBZ7yKZ6Pf/bbUn1zBWCkE/Fq/le/b28CzeMVgG6+0/g
9kbo545paRIL8n+QZ4RluyyBKh27LL3v1nKxiNGiwl184ArWmwqdthyAhiBagVnkIRmtj5YcAqGH
xtpOpnsJ/rq8phKQWtAUK0w9bfSIUawV/vgNwgg7lOcLhuBjaoEh9ZpVT4Muv5N1JSztih1p1Zv+
3TtJEZqJXpgC8ZXFJKEb5fAhXHByWHd3JA/oNHJlpbVksMUGrPXVm+z2ZvSsD3dYnx2XtSLqDbLt
UrT6xB2nRTrYANA765FjyW0rmqYIcNqh79hDPvPev5zwlJt+ZkTr4y4jNVgAanoLhsgIwLfx3vwm
9CArhmSRmEaLi6mULFRlGTyqsDN5LUCIM9QYmjjvYiePuVP4zAjiwNeCJBj5a47y/GbkqKG0iqFc
ODXTnbq348ZwInlDN3cDfE6BpSuNcsVjJWm2hEWemPF8R/pbB1TNJ9jSCScNm/feA+BSeQ60UCfd
PtiYB7s8x4wS6CM4NfdwogSmO/OqDREoFEeAtkn524/W9psUO0wjjsyHAAe3kHnGcqh12rbQ/4fl
cB7WGzxxVdHjlY/rvYxWLZvu+hqUpDciJJbh7c/2rKCuhzSx733LJAj0zizLSljccOsRUnQDfo3l
oPz5jr9INvuvllCihjKcvOzqWsRnxZwFzZIuvzMMbu9ofHjl0NlKnntOevaiG2q6JK6IZiA1b0og
LSIyLDrqzaZ8kc2hImlIdN4/l78LCqGGWA6gfrmOnm/UPfoNDRrcAfYUJMoqaep65xdyH746Zclo
2VBWj8p2KS7EGNLcEuHnzf872hBhG/AsnslObuk0gRrKlYIKsnZ3i9+iv1eaapM0Pou45fHzTT+b
HNsYdf96S8pTWaG4DVmZ1Pbv3VHXj8QsZI9eDmhKDUg8O9DwXPgFhdFjzyyXxXKw51lfsMf+qALm
EqI9ccUmV9M3rSmP6OHVtAnorke/4HDm2yM4Lqk6QZQrhCfh3S7MAIBTs/+R6LeYFFV+QzVxlX3P
ht9uUlt+plQG85/Kb/YZ4rRhyHqdaC1MuywdGplGzEMmCpsv0G6xigNAmE3na9ObPtKWxiAIrJ0f
GIFnTb/jY4cAd0fFUpBW/3gbEcJjFlrx/YdNyxWpl+twczJ+QxW8Wj2cV3eLrdCD6mnMVAHdIiXE
HaGFAXEGf9xl9/UGZFQC7LaREVclUCWH/XmFjp8ZBEvL93OEx6QXQFkUNVyXQTCbzxgQ3KrJOopC
Q/QNrXP+crc1x0n6qAGGocWuVXZYjRbdj/024Xn29VRcvK2jEauUORrlhGTOt3aBEZgwpoMqwjrn
HXecmbIXngcGZM1l5BORRDzYQrTV0QYN3ul8iNyFoKfAI5pDrGV7JXvwYGiE0b1WGc6KFAG5xenb
ett/n/OnOyDCcty87bjyGTuGw1Ty7bwYUJvoWZ0Hv9dUHPawCdiuvlFcJdLeVO6fLQeudnjf+ZX8
k6PNJi8Z6S3EHc0Rh9VIp/QBlDlAifKS5ATaqcIfirTN1YM7+HuX/jMdbaO94L+T5RvztYhwxct3
oO4pu7PK2F+d5pNnjhC/zzs0wvjkznvGKY79gmi8+QyQdPyE8RqFYHXmgbZToiOvu0ue0oP5wcAD
PPHBBHGRGiWdaeuWijp7opiCs15sIQc/0x7Z9FYlgNp8pB6ITVdukGZWVfXyZVnDlsDx5phHKxYO
yIsfVmCKUczLtJV7gU3i+qVItK2JWBZoDapR2NN7pHY7hdD8uZ6nQNxzUJdtEXdu6a460Qa5v5Ct
czqAh9uHWI3HWBZb2FDabRqRRfLZYV7MTto6SNOWZWSeiwNXnDyrggwWhNh+wU1MPz9u2Ui0IQKj
VOpTkcfn5nlqDkMJNDrhY/EiVMOWEQw4dF1AdGvBJyLcmMLG5m18swTfG+1601q6w81L/pTyHyF2
fX/FEj7hiF6wy8Yq5qTww+eAeFlJYThbX187Ax1WRZ5zS/rVccmKgYsU/d+6mz1NAsnhd1CdhLC5
pSJ4Hd/eLe3rpG4CJwywU99q5pMExp0XUsZgGBST4LJhWRl7HeHqhcT40vKEvu4ABW7ZXYfyXO5Z
/Rckncws5O+iMYu5BchxIUZZocdNyM7gRGq+mUC48sEWDdqDocTnBlc0yiQEAy+S9OwebP0dSbSM
RtowQ3C+w1/STeI0H4dP2ZKkSm4jxpsuTdL2iF68XXtPBCuSmFXVkvEJtJvs1yxw1hKAnY9WR7Wa
igV4iFIH7t+d/HrtrZ+e8IsFwvVYma+nEcnsxvELXau0nouPNgaGJVmmq/9mtZkSsbRTQUKE+Yrn
pKJ+8kV89RQtFJhOx/hYWVM7Ufht9JGXt0S6hi9+O97YhCZltuF/Jn2R+U49JCqfvGyHYS29kMGz
a5N3Tm0766wrdl69XM2b4mDsqTuvk/vepZgCJu3++VefcxGgIWr8MY7hgkF+OojwQzLOkIZ/DTY9
n8Gwt9d3O2hlw7u61rlnX1Wio6KPuQyf4AotfoFrvJGMHFA5oMnUV1VX6qAQsDsf/Edfu+ipPEp4
5b9ZCSKCOogI7b04+r0SWehfZ530dHirxgG9fg43iLI+1KhoA/6lOTG/6J2oHj1ahRJ6OGod1mtu
P4L/IU/dWqJTbN8swRx9PDGAZ/V7k/6rKHqe3xldejGoJv2vp7AZTRl02EhwSHg31uONKEf3lPBs
Jqo13FWNwk7FPx+AuaMbsUx3b6qVbg6RkxbnZxX9MYhsruT6tIF9cFQI8gJPPcZWUfvtqYaIeam6
7l36+0sYEfwU+5BezqQVlvRV73iZ2mteaainR+cqED54y7epJkz6tfpG2jZ/hOugC6CIzUCs5pNJ
KjVFQdQLp/V8XYLRSnOUeGf4jP71AFs6DOJVmV7jBwwY7ixGiAk0cfzf6dKkKwmqSj2TlDzFigdP
oA0CsuA85hB8YyBA+6wkpiu5Azm91zEBo02bHgE110lz8biBKq9dckqfko8bYBL4w1TvwvQ4b+vw
6IVINBbzhPbCikiVovR5MFj8S1HsC1TWZOLMu/4wKY0hXTKKKtqyNHVvJkG4KVoZto6UnLti7OMZ
MBbOK3yvD1tqfQDEPPOK9qDCPn+NL9QLHZxwvaS4/gk5Nj4x40ElrJM6y2F52rlHIw+b1NOmZEGA
DHsU6KE1XwLM9K01kTpSH2aAVhs6KoMR+YdwOixSAXoCt0rkWIsngdleA51IkAMQgnjijEoYbnOf
dFov6ONKyEDXv51q0ru0WMx0/QdKPFPAMqolzG+RRsdvplTe7WROMqGBMBORvtc77BlSf7Mc5tEa
4BXetrg9IsBvHHqtrIlJFdGSDBuqR+kN5SClY8uBYbkATR630Tb+rQhy+cBoUqrLDxQpXDv2SoBW
FftVEv1XsegbJM54ESSTIg0e/ifPhg2dqyxYMq3rwN8bheozaFkunnOKc3k6GMCPgU4m0PWLauOn
5Urpz9DOTAEHrzbwNEBY7jmCzCU4wP90p+cEu0NFcO5h/6R4m6BmKiuTiO5jJ4m5X5Um8iEb9hAC
2OHS2RhPlNSIcyyTWn8g4DKUbtCI18ciZ9Z/5YvUjjt9NdZU8SzNVMIXNQf5tQa55kBlNvyifrbj
roo0WU7N/Sus5sNAENFuXUpxl+wuIBUN7h6r9gU36QBacq3wJPnf0N5qKWA0r7yoRREa4Q8fNjmQ
wa4PDDduGzD0+KYoyHD8IDV/7UJMcmPmyH+uoqER7HddwFEVoeiL31iHFKE2AtMS885aAvsGkTaR
3NERdddpDSe53PeDhMW7ibMEhjivi4zhzgofjMvbn5+C0KgDj4AeS02JdXGz1PGb+pTfTiLlvxQP
v5j5XPeI7FkH7P4muNgOnxaWNThOZ2npT+Fl5T0l4WHxt2mhWYZGdV+bYrFzZMVqytHLvVRavGao
R6/fAVvP/RxZzW+04p7OWKugWYbmCPDA5AaGAEuUTMlZOgN0DLmEvUTCIhag+t9//DpQ4qpt9KPZ
QfR4eCbVJp67z8eQOC3S4WZ6cq6vEBu8rkYnnckl9XUCArGMCElpwBGYcRvzHgmyqoQnmBxQej5P
quq5m/MpQ9vl06BX6qq88HvFZ+FQgW98/3HODgo2Az/7zNXMn2FLQ5/jae8sv804S22RsQHM9s0A
C3OaVthA9tyeKr3vGhGQiJoSRCbZFQmTE8m0JSUsRkoj/FyhmY6ghpbE2G3MXzrVslbcu//z80zR
MsvtYpue+qogi4s6yQLD3c276OKNWb7dreVXsvJ9CUXNaSJtHXLVkr0j9FCmz3cELoOdRpoZeFFo
6xaVNZSMAtHI6AB9kENXF9iX+H8BZbu14KXfmtLVsfg6Sbg6L43j0XVzWgQzeg7Vxx9A99NdL8tG
gYKoPsbbcnlv5MQCQY9P8MeOivIzd306wbUQCSsVPmH9k1aH9kLE7Qiu4sZUzRCfAv1pkmjUDT2K
ihBRjvZju0A4c0M2gz9rq96fqLLqw8mYHnDSMrIoaPjLwknM9PxSBTNitdgCo3mibgePLKyaOAll
XTTHi55oeQk8lSczx1L02B65r1uNVcD1H/5IfU9fIe6cwjNH5UC4A2fhdHbsfIj/0KHwQJ9AtgS6
sqL24jiuGRi9CzSI5ytXJMEpCydN7fWoehlECayRGDqYmSePVf1N+/D6tHsUWPwqQAtEMp+Borqc
FqmDjvNJJul2lGRLrMlLipCNtW/DkE51QTHUmev5GTM3MgIwT5KwPj/f2fa2nS1TuZgnr03zMibp
SVxpwSqtaPZNUs4lfmXWUwiDdVeOplAVzzoEByTZj5pe3M1R8VtfSSN2dnoPkFsK8baw2ovXRzNg
m6JgWVHStSL7x4ev2GZTlEea6usyp/StwxMDpxdptLnd+DQA1GOb6/S1nMelobsVem7inefzd7UV
vLzQ/H++51GHs6LuQ6NChODCrBCS6RgKi8VNwAsnc1wSkGqxPsbVGTTsIs00lp/aYxpJDy6S4nEO
kfYtcz7vFVxcg5Hhu27ACzmQzlJbqL3JeqM5SPQbE2kWiv+onZmWqDraFC2N6QwN4h1lckUtYG6S
FWjZyKdZ9pAFaKwrfkkJptrMzPm8Md6HLReFI5edco4bGGI5kjwLirtOM0UHpNiydqIfF86dF8UZ
TlRHLRYyTfsnB6pRlzz935XV4YUt9+wYTjMV/HJuu7lpB9C3DB+WueSytFBWgt46W8jMC6gtyExS
Qdv/s1IlKU/QKkpSqXUAYcI7TogOmOpRmR61jiKoEzbC/T8U54YJh42Slxx1HDGYpc5XhsgwmFLF
H6HT7Y7tOtuFmrBdhrJbLct97mHAm+evZL2d/Hs2BL8L5lnQw96qnrFrv0G54Kq9m9fOV0E/Od/o
fq/huQHC+l9nu2CXgAG/JK6a7mUW1KAqhHHTb8NjZJKpA6dThV2YW98AsHaDnOS9alaPGqzsiY3y
TLqv35sfJfGGghBtDQYh2pu8XlM093C1tR6cSf3l/Ks5iu5uJvIblui4cPVeCgphwp3fIkzmu2+I
EnWWtMmKGAWw94aWQs8IlVPFrhbhJIFv38lsgv4BpGeRfMrY1A4ZBcTSohbO4QCxE336jgCGFHhM
kw1nxa3marpBQeR8FKn9xNR8ZUleyy7PXrALuw4rW9rEkHPQgQtqtijazlbCjJ+4hPVQKENEjgDr
5ednGViGdKtywEO5ov+CoP1/fqB8GMrtlM0za9rQxw/5zVW5NE1SS8XWVOjIkJSOpUhXXwFxClAi
Prp/162isad5sc5Z0YOpNHzZOXSdCavSwrkpySP7QH1jmFkqlKSVl6W8AEacWtTwz15/xipKIPJC
0zUry8v1NlvvmN6JR5MyF8XyoJGcJ8j+c59vBYdoU1sktf1sGSrBXMPw1xz1cgNza1ACWEZG0tCC
wlftuikt4bnITm55cFDBVz0ALOs+ANsldtZiEh1hWComi1UlZjoLQFtPG1oIOZjFigvQqtBmQIfu
txKPKWTG6F15sDCDUnihomeBckRk1CSL0e4SPylP2scK54b3jlJ4VVzjUCCJfIGjFzIVl2qYVawy
Uem9/sCt6d7X9Yrrso/SmPgtn/V5KNxQW9yMFeAIWFnIGB3fu1fn7vLSk3jIEba6zBX+EwUEpw27
zAkrj4E1aJCHw/mTbhkuC7+dvLzuN9w+ozkenHLSMidIWhEDB00hWlFILsE151o9gCMSPgkGWzCN
ryjMP1eqTJlxXQEiPfjgS3EO/y5WKmqowL4I7e5b95hlKZhITxIbsW+zrYhZ1hR/HU5E/gxbYL5x
nPaHIQOUPtmeMBRkAGjjpAzQDyyptxq4FtyMgguZdRbIT3BO+AtUaDdO1FvmY/Z++3j2OFcdEqkl
ZbHffmh5ARWURy2HPnsDVolZ8bKqJH9OE8/ZKDXsbkcJHddztMAUyEj7WQAShzyk5vmXsCyo38bF
Jb/DdpcPMBuRrpoH60SwwhbdsfcjjfK+ogKBKe6O0c5juuFDpWXwX5ki4lDoQ5p7XUEF/D3mZRtE
SZdTD6X0wG2UKgqOU02DN6Mqw1VQVOy48k+plWNollJ3s62c2N3bNHOw6jzUZvIy1090Z/JaG1CD
3KNw5YSEPmlS3LuYQ0LSV1GJXlm8pf7Xzc7Aug7wLnUrqC32fx3/rlGWR7JXvQAyzd/7dqqKxrrd
uEvaAupEa3fn0aRs/30Pv6jh+uftkxHb/WE5H1+xjWhwfHNQZaWk2zqKTtow0heKzEV75O32MFSq
gwOJ5Ot9sobJmNzNVj0EVF6v3EwfM7RNyBnAKE6r9PM1QrOI2xuIUJWowKiJToynG7m4oCjqHYTR
JMPCNX5G/cRqCiWzRvwlkSdxY+7fIbkw2967kgK3ExsAlpqLBeiKBntXIM6SCAVzlnlJMQW0NgBC
vDiZrMf+F40vzlQv8lZoqy1vbLEoDxr2mUGVA5y0YJKoTPlJgNgoDjVkKI2evBvmrA0+xh+rCpYR
XwNwWk2Ehlnm+tdy2BH5tYwrgeuwvOIL5ab6VvlZtBFn0sdfTJGoFfMr2NsElY5IuYIfseGVbx65
RdnZf+vf/v6EIp/beM8OAUcRvmozlMBERfkJPgIMqEEXCBpV1r2vsrTEfLrfAE6Xt/UMqAVbLLbv
CosCiGmia+D2DxrLpZ6m5gmNi7Q85FET+exG+/Kdz4XxLktschnZiLFJ3Jd0iK52b/ILfT79/oko
7q3N4/sEcOk5f6V6uoQfuUfZ01o94pA/14Ctrh6AhAb0wuwYcsPaP5gT7ttnEhbQLQ1EEPj+CVdy
h5YtAPSep6ZBcHTZxriZs2c20jI2U23v1Kl+i3nNIYnDqcTGCDVnCb1q5BXr9eupvBNxfI3USKen
gIruNigk0B5tU6q9hPAvlX3riQ39Ae9HtiMPRyQ7vkH8Sl4qk9qjisTHEcbfxqPx//a1CbUcFenT
yOTQ6Ddaer/iybBCHnm+nCE5NsLkivDpDDBouUNOm6XPkdF/wIS7ZbsdOr5su0qfyqc9UEabxbts
qe4UBSW9Da4fxxV3mW+nyskP1Wfz3BJZBgaMYzdB8TI/iCG7x12oeXpDOJc+JSuIJoW847AIiVt/
jrAvHciwBO7GXUxAEiAk9u+iAxQqKT5mx0z3nOwlHBo9DvfknIr2wrY84MpL0kMmL780ifV5eNCV
+GgsvPDdObolFBZBs1Be7P7ydv+I4tcg1PMiuL4R8dWxEtuc1UBLApH0lg2B/qA/0Kc202FEcGoV
L0+11uDlwLGctYH8+CyHYg2EzSNSLYWh+BcNsfAupnYkN8ts5PZv8fmk7H4zGtoDwZXMXx/yRWBc
9jy+4bfRCDwXwYi4qAxIhp6MmAp8Jcyi3sMKirdz5Mr1juVUu4vdJOcXsyjw+gx6V7f3GVah84l9
WshxZoU/A2FlpHKwYygDAy6Na5L6v/STA7vgOVk7MtR2wmkVOIzhNXdcUgPR82ZCBHV7EGrB9xYa
ATSs7x/MfCTKCKDir3QYcAYETGbDFNQrHJ62ajPd/JeZuJlRArQNLzX7ebJdxKau8hmw2nppK8zZ
4dTx+aXnvb6Hd7o+ZKdFH9/fW/znVNIZ4bhoUm0sf2q0s8Fu1NBL0BhnUDZBoaXS5VukuIJOI6kF
3L8e8WfhhFEgSwGThuav0RTPBayQO4VoDhe0ZQuOweZDvxlZWKX3pr7I4i7QkzIX8OOLHbztzJnU
UD10v20b+vX9b2+ODrjpZU/XQfykPETI388/T/nlsWRvBemj+FcTydZLR3vtqf29un1mTHl9gEyl
vOPcBx4DRuvRTBzNi+TAHUMJuaG9xsXFk2T/G6WdcN77KbCfb20lg0Mrdgo2LW/nw9TkZ0xCbFZI
/GIlf11huSiH5r8191N80QXhAgDk8RdnOytPYiy4o8dlFcJWvtseLGFDK9PlTo5KGITPyyn6uQ4Q
N7Feo9dCaZkDAXxKGtvoaRS6aidO/eMn8YOS0OPoHwgzoupoXZxOxMWOz1tBzKtFKYC8RbjGvu7l
8P/twr/a15jGryNzhJNTDN0r1HHdmq1zq4tlkKnVwKlrIS5ggPDNhNNI8TJfYfmFX672tJJ0FEtm
ZS/Y/9HPQQUNHisl2BL/DKTyYyiPN/xCfveeWC4piqGVn6BgUWxiuWTiJoCdRmhdbrXIKA/XO3Wm
gPvkA+ak1Bnzjlu4c6J83SvAMIgJsvjlHUH6zOy/8G2Pjh8yMDUpiFIBiVcg/+lbOkR/yOwqRYUQ
h8Ynq4aayNpldKntjHvnyForR1H4G61v3+JBTQ7Zzpc9VjVCEP+BMsHkyeFluhGrpiajMX/X/wKw
JD/tAF71p8J7zKT6stmXJGA0aK0qp2HKEfUJR361NvBS03bbNvxODqZQjqmb9t6/iblaCIojWONn
RgTzvMw2S/Kib7/oMGy12iq4dmxzP9vWrbqgU51r2nNA3glDg5tG4G9fx5S4GnV/42GRPHIdz8lG
T413Xu7NU1JxRyAa47VW//aC6QERz2gt7Pq01ZP/sYZjKDiBwjsF4/es28zsFJ8AsyOJPuck/9Zc
dj6v3+1R4PT6lCzc8gRXY8KffVfPIW/jGefdcSTyP2pnoAqz8Cxk5EgJYL9ueuItjJyirXRdd0qz
iPMRgzLvPbkGvHclKyXLZAv8ISwnR/uD1pKD6CQBVWGxMi6N2qiw1Hn6euOtZoRcpN/QTiLcIQoZ
zW6+qZZbviboXoe5pknpTgn9uB+m9bGdJiQpbTywL/nj3hzKDdtMpH0kJ6HQU3PY8pkMM4BRkR5r
jj9x2Iqomg2xMDEPj/DCW2qLuRgLBJtmw98k83ihZGplHQt+OXN8bt5GVctYVtzOT4ooTB7PyP6z
X5lJQ/3J0toaYJ8OPjTBkKG0y1bUts6W5XUoy39mmtrtGWLH70T+AMRyKXP1gC0lWBnADZbWqSq5
9zrBn5BPFQLPTzOPyOq6Nz4KOlfR+g6A5fmf/Sq/iYksZDIRL9d0yS0MZWuU7FBBXZUJp8yd9C46
EWswboRi59E4ELfbS5nhF8lUGV4Yu5xYG86qL3haTEngWTqryoSZJc9sABo1wiX3pgizgyGS5r9W
Ag8Y00QTtHQRPmXN8jlfm8DeDajhIYWfwphQ3YZsLmpjt3fXkOUQKFUSMmz7QkS/SpPDu14Gjk9T
MK1YsfMt1MarWm7vYIJ+rS/jUF77h52To8fxpO3le6D+VVY/XP5MDIBw7SuiDHcY1Z2jNJkchxBn
MHiSzqaf4eY4O+aux4gmpn9ID1Raqrq1cMlMyDqwPkc+L//KHGLFKt9VPagH2Yfk+49TUnElrj2n
cElYRZ2F+eBDC3em9BpOPywnZJZKjX782DlFAcfBaiIk2PHlVqZO35f7muXMsCMkazH8Mi/bB3ti
u2yaQXI5L9Gro9NndXXZuY+LoKtCHw1ZjJUcGVlP9p1kceOUHz8I/KbY/hvZFE4b5HhP5/2EmXVY
tVgw3gs6gerJxiNt+MWw4xVYVpzi4703kBi+1XbOyRPY18SmjFCIRPI/WWCvJ/MFumZO55qvxlwQ
xGHA2IlGEbisXRLou1/oqNoGL64sY9ZC+XfpFfhGbQS7t+l6kqnOH1VJARuEWTfdNPfvFlE/XIuj
NUayaXIAw/wK9FrPFEdX0c6QmfhcFyNeLovVS77FqX3wvlm6Bs/Sd1RpQhIHxec/5H9eM8ANq5Qz
ylTUQM9I0iwrg4MJX4b0YAFIBDYHq7CPFfnF+eDceWhNq7XV+TkIJZHaB9tDJk35kJvRT2ijmU1G
ssayv/C4hpbO/CcvH32Cxr7CWahL2AEQTDDxtw8gi95gPdHHct0l34Y5s57M35Z11Wy4LpvCbmMV
QIBQNt0V8CpxkpVnhuvAqIJv5/k9hC2CnxQQNmGCub7lAhn1nLkmzZ4NHvVT6IGH6TAP4dy7dT6B
jdwJqjxSfYk4OSmYXwPdRFV5AW2RJXV1hb6g8AX/BhJrkLoUGSDooj6KB0pyuwaqcmjPGIePrp9Q
mWs2RKaOYcebO16BJU3uNSJd2ei6cgcivo4Jn4rucmBYNQkQakS1Nw4rwHPxRtLl4rC3M6oHYrSL
SVBjzEbfbToqSQiSRX84oFmoPaX3b2iBOoX+aDGp+oEuZY+IjmuJ3KIa3JO4xpc/SuArwbHkO4jc
TeKvt3kMNCbXNICTIKCY39hwlkh4woXxtUGai+VulvR7I2VCm2ndxZOn8BveEb00xZgJBUYDrdx9
k9RupDDVfGXTxN/frzF1ZRzuXSOZW4m7pVRUp9y8KSiLMNdisZE4wCGOi9iySS/YDLeh6SB/Cg4x
zgyoHkwzA7EE6cJjZb+Hgi1dSDE3qjhWW7H59dYEhpDQSFb0Vf3QU18FxmnTdWWunN3yj29KORcl
9IIRAg2oSFlLnS73bufeYMg4iFXOJYSSrs5p4C4uCqazvwdgKGPqOqUt7wXKs7W/VF8KfhwBgtd3
U0KJr8QYjmgagXdYakM4fAn491mysK+osZgoHeaH/VLXA9iWtEi/yX2aOoTpFtwdGdYMb1yGy+ts
W+kLS++o70xy8E1F5pI7KbfrqYuaV9wYcZSl2msMdyzunb2ZRepl312eqXgg1lecOiXwYPF6b1Nh
wsPWJSOx497e4Nmdm7JAdzubIxrr1GI+hBJoz0sOwE1F7ujTRVHoPHzc35npn3cEcomzMZRqgyot
TvG4EId/Fv2ph+lqfo9TJVWe12XqJ5DlRwrmBC5eqyYt2FqliwCU0tfch7sxJTQ3O6eewOjJcTL0
07zeIl5du6xL8yMvwFMLuUd3VR9kVf56UGQCk1ysJF2kYNJeF2xuzewe5muBXTQcEECXDvMRfwtr
IIkkqMMUgd2/IkTLMuBwpAzb+/ib7pyxHi/7WpkFDje0eOAZ7KsOzyRsiV0XTPAB2VBmCncFFe2i
Q8VEoFDWvalcXiPNXYCVvHsy7EiVGiIgh4bwcn6sKhywb3Wwa8yLLMoPUb+j40VI4k96sytFuh34
Vj6k7lSWdEdF/ro5TXZMfi2WoHd9FDwSGuORCXG8pVA4LOX8pXmASTlrKGpDidIjq7uqqE0nsw/k
zfaDriCgWEQxl3f1WsxGGruFAwaySzIkt/9I95LQH1I1OOW5hRn8sK1uoUrHBQr/9k+Ltl6gW4bd
UJtpEUjoTqsVadi1zPSS5UyRQ05x4kOCcxK3jDHdR9cESShhHweGQKZWeCTrCQEy9ZcMl4YTSHlT
MVM+JZv52UJKuU9U02zTd3IHLdAKVEummzBPSN72qzLKRGdATyeJEsEvgk3TKbj5m9tMnhENgnNu
h2hVXvgybjBsXccDs0uXVN68OiJ0axqIVkrKFzzAKrrbSrDZ9uBcFirjBQ9KuLIZqR8AxbN+wnNq
wR+w8G3R+M1YHs78YQYVj8ciyKr6Bp/shPHb5V053AfSitv8anFpH6i+45SZNRh3SSKOLK4Dvqfn
rdL0TCTugQApuRAd+gcytg+S0H5aUdAu358IcYPbO9+wS6sp4C3E1cUfV/VvFKr7MB7eElSPsRka
KJoNMCmSdqbUDiQkqILeYrWVmqA0WsxK3T1bRb5v/U1lkFYeHimJAPhlaq0z8Td6xtFLjTA0CPI9
nAEFmwZp1URt/jqOAilEBskViyzvsUcL+VSVzgR9htIxT/2zvuyM3Cjpg1bj3sYLLM6tvA+oR+JS
jtU2gwh6WlyNIJrus7SwazEyDoFOKh8Gqwd4ehlY2uJOyvAnFEkRIc+GblqKlFiWpJB0RaBzp6rM
Sn/DaNWXsDoinRLzFeagafcCjrGaSG7cZkuVDGuLwl3YdA7D7+VFYeCyrW3YGRqjQ4V8vjyBvw8R
BCi0lwTt4EC+0+79BLG+wcm6fGdzklqKfv91waCsNLQyd1BOrTn6IBfscXxuihai5FMBd56MrkVr
sVn09zrlpA+tJC/510RhBAFIUJnIywgdUpXk+lKDOmGFce8a8v3kTmRrG76uBOJG+OjE+IO24GbT
AInHMQBMtPbAkxdyOKBtwjHHqK+lILkUZsT8E+66xXJMrceon4VoMDmmB1rdCvQ9tebR0zMY3w6C
6FroiSATa94oOUN8qfyCCXZE+j2B3IZq999uvvVsbUFKFD4tk9CQHZ8Kpm8IqhBYt3Nh4aw4BzHa
x+/mZ1/41Wb5kUgGmoVk0vVTMZqQEcTXz+WhQIMuekcWieC48TGEir6Umx9keR5DtUXmv8Mwqypr
m97+ncIqJs7B+9HEmSHj+s3QCrmU685zDdcPaKUoXqYJsGySdx2vy9+oJflrFuQYwdlEMjqlC1Lg
Aaqy/1SA+pN6G/QdvixS7NIO9/nP+zpU/nrfZJt++26zs+5bRCQVxtCcbdwRvKK1IMr7y3rtC2QZ
/1yQooT57wEYo8pqSaTnnsyzIKvcKtZcN5Y11Fd6GWv0qkCtSa68IpaAcUITbS/GsIUKQ3cS0xC7
sD7DtO2NxvWRhEgwQ1E31cxXedQ2cCyX9fKBcJ0VNPli2jwDWrlaI/w+B04GiOdJAd+WdTkrgT6b
Yewk/Iy4SWhoJbEcj8Z6iYor7BRCfeuxpIUk1nJrEmRYt0UfPpMfEbZG4fHvjqspkRj8uirfPCvv
BG/JyhgjwFmnwtrty128ch4c5iVaq8BN3XNcZuscpnd5EFbrdb+5rqpoNg+GLyQkzjdS6AqCSHmp
XT7nh0B3wEDAJpzcJ9ZGf8MDx2oYsWSW4FcrnURnXsN/MZR21mLeoPPnB5dBbMABERwAn1YFewWm
rkr+sG0LqXxfiuedQvJA+kt5ZoQuLoUF4KK0Q6XzKkHH0f4NHboVOGP+CoEKqvZjNYW5G0+F1qRt
tiKapWgjG/DjwDG+w4tDmvULWNdAAUS64a8xDvctglI8GMVSTJZK2IE6A/vX+BlyyAyCAIM9uDyU
gjK90PmiHD7l4TSiGj6N/sYvg0qXL2F+5iRv1AlQIAAZvJMk9ILCFI90Aqo1Qf9u6JBHeYWHoeN+
xYDqjLrtkQQK6PXLzS5lgpi8jXLYdiIA5j3+pjrw+XrE8LuU8rtI1y9Hfv2NDtg+NLIqJn+NTWCO
4m2lk9x8dCBFmZjFS1LGTfURUZAT95NYQl24yNEkMmgqA2bn3vuqWDNX10ODNC3zd33ysLa1lQJ/
o3GQk5rB/7sxxGCPBS776i7v9V+HR6SOUHMzfvFTmxTcUtXtTkoGXCIexQ+J9COdBp4Ywe3ixJLE
9JuLceVkAglksfM8siHuH405O1fcowWd4zojYgcsVXdKGue6VomE1w7TvKR7PeyMI1AGNKS8Inp+
xniarxhH6kQ8qZwL5NQXmq1vlou1aqJP71/jSP6NB696MbWFnrRTb9LUmyXJtGUMI5+QHgqoE38s
LgZ32iC35B5jArRlGKX3PrltKRrgxgyWMKebsFdWMyNL03rsJTOgzyWYHZkyCVrALSIWqy6P+e6V
Q+jDIWd/99hID9+pC3ynlwwJ6IR0V9rspNqVOzPrAlAfe6aXkyMKI4VKhgIZgFxoUdH3z5zzKe7j
pIK0CR6+Jm/pJtxiw/PKKjfTYmeof13jYQAc2rOytA4oil8Iadvd2eomuovcdhT8pu71HdW+Lb39
0DJwa84TH7IMq7t/l62+L7+djy8o5w894Nd+LmsPHFtCex44Tunl+iO/gdKRzSOpRpe0j3B+xICn
QIC9n8ufzzLbzLIe63TKXAkHob2ivhLDzmWvF0Xeo3J77OOOl7ot485onaTSSjItH9mx9UKbXm4O
scLvbtI6fCw8TYsBjefaF3apflBs4s4dhFVdHD7zsqq6cpROZTNQP/B90UZEKG5NtFzDhNx+yrmO
8f3Jc7f+gGeWDmnLtbcwg3KlHFLxtHTxA3r9VYhfZvuLLS9hRRU5zU5kK5B6hCMe9HVgq6jqaE4L
3UOnfvUzqO0bzsHkSyYqT0wCwvv8QDTQHOqFhCn2/iGbPFXw5AEYEjRMREFakRyV4QKFNsX11QnC
Fdx83rBRvi4tA18bEzOulI5UWEFmCgeI57v6hzeWMuelIISaNSN34RB5+P1OJIKtzyLl14D+HetF
gvDCNYtfNqzSyecCdkj9GVZ+FbDzYNoUM0+/V612IOynyThqQd5QznY7JiRgjcElGKXVKRXaQHWc
P9rUXAn0jQIS1/Eefn1kOanT8oWqm6M5wOiUeG696mhG8/YIna8wUJRj1WrLnxxvfDuzNeweafRf
4TiKFZusEjna+g3unecm+ZRaIRB4S+7T24QHjDa6EnulzK+XraINt9rBHnf0cf6L1zCf/ba2n2Sh
ACmQuEsOjsYXdVZYhnFMisjHFvOKO5fe7JvmkHrke2t7kihPTF22IgDtAJIAuoLHrMUD88t1gn6Z
6TR/3rxw8ED56bHtt29cHm8op7fRdqXXr3ETAn0XIQUzuTuTiQBLHvauR9XnpazOZ+/dtXJlO3tX
rfYqcqIMAmmg2RGGwRdJiSp4Y4D9Q6i+ZDOHwxA4Kcs2hdnb2QYCBI6tKxWKsSczbnIENrqGNU8K
MyatGDtYkaiw3x6HCw4erYKWq/iF9DmvDdD9YFmYR7ObfgqkU1Eo/THYvTozgADUDum7s7RMsjNn
aCeUrCcZNJVrmYAPWl7wdqAi0njpd6dRnb1dDnbAKtoBHV5ZIjbSScAxDJs13XXDbhsXBIpI6NVm
JzmHt5CbJl7xUZ7GImvOITDMrZ1FAC17vaBQ80eLgehpMFJNd1B0WPb9cHnczbwkEp2vaCIj13zF
IGvC3pvaltwuSX0PmPXpyFmCzcLw01UnRU2h5GeELUekao4JzFqQWEP7YPmYteWmBazXmMhI3Tuh
LyRPvXY4TPIH2jI2Glp5al5xjht2d7wM721H/6Rquf4kn3Nz1sXttd2bzVnVvrOOCYu35S0B+kPa
7MUig17XLTh/EDMAZcjyH5AskUMVQz0g1vd+NZr2SpirKiGsfBoP62VjK1JGtgRnnYXRdJpTLgLV
dxShbfIMmRH6JMLToPh1L/0DaJab+Boejma07OTnKSIreIC68eN0nHX+AcgLIN6bIIv3hTb6euF6
hr1ulWPy+7PqBpT9Z6uwCu2u62ADmTe7EYCs85G81qSjrrB3+BP4tb0SGIg0nPgCov77DFrlNcXR
HzFsegsNb9jgRPru7kwZoMmxLMUHf1jvLQs66Q4mKxYRs8EvTQokwXTYWro4yHRUMJfPWwKa1Mog
0z14vXV1q8Z1Gw1feh2nNVpjDESDl7Kg1Y8ZG6ZHnVzez6hWlNztVGZp3CPGB3KiZ9IO9lTtnpvd
XOKGyl3Skw9ltgOP8fjGaWOwhNlTDkPT+NEfThv8f30TVpb7l3mMx+8w+SsA7omYohXWtUUz5YBK
EDmvWlP3FrXzeS7Z3SLg9Saek43YD76QEXn3t5cYU/A20T+Y/i9gAFWbE19IVZ26ka9oG+/19fG1
VvY9z9AoCtTE7fc9dP+nuCYzfmMiYdADt93ToA2IOOOzcBLF2mIyoSGZTP7U14g6vXzgJJ54ObR0
FaaFv32yzEHa3Pd16MFU2GOUWKanN+4agIxOGlQtiuuVYRN4hVZaT6Y75+6koXLQgnxKqPcknx5q
W1HQZbZgzV8j3M8A78RBMMzfVRaLrZBsuflXD6JORrS6vB9Nz9UHsmCj8pTbSdSBRkjbbeWdhcr9
2bVj/VKTNtmzW9Sqsb/0ganumcTfdj05zWKa/8qh38kX5IoPSg3UUdkgkAj7eXgwnE76EDYacK/I
R/TPbCgJnQoJ5Hlp1y4gHjFMP5pJrSl56gk1f1+BHysQ4Q66CQ/KbVkqgiehTLeQ3Po3f8WTJJB3
92mQBjLhJYRd0hlExIpUcQYzgRGb4Q55dg7Dx2E/cUj754sIrQ/r4ASrNfXk8r/PaRaOEmpScwmF
ozulJLSlslgKXudvxaHE2KTNU0q+ZIJFO9PY5x1XKz/nRtVBJQRw5kPtVobnuQt5m+C04VCAaZCk
LntRRQamejX8rIkfgpsUJ7ekqnaNBt02YtMAlb8T/pRzQ4qsVuCH0vTK2zsnHwLc+hE2dezTqRxn
ZNAy9DiVPhYMFNqseggC+tyHdX3HT6bRlCJ6zNXBZ+bABjqrGiyxJwyWsDVbhHITZ74/s2/fMMpX
k9fWJ/XFReZ1hDadslnUXZDx8A/euihn40NUpuV2RktFW2HDwm8tL3iLcVVtNazdUrB6JUmLXGia
6XSfET6Kp+yB09wmiZUb0ZQG7FQEcoYbinqJL13/EjgJFxRuZNiUu1N5l4rSuJ/14lsCbjVP33Jo
DLQly9XIT9sKlaP4qd7gPJS0VbjVtoxHxzOqT95CM6XFfT7N7bof/WuoHTlk6XMWl5aw9lZFykvd
Bu1uT9z1uI/ANBXOftW0FjJDccNfUVfYsakWo2sv8CpNsJA/aY3lFD9GQ5pT0qlcRxmd7dad9tQb
6hTTQirbyyStcUdabedrjcSLirr0yumVycpIafTjMpPZv4H9kBobw2IgkAMermbJb22enIRQzIod
RnEuMtFHTT6tEITIFpaRw8ckrQLNEUMNNilk8UQYo6bsfsNJsTjjavWdAJ9115rVNNTPPWipopAj
4YP2fgVQwA6QQ6c/vv6MvXs9PwhapzHdecfIXzll8JN2JpWl0XQi1uUhVnXQBqaHpHRQgpwK7azv
B6RH0IH3pBf+n5AZyfR8Vqn1zy36nOAbTxMELQY7yBxagLMNdQY3rvr1W3VVSYpFk9H5mD6+Nv+D
u388zC+AUBnaVAsJrt2rPz8bw2oW/7T9HDlsYoYX1/SsRhGyATM5k3Hl7rYS5322U7HUqGxFMJcp
xAL/7+mWvPR//ealEvf9CpryLsLEN+jb3a0LL8qTksc0IKfSe3tC39Kh0jZcyttSohAXo7NLO/e5
xD6/oEi9EFAvnPhCoRIu1At+rMSBIGvWJq4OzlssiRdr6lR4bkm2F/n3U+1qd9a2lg6hH05iMgEF
LdRunrdVkaHi33xsDdk1OdcfgLWwrFX90XwPYfnmE8tyHAvnAGrQ2tjHmcbAHsbNIPYnkVZqcC2s
6HRFKsfxtcFc3E9yRkgaW6g8AVdVFIMaVvPBVEB/haC1+iiaxfVzeB8BOKvugJe6mv5BBanpFmMN
U2iLlLLVRr16CxZn9kAisd1CHm0V5/yPam/bDVA3h+RZVn0tJQ886dmIz8GdSpQrU6/Zxx2ztadv
y6Zy1zF/1qCf5c8RvKpL3fxehZCHwy8+qHR27KvnJgJGWKqp+3v7PHxNLDBQF7q8IIuS385POkfM
96gduJMzramoWrD6llh4UapUxYW+2wMjFdc9Rw012ecySnR+QLICTIfpLt0h02/JxgZF0WA95XLS
9TL8sFZsYnaPyaQmfcA4/ELu2nDrAF5YCPRi4e2bne81+Ic7q69y4alIiY71OUCbu52Id2BPWBUU
9aNOyA5pSmJ68XLiZQdXnb6y+c3lZGWJkqs+dQncDNLD6oB885mvXMbLgevPy312T5m8TZgv5bNe
RCzXgS00a3ErLIA2ixl3TILmCHkr0i1UC9n8/Xtp1P5BZci+aqhc1JoiXk4OiXJN/D2ArDT2Vp0I
b3RMBHU41Coo76sDUhecdnUDL7w3abgNFLuBk2DE2hxhsen5acsmmjDgBt/D7OpvMP3lHtG2nkt0
cOtyoG0iXrWwAuAdaWY1AFPCaGmpXetJLCUnDsGIZprkmrChEnqjB5+cBw7HiHXi9W114J7h52mi
VbBPLzxpnuxiFvrIUW1mwNbejtk7iK+xOxxz5SiQXCPq96t4i0l+6imiMCJ+R7Y4/iivIYRCG4tl
aCRwyw7OMQpuZusbCuj4RhLws7cuB7s/vGd5P5SGdicqvGEZeMYGlDo3xSVCFWz9yr1UIavsrlS5
4Zhn3079uutoqebwJvBZzzvc3Zbey1zePEqbIJHrpH5J+q5Ps6NSyrcXEDUB1I0des0GqdS8pB8t
ducxAkYrBajtF3gAoTN+jUOplxE6+lSxP84qjuNo5FLTHtID3PmcwVAOULcXpjrAOzd4b2JlrKRH
rzhIqzdB1U5/9GJDybw1BoV0NAUuUEXKjVB/n5l92DLlfT7o7hshh9D/AMQ6hZgOeRiH3hzKJ45p
nQIqeTGrgaDkWVOS1Hm+ReQdS8FjtESqtrtYdsZR7VS8oIxYjBO5HjLkxOlMFQQZk0dpR1Fby++N
IaeIgDZpZkdbJZPhllRwnQdnM4MsaS41codz3lw3dwBs4I5Kl9ycw+5BHlbVFD4jdhvTgBg256vJ
AYl8KtZN6WcaiNVhdS8JusXTOfTWUcb3iJhbqpC+uSShETBK9UTkqzQQX2XVZAghmT5d7A5SDbKa
1FoOkBEfxnX34MhUx5fIlch5uPMMlOhWJboCPZ/DT4v2xn+JsJ/Ubpk54tDpZSdEZe3WIENsONaB
HPBb2fu0xeo0wUCrGU3FuPiZHxE0+Jsq+O3yR6XiTyUe0saRNyYDE0wlsDm9Kzsk3XazUXwbindX
2jyVIgX5E4SNtw2povT+dQq0pNJqaDmKZB27eMI1oXf0XeHp2epJtCddOmgIazONpmueZ/PHaliW
RQNpuzJQX0cFUSC1TSxCT2LERgbc7z64cEw7JO1HoK/jL1H7DtLHUESzDK6PwGr67SdgPePLUwIS
HMl3R4qOpoAydwaBsriP85rTDNgCWxOrxR0Lrn0R64YF2XuFvCJe1iwLwFpUnyUwtCflmC7Lx82b
doRdFD3DHK+OlHHaWEL35elvmEp7Wg08TfYWsGakmJoPZkTgaOj15HHx/jn1RlRfs/PNyM6YYH1E
/PMWAQSOTUxWHNMbNnwVCfDsRcTRwLgvrLwnOyPO2uOWH1zLiaBaUF3zRaIsOAaYQIxA6FSu6+oQ
tE8XfAJXrTUTQLMZBOcZK4snnlvQuXrAuPI24GVjgVIQeVS2hKOUM9gM5iKLrYEEoXmUTbdp9+dw
F3HI+5QfjzY1QZP9/mDjtt8CEIF+Ltq9XbYg+f9JcjdCFm5uTFFLAzeiXnysOs60ETpX39CQR1fX
SSnz4Dlkhhya7dlpvKLKWkIJ7ghK699dTC++8gASukQt+/UGHkKygQ0u9pkoGcf4bFY4G48e9hH8
Dx1UeW4XmZrW9r0aDLXFmswoQt7G0X5bjZtxqoOkbpXiry0AhyLcJZmApnN9Jp1L3xIoNH4WCBOs
Ek4yLXAFm6rBDZ9bfanncpN5DxqLeQ5rENRIoXlq/y37DwdStM5vbLapq/f/5pSWf0cj1QNTa+qs
q9VV9hiGu+mIseugrvhtoFT6YKgfsSQJnXs7B7GceS0t85t34/snc+VzSMd6eWpH+9gFxWPQ+0cT
hrVzHBQbjJVBKwk5XDqraezxKd4b9ZYqv7QrhUK8APnz+tJT6k4RB3mBpbKqX9ko9pMPXXWH+Ea4
XIHVNGJqj8zdI2kFz/fRIV0xn3Dlo+L8jQjn4esjK3qV7ck5cFpZYN5Z5g7TyVsqosGrEScDv96z
u287P+v4t4X3bo/nvy1Oid2VZkaLYixWcF9zjUjA48SNoKCrh0RkKAci6NMuqIxSy4qQCtTVh+Uz
A/qd0y1FU/qDUA/LGU7bPv4vwQh11VJyCaeU7kBtiURSUOktqgR1D6RymnIYRfftcGs3gX7WLP8J
eypAYsMDjEJ7R53RodXtNSPoyueC0lJAe7wbt17oRYmtNbsD9wzU81WMdhVBKZQH7tQY7ek+uTGU
8HARSjM+ZGKfE7cVBb2p60A9vpvYyp/D5/ICDuMHFXeqmideJIPOu18c3iiIqm3SGtIzJr6SnNWx
9NDyvs0oILgcThnlmGCnUnVJYK08R60CnBM0s/wDGTS11ayvD7aYUTqzTlTfKFt33PjfxdJlUPVY
Db57Sj7rxSRzObtQ8a0NNZlHrBZ+y7B4AlMmqKPkIJb+gsjaLbTOyPlRuJFn5ObbHdk2bysJRugL
dTief/2pDDih3MiUJTtBl8Way+v1fLlvcAR4x0IcjnOcLz+uSe1avcyIaMMY93b/vUHAA3wjY5vS
r2C1+u7nm2mcd0X2ElWPLA2l63d4ahh0VYgWHXjt12du4gx66B1ysZ6bS5Nt7QC2TPquzOBJ7RF2
Ct/HtlUkoMR3VcNMF30KTuvf4sTmie1M6VaNzMoDLGY6vNbU32RgOVPoLsCBnsQCrjfO6qFVYDN9
8GiAneA7pXZu6lV0UW6q46SWz00pgrucE9TRPCGb9OsZ6CQktpKyusXXF3GQcTaiAno8c+cXbfo+
Yf5t5xmhV+v+n6FEj/2bb/zykgMdj5EHHfA3bDDvinkbcw42DYBY5me/Zh2tPYRJSPAEbP8uW/7N
HI8933oWhKGvrqXx04XYYZXuYCFptVBF8TaQ7Le0AxZH/iOFPdpuk1nS42ZQYr706sA7fn6/FVCR
/SEg2AZsih+VV4IXOgUuFuvxrz+ktHM+vQSFCKzhACV3Ey5nNQOU18wFzxs5n/OT5nfP6fg1hNoq
m2NZq+X+s6m1roTTl6tI6AVEsnl1htg1OZlFYkJERHuVnA0yt5EKHNWLpQ+yCVo4jvMlepcM8PrV
nuH6XuABZGDk7SpXkl0n+oS36QnbhD6r7Xj+IwUczQYG0Hck1jtWGqN04f/RQ8knjGqnfxlLxpGL
xZ4FPNok2IGLo1xTHdahiIRKh6NZmiPF6AEzNsz/99G/5KqO1ps2UwHmlBShmv0QGNOwK//p0vjW
og6yYvFx7l+WVEXqEJyPmy5oHLJAAQW+oqj0Y+JBZM404twoDRQUDNZg8BXepBy6FcpTTH5cDlqi
H2sDhzO7v0hl0Kvy1G87HIspimGARvyFxPdsv1CwLYmdANkKOzPE/8H2ygLBm6OT/mznoYE0TAgV
RnSBDcyl6+4rPZOrFi4KyOBlu/h5rsvIGD6fPb4Q8Gbki7uHY1xdEcc81oFYLt5JtSTTnkhHjCsG
aZQZj/tad3ve00I+wm9Mq5DLRnUrwSkg2sfhXnKQvvlZwMm+EbWsWu3i7Lqiv1Pe5VqQD17SQdlh
FNXfCP6tqne8Yp6NaVwWFQ/VnIXOBhXCFUgofKAF1cM/uai6EBIdmWxXgwtt4cEMud8T4ntfGU5K
ReR9nI12vjy+6VH6MPgMVQ+OCxvDnx84dEnOzmyY+520hdZEfwDbn6D+giMYnS+wd+5uceZ4sGMx
Kl8RJ0VSSw0/Wq/y46t7KOEpfEAZNpfViZTnjVmqSE0wHuqxb5wnMQMiDnm/QkSuYY9aynWctzd8
VLntib1MqSsBqOz3aZut9jLZBWET1hz++7tLchQnIgFPKd0llHME7TbFjTIce6ds+B0YZ2UHIbzI
ibwu4TfLuxcUj663e34EuQ01EafWON+oxtE4x9I3abalA1h1Yo2M101uW45Q8eEpWr362GM/2DAG
o2ppqnVvK+uKG00EfUwZRP/1Oigjj+7hO9E962o73keFCz7h/gRh9RmNl2PN/ycq8DQ+/xO3X6gw
lRgLM2JZ1Q6sLX64nKkn6EwG42m/Plh3WT2ie9/PuV8Mtf+eysCIYJ6e7kpjG5kAfMZ8dIF3F5DC
RTY0gyzFgli6DKkCShc0YcGRuVcEKUgpDI1OpYoR7fJH/JHRVjImuoy5/fpbAXZZMBoI+5jqr0QF
wZkVnevlklvEPeO2QI5KVrrs/cJmD7Z6mAjQJW2cUoYK2v0E6nurbldnGhI8DxBjrK7HI2pfboF0
zSXevYmqTjyOg5oESc/hPaFIZ6YATItPr+Xb9eSz3E4kBJO5nx7oGix3v8Hfds/H1aCbDfBobInG
qlJfn/hL3sYceGG/AjJKEegDMzddcQyGWo9iicZ6EwxpXmuhDVARCeirG2bjn0fDurVx1eIv1V/N
PjsCplD/XT6CTud4oi01N67mTHssI7sIcBWEioOMsFgNaD4SNUns8EfH7eGgQSufaglLkWO56aWH
+nLFH8rjSq3bN3GC3YTcKtV4Qs+oHeFO6Yn5CTXZXffBeMpbpUU1X43WE39R39FbeE93BOoIxwtx
DSmACojpTRfYpoxmCAw9UURDOsEYqnI9EiD5s+nqo5x0eNh2N5SDzy57PjM1E0KupBehfELAd2Mi
sIZtrxPmRCrvyP9o7+Oi56QD2FoJcpYgsHPbQTVo9qEk5Gi8Pv8TEzmAaMfYPR0sox+4HXfWVfbQ
CXNcAYaM+0tPj1LssRzq9TmI8r4ZPwY323kH99wkm4TmeyaBbAalNgpfjM5G1hjis+6U7NOtPZ0u
m/rgQ3rX1UflTUrbWZs/3jrKsZDRBK4oqThwY8px5+w6R3sizAnR3FKkyVpX1rtSSJWXhnJAygHO
5bTdHyVSa/5BP2kI3nmtOMSvSGTCGub5y0XEwnPNLg/UgsR8q4clBzogAFMnzs9nDt3bkXU1A4G0
4wdovCBlJXjqFpd51UQBweU5qu9zBYiEVCvsyJWYvwZkf6BuGxaCtzANv4rQqotyC5eScKS/XcOw
g0CgYK72gHpB4zeUlSIpp1CVJegV60I3J2ADlxP5TzHcgd0zoG1J8qKEfYhrbggCc9WpK24U+47P
XegRcuOOpbFWRCuS0QVQFHbGSSyz67umvy1+8iPYW8wG+6frKUO9nfvK8wNvYigze4eUGXOkLT7B
5q19EXHkOdmw0goPF8ZGLosXyS725+5iz731rpjIchdmprXjEPPFz+YRdkC6AUyBDamk6rP7U617
F6PRgQBapFPOtFJP48WiZSQCWroq6VTpAT05FYb48coarxL3rGQtlclUT/fBvoEqSmXnRIwN7P2M
KAQhm2KnQMvY6DWacWRZSUibivtal9m6/d/G7DmzS7nQo5I1VCFyD5XeRlHVie7DsbQuFV5cu+r/
rEu141UMd7HrU/94xlzKgRnjRekfVnnLUxsd5+ZOBDNxgF1/rZrPoabiLOkZd+3EWBGbsmN4rupi
HSMEQIEvOInrhu8c0F3q+FA4wEGtHOwG1ljtXtMJPOcD0s70UzbjwIZwJe3lRZTE600FQTVZ6K4T
48lvnm3+RK3za+LpC17k5fEZlZWPqUz9WCd7V71XBp9ohbWEAnQQ3khH4IqpugYmDynVBbUihIlQ
0fARzTEUT6omekANunvTkpsu1ENmMRVVJfA81fAfDvX5v3fJO5WUuAuqYWTm5138IamUv1nKA8uL
CB164NfKtKiA8sldyH7h9x58/YlXxIK4FNOuhVZIVVa0J1McDspzVFH3LvfsLVMbMCKANH/GL27j
YHijmCNOJ5mX5NEnajwbsxDS1sbNl03mcStG0DS8ACXwtAjlKz7xYmXN/JDGjmjG6Sc3jvh1dVpk
1KTFLrzh6MC8c52ANGPbBOZ8XcUCjJrsAhPVqT1BmjzLW71vLt55shF89Smc+QwYX0A12W3HeVTn
ZzNt20EOLPLOiT2LEQxHH5APelJUqpzcElwWzVXp1Ghl/r6f8QniyCMx7bTLYy858Y0Wdh4zMONl
TmV1wVjvBTDMqjc545c5YzrxJZL3UXm4tFhJVan46L/AlCtg98UCnY32pxh2A/PNgbJ4y6VJQAmk
n5xc1cU9dn9L/3zy4mcofXu6yarpkjxFwdjlKnYQ1Eg4QVqLgCR4exMvl1R+01Z0VTRcKhToFx+o
DuTr9fMzcpho1Ma4rE750iAz4IUwH+K2UfL6lUPf8kkZ4wGB9KinRpUP1FBJhmvd9+IkXTNMCCi3
iqqbAGn1/mX9oNx2Dq20Rh0lUqKr0eguXSnGfpUVa+Euj9vvUGG+jaXyAuqH4S9lI3DveZxnMcmo
pE9c8y9Si1tIuK5g2gGzP6PhNwUGU+t6EUbEg0igcJSd5JfzBc9p9pq4Y1yCAOMfI0/AP6zLjCir
xzlybw45rspmvC2kEkjB6N5FKNhoWEdtietQCZDweJGaqm0OTBz+C4rov2tPdJQ51EG72u7aY0GB
tmPHipx+yFybtZgWUGmlif7abx7834z5smL3bjNSyaBAQqqSD5qlUzXIFS6vr3RQD64xP/IhK/kQ
448pCHW7SQTScqrl/mrWlFxIjPUx3wogqWDGw8B2AagrIhcF4wWsnA+zmBCjqGT7t2+VrPdymQOr
zuQKgEbmX6pgf1WLOuCO7qeaSngqy/GfAJ0X4GMSx46GsH8sDCmvE7yxVAjNAwN0kc1C8mRjvuh1
YgvMgX4U3abJsNc9tSLRbecc+Fxnz8mUwjTcW+yVXVv2xEyhH3b4++E0iQAmnRBejHGQ6ehr/wqq
/MDXOFzZYoUM03bXsWeLmyBuKx9YiwCiknblpyNgHHmiuK2SmJfCHJ9ezXzGeEO6U+DR3APhB34i
lEyQrLbNTxmUU2wzNTgqu/TQwRrBDf4uQ7M8vIEsuMr3jlAXyfJasWJuLs11sG9Ehd8E9FcOesJK
1En6NnJOpra3AjcOOJBJzscSPvOEY8umwuMEXUpU50DJ1XB4BidV7EdvSUJnOR0EyQ+mqcQGISc5
VPG3bzUIT5AhZ2Ap34hsOLkOk8+pqSmI64nha3AKUdJPiOnjWCuxEz6YZWyme+taCDZDN4jx+iJQ
fkRRHSELGVILtnTZZ1oKRfNVJAyhnSc1my6fyeufEFdweagZO4vsy73ZVZeAsz5CoHsHl65hYB11
fo+JIvXD/eORS4RqjWpexCU4sr/pf8TbdwEBKkW96WTIVYI7cVt7UkgigyZaMb7+8QoLjbaNv0fb
pg08GMW2QHMjmfO+dytiQOe5wZfPSdwl0uoepMjS5i+pDEPaZxz73G8i4qryso2pLZkjTZdnZx4/
eSu92pGZb106AJe1pJhMUbVD7Z+fuDuv2AcKbUlUuqid6kB5MaFCE4hP0mOB37lGqUrehzlSBhex
kibLid6zi8SIPEvKBSwJwqA25IcRt2HP4yEbPyQFRbGeOhCaSARJqNAJ9/MpA/75uXhjo4ZNMzKg
TDMcS41J8TdZBHl2Y3DicwI/6erUlfLO2VxxIKJ9NTQ+b6r3LsC80shXzJ9C23c997uWyEJHsNQA
op6S115UyjaWzEvL7Cqj1mK8b24ZY02SyyQEwyLR5E2LjtGKS4pi2ezqPmnQPPCgVcZu6+8aOWn8
ANrHfdpRfZTDfncWdiA/Ij5HFTcR6TVoPM33GakoCaw7VnnnhmNGPKogtGkCrVShboIgn676+2Fv
QvtRYY1yAhR5Ot8GUlKjoNTsIXcCobnH+y7wd1P7lHzza2/TieTfcPp7Snn7aVNjXGyoSeaHFljW
X+7JdHlJrXAi7dhoien/8wOdoRyiS4oZKW+IEk1+0DnsT1kP38U5Gh5e91u42dOeU2E2XZHznrbF
X4WB9NUHf8gqiXPrw6EqoSZznTegbgUSTOovzzs2RngxkBkRTLKTWFoEYxAuySpeZEF3nv9r74x7
a+cPoH21lkcU5DtMtLaX2TUXtnPAddYQlUEClK+JWWYXiemwYtaSh5YDOw0O8cDiFYum6JDAspbf
khXgwbMzvtQjMLBfpES89zdWJ0r5A5VZEWUXmUA/YCLVJjzkZbFrIUnHIHtbb04VpCnxAEQJ1BIW
CkAIINUIQStoUi4Ah7Olqaa4sV4qlxH1bYdk7Sig9PacOCZYMFWj14Ot5dBlVTlz2PX9WT/jg/7w
XrlILdkcc8qdr5Mxw2XkXHnDlkzpY6X4f8lnjWJe+pXXyWwlS/C28czGIj9KzowYrqkZ9FJhK+eM
/HUT05t0FPFOdjJXhxsKgnYp3551HFcX7thmrN6jc3uzv/iWqVHeTa62flqoTWf49Jd6LGukN13S
jE0lN8EfzDJjqCNEzI4GBaKCSvD+txzRRyb2UzfSgChDtB5S+ef+AtdjK1rDuJQzlOYGNMu+OvNw
F1HB0cWmwZfT6dNqj8mAiUOvBmS1w1aSpBznXfLNUZaUWD/n+hTJe4d1K4yOYmHv24Pmv4L+cMc4
J3IikO4f1garAru3K89hY2P9NxtkIhnsMRhLIYg6B3b5Jd5y2hwfxgquWunSFfWAUTyBJ5ea3weA
Xsr8tpci+jHSvCUrfsEL+BJKThqDSVKjDoHV+gTInmDZ3kgg/6g6tYwKKXML73zi0rNW9cj8XhR+
2r5iqRElAnU0zfTDDhWzJqgvONnmmZSNQmv4It4tGjHjM0bOAbO+t5VUEOAxjmb4WKpSH2hth9DL
O4SUQbnrV5y5CUu9wF9bkNAQ6YRkyF/392A29lNa5NR3sEpeG5NqImOt5JTWbsro7Kj9yuOuqeWu
1eNDqvK26B9QI2vgqx4SFdDj0lyeblIRvM9965wVFbqDP0T45HDhchC3XYGWHKfoN7X9xd7IAcal
9w17qNA+u5PkMphBpTOAWOZvIA2wkgrSb6TEKGb4tBk9dt7i5l2k3mPdVEcHdBq0NCsPgYc37ITY
uXmNb551Cyo1Nm43hpHTfph5X3y2HrD68FV4BONnNRBVS3Vv3dOJO2qNPLFjyMpRhpEvS8vwY0dI
A/r6xYlEMw0iFg8wVBqLpPP959WuwULaAhgTEfdJeoLKxyB4jyCYD3UgN8pagS/gA9ysYRjHv1iw
LlUaA/VbetpZN+esLRlahB61cmCqIrhHLFD4EN40R5zkjNT9q2whJ2rxfEeX5U+asP/eZuBQ8iUT
G5GMQTc6YwMRwSQvmlp0OLwl9hppYcz1CDipOzoaGDOOb3xHKbF+/cHrQt/zM895G7RtqGkKrKc+
hLP94fGaZ6grp2Sot2OWZnE+dn3DNyrfEBXu0tougdEamL1R77Y2YkUAHz5wSpP8tQeFE1dKMCse
aSiJxhdOMsOqQ+YifZsXmP7CJQ86buEsKDvkACZumXMccbfS0tESaAFASCNhFd2bLD05DYRffycQ
89fqTlsQP/vVkDmybhxKrK+bHFrukNa+XGrCqEIQTh+RTRnDZ0yntMg5MRX8+e6T75iI/krrt2ec
kz/rZs91GZSQ5GOCzAtGCdZI40B+lpMG3hN4rklvIIBgOdSDY42lDquwYtdgxC8cTeag0jlHkfOW
VyZ0qobqtgBh48et1rLnNg+2wEQe3GjfAKALOQkxmjqASMBGpBQqUUrWxmcvvXqXGioK3C84i9jb
WZAkH4CJWDsuuiAaE8sSCZs8hFnI65KRUK2Puq4cZWI12hllBMvj4BD2dWx4Z4qqS8sC7uxjy0FB
JT6hPq/hJlkveZ3Cmk7arxbA5mW32TDOmn3KBd5h3tLaIww6LQdqoG4vOAsPu9tmqiOHrZsf1aGI
8HXtARFtxne22b3RB8YhOZhQ2wb6JjSgPL/nFRnFfog/yirzXKloJGwezROjxzooFUDZ9waRjGbc
UlpROFtYNkyDykbsP1eZSoXkrlWgZJXlN8V1GJxZ1R3B2vf+A8iEURgbmyvbuQnR1hAkS6vK2Ip0
vz/wYQ3X89X7slKNx5cjC0WG2s8+8JlkQ51QzU2BpBWiqQAKheBWvEjjLuH/EcgqhCkcZslL00eQ
vgTSuISW8w9r4F6g9gZU06R+dMQUnomgBvO/5UiBI2kVrJUYxNXQ+A03in9yIelnxROoKehHk98P
q1ogFofVjKI88Vm4YifUJ0IvzJsbzusgvDKzohTRk28LMuZXp04KPnf4Y6ibS7eBU8lwmYlTzXYa
+pSF+Ib9vzH6IkJ2VtPrnIqomdJQe/MEab03wujM2/Llh094KsDuXadz4LTmWYU1Xq+GIdv4Pq/U
9yognHkOn9XLPRzpaoPLIC4ypzWpxgYKZ4N86w7VYrsEzb19pe7RLdc60iSdRYPxfWi5+MuMq1zn
Qo6us3q2lY7lgCpnpGgjTYB72OuFPXortlp3CMzxL0eMaBA8cUhs84UAJh1aXpKz5rFcX/WfEd4Y
po9l687HSaPNxNHicFvQVvg21aVPtSUOfZ/6I8sDiAGTnHSo6NokrO5hglzU2qd8aVpBATTjGDLS
eghxk7PHiweA5J0vDY1h9pHAB/sYbweM82q1/sznzThIJD0r3abjeajWpc7S11FbSXEZDbfTiZY1
MmCcylBuGxl2+TiqQtdznOcCKzlF2uW3j4p/OtEQDH13YkrGEzSkyCRycOHMljtp0/N47WByQSVG
v2cyYsTF/TnbwKW7pGrz8yPw9Ysox87IhirjGjJZsOpTcjBbEu/bRQdxhvNhQ269QTZZbdCRF2gB
N7DjpWma1o8cseLbyhPdu8cvySSplIPNKAgrkZCgFq+wYOX5nJWtqGjWtbz7k1tKzNGigWLUVWnE
Z7hLwMBluYTWKVvhQ3xNfKt4+K+noFwTHNyhQqWytX1lHF/43TMEvUriIuVOmLUcAZj8tf5LQcdU
NoyrUmUxmGWMu4d6RFqgbtstBOqB0dJY5u9yozPit+PAVthLXlsiHZ9Y00VjdWxL4KHOpFDlTAOR
9uttWH7XYM680Kbyx8PKAzyUx4JuMEgSS643yS4S8za5ZczSuIe0PvhUkj9X3FqQvF7jksMnKNMe
a9fY6vGOEbkR09G2uvwhAznRWCuWKEMHSDVqXlVqoFMQB1H81sZlFlky2vVi/4JA0gTDyZdkILmU
dtTFriMX1Fqxac95n1jTdQznvc90PAXAVZjK9i+OQU4vyfWpo1AzuKfmZllPU5IS+xkEv3l4gGKt
+JRQmxoWfLwW8Mwt7XRHWfoAwqcKpDQstTuvkUnGLvl/0/JendYpukKF/QUglufv03kelsf/LmCl
A0g0QCHRQRmplDbcwbMqqHPUplS/zNpfk1DL3r+7gP67OJgnuR9hrTvADmmbKS9U3azzd+8Kq3nu
E8DjLOMyOIUDMReBguXalcPyd7fszrAW0nV1WFlQ1FzLkP/bjeNlDt+qoyJGjeu9/UiJIUHipLUg
AMmbLTd2HLQ+u1K/tBJ5PcgPqlhwI7p565o9AsZLMjXqcHLb70hJvOLVZ/kISkntl+eSvyZMKjAZ
VEww/eWXLQWXkpgfQIPxJgIwAcQzaSZtnx8lB1C4h17dimHseYtKAt4Hwg9mGUSnV5im+ji9dVGa
pc91SP0DQYfOvJZ9yK//wpaax8k578S6mcdEwxqPqY10O1lzKRMrJMiZXDYWmyGsw2bntobM1INn
vIu8X34ozPbo6ozdbfX266PSXmovmGaAYPO1A0hiRFCBSPYIdbPj1nWTzHCLNVNGuXowXwVhyCfd
ZKU33u84Hpfo5jCzBAN7buHlmhGywhMauc3yHozPbeRdTfHZOfvNCLl3QRDVgtAki4UrBPKPRF4+
zwTRZoZJi0KxLNeu+owQZc1lysX/o7FOQ0BNDXFHZHCCdfaINoAAI66esd+REjTbOWf2i14DFrIB
zeJdev74NnLXDvZ+EDlhxoFqs0FOjZm0pnwuCknrQlGjU9l5e+VNwPtyEbfzJslBiVnl4WMTL0aI
umKwm6DXMVHTlFB6MGsLpQmAZigUA2EyYut+tX9vnbV9ElhKW+lY5DwuKW/3Ujh4BriafwvpQkUS
lRfdV1+KQt5PhByQPhN/R1KLPR6XwqMxHtnNqrSG3B8DduHsKUlepN1JzAA1gnG4gU+xYXmehF9F
G+KzVrzGJy9OzgVOF1aLsV3n/3YLC6z66xiY/ALEc3LdyAfZn5j8b4U7QT1OZzFeWut6ciV2UYT2
4/XQ985jHtSfP2AruPp4DKbEBshT2HRx0p7vQmtjYl1rrAt8Xv5hmfBBuXF+QzBRuHbeNv4E/e1h
zpifXjU9xPvbZuozPl0a298/fBofgRdOiQnXgyTkx1KNW41U58T31gH4LL6dISg4PWZQgwlUC4F1
1DsL41KA0xI1jCde02zIQeWmLtFcIfrhybTP1RvqeptIqJalaMTW30iRP0BsJ2l90R2DDi1mIZzE
xAYkRoXvaGrdPVRyZ5Y+Sp7gC3HLiJTnFi/v08l/+60fm1uSt3P2o1PcHt5EZQc2DgtB7Z78Muhr
9RIaERLsr3Dskuu3TMJ2XHs//n08JzlX022JJbRsotv6qJTH1yFH13tDx0Nv+xvZ7VBA/imifKdG
wzWXr3364ABPnZfMYDj6MeWTi1wE7sJ6sSzc8aTZIm6W+O+3mGXaymXuRdZgcB8xP0JhzG6/znBj
IFc0s6O98bdHZutD7v4DN5437xzbUYnVe/BeX49b4ObZG5cpXDnr1tKiOD8k1DNvTSO6GjWCFcCQ
LlNj7rdWtukKjlNEBdrZPnEUJOGdi/v/KlOIp77SN3rEAujLOi9o88+8di80fNBDi/rhtN+pHaSI
3FVhccrrjnEFN3R4dlMdexAPMxbXlJ6g7G8hPMBXzVsi63ET5wPLCtrWD8bL2Z5U2Cj5Xj2IDM7+
DFgRkjZ5ZT3kMLHVE0g8O0NthvjoE4MMXYbLmg/eqkxzalxAeg4uOBuZtKbwn89QWXAJskd1SlFL
Z8Ajutai+x75vWeK43gTRTyfgDKp6zRRakwHPVv/DYa5F9ojRr8ARexmJroEbcPFh+tOV+GHlVEq
Dqe2h1JNNZir5apBYLGXqM9++QHxT0oqBFhIAZh5xZaerv5hiplRkXgt3eFgiTqa/AhcygHGQJBU
mtF+HUIQ+lYl4UFX4KVKnAAyHgbjlcwj7sjSXlLEKPBK37DEDFShVDi2hJ9qKpmbC7tMXmt+MTJ1
01Ou/AkehMNH5XfTYhYKlPQpIVLlAlJrxNWo54HuejfUuJYH3XyWjg7mANvGYaVEjFlpw13OA5j4
IDVVqKThx2XpjglgCa6e6G0mw04w+77+7C+3k7o4nM2/VrWB0jlTy2pWiHQj9WJbWyiIoYzlyXS5
vlsXJa1bxPqjwlV2OMEaUEP00/tFNG8n1MjMTMHwjgtn2xmwoeXBjB2en5DTTSwrLaXT3r+88cLc
1dAyFYpfABDVQOZmnB+pGqdYLK1jLCeIuYE0N/9Dg4ciWB26DNg427tElwLXCl+9GdizUvw99d8a
E9pxORiyV1OjOlF1vXgyMI97fGlmgcsm+Au4RLcrQzchu9gg0+l6RKfYtLDzItuw0J8CiHgAOpdU
B82MmgQa01IQlZattu6vpyKg5MdZJuDBQ27wVrOGVZye8wO0F5JuRFNsyJn11eOuecUPkxneJg2n
FFDGdpwEEK+B1r7tJ/0GNpBrLoam1SQ6Pb8oMfMMxWCdSwnzV9gqcI5tnPYMBdT/3NmUzAbWt7tk
f/9kGBsjtT8XOA2BWevzmdYA7URPIU4vY1AZ3xA8nz4GCWm2vVUpdJIRMNFRtRej9baXhM/N+xZg
J82M+pSzdL94iIAQdzDrlzRuclsN21QmCgQUq/C/dr8lY9BYoyFHiBfQYuI/E28fbEM3BknDAQDD
c7vZLnwhvtSSOd1Sb2PJUHqYblnlHgyxSQdUg2OjlJ0yHfDI+rBl7W4jYF1I4J5dXa5siCsalRwN
eEVA0B3fwpJxibnVJxzhlgUQFvJE227zdVNesoGZxxsgBYEIr2B6Ru0NMdDu98ATkxjf1ZKNhy0G
pBWRFKRULf1UNj8y3La0QArXFbg61jEZBppxKFs3KRa/zDrVDzqOEK0WxNDAadW74GeX3KYAe8BP
`protect end_protected
