P42407@HAGNB260.13796:1641828461