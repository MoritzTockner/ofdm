// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std.1
// ALTERA_TIMESTAMP:Thu Nov 12 15:05:50 PST 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FQYHlDGemvpJcQ9eiBcvQUnXpnSvXHSIfqKk+1Q5hwFvKcw4H9KsVikeEOLmJtBe
L4LcsfYJvP2NZPWk9MiKwJgz/knpOZwWqSaTsypV31mAJkzdx2Qn16ynaBChb1S4
viwOe3g8Tb01hybi4kyev+tmgUQX+GmA0Ri/j1xIC98=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11200)
r5Rcw8apQFv9ATmWpFQd61285T5f+dqX6ytzyoFOm8YX747Wb84FTjAKD4oGvERs
++ez2DZBUP6thnpLK1quEBSYFPZDuJ2dG5mQSS90qAf0ACrW5ASlxgZUIFenqmyg
r4a78ndHuD6HbWSiN8TX9MDM1jLtF86e+kviA1fLV97INZ6CKiR21ACeXgOKqfDt
0J5Ubov9yK+1knPKhWgW/uf/qS7XpP4fbtWpLzEybDbcNdkJDZ37rhigDwx3USgr
t+mLd3+HyKikhq96XhMiwC6THsq8CDf8ylpnTaOIlvRtrnW7bu+2PXViB+IU6jIm
48Bbun8OVG9NM9hNreHRfsi3zbrwijFp32Be2Ne4TRaEVPfEX/LUOk/a//82bx9e
0Qy/FCsduOvfanOH0XZ6FnbhHHZBKlNwTnp1MXams/1KCplxMq1zB6civlnZ+OqY
cLxAdcRydujeVRICXnpcFFPZQn7vXCM27wc0i3kSYcC0po5tpd3ww8T1iUAekESG
T49vu4RUgGaW6KKVTGP83anE7k7Ph1dye7QYwEVQUFnGPYqks4oGkSGw7sqZoQFE
ggxs7LiHv+4wVuJv5vxCrYI1JePHl3EXbPSkvplyLAkxe9rX+dGL+Qq8ZNK4L516
bttmJmgtCnycKJIaryyMJ/d+HLO1mpKjEhG9h1VWG1ZiuDOgUpjLTHDg1ItzcnW1
QPn2MQCFLhYcTElk57ps4ytGozmJ3L1G6BJSK5e92enjb9oGhBeZSHx7c+y8FCse
eCuJH7G2Bi8dag5j5t9gTvo7cGl5/zbKXu+63op6P+BEpk7NMdwuziFCppy5z935
ZgbXk1LA07m1q4IL2vvwMtv+/VCIfPx8lEs12l2e/RD0bkHTmTCPraGuhlt0smKV
XbjK59Bwkwss72G74NSwjRIrQsyL6zKX/MLSz40Su6gvonlmQaInBV5yxi3oRk9y
Mp1KrRPwf1IuQA+V/vE3w0Bojj8syqdmHH82Y8qkQH1HKxlev/tNbh7D26vzSshi
/H7mYlsl9NycxRZpHQU7aI31HQ7yaLpgRxgRjRzd2SdYq01rnRuK1Is/2JB9BmXA
8E9dvihFaaz5hF+Gw34ZDQqMvsX4tWqaJM8ElW4njzLkngIzoKrQ/5MiStw1nsvR
I2MUY44MlzhWDnbeaMh0kJG2SI4S3vZM+q0cDE+pDu5d92NKa8RqKXbCIUhUaTKL
kuVwLNAQ9ccTMVoL+zaSO6C2h90dHjXNLKqzXJbjq+cLslHflNbOd7+bvA94tTx+
dFKT5/oN3jypFdEY2Mp9ru+RFefv7TSs3IlEQHRiYQRpKq9h+zCX5wVqwdTiq3Ex
Tu9nWQju/yWh7zvVOZRbfx5U8mjQhUwtwXu0pRLinDCM9+4J8iNqGRzJ5AzPc+CN
1aJvmV35NFgQVowtJAx/pNiXwwX2miHv4Fz1W/lSxPHVxuHERhzAAmWqZLuGrjqV
S/vixFhO6BHJ3zmx99dCVnxPMJgRleqwv8ADLoXyRwq/UqKKtlrhSxmyjr9catgj
3eph5wTVdhJIiejR/NMT2Bj8whbLF7HAHKLyfvmyNRy/1DastiR5ACvYqEy46qsx
7VXuYy61eiFhB/MWDfK1cNFi31M51iiiVLMhpOgVkcdPJYKQL2/Epn/P2lE3szJ3
G/99NU2Q5+a9vsoPErlH/zbcz3nYquJAJtaVTDgCqqfp6cm9jh1cJSrCldHi9WdY
LcEV3enAO3swGKx+k08lCA980E0hb/uRll/NWRZX2Qf4D1So4KBCcx/dd1KE2Y4g
D0moK03luGAxuPLC5pTfo6aom1ZETBIknkqDfPw+XhnVZS7ebsFg7rjJYW7fVbvL
g17FjwOIOhSXspz8916IjYaHz9g0J2tVedt9KWh+zbdD5J04q1GsXkyU5XW+rq1h
89zn3bJBwxi2v7NEQ4k2sxpmpZs/WNIJSNkHUO32IN2b/fhhP/IngsNTOKzQP7Gf
nziQ7LvBn2JIe9W7NTBOR4RkOkxz50NZJYmGzFsV7fdYi9xiL6UBb5vtVQOhXjO8
UzLApQZTqYm86Y/M0wFEYB3MSpzz4+Gh38Oh38p8UNy+AY4qUH+0oTJ8RD9Q5Mvw
XO0tRe1BGYlV7CS2dW4JNDUXKGLRfHxzLuaG+wDawNiNBcj6Pfd0j7gplySfbQjd
o92ImI4eBarV3e/FNOae3kf2ccY9B9oSYaQQ8JnM8LfLJ14AZgmKTmOs93xqNLWA
6RK7ZkfhbfwaMT6IOJwPCbddBd/Af6ky+hmyH0NDEni7bR92csoDgVybUJubw6UX
OTTNMqwOfCUjq9x2Aorxy4/Bzf/b0H61PfSl3yEXa4IPSCbKjRrTinUw/AezhsVQ
YmXBXDhfHZp99b4asWAqa1j/R+SqPGI4ELK+8zYECGrU72SLoW6JzBkepldvlKWn
SHXE1yInDCPspJ15bcvB7P7qyQEAPDHUp5zvR3FjBefHjP3Mcueg/rmz4aH3mp8L
0emBBgAQ8SsB7pwli2fNIh89zdUxNAc0K75vSgpQe5pxNASapyF+T/ug92Bb8nxl
M32lnXl/jfWER14o8sNApZoLJkGj+pAvhO5GJ5YcOTmbcC2NjIZJS6daYuKTWQnE
voRr0qXL+BvgAjE3gsK2sZao/XY5uKowE+uXxgzrupItOgxA27CTg+kabLoDRt7t
yRsiSH2cZcAVPXIwHrIk8NtNYjB3uhyG2pSUpnvL6Lqi19qDHP8HnocUGCkM+W2R
8DJK9QmPz8uoBVF6Lz3w6bYNOAjeB6AYli6XtvfjRyvUTizxF0KqRRnfnPdQia3Y
fNR56cpPZAELvZZUArALoUBiCZX23YlXeVr0GwJoO1kHE/1tgAwDW0ZIIxJ7jer5
V/NsQkE1PcJ6XPCXsXqbqymw+BFA//0IQt8XYVX5W6ky1vk8GhlE8NlRfWN/m7Rp
1FkmNfd9S2drBdb9EcCKU8tDfaRywg3Ju+sU1Pc6Ov84bpjcTU9XRUxTkEQk4SW0
r/oJq5r4SvFHiyUy7muzim5zy//5D+gqT7E/merdWuk/W51a6eEiGO9xfXJp/z0K
lA1WODGhpz05RJ/bsfyfYVe4wI4oSU0waWSqO3+jO7224rIL2vU0t/gPXukeFBZG
K5EGBKfsvjkWEdNMWNM+aTBun5Y9vt/u9QFZHM8Th49ZXTD1VtG3vDms0OEPlU6v
5uk8ipKUBWx3pE7fBkNFSwKNSeYJdTzZBMtnwqnbxa/yroZhmeAENTi/Z6lF0rJV
x+85+4w/scvXetWQQDy9wjzon9zLHi6aefMaWK37oEVqIaqTcBhjS0dzKxPUtZlb
ZER695nPo+Mv+bvgv/EENito86OQDzevEOc16qGf4gHf09peWINrRJWZPdHcUmwp
bb4EjxyS8MHe+R5SwIXmF+zN1+sqaDomBa55ga0wKEbLBL8XEqjthYEJm/NKdSvx
Fa1uZPGdjw4MQEll0JS14EfoeUpgco08HbyHgZQOiBge1jvUbODQlBFlnxFNznXF
BM+XK7MKOlkmuwRIcaU/SVn3ts8xkHR06ZKqqLPSRj1dz48/nmPsQdDExDoawaMS
IMQZu5GtHxmQmVqNDWZcaKGTEoPJHyRUWGXj8uzvw1zTSrgYXyomIgYt8AbzcvbV
5Zy6JvIVcDbVmxcc7u/lfGIVkgfpCLSo9VtPtfDVmEFWbla96igEf3SovAU32AKC
u3zBAvJRwC7GVO28AZLMTbsOj4PG6XHfDZQc/+YwL6rPgqTqnU4/uDPlPjaN9RXL
ShkC0uczC1lpCNgY948UfyNDeEd65i6400jncmT5Sn3tEgoxgRg6U0ZlNuE0FXJf
ueKhM2hH/VbS97nfEebJ05edw22cDKBMklopqIhEzvn8XC6QUtj6nygVNoDHkvRM
MaBQ1///2bIseGTPrbpx+wdi9FZ83D9So6cHsDscL8MynpgmsheKEYqcJjqI28Vs
r3z6kATCijDfypCJ0xhXL6XuHQ18FMIg0z1hMdMnWKMy0xH2nTBdNJg5L7+mtaiD
hs/Kw3Uw2Qn7yn5rudbNsbPl4AngCeg0wcmFDkauu8qRNsKUHLWYMnWt8sUsmFYL
6L5X2FXulcC9z1FWL0dPwk98poC7mr0CbUdgL+H92luPLhSSrOm57p5J7JdrPo/S
jmxwyHAmWUNMJN4SEY+MDoIFnB5evMrF5eJgJ6KUeGny4Q6NtYUMuVH1eGYN88KG
e8pGXpI/0v8xmFpTUh4YCQg0yfjX0nWnlECYm6HkUvSlPKyHafyuzhA9HvCYLfzs
jkOVlfmPBvWz9YG4XRPq1kztA5ZuTZ3TdB3GgWjDgIkRI6wN2xsZVi7I0lAqKs8l
M8TrefPHqXzQmjKsg88dAVdyq2d004vzjDDYF0iJTKNo+lVqX/0ZknYf0h/nq9GG
8arSRC2zZ0Wzu0Shnr8Bewk30yYhDKYz8uPU8YjqTt8PrbLuxa7gEzW/bHnji9bm
YiFMXOdgynTl5HUFyHMNu6LwtMWxI6kYf/DTuFUI6imUcW7TGpQ9mMiLuAj1yPvK
LCKtW7dIry21lOk/If7x2Rt2t23kKvdwI3JXiAvSRc13XxMg2tADZ/LvJi4uEyTf
P+R7k5J7f2MF53/9+hS0jOoSD3zBrbVZ8q2/BNd9prj90d9KPC2/oKy80OnA9G4B
6O9pqemfNI1W1rscLPg/W5A/o1SpmUmOHQAhHnyLIfPk6+eInCN+fz6inS26ItHK
sfh28Vt5iwycR6oDBIp89Kxq9NQEehXyWYzyFQLfX9qUwifvbH8xfEz23ziOLmZK
NcvmAihfG9BEYqxjKViwyZVu5McgqK7Ot4g1+i8EJc0GLWOdyI7VCd+eSt+YAZ41
83OI51a3LJGtZhzcKd4+XX32gg90zTeR2TryvyoG3vIKf8R7z25DVQhgUUPqxB/9
O4rsVpV1Xp0DytNq7F8oLQd+xCydkBsvmxtUQrHFlMuKSsnMF1Wjc4LKfqa7ZlTg
1oxOoCYhRq+Bu7lmuppCP9+V3PG46Mfe7rjGgkc80Dq0ICyd1eoFxEtfvoDaL7b9
KjagwDFP2ybA7vSYPtjpmkrnGOp2pjHvy98NY1C6Ez8cnyhCArgsPzAeJ8D6JvV2
8SmVcH7p4P1zyMux7DQLAHksGddcASZA5oFt9qSUFnsv17omJzF8DztVLmmzjOb+
rdrBuUUVQb6wkyj8Q4shHll/smD1Ttbx1+NTwuP1CfQynqX4aHe6b8l4htazd4aG
Kr71kuAUZR4MCEJf5f+CfMzzwcuziyaGbPkoeGE6rsmG4jKRH9O3C/D+b8GpktC0
RIZFqcHtskl8Y8KVngDRT102iZqnWrC/z3zkFnl2ThiCdTfUgG9KKeXcQ/mCgWxV
sxBPoUrJGgm9/Qj2JLBn9ekZcz942oQ2xb8F2kask5sqzltAPn/f+wuJ8Z+eQmjG
zX8922xS1Y/Mm9WC/QPmKBS/TB2ZtiX5UoSXABWF3HpOAuJpZlx0GO2Ty56uuCST
dJLio3xrNz9S8O1vKXI8c5pF8uwBAB3eF2Tp1udYWmDkf+xJljDQ3ch5Dd9FzsIl
qWHiTnZmb75AqM64U3elAZJowKIqmOU1UPWRLgsoyUXIWfq3GL5fAJ90E2Hxpgw3
OMaEdkYeA+IdY9FYcMpvdmXsMclY6DvQxWW29jYxUErjAhnQiM0IFnfhRyKApyoa
LgngqwPXJIgKONftiMkcvUbcWQU2LgWjeL+s5onhrayS4rDn4ob5SDWBjRBYll6/
irbrtT72wPh+CnIYy6Mf2J2QC66ERKR0GIWMpmq5qG98iWOYKwKE8Ocs9pAfubYt
6QtdtFjC5fqIGKJazWA486fRyFOnh46pU+83zBduxfp9iZAUOVCxr/pZHithCLmM
ccqy4RhOe1PzDKZGekA5f26jySVt+LmWxePl6QQjKIbg+JnDSLD76awjH2R37E8C
KLQK1LshwgGLZA5RK64SAV69IOQFRTL/7T0wsmNwii8IlM5wliJaMjaVwM5s+xqd
gcA+BlVv/q7nKvDaDF+qEXJPBPUJ133l0q98+X68EIYzXrOzl7VDIe5/jLrXR3KG
C3a26DIfnN5SEuRijedXqaLNtGVdjoZba5lpppkvThnszpRCehBLrEKwh2Dzbqr+
Sa4Irx1JIh0AKv/H+Mnhq5KDsitUi/LHZv50ulKkybBZ4vI936puyPTuQJzAJlpd
OArTzZwq4LU0UiDIizRdJ+Jz/IavW5fSZgraB/z+GHxpbzM9lc8UYyKYf1pQbWqk
H5/H7Y86RZIgdNg8Y5jdkZWKSsk0sTtLMLzM1+Ujxp891YOfvzElM3OJU0svb+Pj
gQozMYpsZmrL0qX86guVkRZPoXlDByFG5T+XGO6SFOhKwVdGv0VKn9jW2dQwLY8t
u9fSwvRhdskZmj7UJjJZzrvoRhT9K2R8TB0eeMzo0vFjAMO++MdKfnAkVvLFXmNr
baxVwsQD9SIhy0KVqqGB1YubnjMHzDQAzLYl6fzWVcH7YPC1u1VUaTTdk/RSE1vr
5OmVyaO9ZfmuVPCqMqbq5FYbEb7+gW2nFwOECFGQCmplzcX+8EZBkhdvW0bYNPXf
imQXv7SaZRKhX60fr1nT2uaokOtaQ/+MplVsQzbeGC8PzP91GxefjvXa/eQVPExm
GjEYo0HXU4r7MVGaUI50b9LAzT+A/OK/u0CXcdXZub2/5irYI0r9hLsCNsz2a9UO
7Zzkl2xtO1yV5+Sh3BF9VSXD2pSGNt73O5WEsY0RpaBpUxownShTmWb6agJrGtt8
tUW3GsoxZTMBXlp+Pa7t2ydAFcQDyzFsckzK3SLUjAJBwXFJ3Ckpz7jC73tmpigc
5HE5lMTX+BdOCbAtEnjRu4ZZPFV9yDfGVrUluvbcvQ41vAQSFbD3zZ3CX6DyuBp7
ZuTTci21vIpKnXtEHPhK+z/8pX50MguTsdm0/cP65raiaLedzCVHm2qFmDbXNR4H
lVQiVk3iSFEaR4axHxJ0smH/2O8fX88aAcmge+Psx1zgzV3iPqUn02OPDkmq9URg
MxNO729rTnRh5+onwlwPeMzXyyhlVizGttrqNoLApFySU+nIFC56wh7MoFfz26C8
va1x1fDar7NrprQnaS5Zly94VP0t/i2CWV6qwewvwYLtZcSuKWcmeNs05T5GCJbE
i/9zYID+MzCAa/CaUVyqdXRQpM0OD6+1vivZwCHznuxh6uMLKXh1m2gU6ihAMuLc
YkDZTl+rQ4z6I/v0FsCpkhA9G2WjOvKC2xrGlT0/sSGfUfvbOGDb2CVxAMyDJ9dZ
y6Wd9PKrRHuBJH/dvsVV+DTVVDqB9YRaQ7cR0pRVrpZ0+9qEe9nYDrsfXApGFmrU
kXb9JCw+4jdTjGtxQs5lbuem6aden7kBFcYXyHYaXCvxFiyqyzB1l/HD+3ZCL7zj
baBNCRiQPv97Rhd8bylDANNooateEuGNJ0SXO37cSz/Tjk9N54L6ZU1NuBfXzXTE
2sP8Uk+J4Fpj8jYE39O2X7XoD18n+vjIGgzSrKGEYltudQbPdkDY5MHRiwbD5PmW
BWQkMHzOaxWl3/0xhySG3DKjEo2Z+mL4ttf68qQZswtrEiafRTkELkhAlFjmnzVN
7SM+QUENFKhe+AyY88qMrVpRD16Ce072ZQ/42UASoOxf7+sgDGCWpOW4Ja+HA9hN
fv28Jul/BZMLDj5Ryox7FDKjIddKTicRRt9X9z8XbWca3w4MXrTCJPC+5Otf5ps4
jEPsuVSIhhsUKXilfrwcd3wep2mAUwAQwcn6BVTbYYIuUwv6oSojX/1xmGwEs4Li
O9kP9uWJVzf9FH1Q038pkHcA19zCAWjz49pIKXOBDmRLRkuEX4ttTege2YTIcGbx
IiigPSZh8i5up6ap3Sh44Ozxa8TgvZbfW/vLVgD2AGMuEzZjG2iOrIXV38OfsYJH
5szMVju9UyuVKo59FVefrG/9ERnRyyIabwpDZtLBW7ylexJDWq5ZVh44W0ggmvwu
AuPn5XxRkHTM/MGO8wfJAiaV4Khkgpk1Sy17qsAVTZZ9QTv0f9FJgtHXARCe2+49
0z/dZe3k7OfPCJShsiswOa5ekeykj8xQzYq7Ksqw2N4JTWxMyiFTjHbQGuMpifp0
wOD9gOLE9aVctxi0xgacU6GXdioCuN/rD9/zA+b59g0tTtF41N3XojNzuGv0tCiC
KeOA4rIHLm6taGUHcmTcvCf+P2FAjOfphC1Xyk99w338NzrU54QPAi8iu15M9wXs
kihh5NuHlvR3RK3Id5KhYr23Bw8AAsV/2j0iSo/QahUSbLKMbomO+tbuqiyjhAN5
rArw+7nKKucM/rrpMR+9qkvEqD/X+nudvotAXrRKdud929A9BSsjr0oNU0Mm6HTU
DiBdbI2AqI+oGvOnFO0JB1j67BdOg6TuyMVuH7uLXKlky8f+uCJme2VFHmbWQU/4
qsIAoT+VoEdFtl75l4TxOEVUq05RnIOWXUZD01Vpms0hCHCk6ZkKOfyK3XtJlpeS
cd6DTrmUeXy8FTmpcKkBkzoA2XPJfxFtrYgYJHlu0w34z72cvYL8lGhSPM4GuSrm
zQPNw5ZRlU/2up87lYUuic0aS/Eja2mdQWiz7GVP3pcm4BhZoQNkHVm0v9FEVCu/
rtpG9dkjwaly3o+5vzVq7RGY65WmTCg3k4CaDIO6JtcZTiLAcnJAetnYYxtm06sk
ui5XoMXrK+W/BksGEmXS/3ldwz1QmK5Yrm7H02a1go0kdQ0KHG5KbvOW+MBA7Gh7
zY6BSrbvyoYpyuqeMBzs8Z2BgR2yEoo6jg86D78vX+gCAN3nza5EZbNfqR6kpBF9
b/MKmkhNzYdmCqgr65arGUnTg+Ho4n4aUj33C+2HxO7jWyMmEXEffLuCZdBOcY9L
kibi+sY697qRy3hLMGK6vxGQdvOQ9+k+iKQzAQUmemHSvX3MI2SeDkShQ3v90IJF
vRXcHZkXNwsemG/L9ueyinWHnd2ZhYptxedUvN77r++W2CUhg99UyueZHcg3V/OH
v4ns8lxF4bK349jimYx79pJcEh+6HO98f/frcTs2iuVhU6Xokw6Nq/5BZ5zU1x1q
5H+5wtaAsDSPlOhnzLuizYv/0lQ0lP8sUJNleFLLeX9y0P8xcTMUatbcAOjpgqsN
O8VZI00vVwkxRdx7fxOMC2B5MNkMWsDoathuZxyTS7rdyKu+/36jCBuNdPCV3KL5
3fuH/PwW4ti6hmEoTEl+MWbbEL3mVyc3iJ/TkYbLv+AmCmEhCdE6JpsVSXnST4Xp
HTyrkUr4bmSMH0A3MLcX87/pWthoZCRrfTsGE/gj0TTxc0+gtv3bB5A4LRXOxtzl
fhVLEIy92E6aY9AgZKlBpO1BDa5zR1u7ILKs4k482WY6QrRzcKd8Gqt4oMdhD9ah
8TtckoXnC7uesN9g4o/HqKU0SA/kV9vjHNF2+Ilw801fs5thqhXYlyZmelL+ucdi
dzZI56W7EFt3rMSKMDdkht6DsNnb9EKTq5jbinwp4SIppghNLDa9w44iLbzD9kzw
Tx7yyaqGJW5rT3EWUcfvBH1mGRGynKa1a91hzEH6T42L9H4M8YXKytyv6caO8z3z
Ke3+LcXK7NaQDySih/V6riEeji6LBjSDaTXArGNgVvWmoG19IkExNFbqFDSc1c6X
EtOAtfFKnGeT6ao8SnKgt/5/uBOOQQNsvniCxibt7CeCHIVEDTZQPJzIDTudbh94
9ydsiN0tsNsswmjtOlitv42WNVUnVsOpkr2Ti06VVeU8bycQo8PCETCT+XlDaucA
towMTXGH9pI0GEVEnSUpwSYZoSUv1hAXWxUhdEw9ZJoreITM9nVhgYZZfQR2ExFl
FDe2tTzcGNVCJcgbJM3VlJjE2VMC+xQPHSwK6KDDoBYV9vb7PBOrbRGzFA4hh6ph
e12N4t5Zvt+xn0AZm9f6lkUEF+cuWkBaPbfPrCWsBeNKsVP5J2tpbVu715P7dEQK
UsQTlM2cuInKL07AH2e+MYrr8it+YpWS3YLJw/+IQGfi3xhT0ENQROdJdQ4J0iyg
W+DtcqdOGHo8entmD9MdKinHuxaJNSOKrgIcyiiIrm7N74UIBfCmiFmqO9qUM7gj
NSbhQKHC9aTjJRfKwmPTUugQc2SLu2efCcQuaWkiemyjvg9ZnFI/5LSf3DRlTZL8
F22fwxqpZuVOvKxGaVnR1fKRW/NxBSICWlY2iKDPDj+EITSjdUlMPD7azf9l0DfR
nypigc0h3Kwi3/7gw7f93ew1JGAyYlOpIjlGpbSHHxL18J/z8QRlJEwsziUgyKx8
t7YJUDVTd2DZL8QaAzs6+C0jSGOHBbI/KqoXw8S2akk1DqJRelZnDiT6W+JpnFAz
0hk8D8HbthiOmpNxK3TUTvxkbAE4s/EeTCdsWCdcj7WwJlvjckU+ObzwL9ujXRgl
4OGBGAhjGVShxuKHXGnY2dcNNeXbfDOo3AwBiDPJtC+E+Y9z69Ny+7qrFj0/qiZ0
T3JEcJ0L9HCpM+EB6aOFiEpKgHcoWWYFR1O462ImYfKv1erqEax/K52444MjnD2D
T7uddY2Ei0XGQ3QghtPFn5Wj3W/w5nQKb5E5KixBYICzJTMcbuuS18sqvCiI/9gy
4yo8CheQHj5Djrd0buoWTMny7+27HasrLKET9zwPnGXY6YfOd311GfzhDg40YWon
nb8lLWAI/jI0zF3Pl6qwFaEVHYAqhR1zAcpvzi1pSkw5kXxSOzBZDNDlKZ/sfRCZ
UazVvka4qeivJT14l3suyxZa3shvGYG0FWZiLZftYsLkQYOZZuMjqtcTe3z45M3h
qai4JrScMJ76CC/leLEoFio5OqWmRtr6tCVVsT+hfFqkr76dcVgMR50LLuOETz32
zz0a0qRMsPmQvK0gQq480/xzo00JTO0YBsWURQg0DGsib87IA2fHGTOzqagG204e
rT4IELrnuyu1Zc96Dp7fWGRAebSQclSYeHSn0f18g4ztvHacorEAYO5ZoSp1PfjU
G3OfwG0Sv4GbGoWL7a8+6Bu6FFxTI8LBuIW1yc2q34NBRxHG0pEJZxD8V+ohQUoy
Wo9ov43yHFcyhd0s1DOJI7MbZ4fPdht3EsPyygx61Gc0awlu04OVN9ttX4uOThco
3DrB2bqV79TaHz7zSDbSu+dD06x6WRs07u8/BAN6xHUtSbxL1BczvrOJUVKdKqAd
hqkShn+Sfhvx8RB6acwlxtF6m42RnkvNFBWk8o6N0WvWkg6LZ1PqoYdRQsU5dldf
OjIm6n9/LAXPb50k615Kh1nFt7GAqbtrONqaWol7LWvx37j5QSecGa5qOOgFC3Hx
XgJCNU2MLIOqHjems23uZ71JD6G0QWSTc7Sgy/Duxs/dM58ggh/IZju7tYUZxd05
wj24E3P1BVQhw8k17cID+9WMy5JTthvOVAVBfuLpRCNUxvBIAU6FCxceeo2pNN2t
xG7VqHRu9vz5qbzeAC8PUMc2WCqSbI1BLU2KRtKk1RwGA9lY2c5nVrAyh98wALS/
vwLV9qsH5s3jdpo670gQ9XdIzQNKKzRQEucJMHsXEG1Dj7A3aH+hlRfE7AqZRMKx
/4mNgNx7d5E/fbl3Q6k8e4VCFH40yHnr6Qj2YmFdrj9pqHf8cRp1IdKH99FNv+lV
i0u5qxM8VtZLaHbEqw48rtUCf5Zq5Lv1QEXSMlVvnqFHwpupM56iQ+ypnJ64yXbg
oB+LpF7TjmLWyzVzdvi8ZxCeW6hTiCeLrRj5tWH63i+5anSfjjiIFcmaLDIl3utI
BXJTffLR+Lh/kN71IdEj9OFe//bqZVDIXyDpVSVb1VUzlRhG/WqY7zOiZdlx84Pa
abZk306P34J6JlZpPul3Xmhvt5XoEM1ytjVyIDdlOCo6g7MCjF5perKlm3U5Za9D
F9qP0kKVcnP4BMaRCwrsUBIEr44CiNBXOp8SkSRkTPvfiCWlYjg1rSAkExZ5cQNh
+4Tsj2VjAM8mdcAL1JdAm+VIitaQdPd2zXrqt+hg+QXVAr+bEJ0+HOsjXv+kIAgW
HS5FfxGoNhaZdRHeEPXMF6A2wtVvYR6V9Bo0MWEDcC1G09rqfKn/7QlzkQt9n5CX
j1Hb6hfGEZFPTxAR5CWefCECKsLcoXmdvYUCi60GyILnvgKDMNzvE9Wlx/1ReRzu
3hgUO/o89VdkN1NJdPLq0d+Yz535JNNSesx/LB3b69/+HEzqNfL58S302jIInby0
yMlC2lW7VevBX8zHU31rnDdQezavzydoJZvOPFi4xtfzj90kudotO3LgJ0N3mRqi
4MXVk5zAKgQ9YIKNYwN4HI/0RN1YTSxhdsHMzQXqGp1pTC1zCG+wbt6kL4TIr6lM
WWazMk4eQP57cNw0HpFXGVnAxjQB/cRUrQEp4t7sPC+xmS08wFk87N53M0d2JojM
hf5JdDmCQgqSQoBwuq/8CtoU+io2K2bbXdx7OjDSDoZ5ORg3K3uFXsljMJxJ5z0a
+LPk4kIQHl/8vyYmoRZ457oyttTMH0qwZznkkcozZAuBJjBS5Whhu/UoNOYICWEr
YIwC2Ptx02xa+BdtM1baF+Z8iYu8LTPixpRXt2BCiCIi1I7alBkK9cnqoRqywJnX
hpPPYgt4FNIraMBhypjTWPfDYcIUzURWoF8fnwUnIk11NjLKmeIIbWPN6MYU1f5g
OaI2ewfxV7wNOE4YQRJn0uRJWJpw/Y2s6VsvhHefmJw6TdMJwRXtrDeiHjiVPAat
MUouyvZGAffhKkAWnL8c+gssuihRAImDZnvfyMtDAz481PBIcpR/XF5SrWI9/ky4
qr/rNfSR/4pJHIBqI8mFR0lW7ERuQ7fJPDXa5/P+kXTf3VCUEIDJO/KJZ27D6SwZ
c+LQ6Mq1ttyIpYmRafH9fhlJ8AFVtaJ2VcgooQrb6MNkIcgIIwoLyp47pMoceBW8
3FJQi79JcsN8QTO9CsSztQSXKssKkKIQuFoCO2atdXHaUEEnJph8qERCpPngLn/V
Mzvqhq/dC5Kc41/Dp2lw8yBkHxdSdLPNQ1CY4czr51PSrUzJ6g3TQx5k3UGXPhDi
AZiU7VRqwfRYNgWcNxDoGeOfJiaKDQlVkE5SrWjrL31h2nKVDAXJbujIxGgH5Q9z
GN+buR4PFDhM1hxz4nl38q16CS0JPrM59mVrZBeBxMVZNn8rAi+cOY+NtFE8P1Ld
/du2zLntOVV+xy5kdiBcEQ2k0xoS1qAjMe3kPU3W4MEdnMKZ+keDrdOdTp5OHRi2
04pxvt2L0GSXi7ZPbnPn8A0ARH7IPY1IhL84zxJYFQAtRfQ3HDTmpCfIGFtFuQ4C
/OuROmC6Vs4wFa88r1Zbx2NGJaBxu1NGQPQIAei7dW5tf5jfmVSyIptGTnt7RoHy
pWHv+rxtxzJj02Tq9LHGaxUwFiinulFJd1U73GEiGRe8TdSn59+5GfqgQB8Vip2O
lzKo6DUaJMBu+PWYs4MBxWycQeKYsOdtlvtfYWFQ0YOKavzir29qNl0pWou99rvi
E2GLCglkBFpefrZ61SBkME0pGctT/jITV+urAiIB2UD0H7J3m/qJuzD2W+BsXwse
nfZK7VQN862mW9v21tn8LTnE3zTRAKV5e8gxd++7YhY3RL+FwhcSEn3x6B+LI1DW
Io1bn/LPdyaNiF00K3jIPnPxPUfzd8r2vbxT2ldgSMTuERm22wJGM/UDwQjGHB2E
EHa0gNyPTomp/2bcyV8n5SRHV+zM0DTpm0gsqaFoaaFirIQ32jzNnGzVw7DpIf4T
ki+RNcuqkupxd8Pr6ma71cPnB4ou8ofsosAutp5pT/70H9mcxcSlZmnIOwQSba0U
VfoQAQbn5Z3NuCqZCLcexDmhUXAo/ZC9/DxZLxYP1+5JrEdyoe3q58h9GQ2YPJHy
S6Sp6Ro+87am9VvpQhgXoyrk7KN+w9+Hp9iT7udHewfpkBPv6NmjsLcU5sYMECON
VSjgykkeB5sNF68IYZ46ijwcZNaZYeVcOBEIucE1w5iwXrCo2swUHCgcO6zkGNP2
fX3Rdgy868opVNXdujERK/xerwYPb/n1/p+6NlRj/AoKmAqJbcIvNV3qULYUPMlG
ekhW+r1PKrQwc+PqJ4tcdJUFi8sRbekriQtrMuscVr8r0P7yVz3s48wERVuSHfy4
eRBQovSTcoRoBRZDG81nr7rmthrb93BvtiRScH3jTrDChX8SvZLK4TsgTJAQvLdT
Sm5GBzeCh+/kpyGHV6njcEpgz4Z1sZ0y08F3k9qAfnUgvyB1PJWBNjsY0CtGkiHl
AKiNJaVJ7NICNYIqGyvX7WB1Xu6h01MKfvSgN8eNKZZH2Nfm+75PsvwNpFlJNf/E
OlfY8nZ4BmRdIVgJShvlNPaspynHZm+G3eGEDFX3Yq7OmTUT7vS9u4kVZ/opijqt
ez7p6vQ1svzuADuc4fVM0j0rLslkrCfM/Cg7oVk7inzv6VecvILzxSnCW+D6VIrH
GajoGRXwIS+JcC26aYlX79jKxfknogupF39w/4UZZLtcpFc6s+Q3oFIPRm0hS9rC
lnzr6fveRQwkdDjegQfo3DizJnJGeTW1WaEia2gn+3HUBVV2nRaWONnmnVeTvvIL
LlPSHOa8HTyLai+RBrskq+KZ7RuWCWn/Qj5VUGfheB8L0alT9NU9U7n6tgBDuc4l
a9NPigdAhvLs/y6/bk/zGzUBTf+R411eZ5xl1ZK07ZRpauOdhnLljHbIuRIFudAk
iYG411kGA/LcCmIbOs/UtMRV3E4f3S2UCEjm9MUFGFrMs1dNTyPrHeFTh9rV0dw4
yxB8cxPBOPX3ukuJ4L82BP/0cmepycfc8uYHZFZR2Vw4iY14HdeJrKw7lJr//AXt
IpbRix61VM/H9Zq1vIzOhp3iN/EhWYQOHNmZ7iozWLMrVlQTKsfsEuGJMSIqFvlG
JUlJA1UPOTzWdI72fn/EZQ==
`pragma protect end_protected
