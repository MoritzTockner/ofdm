-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ByHvy1oyJRK1rbFpBwP+ebQ6ogSedRPRtBvc9cvCywl8DmXD3XTJPWZI7NRC5yDz7Gz/Sa98l2YK
bGiMTIH5bSJNC9YCAmohK7WBv2+aT/JFqkOz/dQf04qJee6sAl0gwgmg6TuCRD5g/YaMtxDcCKJb
8mUuiMNprbf3fNkJTWpYQcoDK0ozZsUqQ3TozMdBAtHyYUC2KZ33u2jqF1Unpe1xFe03Pw+7+0Jt
KIyAkbdljlMUFo2bozC5xFY/4XTRNFo2S4rH4s6hDzQp9bAC89M1/yCUSV4+AiOPYIDcidOZHM6R
DZy7RKdwne/Vn6WisadADosDAIpaEmNk5urzeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
97GfWRNhrAh0ZKnf2VFzE6L+WdE0cpzMhbsjcUgJjWAzI+ARThqPec5XPUQBQ+OSLiJqzhSD9iB3
diI+AOkAsHwgFivBeOGSAX8WOQ2YPgPNM0z2p/y219o5crU0yYPbU3qZAP1/+M5Z3L809BuWwFSp
I9w7N0tB+nX0rqC3w923KYEPLfMBlVmMF6N1ZhUg6AAz7q3m6izJk4n3l3akYiL6+qzbK/S2dqbN
YCrzPzha1v0dFqmMcbi2FwEYW18TVbhOo/os0xQ7vWRiE9f3vfaMi2KkDmmLzJgHGUp8qHatVwgt
ibQpXpWdrj1R8DtfY1bIcvP9rhEiVAwhojlSU/yr2xoonGYvND2Egd6wDhKNJAlBQgNBb/7+r/8P
XbH2Ne/M659E8kOVNVB6SKIbd9Nr0PKoiaDFNsh67vpPCcj7Wt5m+wnwYi4p4GNuliJK+fme2QPZ
F/NF7T+Eog0RDs+sZPy3irbiAuJFOdgfUrOsDgIDpWoKHzYsTJtAg/xZUAueE41E+elsjOFY1OKT
0k/nMix/EmAj6pW8vkpHbonfP9ZFwiCs6g8bdKs0LH1dKgQKobIaQ5bpmgNSEU3E3shFEtf9accD
rF5T179pyhtfdNivrcUeoGCIPEvE4oapamRWl7BJKCTAWgWO0dWHU/bmprJTahFyqpdKcbpBEHZ0
K/lG2iF1nS18YtO2+ea4yJVos9NC9LwPe8Kw8DrbyEKTf6lbssZ9Shk5T0NDuJqqecOZhxygyTNO
Id+cecVo2soyMg1MPSop9JqERsyJQp3K4OVwpyF4cc7jyH5RDmn6mpL7vXG0Be9yuEhd6V2KOpsX
zlxzEeCEikbL2KXYnuop+3ItsMpL7TsDCPbD8qFrGDc+dbu/XapQgxiwjpvgLzb2IigW4c3jx19G
ko3+nBQBSXK/6GCZW3xKzQY5qfopARYUIsFg1mcTRmvJrk1smPD676ExDTSG06Niu/AcsJ8Z8jSi
QvU/bwa0vlOkIXBtZiNlW26KfcgoBy7rg0UMeupBZjuOzyvlQt3NV16YDh+TtpH4gW5hs1oOmJS4
fnGafmGsdnJjqnZtiIjVsX+YM6sOPim4kiy0tbxKLwk17eitYwA0QG1bizM7lptOLaG6gWjrUYim
Pc+vHh4Ycj68Tm6JsHk4PAv8lCVmLeLW34zlxRwiGtwNNL3PR7FJM4P5LgmXBHOMPZxagDGasj3+
S1h1sRG1Zk+32o+Bn/ui/ouibTIXxd3fDAA9tRvZYpUeOep0VruYxxWx+2m9EU6I+QCNfIqZ23Va
qq5rdyic3K24alTEggSOGLFwbeRGt+QB3C9mn02dby47QUCLX3kmsD3opHDh2JzmGe7ns/Pc6W+O
34zon098jmBzl5GoR0hxu0L91QW5OMwOR0bo6ZgOc/NndaW2lu39hfU/5qDgKSA6dL9YswW8waMb
3xfQTncVrgslBrLcMDyFOTEz1Ja+CRBplXo/dYbc4RWHutFhYQXIDLHlolBnYstpgfPppzP3uULB
i7fb/YqvR/+nByNHM+B3R/wzsCEG1dYKG8zEpdGRrCVaMJKU54F1IPJy4wAM37v4PEL9f7UqO7yG
m/2+rrR5fT6WxAweTzgR9br0PIX6CiT38SGbdzYX11j1pqemnnlHaW9Fv6SiGLp2+m10o6V1aIGY
IbNsnInSR71hrdD/vRj1Vso+yCO0FWdYd/S/erHIkBvTAqO/Tl5HY+xMK7Cg9wJZQIazmeREhPAP
1NQtK2trH+7LB1wtL1fbPW5IFiv1v8HUidZ4OJSx5SVoFZl885T3KzL3QBF9Q6Rg9thDFhnooIqt
5sLwOA+Ekt8+2rU4cgCNssIt4W8qFBHOW0zgpF9wRI9DdHv/eofDKcvXVX94G5tnI3AOvzL4SYl9
M4zcD9w7UUkhOXCyZJ05UP+/xblaiRoUrG+j+iT5m5uc5LRf8p5prxQw238N987RzbSUd+2gsZGF
zJtpVvB0NOO1NJ50KE1NCoKsPlYGglcO7FWhlQIargzZJzNmclUKH6v9SAg1vRFw4k/Bj+PM24Dn
xeip0kH2MB+Ep32Mm6Xz0w2l++OICwhtBM51kiRkJcqSz+Juh273cvmkP9go2rYZ6z2owC5DVT++
jtAKj0geCkH1myUyRWgthxdaKMt2YKZ9fuOZXFM5TVc8cwmNXDgkgi8nXyU+UinaTDDnpaWI393L
tpSdvBXZjVWE+hJqqDm09vqnWjSYAX8+QxZ2U/YzVsY7Wn4Ta3A6k+AoXZdD8KdoJE1yl2ecUlOO
EI4Hv7E3C5E2ZtP5wyTHCH+F7S/ZRJugebeMMbJh8xmaSZhSBCVIG61GvlEup4SHQNVY6zEiRLyu
yJlUu42fZJIiRsf1ZRfXRX6LTtZGy+YANwzfnBDt/dOUezdmnaNUyyjXhU2NwYqlJt8ob6ArsNYA
cXp3H/PUXNQn+oPMMFJmUIloWY5/KH0kPiC33UY78z9mAvDwThAK7xxiNjvYmK8LFTjmmjWjOsOj
hXGZea6ZdyTKVLKwC7w/tcTCz4SP2wh4TDxDWkMF3zq7fjQIEkSpxFbihmKIOJxzLfrT5ZZhg5IG
mRT5xgh91E85xm2SzoH97E7adaeFqPao5Lzc3k8Kuttk/+7srV1WYZiYXVTJmorh1Mx2RysDzTD2
4qbRa5lFMweZtDi5KKJHzg+REwBRpwOtUCq4MCBCnu0wfEm2laL73zU1m+b0NciCfngbb7GRe5NW
GuJEAhdeM+mh1XRqdLCej7upr4zLvvMJttlMxhqb8CVytVj4dAe/nO1Yxm8RzMGKuB1dZ8jUastq
P2q5YAzSzhT05pviiIZjgSLlF17gy7Iwv7p0HsQ9+1Cxu7EPdmm+eOS3EUdzWBARiqLnyKvq+54e
GSgPWUfcNJdD4cl3GC1A5FRDRWyFW9NldHcG2wmkHxj6yxHqDfVXGj4+ahZIJ7ol6oNwGSXrsQS9
FpAafIIt3Wz5/tZgARp++GCjUjz8GEwUOdVf/ptHz9KjLoajPpGx1VsRvuuEHgpnffaYMD+alM99
l12sn4DzkzRasFNhwLiTuscmNbMJ8rQTiHlt2khd4J4GFv6NVQA/0zsAe4BLbl5GwIYN0BFqA8x1
Q3rgG/JCKOe54NnnkC/w20v7vFOkBn1NavusgDiFCkcTkf2CdhL9UTZzuCd8kZasWgAGNMN6OZOz
WmzB09sH80JUhiOgoNaaXOSkCn/7IgRn2kE90bxL7A79jBuBDxjavQ+XLFYjVp7b9GO71do6wBz3
cBtK1xQxXBZ5HTp6WnWqUKrXJLaLlf+XJJfYlUUdWCgVGpRZFwiZeIB/JsE0PCjk7ux8lFTu0mo4
zG1Q+GowXTsVbbg6Vpr1nozOJ52eH/3ZfsuXlk23F+4R95GCMxgHPcZe6TF8iIg73BEvpvWD4CmY
aReZeRUGJRKkbdZioRH3P7oaTe3ws7GL+OGuiefD1GaH3oqZ/EZYxJQMvm8UlXJRKXpn7quv7rXd
xHThmG3iJ+dpG7/94Zn2ZRDvJSvK0u5ubSGbCrB5z0IWSCJ7fA5796T8xwZMIl0gJmLvr04j7qyb
UcowzZyZVs0HZihPNlpxCYyNPMS2YF6IcvJekhca82733W3Ee6z7H32XuIY1huaVFJ3Vw3J+mH3G
ZsCFfZm+vBNV/xnVARBWph91RkcwVJZS6BS9RkvxHjHsUMLLUguuujC5fkiYJ0cRei4mAAnMboqK
+HA4Sgk7C11vdhpRoS9hmHaJsJauChaovyIf8iVGu2aMEM1elUC9TirR75JnhRcqWmUfKC49wXa7
DJAgvZ9YVk2uktmBXOL6x8RMjgTpVfrsvDubeN5C+PlWsXrBdYpfgAeGz3jyfrIViE6sqTUfbHBC
RSLEemFGKWdmHoXdt9HUh2bTrMImvVwEQ0sBUrq88KXjfnvOMekzWIoBmIf8nrjra2WArRUT7hKN
Rr2sgtoZP+q2jlOGuJlhobhYp2+jjIXF9WY+aXu5s5OW69redNLLaQgMRrXWN0cMgm8zyHQBD9Hb
BQ/bgiET9K3wPtKPKGRrLI4f1K60HtOIoqt4CzjURChOkNcMFLAg4SX0v9EXHsGS6vB7XgMvLZtP
TlIhEaCifuGtu1/wL6DyId/6omWCMavYKM2oz/OjuQ8crGT9Eafq0D7InDKfOmrOpBgpPjQf3wa7
iyzPm88gGVYShaqR+8tUgjQPQkYTz6WZ6xPgCTXJ0r2URvId43aNw/Ei09Y8+7JbQZeKncczof4p
BCMKh4RG/itAFTj65PSzuxWfExJXcf9gHzWqJFP8YdonNmS/T50pjmYVcrZVDgZm6hpA3YlLCv/H
7XZbqcW2ESWkLor9CtI79Dk+eWwdqCGH3hXI+Y9RyOfM4A+RmVpcopICAHWkLx8EIWAd4w7yRoSY
6ojH3T8a0UcAzTdhXTDrD0aWmuBo3XXywCxk1uzcPcOGQwW7dP+J80fDHDbdzUTEAxhDKXXpOUVC
yIcq2Xe+CEBA+MfvDqT0lQdcC2SnvoEh5HVfjB7KVOo3X3KLwugwUXKOiPIshA4x313vgKvkM10r
Q5eGMA2PW0XNnQASiHFDQdwQAOqcKqaJE4MwPujrE0SlipjpfUuVTbtnFup7F/PRbwoQz3nqVc77
I4nc7mka//XrsCHufwrhHWptHNLvOWNpuEA+4IAD1RzJhNnvYfQLUqubugSOSkLMYJM9XpUYE8WU
+TW41LPyhAsuVhWZ0LSIQd9lX4Xjrk2LGCUIdv4Vhf48TOf7OcPd41X445JHi5ofYUx7XshI1N+p
YA+KbHbPktE/T4qGiq+84wo1dCnkKtY4rtwoJFPrERCYTTvWyDlHx+3rfp67J22j0t6+a1Pv+9cb
I1HNm3UcVPQIr0qplhZ9V0XUxZge84uYz/kv54M2MPU4kxmaodX5DHZxBcFf8TyooDBr2WlnrDy4
OzD7zTJtZVG7dp9vStnUkfHjLiDtyGtvAmVn2Bft4Viqf/ZxMf6ebtveS5wdFb9qhnZDbcp3yLcb
Q3YTvDrsGfynE73FD7mwhjmLbJEavg3cREb9BsH7AbYyojvT+dcas2PA9xLcvqEvDoht9JzWd/xY
w7O0SlDEF88nqEmJlaG+q7WTxYqLoyZCp19hHO2UZxb6VSLDB0WVt7aDW5FKHegOS7ly8KA6z/yv
v/m/evaq9heOqMrRwFQqU1h/yOWOHR3C/ecwB9Hzu8cDGOo8AB+ZPD5RqiTgbynGtB+tGi2S/JG4
JlXrhFcffcAz/9Bh5q1N7/JMaKGy/uTs6+Rkkq7oVOT5KYStm5lT7Bx8zf83EzZtqPdZHRthJfOw
vrr6+Y5E/0M1g3GdEHu/JKFXysHn5ta3W4RXsHwUIi8eN3+NgbCFHlU7WEP/4X9tAaH4kh/57T2h
RIMAYLktaae/QvYmfRC/lp8/hgFlafblU/2UjQfUhEuu4cRsaTKMkrIgTg2pEstKPzngA6SHgbow
K3bTy9SoQ3i6mLt0kbnx1mBAsNHFAotEYoj+AfcyhXbQUzCwW1htfy+MHpYdGthFRqaj0sQYvuGR
fyYeilvqkquOKZtI751kFDkEmTpKnV7HHwCBMF1KRDooXG0hWX4TKqSjsmDRVA7JDBQHuKKfYi5h
Hf9htLsKsOWaSZ+hXh14tgFdXikPRCHt0QkK6C/xQ5yrjl/MPTcCVf6C9O27e2QeNwwSzU38e66H
HzRWnstT3+EPPWwTraji33MQt1uDffitKwzgjI1kBwrKsmlTXIGjA8mOwdZVVtU2xq7nzPDulSL8
pnEEV7JTjmBtkwAC2tU+x4VpOG9ixkkNR4RvdBYI8eKZmfclVWCDwh9SKPEjO4XzEfDF63IheYTr
Oww/o12gXolsqrf5xZ8hOZFaWf2nf9HpgEIkPTb4P4ZuzIs2EpSG91qwtOuDEQLqmK0782uj990R
S+azfAkWeec2Cr1mQ2m7v/s0vaMwksdI0JQjUQC4D8HrXXHkxsEffOSTyJPNIjVCagE1gmgycSE1
4IgyNnrW3U8TEqNvF9fv6iJuG6W/ZuVZvkjMHrG/Q8gP16Pq/Y2Cqx4lMgUi5PnWXTYyKi+8GKEE
ZtkvGPB1++E5W06GqXUZz+JjznboWoCo/DcdkSq4/7tDWcq03RclyxdvlVYvEIEDUy+8YivFybdG
Pp2tkWtqXxmPO3fwUCXvIR5YnFJTqc0ejdekCEgKlcBzwdzyixerG8jvQQNj4lx6xM6/cnvmSwBY
YQtJx6vmor9VqOvAq9c0yc2vzKRevOt1G6y+xYGdoF1yhFCNyTDYyqMIfl1yb0pqBA2jo5Rirxrp
VnDXNjgB1ktfionCk3UUXfn2rLlJn+sSVCiEpdwyz/AlY63SER4CXdnoB9uY4pjJZ0yhwJ3kmpc0
5uW5DQuQ97VZKRXY675Bfzah5zkvVFvaLvzm0JwMXf3JbpX5EIkrp9RPudXOTYC8FqUo5ifKbEKf
NycuXlON+V5fjXAddgsIUNiGCufmJopFKtqFu5wm1NdgifucRlZdtIh6g/uD+vMjeOM9c9otuspu
/Ri244KA2sBg81d9EM2ez4ZJq+auK7j09Vt1CBf6QtnhZHzipqRVo5zgC6eA81FP2KfLP9aztWKH
KlPJKh7KLzRrSoCIgDosVLd7zae0/llEy24VyRWMbYDRTBjXsibUDtQ6KU5EShTcdUaCUOIQ1iv4
3UqZBliuHwSDtdBCEXPNtLLkCkmfSvYHfo1oqhjE7vKYZdAhbeNssoD3H2IlPKeVyznWUd5Ug1No
jB06XJnKIF+dEIrOZOjPm9wNgpDQwcdNaDfXGWk8Y+oCXxjjMwxHYLxoRMi3z8sg10CEnYZCB8nQ
K+amlmfnkJFR86cRwRsxCXf6A92WbBRviuTcTGRDYL/CHN3BV7FPsn88W/LB8uZGe3UAzU5aNWn1
8NDAYi4Iwoqbgb2jD8eWF+8rysCh22K+nkbd3+cxVG9/aG+P7unBdKzypuXI9+qeR/IZc8B2VgMS
xhN1OPVBp68WBtPtWrnkcNv0h13CpocINEy3fuYK6wzr6c9tPUbc+wEB4qy1b5D/H1JwzmNPOeEt
BuXvgBJlN+6TLrY+ba8PnEdJI1Z6JSE5TGZ0FX662Ljo8nIvifM6TEoFjqw0uEBzIcxN/1uzJ31f
iUxfWbe5Wg67lusGLWqRtGw+0aphPsZbArXrfQuHBflvj5gJCBd8PPsOlpC9Nl0ua5znY3dP/qlc
GKgyQjL4g8UEvVchgWhq/IAWUUh+jbktjTfPPB96PayrYbYCO4r+GruZi7Xr8so1iQ48THqEdlR8
Lyjby/D7XOdMzndGChMoaGtVF1hdT2U3yUJ6weYHN+/cCSoKLM8ZpDHeaA49h+7QnLEAkrtoI/dY
E2mV0Wb/wC+tdEVfUcecSC3SHev49/6CjAzbu30HqYRgKqvZIRSKnY2iRjWBOosCqsIUn2JDzbCp
GYndY9W/v1fDVNx2cm6qfaMv8WosADNuZiy2C+yQhGBqkAu+v+MVrW6XZiOjHh/bAq73paUJIwtS
sCkHxG5k+m7efDQ8qe2buMYXTfNvGkoM7D0WE1y11udI1FQ2XImNVHc06zcaBE9srp2h0HkkNh6L
dQUlY0VQRZyM4o8KyIMshwLmPuK+Ok1ur2J4fwTkOsX/4BXV0YAB+PLMOMpp3B/VUsxNKFE3jdBb
LcegGivKVyXVRDxKtdY9auItmnXcNLdmlaz/UvrhrUBNjaBuJY7lOsg35u/d6C+L+B1v794fMfZU
359FxULzAW7LTEDYZFWtAMo5Qr56Jote+w+TQDSNg4fxDhmqSNdaK1nryfTAGItvEoGNAKLD+SGI
eUDOwQzPASkLl8lj0UcXkrIvKsCaGH048anJ3NebqvgaEuHn4rmqLAyS8YmQgwiVBzFYgsKUab/A
kFeZpZAxI9gazSKJhQGemvYf3gIUL6oCWxxFI5GOKgHXwJWTiCX8QmN6yTIN2OaR7N7/HWUftQb6
mN6WYb+o0jnUV6O74bF4t236WlhCM7soBx3RhUMskVyob8GcYLEOu3YuTqUHSEI5CK0BMgHVrGAt
7gsRGoAeABJ4Nro48GoqqJr/ffhgzxGo3daQUNcPnlM2uKfxTKDWq1wniG8BA6xlye3uhj+uHBDJ
rsn1qYiHx7dvhLW9Y70BK7g0WRAYBEySdm5f2ZTJJUytE4f0lZeHsOZxhEezjW6vmBcsvRPvsFtm
P75udsKPKJS72tdnXjXuUecsV02Wnc4/KkJpYdxAbxw4QAtXUDimyhbk033dfg2pJnu0vFZyAOER
7SxcbQTHDNw9u4FGfnoiTyNp2MSL4KuY0nA6Wz2k1lV477VBQfrCEl5Xczdw0mWh8TZcSfewt0ys
ozMF+lrKdxhElbvPygRdtPAfQLP0V/kvoK0H7flY0Ki5U88xOBe4RW10/Nt6XLq8AvSpN6FAhhQb
WSrLJ3i2Sx9Ecg5S++0K2m0wRbL93LgCdPpF9GweueoZap2pr8LIlEQrYv5NZkhyjx+Hc3eKz8mH
btxp1Xhyv8ea4VvipnwY5CYUYWLl4lm88vjcZsuZxE3GL+uZ4fft8WTlW9yaSNVfMUrqZfiSRDG7
7TmigcqLcx36hXBRYVU1NUzKA7d5070i71N3Igfvz7RD/rxmS2lzA2uuzpISNDlzft4J6CdAp1Xg
d2FEbH1wHJoSRunfozuGee+8roHA8pEPQ5y7TvyzFbjhlvxTcDs+rvnhTLgTTS7i/La3hgwS/ipD
7dIcV8jnmJwCKWbPTbm1mwyovvGxgN6IjIYbFVln29/VjnSreGHeVELM8Uh7oIUd9imCarTLCzCm
lI0OaLuBjJn7332W5+2rdS5UbpaQv+WYqOJv1cJiMDMZCCID1Z3sn4p1ueUUlhD2ZFfq1TMvYzFs
tCPs+4nX6rTWa0hm4uCXSWExr+vkAGPE6cxw1URQex4BiYCXSj3cT/tkZgtAQdOp/cxgYx7/0utX
Da86X60Y8SXK9a7SZCYeH9JRECnuly0zu5X4eGrIgqWYmhyUQ2Mpf/d9ZiDbzDQE1Pej/SrUKFOz
u0Drl902Y1/+m+YTcJPW3tPQ5K3SQ+MxO8hU/Od5AWnT8xxIF9fnkpPLXlWx7dAd6E9vWdi1IYoB
dMqITBBbFZAUIfi6VQmkBgK40fLMh9M372nwA8zADqPNK6ZPnvGDm0L0/SZjsJlD48GSXX7gdAYU
32jb3AGt72Fy5/nrHecbloR1BG/lPl2VNm9vJiVIYLh5f44PkrorwrdWp3WFMgEl0kc1d9TLMVMy
INyS9IFTICaNNaOszmnjt/5yHpGw7pzis4rF+VndXDaON9O5oy0yGyeRmpLX9bMkLmj4hi5nWmPY
sqb8frqyH6QFk7JCpCat99mNdcYnt2qGY/U8JLiJw+98+xU3vVRX/9qRAajrEk62Hvvgm5Wqe/JW
qZn/zf6g9ofQ+vkGYy/nrN3suLWx1GWL17Hm0b9BxG8OJrRDD6KxJWCUpnIVN/b1yEeR6mbfuA7l
wYXO9ov/X3Cz3jItotLCwx0895BsqxRg5tSv2SdUrkXKjikdLMb7/LkkKlKoNK3tKlneNiRQtWH7
g1nKj/3IXFIjH8umiVO+EKgvHq09nZxo0f8opBCkymNbydG1AznM5iQvyfts5XsvXwiu4fqU/t07
iDqB1vrAXNakCAA8jaBdqOkrc0/EtGUzuefuFzi2qbvXeMiKrZq+u2+x5DWAo+EgWj9aH2AHwGS0
ADAQ0w18rO6ouphv0Pr+0PqlqqEc/bujbj8E/nE9o7R6Vad69VH8Pwxk6hi1jC2bzGjXwaWM6CJj
WDRhfFCyexij224Rw69oQEeH/oO3YdwrZWCTl50vQ5fth9sTirkEljSWovMgYwyimNiOIgEIDNOb
hCIKHZ9Tbfo6rVvYiLLIn4PSwjQ/I4SEbU1RdEzdqz0N2/XUldPR6ZX5YdtaVmYq4ToHuhED+uZn
9ENbKZj9CzU3SyhUqQEfiQQYnpZwp915N9ucSd7xbpRCuFDGlWf6MW9VkPJlFJaILXMd15pB+J+/
jdv1OpdexhBRJzHhjYfbjuSb4o8qMUfzPzbPiqoUC261a46WnpkP9ThqnywqCYNKh0Kfcfah6D8l
kyVDBlxu77Z2yXQpdK18K46qReyHyG9fueSYE0SiOupalRZnSGFKsjJf0EeCQJG9gopffPneBnSK
avIf9JtjEzbvZPhLZcWqBUCNxqQmu+9ACZmWZBzPTs4LJuO8nDn2qrBy9EkabK/EMunlZ9eSGMBU
98DcTekgSEOqoYLKBcyKnsei5k/6lVnVQ7qkw/aON4/IpM/Qcg5+adw+XkXkn96KlT82SQ777OUK
FU+Ig1Nqe2wqZs7ilFR4Ms3g8wK/P1Nyph3qCGWKGsHvg6lB++iNDtnklTsJzQ2SMZcjc1LjeD0s
WGBdj0I4rxsUSqf3oR2oDSPeML0kZxHT1Gub0CbpWa2vJUwpizUdpKAxa3rXyXTm60FYb8Rw1fTB
nonAPRasB226AV0mCvckOdiW/3hJGiP/e6F83AcZNI6eVLNbEopAwL+oHCWUlAyHEJMgSlFF/k4j
RSXJ2tvz1L5wL94ObrIB7Tqb7CzCKgl0pgFN566fCSTRS/Ex9iFxOVqf4qtKhtKkCsyMYqiPMnHm
7HR5/lTPR4fWhwNbTls8GvrPrEUOccrENjK0rL5xfrZIEK7ZkQ0MFnK13svnCjCNvFnvyBG28nuK
SuecDU7uX9MxSIAag09w72oTSRxwnh4dGTZkFeADc32XQShebEKGwIhIOI7p+FD9MKfeEEjWKyjI
upTsRamOSYD+5vV4GvP2OIsrrvgZdYv5D2mGA1Fv6x+8CPTHVpXIlINadXcj4eLeJmtatuxnwyqh
XC/+aG76oDvPiJdYPlEvzyih9my9+vWxWDpVKEkdQkmqPhSBu1me6ELGibaTkSxb2TSER0CfxL+F
zjlFhKu1Og9q52vDPAoTVeabsLQxKBgnJBZOxXo4gU8Xv7nDZhU4GkbWVm2Jq0QW1c6qq0EQwMM7
gyHXDDw2jwyDZL5gEZOhuZdTjROtMdLy0wmwCUiNUOniBGheMnUKXAzzxTauNcZ/LksNukhWx+kn
rHdbj0xoJ0G56HhId8hqnF6K7X3kAfCjcFYpBslPbJ+QMKUPcDKMnr1OiRyJiNaKXbP6ahZJIuhm
NK/9Mqwwu9UWB1wtA/+FfI7SHg7gO7LvZ5AGVqWIOjX+UVS6v3YxSERQuB/wHTZuHkAJtcf4TdgI
aIUufE4FvxcvgzaaHCopn+DWitkMvnPCJbXeIHoYg2hIHwuxw/L4BgkGaIfWHKhoQm399ZSA49tG
5evgcc+3jBxn4/J02raVEhjgrRFJRoM4sOoE0awV/xp5dyUFi5y3j73ntlGDnfW0upkzR2W4PEvQ
b3jGmRLCJ4UUZqWTAhoebCog72xI8GGy0bXox67t7tSP+Rb5GSofasDB+/yukrx1hF5efq5JHOD/
vuC63qGQs2Ea3eDgsfr6SM1Qxm7uLCsOoq0tPtA7KAPJyXzVMgpy4le2CSZPASA5CiBP703aBbyT
HgvLe5uq1V+3T0a2bgrmOangiSua0108hJ0SnAAXDPq5oZvosfRE+rLMLjTFhfVUqrjxvwCiX3CI
eiCjLccvR3CYZv0AgTa7AdKVISL85hurvDpuCryAVNuL0FLrmpuMkVHOoEjbIpBQ3s5p0+XOAdOS
Z7CJhu+LgSpXQZ+9p6O/nVIZDVbcSDufjIZrDJ4yNLg+bkVn4miU1LHO19FuU0DeL3ltiDRTrwp2
TJlpC4VlXCtJjZRfBZkcyV1pnl2l4F60BVKoMbpiBLBUObLq7NllGGm8SbfA+EU1HSoqgRkFNa89
4i7tNPjQmplpgatNXlVavy5ekhd0K8AFZvsUnxUau6RVzeSCoqHVQoPkdn18zFO9puEx/dj9LnfV
CxGTanMPVAmnDBagew74LY+2lyCccvtc9BK9Nex1eaxHQSQ+zTE8iwZeppRFFSVFcBUyWa+JvpXx
abfMeFoK6ruZXicRxd3vQOKR7P8ElsgDRr127rRFDn4S0tXvzKXOeMRJKgC7WRtGL/XnTfWxFotk
AUUvtKw2QcOHAtMDODzaxgOytxEYfSoHhTbDwNEo/eSu1A1blPUPmGhYrOlZtYTsYgnox54qRsXr
BVNX8NXxRgz4dl0aMSGD78NjXp2mqZkh/9is+rH8/eA7zpzq58wlER11D2XNHvvfRMEWi+9VcD2k
p/HMdpI86qx1J509wvAjeNnMwaIZ+/maVTjtDnfunCzv05YCJJC1SDaQo9qTzC+pTbbmI6gX7Y2R
oY+stme+4LDIelPYykuVzbAeKUvedyRqsznh59/ieRJAZ8WAXyR1GLuGt8hrPDC7HGn3xuiEWCx7
zWE46JgsExoKrNnOqZk3csM1qaeXlq+eroIR6Tuhch0gAt1uExkjpfdElAWuqvdU6Bwa5PG1ze+x
klExo77NGZe/1LKfZ4fMApi6LmSsy010GydC0pJXW8SOxDN3ZKYT5kDK2iVDc7aOKIghXrI93Z94
e5T00xQJ2qXaeW01fnM7ZAqRT249XYe69zwITq3pEKU0rLAf6s4xObFlJXQ3buuhgkS8Hcr4+Owl
KZWwmuqa2/j6nyPNLVFubkrx6Dlb0BoqTuvPFcGAHDQM0teAWXYHjHfn1vV20W1bGUQ7TaaD24j0
NozIDKtkJp9GmW63nxMK+Bu4at4XB5Wzci5eSxnBMdGGWoon/Zq97c+NOn4blJ99UCHZ2zseUYbP
ubowppR3S44ynGBfUD93xVhbcbVaDuUo0zq5nQbpqehego9ll8r814HNYS9zV2BOF/TjB4V4Z6QA
8rx9f71XjEO63hxn78SgRTjjcQR4XzZtmMXJz5BhSuGR2L46eiOszyF9WectgOuEPdWbpJ39aXvw
i5rz0JEGTutRlt0SWw97la7pHqpigGmVN52SPaz1OEnQaJYZ7hjqLBBGsJokTuAY2HVEIfyu0ux6
N54NjlZvoqSl6Bl/893S/g9oRSgfY8Am+j9PFeZStBEy0IPV5dXpla8zuLZPnkEJzzdawgqe/s2F
Oi4n29g3J8oOUfNE60IRhCRxAPm6bx95mPbrfle22LxkOzRr9jXMYkHgoMHcnBSze6r62LjqAnXK
mslayR5bxn18cNLGQjtCmenMbIDf66l4E2LijyOrE/Jq0L11/fC01mqorZ8+70BTTZVW2J2/Fyt3
evw0fy/ry+mR83neMg40/5HZDSGyuPZ7TfDJX7ev/Hs/3Bx1vpe1B/HxFBIE560uiF3yFvPqiNpC
FqANPOL0Qg8jyoEfsaEkBCnOBPe+Nmm9oXxl5Yf0C9c4Wuts2/5o5jjCBEtPTujowNcbXx+WdTdF
nE/v9MSbpTi92M9epCaCh2d0T+TjMz8NnfGb6zvwCVgHv24QG9GgVvaY42dTUQCUxhGzHr8Y7fPj
/NmJBNXMRnuRS3t2y8tUNSVqaq72MJI7BvhrGFgjw5MV/FJNl6nXDB96ylltjQ5esav9EfRh1PaK
8qpyZiIt1HR68u7BS8HxYEYqBb2dX0xAxwkvOAfWnI+bOF6rVw6fQ+2MBG5EP/oJkJEAYTl7hAmH
Abc2qBfi2iRtPWr1s3aEvg8fLKxtg1lwB0suE/6onORQ8ssPLx3s4//Qi52+X/zrNxskI0WB/RTw
HDtoNt4yu0F8vU1YHyLnTkYIe+OiLce66+cS50FIvrOIaqf0Dl/mdUFPpu7IDdgDjiZH1b1lsUVA
NCJ9E73ysaRoiEDVCvlIwe/MGrcynJ77uJTcyJr3ikr4rvyRRGFWQGUgFUoBG4AdEUnbLdppPVG7
COdr7gBQd8rgyX7eEB/GuSfEQXCRN7N8vUUXmqlXEBYgYHxR3tz/B//d2ofiMJ8uk7TTOHgSXazR
jWIWTDWh6PtAnMXk2qjC6rBZZbHdgZNCWo0fjhnnfcLh7MyOPDyH5vErD6L4SBA1X7pyGruReHHH
KEEfx3pYHROEAdueACOSkm/MbXte1vXWOdpHhWicT4GoV93mOGE3nAc52f11vv0UjLjXqvfnJ/Fd
29kg8rPoBspGGKYCJSrfKTQZw19qT8ORVUrGJsii/CwFDR+bGlBACWJSIyeGodvMZdgLBn9s+hm3
PSx2ul9ykNQgxy6/0bAexvdPpswbJlFjmUOzl4y9cxpvhNKxjKpNA4X3ZmnPkCcbyPvRfUOdxV/X
wNNGjcQBa/sNr/aV8L0Q/kqqk4eaWhYAonbUMsc9LCfcMKZa3VD9U01EQDffxe492Lm0TbefLjgW
OEzudh6yos8dvfdJFFsbPiKvsWGsyiChHMFk+JOC6yDmmrccoQHN8foBcTBmYULbDvBwrf9F7afl
9NdSZ5ZP2Zpb/p7jhd33Lvd43FVpqYo8wXyFO6JYbI8W7B3ntrVroimW8492QACJJqodBbcHV+05
tJtpdAaCWK1e8WnnASGJntyj0kSCdE5sUi6E4DNO1LevBBW0DrKXrBFFd2Y4o9Ju4UyDr9vgDEG0
He/G8Cd/BsOhGpyZYLIh1eBj8SGf6+sI5e9vT+9HxepETYj/lUUa77/xVJQBcgMVtNaoledlHKs/
88gYXCJF85aveaeODtu6NbRX0TpSc03sXN1iKZkNHi1nW59TahyzkHn58hpsxp3dLE4T+VNOO8ro
7/pzNoDtiKnbklfnmpT9Yo5SauAxQXHza/JuOOqj9LIyJkh12LfO3USNMaia1kwpr8oizW5pLKrf
2G9U8rl/v/KIQyphxVtlRWsaKLALk5fZZl891Z4W3MCDc/d4IjgfCOpz6gcVvbEMfltyxqUW4zDx
KuTG+Bz1xXP5deeXYJ8xd93zm14uqgdvRmpWqYgiFiPeI7uvqwd9zKwiOd6MawLPOyC2+jsWO2WP
OUzPJygWN4AYsAreY+fXd0N5vdOTDU61X2jRi4uWa0NA8R8gztNFgEUEfP1msQ+sTeWMiddadU5v
tBecZdMbH7GxNihzn5HyrNDlhVcBlKVQVmCYzIqbkSf3TfNbU8R7pH+Ru0xCgjQ+AxVv7++of/sw
frV5cp4P/euQlOtX2gJYg5h/3ToFYfTA+qN+p6SC8j2VNwQJMtcFnuiUhykeH+c6csmjcD7bvcDa
lYVNQU4V1fiHRnLkZXYklOz6q79xMWc6ti8DdGnrInBG1jU+TW4PZvcax2DxtGqE40kzUBkmrcnG
ed4j12jpEWnVsZ6iJa/gBjpddszMZjX1r91ERcMnXlVGbxyDrynaE+RI3BVUo3hLaBGAWs6DhAdu
ZpP/tIDbI3Bz7JHezptqPWK3WtC35+yKiNY7+0OQcr8AxsoF5eIw/2ImsnH3IGkxvOtxqWZRrnBl
l6OI3Xwq8snxKy7OKEJdxRNQNoAFgvpwUdIrvr9dZ+oOyBvf1ekycA0rOZEI0SWkbcWcuz8xsrSs
XQvCYPjB++4haoSCAKmMVP2jnnUvzvhcBMHKM/+EQgIiniBVIm0LHkNqeMNFXImwI8Yx5JFapRxZ
2Tzo0nRd70K0TQZ2X/wfeUv1/qrjFkmfaS3JMr/gt6cKnHpjzmt0Taru3996T/bDeSrLkrxVhQeY
1cuzPmap9w1oB5JXNH0kgpa1KPCrmCVCLGHvGi9M85aTsKCp37cO78v8ALcLnmFcxxqsfw6C4pac
I7M6zfw2KRO1Twrppad2tYkPGd35gDMY97uGOgOYqm8POM+3sve8eOGe06CpoJin1xYicwp0CzWt
muLnuMfdr7rPzbBJxmBWkFHwq42WBAahh7mrmD+srlnQthZ1FTbHD6zMRy2IRMWlryI8CwO4jR3G
YcSTQUBMi/GrNJBivUJ58Vryn5AkPGf2TxK+eORDKYCSbRMACdXa/s+kZjO0V8rVFN6r4bdN01Vz
B53h/KirH/4Tnt37b/qfHVLc/icUyi4I/BTiQj12RBAtP+jXnNR7MZ9v+qVLA2wz2bMQSuCvmZoA
GgsZXoH4mqqo+yUluAmr3CSKJfh12gwdHynEzYu8Z71Abo6nKAictLb/SDsHbpybMURbaG19BGEL
0D2NGCTKuAE0pf1M03flQmQT06Y1EbZTK5CCWdSjuXNp1YL6CYmd5ZD9fn2Ba6fFKW88vgARG6Os
zdUs1mUjMdiHp9KeuOQxmhdGAXy6DR0Ah1RdsxnP1TScu/G75W9zNrLxHFkprWsDOa5gCXhqHiwF
vJncH/8GEdd4FvT55T7Pt+KB9BeeUOKg9DS1VPhVL2s1IJpZGs120hd1jvqRF4GdStOqgJ1V02hE
bK3tfS2+D+mfds+Md7/regJmYR4hileXAbzajIjCp4AZPsw9HOJPnmmgV5GZaPyi39ogHdE6UClj
nSP0o5yEqSoTbrhttK02Gjq2WedwRIVbQD+mnMDf/5wiW8rbJBcgUFxJjEOe5HrhkiWNahAuipX7
iKXqU7fSuK0AJJD/OqB1m+PbjBdSn6STQ5scUyV5lMNof7Z68NEIeE7EDX1d0TpqXpUQ+/kyhiNZ
loEOUBkE5U2J0AnrVcYvMTQQLKvkIFI4A8XuKY9H6NcC7BDJz9NMuCbo7DDXr+4HVWZtI/L5ISDN
tX44w4c47bWOJ6QDyVMnGIrm2yNIWFhuEfvPijDH503Fu4ehRKloa5aYaLqF33/6bzLYCH1vH1dQ
1naG404HMV88sDbTU3KWq2zR7/JzVHL/J9OFAywA3rHepS82fbq7vRgsBTTW5ySgxQclnA3BiGh+
P/zHn/UGLbfOd5cLa7PAURIJJxKmvK+JgvlmKR4ScV25jbFoTr/Lq1vJnIIzlhwlh119j+eANkJ3
zedxkV1EWZAXULyRhM5z5uEeLUdxtYvETpsvIQL3wUgrObFuRBey2FLtGlsOq6qzjLJ0d/yOxTpH
/sJ7J4vRInx3H62Cvo6zWFWYrwAgFIKwlSsTAHlREQHhhRqKyu/lg9+MfgnTdzGIwVHk3BuJOL8Q
I0LI9IGiP0ZT6Y8LOPa2PTLitSKYsAavdeFjyCPBxi75QD2w7l/ORoT0CaTbp5YLyMUxcRfoJwn0
/JSEaKEj5Wguo1h2c42XuCh8z+7SwSSkp6pC7R6R+v3fYnuOM3w0d8o8F4ZaxNIrMDpjVdPkm6Mm
JcAVRPvrnNTyPDo+muVt/kT6raXoLBq9AAvSuNJIFcZRVgydyDVRgjPXMyb5nxJvhf6Jh4lHqYtf
/YQEdzPC8gqHMfXgE0psSwJe5Zk5Bq2BGLMRCoR9uC0vGgWVpxZeVVGgb9weJDDIK/VoJFKAHSAf
rulgV00GkMNQOkiMU0DYxNAGTPStTYep+pvbiZQwiDKs8+e0YOw8yuCeEbM2geNzBOSoItGwr9yy
1xKVySX7+ar0NJrzaTkob7etw4/UZs857t6nBqk6zNoeAM7MVpEYlItHvYkFB9cj/vsL0+NzSm0T
Y79y5XrAsuAUjPbc1qTsJtqHn5uDyh1M250cge0Argm+t2Lhugx9nBpqCnUSTXKRKFlHesoeUJte
/vYUgXpkumq6uLeez34XggzEbdudyntFa5C8Thp57nRD5RSeJiaEzpmSgKHw6yBcjs7VNfcSWQMT
CqtC+2AUJvZpOF0Y52/ZR+aOQdACth2s0vhTqcEcFceuA2GxR7yxrpwpPtswW3h/suz+QIo5dDVs
27zCa8qh5x3+r2XaZqfqRE/5Ri86DxYIUMHrPrKFqTRYmjPKvad/LaIeTosBkd0uAD6dDtZ/eOZC
Oi+1FqQ+x6pPkJdILM7aDPYHph1bNXSlNl8sRZHTykM0ANDDaaeZX0XoFXO18W6/kXDUrZvWFaif
jX8fgzxuoCLvyXRPuhZOZL8JvSbyy/gmjiDiQIedVcHEAIPyPjgrC840nqoyR1gAOB/q/eGm4iYh
M12sDujK5BtNqNUXIrjSwDrLTZuOb4Csp+NphJHRLqwmKaXjvDk9vlsV82VbB3DkOSEmAMRMTmQ8
7nGvmQUYwJw/ZCQiyHyhRnl0dGEQEaIDbP62HIlWUHPPCAzA4Jh3Z9io8Lp1WtSGFiqBl6/wgXlD
pgswThCeK0Z//fci5EDUR4kRs/ZWdGwm7zc4KgBXCY3h6n6Dl2pl6Qe4fHYtHJjKOIXDkaE8P2qY
rzcZxVsiSfP0y1TvvdyhipUXGHu9xtyzi9miRhMgx2S/yqSSUvn0JLZ+z1fp6pVQFIhyUNiXWxuM
kw2gQox7Cva5H+3infgdfQWnV2x5XNtawiG+DjzTz0H2PP26j/DVhnpIk3h8IAt88qjJJhTbl8Vv
IWcBGbY9jWkHatftD01uEVp+cs71GWvxGzAgBiX28vbUzSBQp0PnTGCCC0V+PdV/lsChPzTXFDK9
jAd8OCmAhGGOAhS90D1Ei1PuoIZtUXOx8ZVXUidaUY8SfyUYZMxDXmxvI9TEvFeM9g8KYmsZ6lyV
eEkiVHbmwkClkcMBLtsLv2XiaaZZyzSe+6CcGeXrbVurf8EF2e9nfhtLwN7rGymtdYXNhpn7R+wG
clPaT0Pd2WWwAb2+8NBvgB5y9pbePswwq9fnekvxKeSJ7a1GQ7bC7TwEo1MHreqEvDmDHC0p8+bm
FruATJWuJu/KxfX0jvw6P+ow0k44jyBEld1mP6IA00CqSd8wUptE0nvUpbKV50f12aQWiB4Vv2n5
21tcHcsH4mMfYVi2NPW0Rpxr3JOIzvK1unqALDqKonKw5+cMIx1o07OaiodEIGTek+S93E1Mk18K
2Ow5DN3U4GO+3BfzIKDYPHHxPjOtPcFY3aRjkHSN+E4ypaDpsZcgjtq2ND0dF9+WQZdaXx0+PKDB
NF46hPc8ukB+R3Rbg7i4LZB9WYQJGQ+D0gT0O1uSDL0eFhD8XKiAcqD5y0sLPI0dSM7n8RTGNjey
3RIrDN92KBvWu67VNTuKeVm/0jfj5UvYkZweByA/rrQnDeTeptZ3A71ix6LTpIgvfAnj70DMBp0h
649T2kawYpIqAmBdMcqz/ybfBnpyHcXcgAcNj1lkr939kPNCV7e2I7Dl74RUJ4YGlUFZCMvowksL
ymHYt1JigWyticasIZZWz7UFygiJQoRNz4EJEylYrDF9HBRbBCYhATY/0aeE6mzyRUafbiHcwpUp
7c3yVE/ChtcUK4xoEp0uXm1OJgTM9Uic0IvPf9OJIXJdMxqD0f6OQtEusP3OuX0hLxC86LDJSBk9
Nn/TT6GdDYcoNsPPxaUPGH9smLuWv4QlDz1IZ5FUHkpaSA+WLNLAftFZjbDm1S6JCn/WRxYSxX8C
Qqn4w+Rdb/rwcZctum5cIe45btSiggH5SZ++JUvV+PL5zQOZw2QkkUWB6T2gGxe1Xsxo4G8qjbuW
rD/OsYUcGwgCYi2Ooa6pJz8y2B3YInuS3jsTuL8HgKr3JmE/4LRdRNVEzW3auHYJoVquCb182FOD
eDgDHC9NzsV6faZmVb/OLqCuow079HULtAobNV58D3SyuWukw0hndunukPqI/TAUnS/f9m2zW3af
MRUpYGTMOpxhMgzqLF9g6c4shWNOGrG1w7dGS/32RAUcG1bX/vAddcdYV3gtPYFAdnWvr3Et/VA3
55cg/ujh/lPee4sDBhKpeldufxl8+Rtxv0hJLFpotIQ6KBvRUIL+Kv6d/GyC85prMDx8dgmcO0ng
AuGXWDb7GyohinPxkjy9NJOTRQpXvYsogN+nrml+oqec1kV4DwQOIvyebYuCTIXzwGOrfw3ERjFD
TEQFEQpYZuCE8NwvnPTyf6Wkp/KWHW1qHkgfqwz5IfZJmrxrggYxj/PZJDNYg1iSxdot7MWXBOvP
fRmMGrxwWyu0/mRMSFAFDuBnloPX2z6bDNYh19Iv0kd755LJTwR4dhKK+GHZfj1x/Ec1Hlt9pNP1
7hk+6GE2NC9Dko1u+YuRA6Sa517rVhatSpulJiN357R0nzHg/hvu7rQzqcQXtPwGGE9uSJzp4q7A
hhB2K8FQd+MNL29Y4cg6l4HyBeobtvU9S5wEC0r64bKs9+f1x62hxgifulWa3PPe7L0TxDZmKmIc
8XQA7bOABEPg5V7xzqDiXHuCoEZDiKHhx8mVT7pXMK2GgBx781X77vQZfj2R+l4qfIxJcMLZuxOu
/iWoGgQ8UJN9jqRQwOJv1UaxCHZydk6pcWsuugtNnLjDWTaEDohOoZVk0Fn0icEEVpPfohyKkgHw
iLXc6CkV2gY30NXGMHahU+Wg7Dbx1t/l1NSebqbc33ImRT53pA/nsW4bLJUb3Hd9sgsmhfgOtUrm
iQygI6+Z1RBhG0mTFp+olh5pBm+dOYascz0eYSm2K4Q0RWkWOOPesHqLha7UCXyFE5WqmgDB6lKV
wUivwDXUQn7KlpC3MH5YX77alFnw4V4Pbv5lWMjjUB9/us+vrqOgPBZqW3gecq4Qvcvz3Qyq/KG+
bpQkAbuHjLRJeGaKeYqx5OBfj6z3fLO4FhT6Sw8u2IyKTC/ldK/T8hcgDWgYeSOrkz/KusKDCshH
g9pAAlB2Hpw9eFcBfOJS0j64nfKGndmlk4ZcxtxMQ+uYUvaOZd1vOL5HGv4HaZdiEe23q/agR2en
LGAvvJPMuO13kx6PT0U3IOVAoKIbKjQamrPpyJxABBi+YlmZ309aq4NAR/z4OW+HTs/jmKh8FEEP
9z0oWXY2QuPWYhyZ5lcF4VWMEu655f/GWolyt6b0crW/3Aov27UyHWaUst9v+GJekq1CVMqwapU5
D/hcXGYbo6eKt8vxtgvl0S9RkH+MKU0E/BBYcD3aGNl0i3It0p4VH83WoLiFdGUq3SobNRWTnhGZ
eUYzgUTJmMwUVIkQAj1K472S9dgr5gVjuPvo7JApzsVETBwtarO1p6HpJ5A4zSbjwZZ9naulI6XK
bXh1j/NLzrdKQauExcBNWH+8LA/MJaKT8UVX9dWiwOZLMs/iYkd3l9YjNKxdXJ6m+rXOo1pUcE/z
VZJsRjOiKIdnjA3AYe93XvfcJk2r7QJpBOj/QPnY/3sHDoPEhqrt5w8MSXnJZ0n65+ts+QulDG4P
9k6d9p3z9ZE3b8+JdexFz3C52Imlco90/bnWjKtzvSTAhf+AmOyfH+Jex6P3T29xYLpXos3cmMgi
o65vZYG0dGKV+5NuB+poVTKxetc8NDT6zzc40OWdvsjooulPvK02uWC9D4KuSamMbHv3JpiZECPC
6HlWgJZmUHDYamf+Wha9RKMiTovuE4Id6AQ1aR2LhSWjbKrygncnISWqDlnck9XX22aoMJ5GxwC1
ibsh158usVKNzOTYy8nzOJayGOF+UVK9+14ecz040Kncueu33XSwl4VZN7zpN4xLj6Aer+f+H09P
wd1ub2fh2knxA6T+VkWVAPJYL75QmeTKjpjxzMCHtZ7b2JxqfJatew/6fsAfHpnslKlIobYLx0Td
H8ryfOAvXt94+RcnYnfYWbutaZTkX5Ne8lMooA/o6U2YbVEtU3v3gsU/375Rbo3HXr3ExI+Kotie
spDXzd7JQcHuaqasowZdEMcy/oHkG2oneUPpxIop1DOSIh7f97AUbsX7MattGczJEcN4sCHlj7aF
icCGN7REDPEG8eTbIWLVQ/zNGST6pTQWGbBEKpMiNVo5LifjsfTTO1dwwRHr2vXnQWeuyP6MMqNF
TNh4XlgvjK/totW2H15pOaca85EY5HQ5ZgPZ45FiszReA2owvBJkLtA+LaEXm2fxUuwZ5GVwKwN2
lX4kWdqbWBvE2A1XI0ud+giHcHz6Z8p2eF0P6PPZ7w2PIjWu3+9D9Tk8JS3HzzRjOc8JxM2t9jmi
Z6rdmLs5lGiNI+XpsLE6CJmJrYBKez2mIUZw1RepyE7R56J2dUQp5VpASjN5wXfDNCFxdbQbuI3N
IVHGSilnl+nojWzNKJf5JFVp9NFYUY9bamXaw7xVHMVhlORQxOKf/MNYaNt0ROPx9rOfJw8GT3BK
CehlSYPgySiY3yRn6dYtVAZYW/FXxFKmUbkr5EcLzCje3kUhtEucWeS1uxLGRRrHyK5rzEIVCwNN
2ANt51ViHt3cdTulTSBp7Nx2wtsJo51eG0vGqbZHJkFmZm962hZxItLyQ+/tt9jR8HfY4SPwveo2
0ldVMKfG3iiOULd5sQWVPZLQgeQ2LI8roXBUoy20Vkk5V67NjJa71X334kL/EFo+KUXxmAlOho3o
uaS/lA4xfVoEMC36WxUqSNKPYk0CFNh9R1qO0NuaP1Z5mNVAhxI2TJn4UCSqFGb2qIJ44WmbLf33
uroOfdPKxcMu7lQU3/BgSVuzpi9lrDULsSROl4ToQUogAR1OllvNcIbCSkDWWNFg0/HTLBWoRySK
idp+vRzjBjg70d9dUZwU87ibesew4PsBnDG0SYDvz59OgKJtct2+Mz1Ai6o+RSJ/uC1Jdyt4BWun
3lxxWsgaiIhZMRo97uoErTI+GN3Gix/29fzLZjYtqiWHZ+YeWPYkEkUXZyEg1bADqKpSi+B36nkw
q5/fVhQQ8dvJ2hMw9nnw5F9OMfWsiZsck7Qp1HkbN9lKtXjjQBpCd0ile8psG6Up+IJtcSISzldd
X2dIdt5utk104Wq3/N1eOHBAQUs1H4NoGgx9dz7cK2W5HGGhdgJ/n3Oukpn9fr9UiBcWyUv7pdyT
17dMpcM0rS+d1KtDh2Sxu9xwqV2AgrmvdqrGo0zlxNhO+XK8oGGj3YrDXSUEI37ED8ClX8QeDeBh
H1hBuqT491EIlCY9jSAJCm6XTJAqMl4lAhZ/OrwEJ3WRbG0iNvJdLLDqBTrg/ZbKfRlK0I6nusFp
jbLwogQCZFknwhGLjmhGoHOwGW6PxyZnkidLtyOHIYHawAjt5SclTWVHlFZQ/eNdB2xTf4VPXS2D
V2FApH/aJr7gIxZbuKUGmNi97Bl80q6vj0Ux5T6GJioUbQP3GCiAOKoN3YYt4/BE5hK6Bu9b3zd0
TDlh7vRoZEBDKwgidGR7K4WLZmhB4LKEQMFXbhLa++O5YO5HtjpLHYnVog5W4UHh5TMKfYRERnJ7
SpZoTkFz0qQ+aHgrwXCFwpGEaBhrocGOTscVEjDnIIKO4Xtsu4PtErhIylpPhUlAv3XCi0ucudrC
68tks002WOyAdlxXQ3eOK3EqkU2aLznUAivdbIoNFFgpIR6fLkiIMRaVTqAFwikCzd8wflBNOA5Y
wPrpsLHKbZXJNaiGzeuEidR1PrIEJAXsGVZ/i03TDuzLk+HRns1ZR+WZ8bSw3SdNVlGrOVTIzKY9
K2tqo8WSPB5DYxFizDDiEWwLxxBTTBAXIMf0LEJTwnvOKHggmJ25Z8e4dNyKDlcOYPjiYc8FdKYC
NsPG7N1V/39wzeJSFZnG/Rsf222Ck3WVw3fydAGH9ifq+Pk9khMdYPI0lWhtdDoYIVWTA85KRs+D
ZJ7nqpv+yieMQ+FXIKxgK1fwN0mRzMCh4kJBKk+/qLjTXw+Y92DZwPIR7Cv+SFStAS61oPns06+i
wrO2hmQfja8GYhFYyVRtVqk0niPzCvVvVyhC4/xz46LuyTp7lnT3g5muw0xNVCaf+V/l2bXx6Nk/
/TPuR6RHSxwV4wOilQpbl5VALJUqexbRJvJ69iNFD+drieKR9Dnb05OgiBtGsfeb8l0jZo7+EvS9
uqbYjat50RKYpURQuPxJc3HLzhY7pMJkbeWEtOlLGuL0Hq+FGHEabZy71Qt/u7dMClYA94UlLfYH
9L6hau+zfm5TKmy6TtUeyzb3Sv6qgrrzB4CBCBY2dBn8z7N2wN268p6aXxkY/fMfYUIdilqC7J6y
evVAJEh3lGQjqRgCK+XZic+CaiZ9K9siIi2cqANhdzq2XyAnKFdcAkV8EvxcdSBAtuS+tOSoOoXt
krILL+/KSJJNkPmGSMu3b17+ONjPpeQtUbsqqOBasLQjCyrf9OjyY98MfB/qMkEA+HXpil+Rf/bG
TvOfqWTCiGaJhrMvdth317Wb3bb/2dEtnTYPLdmaP7tmSDrCX6hfnwJfchlLgh6Pi5uSslh3QHfz
g28crfbyDQ3uA/GGj/FLwHeGZsFxD0vmH1iuoAYRoQGDXGlozz3kixLxqFyRucCSQnI/xt4DTvzl
FQYvOKkjkXJHp5qPuB83EafhWMfkV52LP3vyeCVOVQduzD8defFp/KTLG5A9uYF04Y8JoagbAdsS
03lG4nidMEx2dRb3Pfg9Uhkow+6be79nO7nkT2p+qk/SBUMTdzF6AGlXYpUdUJCKR3BBzf5D45+P
Aybs3WtodABIi4VOSt1CBHTK/APFqUH2zIa+aXJnCJ80s8iyBGTW1gf3l+ciO1EsV2cbMg3RJ6CG
XNw8mSE+sJUwyVuRxX7YoW2+XdSIv3EI2UTlD/mVftTMYf7E+e/vg3mX8UjM2NuCJG8L9W/kKX8d
yWu5pRXYG4YSYPPMB0q+CcxrZXQeJEO1QCuLFJS+x9j6krO4Bt4CXhbHEcVff1Kqhcdk5o8PRQx8
HD69qvAUWnTrpP7OZiQOQZfp7HDPQ8oybup7LBzKRvFV86bQ7Q/Rp56dRtZP72e+1WyjOSbGQgxl
Twu2AvKw4ueE6yAnWU637NSdMNIoIEMbfy861qQJ0XawRFz7oMMN778pAn63AAACbBhKLqS8nA0N
zdXkkEoHnqvjoDLLHD36MA53FW4RHUp7pwMafoZlzD1PvWr2TIk0quN4JFo3sEyLnKRRXt5gwwQZ
0ldYR99rmReEJA9wZkXtacX2yxQ2SAXRuo/2sm+807Q26zCef49/7qV/r3vXP5RnfRM3/uca4LzY
uoQTHZKUnrZxAJUsIk6KiA3OTSdff2WEadoeEpAc22soRmPrrel9IKkXEFokziwdFVgiCmUM1nvb
OSzibLuvmIwz3M043PVHtslEZqAA/cwXAjs3MaaJv+0V2b47Q7Pfi00K8DBzqVOwfFJ4vbPhy6Ol
JBiO9yuaFcLPpV/W/Gxb81mvcrOZKn5rT+vwImctGf21wZkBtKewOFCMiiUOqEg1l4lCcqAzI5cY
nuJyXjfS/JtlP0eRfBaP+f+z7F8oMPhSyQYkIU9mnN1E3akkuoNXbfVq00gExWozG+AIBB2aucJl
1G4WzS6ng0KxGZWLMwFV+Nk8fST96U1QaFe9h1qb7P/9ds0D80jc1YmvW4J17X2AhJG0t6lWtSuT
259uBEWnRUvNPrR7tdGKntCErLigIOIfqelmAbGzjp9A76E0QTFR+ystlwZANdqP7yQN2EeL1poW
8ENI1qDblphdaCcVqWdXpNz1qIAbJ/58nF+Lp4TwBKP7bSGZYl6i7dKU11BrIuOdxGoKk0q0JUTT
d5eoHCw0ub2xcjOxS6fYpJVavepOpimI/zMcl4DiyWdbRmJAoadDK6+5Z+X2cd6UJNJ8EidYXXyo
KIkXj+p1fgOm6yXqNVc7ywGWNpFYfAaotOO7OGd0uv6nMZ1uxNCIRgM2enPiX0pvqqEJPyGKbHPG
NEP/AzB0xj4yuDwhLSj2aPP9e+uUuUGU6iO5QPcy8Yr1OodYUWD5WroTGhmvVIIGrJHhruz+tt62
riZ8qNE/A8BUYPPzMFj9dW7JRyrkFMOH4LtyzokdR4XQkpdVlR/SuP7HnCwnOhfthRWZmSObDFmG
4ymyuT6yUvnROfhmg+PBcorplk1ZB5tkVRw2vGITMx0w1brgwihOQcVGd+EQVYKx9GDjCDSNbVLJ
W7NVYHf/dotyf4Qe/CV/KuQ/bq5Z5mikr20vfXvMLsme+1kv4aqzz7lMbeKoG6Oi0lmE8c51Tyzf
ukMoIawCBQ++d73nSb5ahGKikvdvvj9HoFPSYHOcSDFmG1l34Lqo7XswDP+54GJBaTtMZvQf2aZj
C1AzeS40mHzA3zGugF0f8Fn6W6WXS+qfFX6YePbJEUDr+YmtLR0RRomkMiGMfRVAkdpXrRIPBsKk
p9YISAVcqhnd+L3s+dsLk3CXhqP3QphL7+RIPnIic/lz3hWFcl9fidNl5CsSZsPUlOsZux7Sy3xO
XAzdjhiu4CqU8AnmkmXflvbXr82Iw5ssQcyTEbxQb4nyDnmUH+uvoq41n2/UnEoW+gap9eFeb6Cb
wgomtVxrs4mP/1Ga742mkYjyQzli79tn6xauwyGtSJWDjqnjG9R9+JukNcHh31pEHuhH7IgEm3hh
tcGB7IuNHANsFba+layrrzGwJmY79Af7DzY3sNfZ7idpT3LSz7iwi2Q5eu3sm1heRMXhWpNBlGGA
x/SHmBDWz62CIFZdPd2loKryI+E+Ib5qNyubwHGgTBgxgHwwDN/39EnAUvRQFKBN4YCYExfVkziF
QROIXpgRKcdpSTQzPGApmkfjo2eFs/h7A8zkuJa+yNBNuo9qa+hok1IdvKipz427qPsX4FHOxtro
6YJfOSjLCELk1bXtyZwObJkNdzWurcjHUfhC79zYH/VlHwysPUZT9TxGpxoHn16euuOitDaf174z
4pxwskxbDKcHtsz551aPCOfCGpX5/FHBg3nJpbHdSRKbeLYjVANXWDmQSFtSdO6NUQ3zOxfT0thV
xrcbMtevYWH0dT098DNAOwVndA8cNNL/Qc7OsqVvmFnj4bYnAoAnq04U2bAsQrmbaEt67qczlaKA
KXTjT+PN23gHQingrG7cErLfvSF6s4jTo7HGZTn9lFTwPQTgTBt+gv0L6mdRwmA2wxibk22pnCF9
SE1n3djbAkwxLLW1ATQXhX9s+7x7osd5CFcHBwyWHV5KmYdF6tXCbxSFTloNpXDhq1gzhLtSiZo5
62C+rhwiPKcfccjtH7vdG7XeXGjUaJQfNNwmP5X8UUJQ2qbM+u17mE91vVxb8gETvbMfPo58jQjr
9sa3nb5Z6uVO0bjuUm6ZsM87gzlBMbf/IHpR20PRZWVw0pLINpBdwG7fnQtbReRhpoQ7pzPfmPwI
8s2CFOJGULZQijWtQczvsz0WD9ykcjJyCWsqQNCKfcfAQV0dx1zX/ojxjMU4JwBibgGhrIx5AfAk
k7wbfAgnXy8L0fmsh+82UgfKSWfSb79yt+a5dVkdDrljVBb1b/B2SR6rIYW7R8XiPJH//n7KFQYg
JBpCzggkoN475uW/TbJdUtCZmXBgFIKMJyk0+9JIcyeOPHS7W1Fiagg3IcL4vWeEIogD5kyAj76q
VnNIE9LtVhS11NgMHE+P2W0JfbhQNt7xmEYIw7rec+1ElzNRQw5w0YOuRWbPEYSfYv4ObQvs8cpB
+WRo7bLMYvY+GAupY+nfcc37rgIB7uRRepMshjvIhQTN9CVMTTGv5kcpYTAiiTaPFFK/WRAFHUeL
GoCrQhn/Ox3duZJEhLSRRaVFLGzC2WmQsl2ayjqLmovgI0on9LfqRktxh5MqXGuETtDZ2juDUIBT
ju5pnzLXoo20vc+d8bWmtV/1Hsj65b3mmmfjgyVA8WgOW3B8pT94C+2m+L0+7I5MFQATEbwT9yAh
DIIh6jPZmAdV7gK4z5eRGdQwMGWlundyZtLxLqif+T16Bcrde/vYF/Wrh7+NBJkCoJmUBgvDcNu6
c3YdILqUnB4W53mqaMRCJyQyj1HUyIwDVpc26ukmDqhJQ2LxaNsdBh0FkR9PeenGNK4FnEXquRWK
StkySrN0U0cbQSCLQPlNLtBcQl0ChP9NtXeq+MSay5bl8SP2jDCVtSe3NvPPK0GvTYmb5HzvWnmk
lrOH3vu63QnegNm07BNKUMdA7lKpLAloKldlyjwEUGzufSMY5l7oKHNe0IcekDjrEy3D4x0+gQkZ
TXKx376lH91tpkQNYJElExM7Hib5jYLozJL4gfVJ6ggzfZeusLGlAzh0mwj6JqXoyk4pDvk4GLgo
ajeFWP7nWXr2d4RS7Nrfug29LuBs0//kI3gXSEtIM7Wlta9GLsBje7Ep5TqfaYRpQUSaqwf5Gfom
pX/tMVRhyu1fdc4Zp8VmFpi2puaK9+rnoW/metkVmH1sJ8Y31QQkFWNfBzP5b9ov24TOzva0k5GU
bZj+Q08zXJhHOLsZkRFfAoVPN+ZZd09L9VMVGYW0ao4I+w4T1/o3z15RceLI74CdbsXoQOt6Y22J
lAXX69EfHVD2S8/thlyMWu9FfPRfaSzLbqTw2/jj8dep/g+J+2SXkiz3sjhf/09NsV2cvlLCwqfs
kIyjOLl63k2Xt6yGa/Cc1DjaJ1oOL/D+TfTjQzV3vpd8+XslI42Xfvg5npGAdUReOnpuizdyoKcP
z7mjRomNxCFui0/CgOVKWHPFGEwhlL8GQ3unT9euPO7hiwXr+dzb5bwImGKp85zlpko+UYJwn/Jz
7/hagd1/YjU4V9UNo9toTGv/QqxDO5Gm6tw1JDzShzaJpDc5ndxGNqSxjYNzdTxGUkE36qAHE9Ze
io70rzZlvlnD5+RThqK63GCL4dyewP1upmEs+Rg5MrYywZ2KuGmrRB+1L2g5J6Wk0SvdQZPzoQCY
0k3V6xaT9XjVpzpn/R41mRunm6/xbgiJCzNut5QnbmYGAW7iEAoo4q0Ub/Xzf+UQv0ffXmay5oga
WjygRRQ2dfZF4fm9huxEsLOYQ8l5N1aB/5gUrJplNGPY/F3TeBzLQcK5Bd+OQNu7XnD0TZQkMo4/
/2a5dhqwoYYFDDMugsLYiBqSJhsrOHxrMg1miVFOxks4iH+X20lJEfULPAKxiQ8xU94wW84Y4wzW
b4/rxyJX2tzhPtRFgoer1ah5VVd85OPSagzPGObs8/CqvrXPAw161YiHNqIksidPwiMrjffGiDXX
lgCXp9LrvUnBoz+8KBA1+uI7prCWLmJ5YphdljwVaOdWhXKxpu6aMBjTQjWEQbsNNBJ+gX8t/1SI
gpqalMAQRrbji+eqBbLalKek/27BVI/lvTsA3KUxtJqkVayeR0bh1Mh/DXzQVOEYN0LzL9rR765C
5SmsWHSCP5CnfLFWUBd0YoTkonieIBhLmsf482/ttR3rxdh2jV4WAaf8t5RCH/lfzjrbWeE/6BFT
OBWIz89Z0JQkuIExJ4JPpqV2+9R0rB62xWuUrj3JWGYDV7dj02EKYjr+wy2DFaVIXejZjbdi5g1F
I7biOBAoVewDN/EXpoMi+64yxkF6hG/R8i2HHP1LIm3eTtsDU1sCrNncZhuLMnR+5wfmbyRWqKZ5
6FwHSprvRslEkXnecvLTsvt1Uewtdm22QPKNireDHlzRQ4/cexFxfiZcdtF+pMvwYmD2JDuQWP8W
X/VPgm9nnIuX++eokH3fRcLv2S2U9Wi9AbvGqsAzfe7vZ6EDd86N0VFN3ZBkz9XeoxAqG86Px26O
LMRaZauzuX22eHGbFvO0roesTyQNsxC5cVwRmd09HMWpAshdiGGqNzpjKNSp28NEu1GQZ1v59WGF
En9iLZZ4nC2JIYBLoPOncJMVpj2pGYmNf0kur0GEIny7veTC3ZzjmMSGhFEEWmT8lhHrX3AMWnYM
anOoTlL/ezNfKQDVpB99b3TwI51uQpyumUMyMvuQ64keIn8B0YU80l9e31qYYj/VG3rgBMGpos2V
DNc0cfs5YUZbiTY8+R6DSykIz9C+k/7sEzUH77OaHRj94X9WZ1fv7NJzw1S/GVqdiY4J0mWkaEtZ
RBiw/MJ3886mJsyuZwtmTr5mz+uu/y3CU06Eyd6Gs9HZHqQCRuKaJaacbyV2XSClXZRwqC5dA9Vv
FimeD1oXesXi2bEYDN7qEyxxg3JagI41TxF9RvEzVVUigQaG99zTLv1M33y/XPOTRsCsIKgO95zj
DgId0WWbTdDEapD/spd0j3o09g92SSQYCQD4UmIlRd1aF8nGtU0Pl0duTW/a5Bzt4Z9WmitTNHQP
4RWdhwYtaGGG3Bb00kjue+55Qt/VGyDXbqfQ81P4Hg9nOqCDWOiRwDP8bZX1OTmilVVaK02HGYGn
oF0dAphee/x5E2be2pHFL4xXwem4m7odHRkRpXIc9PgLPsWcPexDRAsztITRL2IHfyS+3s7MkNfO
X3oYB0XAZTc9ynDEMvhLthYIWt7xDK12bIXJ6JIHhrBbdkuP67IV2zzZFamRMjoIXAEM75KFruO3
0kvJ/om53w4XXVLU3ZKFnkdGYJZrSk0CY81zP+TTXsoSOhQF8hMz5WTEYgJm/SF/8d6GRXiVn6+c
WFmzZLxS7lxXHn0exEj79eF4yIu+hIFOqAcrgRkU2sZ+YuahhzXpgxJ9CjXQoTVbwjyMGMEXzhYA
UnLRYqvwwmtOKy+joKCpOYhzTRzNZtK0XkmB+xmZxhsEClJ3FX8g7RhAZcMV7ESznoTzv2LFgzKB
p0XH/71WM0IReQ/HoNJP8EEAcokhMKwdoFQH3BsMi0RYo/+eZL27vBZALoeFAVNMkkTlbidV8NL9
TazeEtFPjAeBP4YYm8bu59jP3GsFIKc4BHnmtW/DP3T5bYxwEc7FEJYjU/eo2mju6JXnvxxL7HKx
pnPvgXVkb6yuebJT+xag8d3a+6lJOZLOlpQc+UzmDyerxi0ELjaWkYC8ahtObYcRUUXCGadRcsDf
sOPiRQLRSlMLqFC8zypvjW3V73c/lxxGPOMCpFHUXxHEw7LblM+xLefwO6LA3kpGquwd0W920uy1
pCznNKw6javCyAI1W3qKQycLjrYl8ANft+BbsRUvF5r04XNwWy/2RxQ3QzqkY82FhqoDHUAo4o5X
yzbR1c1uovPVf/85Uuh4dcA5fiQ9BcNBXYRZg9YpINnrwRGon/1ApLLT/K0MMHVwlIwOTNTkrBus
aWHyLjuBl8aTm7iaeadq6n1rXcyW6WyfZN/6/X1x9VounfaS/M32BGldwjRQU0TRSZCvqYVmvASy
Sv7fxyHIpJ+vb3QR2RHQLnsog0bt/FfvwN0FO8pujF5f2xHdUVJVXCQjYCyXbo9WhXq5LirmdrZZ
OYBWhixX36hO8WvMfGk+Pq1CtfKHAk/uqMO5RoZp9UK44ylWqm8bAqF1GjZXBNBs2ixsEPIjayqt
7LQUhugN3K5Cib07cGUrKc64YYtfvY+mkNjCQ37VKL7MWeqdKBPnGW74I8kRKWHHtDI1rmJNU8q0
QaYQe/L7fycUWD/D50KbF3KmSBf42YnASuTZWU2hGgX0/DQDVHUsIWuDzh9S9feeU1bLTpZsRbXz
olfKJQJ+8aOPYf02AF7zcMUjev2nFVBDd1Liynqx2k6mklnuflakldrj5+R9bW1ys6Vg1ef2i7ob
ommSiLOusa2bDE6J4S6J1n7sD7p+KfEk+6IOcJwJlsXQRZe2Z/LImT+ArppuORdytE4rpkBp+TuY
n2PSVM5TLZQIOh6Wz8UDbWp/Xv1avdC6YjztS8/L7Xzw0ssyUq5HbKa6pUHlQ2mEmbGhktfovDOX
5xnfn/aDQxAwAXSGqC90UiJcmwO54JJweqeKn2LW1Mh1duQJKbyb7ZOBtY+hUMZttaQof/3fkHpv
6GjTGBqRcYz8eoGPVb3uMy+PC5RUawxBlM725vQYrsUyQWGWRgyc2i7XunjN78zUDhcB38KyghRf
Kb0suOmjS6jiXPQbtjaDh9zRsL9bwdbBFTdqYZ59sXR4JRoDHIMxvy4QpBaOOvBOadzq4SVNvuLo
TTd42PXuSKCVvPp/CloLqY81hSR6diwWEZWxPls16PA4ZAlHktppsOPyL0D6uL0InbraRbDX45xW
dSftO2+YmhHCKQG3w/QX0cj11QRiylliWTWaVlYmEsbmrwWSq8WQOTeJA2sXIvqoVXcuypJMfeDA
nbEoYhNmfRrcBRZF2gxJEkLUbXzEY+wFmWD1TMjF3IwlcYHGJQqVSEgsaJAoIFicnPX12q2AYTVs
qENsFv/3OHCwNraW5N3Jjg5SUnf8hr34q3PZCiKEz6Yww2vLFg2ANm1SScjBmPM9WNptbfQCtDY0
qmcv6VVSs2AyOyle3z5Eb6mKxntgUa9nLfsV9dwGg976NfGx5EmEa4oK/ANEAqG+GjEqemxVtfRq
mcZQbzc2Ttv5MlMhZr+hVmdESs0WJurltnsOwExbyD1OrRBr15wwKGhRW2Vt+g3d4jvJYXDlhej6
L1ZCOfxFluVDaxuXmC0YMB2rFc9L+/APqA9ZIjrPb2AAuIoQS6Rf+anFNAoWDyL20AIVuOwwT4d2
thYYylMFAuPstkwEP90x0MEyKrG4mOPhI/N8U3latv5ZZEUEA5sCujXZV6WCFKi82LPetbvxmlE/
hUag9jrxrjHCHAvxxm85fClaQj8Gs5zrwFNCESqDPR/zs72hGKzKVyHJY9lPmw/pnxrG2XNQGhQn
04qgh01WpxaCyli5r0/UcB8aUd8i66jESGOTx4VJK/38BqZp9YgYenJBAvfM5MQiBb0GQRn4kzZ8
JU5Gn2qxxEfWJ6vpgZ1b83t0cP96rjmy3rPt3bvtTeflfP8jENdcUVOhxkNnrIzPxXJISCfz69ms
TzHAWRpULMGjttBCxSpoDnjkmHIo5Gj2rTfcCMLgC+O6CjDyXeRefqCMWTpx7XrIPiW/nl56LJRD
cKaM/yVtU2XPjLkGsBIGBdLSWEi/v77QF1JUgD085CE/J3xub685WvSuaWGlpjNfllqFehn6HgTs
qYnw/97b9I6gQ0IOnUgGCkfgpb6aJETgGpumWoPUL/bBo8UAM6ow7+OQ9MGIABYMsDqxiUC+LuKR
F7HyJWULRMsNr8d50xQ3IqVe2yVmGgUeUe1OoBm/Q4g8Knl8aw57bHrnShijd79Z5g6jFVv9LOdP
RDfVzvNTe+/dluVgu49N+1KiqLR6JAebEUg2HfkYQfMKFWKKYsb3nRDSdvrM2ST2eWHtB+XW+MZv
rcLS37VcfD7TS8ddo2NPt+tMsErV/KdtF9T9xzwwwHLP0Wh+Nte4wcRs7LbY4bBbT43w0DpNQgM/
urDh2yD4mTEmp7LMhlLRAhxMwIaEezanMhwHNpUfrcuKEd+42R5+d4XiTnrKiECnk4pKUmJeUZIo
xuv0/nFw7jkZPPT3l4giJMLeiX4pii6IWuzgkDjltnLgKeYSVA14lanGD4yTrFtdd2b9MH9J0QOq
VEDDbyIqSP34xH3xSYq06jyXTpCXytc5sMTuHkN42xFeQUhtLuucAoYriJJpBOa65ULhsKnIasvc
h1z2VKGG1gmmjzDvMsDdboKrvVJhBBH0nlHYi4zstspVQhA+4vLejGF+5TKqydhWbiSwBArcxTRr
Q+HoZ4FM0wqwnwSdRS5DHmCbqxAt86Pb4oZO0S1yuELX4EmlCZ/+a74w3onGAbN3lB7491NpkEgF
EILDNe6DIWfHYoMOriOBOTRlZ9MQLpGVLS+9LrKRyHUYhGs4ER0ZEvZL7Id01uCht97ycM67DJu6
X4AVs+0YNp4SDCCnXtHntTNMARnm6jkp7XnviMsb9JB1GgUFi24m/o8E6c+kfNG79KHsfyzmGUvK
vqKkqut7pYvldK8eOIXtXdzL+/bxbqV+9jjeCNJxVlJ0WRlD84TCtUg5GgPXMOh4B0Rc82DvZdRQ
eiPNAGmTgEmcwBPrlPl7p0DwKtyYLg3ajY+3m4lijV6XKPPNlyBPhCgdly7hAcevniIa+8Qus1ak
2WqItbWl6x3B/1d+8TYp/kaCFYeOKCYY1IBq5wda8N0HaH+Azl0ca/oQu7fqUYHS/Cy/T65DJR+R
j7JlkGm5drzlNjebGnuLspijlCW+4uiTTSor7CNnMmthNL4R1FJCB+L+fnBu8vTCm36NwJ+wQzU5
hOqK4fuGCJT3cuRrd7Wpf3oPNooCK0FB/e9NspRJdewkqSs1qjZg34EmLQSiwL/ijwLPWjT7BhRt
Rmd9l61hHb/yaGQML6vrY5ihxqS5VfO7N/pixRMID1p1R5wvutS4U3b8cr8I3knjmSAcJtRlb9Df
CE3x3Aj7o3qdvuMTj2DqED9nkVpcAvlROFk54n9ATlDkrVFnvmXbPox9a2NCr8FFbMdDghXbPPje
livy51ytmuWkDxfE+aKhxwJ9Y+Po+Ry0+ID1pTlR/C41ixJzAO2b7kVHBe/UdGO2J78rO6aK5rRF
E6/uTIaha/b0Iu3wgntFZPU6yN9kgkk49eILBVs336BmMtC4gfva9LGz/V8bNFJn1GP+7OBbmBke
UYXlQNXcDLckIbIfq66ADBinwGCTHSZBomSxPpQC1N2QZlzTWsuc+MiisesoI+pk+Op3s0oXSJ0D
YCOreJe9SQkANygoc8Ml0h7/68klUXCj8ElmiKd1/KsmG4kWpZKmuvLXw8SGXenvqutweK+Az5r4
QG7bYqB/sUNbNmqzPV+ZQb4Muz7pLp4uwgcGYgApq9HGVWfnflnTYlynWzBS6oBYss+xmMURSb84
PPf7TGgVV9mw6FZjD5X8bt9tG+bZu+wp3IQLZfH3mMTKQpw0fntypQeXdqDa8M+EvMY/6QuaMwk4
Ahn/p1I6OD7R+ZWLepyRlibQHLPYYpqt0abDjp5cacnTLLeS51ouSAcAA21p43eHdV3z70VWnaS8
HcaCyNDUQLYg44GSSXMyqxIHMT0TYO/1+j8uLrAxmAywCsAZGcP7KXBlxz5nkJmAEeQmiKAiK2Yy
3i0cym+F3Xyg7PqxW3mVLFqnuvsMXjUYxBfY/KUgHBgzXo29T/+U4UEexzQvZmFB50yljIp8gKHX
yyG1CSyu3c83FBf8SLDLR0j61KGaHbilhxiV13UekWXgW+3PLkICdiANRN6EZjM/YtQWX5KJYpeu
8LuKf0/h6P4qDW//onTmPOEGFKS76dihypt2IlFJKNfrxd73wXdGIsCkG8fdSX4Melic+gWKoj7o
82l0VRfVJlBw81s1vr9kEYm7qLMiTXex2VUxpixI7kovFIJZUItni4odoplckj3BNCjgr0wtlJP0
y2rQmA4Zw/yWlI2YgKtU+CdjGn2rNGEDVxyOvO6rj1pwYVqwC7A/jM5ipkXA5zoVLFDubmWatXLl
4RzeAE1Knp+tH3GfN15CQOCtu10Nj2gIGY6tKABpMjiiduJSWYH20E9M4WfSArvoJBnMg92LPx9N
XEpFNIjJT+And9ckD76Qnb0M8wlOr6dkQBT6W+wF+qEGvrEj59FBYnXZzEBBJxL/aFnebdEoEi/v
P/aZfshrmjFLC659Jg8HgY+ZU0+T8USMMhDlXj+jvdJvPpqynzhGwlS/z1+4WXA9yxuQVB3aAtDZ
hgej7XQc0Ut7fIbKw1XYu1qiIPkaPPRzp18v/DfhO43IOyokI/Rb1TNO3KLJvEKjVWsXEfP5XI5D
wpgNLUMmUbkYBQuhsJU97+wOYdGPY/WTAnoMQ8zRxb6zeZ2pf796Opa4Q8iaO8/heyvJLhSCsyVr
ijRzBNz0IvDM5wj39vDAKGZZXiRjJxyJIdwRKKCZieQM6itO4Y3FHWwRPJr1zlDq6FdqT1/gXahC
+6BJqgRMpwrPjucNn6gj44E/diTUc9oqubmqdtyO7/H6GpcjyjXmPX10lxT9xadYPZLvBJ8XGWCs
yIyAZnTPOYsirOc0c4JMSH7HhBXD8l+wwoD38DGpSZmHxBc5zHQD2N5ejFox9Yha/L6pye2iucf8
ZGZ+Y5Exbut/38Kji21KEGMsUEa0+tFWtEtY5MBoEDVLQZU/CtTQkLDtuBjFPEgR9wbgeggNrB9s
jnPf96PYf8DDmJIjOFuwhlCtuHrOpiXqdSUMkBAkH9PdCphQwdVijtNPKc8lEuDvD9JMoMlAo7Px
dUdPp4dRoDi0PNqTvKo0xdpvXjGbzBHz6a2Fuv5SrpLe9M1lwbThxIrqp7cjkRkhmHKFsIXnPD9l
AD9Xr9zo34XiQvdw+fi+XyKXf1WBUiZb2R5zhOiix2d1C01IlJb3xAShxzFgrjsiey4a3T0REkxS
0jC5psDa1MQKBDc1cNO1k/aF85jVvFOtdUa4oA+zT2AJQtHoUnUf4fFj58qkg6SUd0sjn+zIFyPe
EDCLndjmliNMmQ3OM8905d4cLwWvhUBnhlMe8T70hvezj4mYOhxzZK7bPjvR/kNpKXneX0HoOrQf
XtL+dO9dm7WGF1uyDICDlzW8P265g33dFUUQ3LfbtXHiFIUfTf2M5zcCLCbDL5r7BFwiGMKM+pk2
ItfyxUZo3u2xxktUDKBn3rpjnicqNuTGxbzOMY5YZ60v8wRJzTcN76P51I/yEZ2X7Glnlu6urRvP
0Vw5M4ZR8RYXYTRjtuWR+9tCCYrxd4YFkA3IxcYjqHY6YLe1Bo1L8CBdeZyUVERN7RWAIC1lTYSE
g8WcDJ6CzLaWQ06fX33CsyigCb8cLG/M21dkPGUlP+vDWu17SAfRWQDYyw2fECv//ClwZ+beNjK4
gNz4cATWw5O+KaM9bGVR1PRsmXM+gD4iGYfynBxFIG3UXV6W41MFiNNQG2QJuX9SeKKlCw99ZfRd
l/e/6RlbVNg2HCJRaTCMneJ6kkgPOY3DiM02PlQnM9T+6VJbVreYkjaB4TlFV/m9wxChEQB/T7ST
llnRjBLwkQUCdKpM7Tki/WZjGEMRcJv9ou7KO7FsLQg2MzTUjx/GOVT1H3PaBOkAQ0EgaL/IH2PP
WdiKL0a5y341Czv4xjlO6Tp51f/zsksEE3uXYdS7fbzsLIhIUjVmz2rRikaRjAWOVF0AJyIKaBgK
UNE5HLxhsNp/x+UH6RgqOiTWnLtoPeRUbL61LhozagSmuRhAeK2UCRayGMfkodx8I64vWTmxCEjk
4sa5BkSjwAQADnT3AeaQwFDTZIMPKIaABRlq3z/SKrs8jhtaIFp8shG6qni5pX8xYpsseuxrB/7T
kGHBo0WxaYKQQNPRvuPSodQ2Cgr+OpSHv/B+yd1YOLmd42oywmkbMEt2k7dJd1wf30ULFqXNJeDc
ItYAybO2q4uxq58wpRfrhIzP+nvLcRJA7ryy/s9mcf+2bXbJfKDmpRwVhf60fgNXKwXvJ+Q5ueV8
W/zD/ewQNS3Q10rZYUpnLv93qSqpi62LwXlQgsK/Emq7QGxzStTZOMo2o9dloqRwq7fhKwm9p5nQ
Ug4cJvyovgMAYpBkguzJ/ZfL40shmLFzKBeK9vGchTtG64d0Vmn3VmFwn7pES6S/DnipujjJJM8L
RjjU3kSW57J7F2eljkIHLhBOHFjCb9fy4j0n2487RXL5slPnE6cVbnnAstn9m6WzUuJjCN5yqPIt
XExilt937slYEc2MpuwJUl25VXY1V5hMnUdQrDvaeEXdL4LGDw2fhM+WozdY/wfa+yiTK4CCqNgr
09r42ds3F30Y+MWi6g9EBJGTZhYZsL0tgNMArqmP9Hc03+FebprqSTah+YYQtvFsJVmHj/0ETjrM
kE9+2Lm5p4n42j84wdVB2ZA/W0NHSDpz6hr+Gm8RRMGTOs1S+TtWk0mqlAa6SM4DpKT8Q3wbshyr
UxWlWmMhUREVRNUceN43ZGd/n9FZrUVmC7VQckUrQzHmYrH28mWAyC01A55EC5ua5le4SH5FcXhG
VgAapN4Rla2KM/GeCoBzl87Ya/++h5mPxdK0jSRnf77CYP5W8yS+0XuZzkW3mQ3s+v2TaICOhwJ5
Q7aBFSU02U/KwgROY1+6SkBPXV8BzXpjjiO2+6P6QGVJjAlemL51wJ4zHglch9WiLUEVbGWzfr/K
iI4l8qa1fDlYfcuock2pxl36b7zHopWAkxpf3ysSXODisICTCb30Pr6XhCqHshAiwv3HOlxfSwgg
+IAVvFOrff2SfQNesxggU/D65x0P3Bw4oCG/1/eiSr6EcY8Mu+5wfLF+seEtvfWaZTaJNFN0G46g
gmAErLuSyJGh40ZgVA8WHs+1KqjxoNGlYZfy3+9l+ekWuzg0JZyRW8YZ/o+hdw8AkLyWVY1JT3p1
UjBSRxiBi4sJ1f5e2d77p+1v4rocXp1KF5TBsB3K1PYvGpuvxefjMQh3Z4oIp5ounjPbCc5ZsTXq
wy/gRnMj7S9Wu1VMpSNQaJTsfiAKv/4L0QqL0kmQTq8NpceL6x7n7PpsO+4Aigj37UHBgmFNfC6X
N6QNIxxmiRQM67gM+kn4Q3/D6Hk5pJykjw0+IfTvzeGAxYPTFy0ss8vl/rTVSGdLEy5NOUAuncmw
8XZZX/pK7/7gKZI7lDjXS6ooj+mwJ848KpfptdagQmHaKnwrrTr/9J7bmfxRW+flMiz45dvIY9Jb
K/zouHThGIiapicZW3vBTWLvsAIs4X9WPSEdQ4bqFwN68pv2SBPGCbYyhO/Xb5y6U2P1MpX0l0a3
NxD32JSeLAi6R3n+MgN2Wpvkc4F+DTBE6K7RTvA9g6p1MGHj5vX425M+CsjUeEkacEicHdpP2/K8
cIRe0GKTdU0WeWjhd/6z87xvu3tmB1+eeSJ8m/yukxNDLYW0qjH3lkmk42aN5iqVnE6ZTsgtsnQa
N0yV9S6FJ58uCQlFXza7JOVsc24+6VE8g1MKDq7WGF+AxXSf0KHfapDhVknEOuXfnA+xud+7FR0b
ye2Ws5m3La3D4QY992F+ANvfCYv/Nd96kN08GvgBLoXXHO4/IEoC5PRgPTvIwIoa/ZaCdP0fONyh
aHBgq0klqTv/lAYyXapeseNyM+eWaQhpuhusMJwr9GDSpip9Ae4VgM5woAAQEcgBhoEzzhaS8V66
wP8QHP0EMzKyrxqZyPSr8prA+kAYJYMa/jtEGupjAbU+pP5ydH2mDfelBjwfrZsen1NISzBGC7hp
m0ZnruHrmxmI2M6fQXWEzgFxPNRHld6OfDkpDyvkmEaQFlaaKYogFBO0SleRv1QzIPGawqT0tQje
dYt6zmMVOMflsq7qCBDDgMwcafC/6uwQDYQwbUanZws8ulGTshyKYVB6tNMqdJurAPNSm5RBknfJ
apdgx6VZ9gEJ2JwtUIq8hz+dvlQAJ8YK7bAlfLxUkLxFGqHao+hhDueroqe8tw/epgEdPUa1ke6T
RRZmdAE9YKRo7Bq8PDXXXrURWSH9MeHGDgqYZ11nJIPMnwkZaNfu6oLv8WIESUu6QlTSj/GDIepT
E6AAv5XlZh8ZDn0UhHVcLuH/BwvqLsSLZqHFbdDVzoJU4DLyNzpz64/ohbdnkwXdw+KArp/4E2Ui
Ywp+E+1u36mC4XbgPrnVm2ZF9jWk352QmsPCAKSVezj6oVClHPt5++OZVTfy0BBpQlhj3ulyRMzj
mpOrG8+kbkcTvgfZZQt+DEhCzHAvuLVWCZ8FFIHC0kSsNCii2bS0xGtpVoDzFLOEWj6QdbQPxinn
L+L9Wp+mTY+H7wlGDOVWIvrjvnZlJcr1p3QbZbPspbmzLQoibHFzvURCODraU/Di3z1ebfd+bauZ
PjO2/cIJwhJWWo+YtsvYnox7OphapkqyScJ+nC8FBtvQ/HVUeKw+zMh4FcJFyXMldoTyhcmqFv77
nKSCGlmKXAWfmEgQuvKPlvtWkBKHUjtAf7lQtmTFguLEjR9/XFeE1DZSb6/Z1AvViP0cERC0Uwh9
0DmjMeR3sflcwX0V5iput1TOf26oDuWlp1RHgcHRzxiSXIlK3UlbjN9LH2qV3Xp0MC/pi1LSgSc+
hepJWKUsd780+QE0+CgRDemC7L1Ofege5VTI/h/mujTMKelZ3N3i73x/2IulD3/hny9CS0aMGShE
ngSUpfmnnmJKebgDTRafKDpiPgsdpO9UoT5KcF4v5TPUSO9k593zamzkQKLlW1ufUPoRzh0AuHdU
2pWAIHyKGzjJX4XnWMAEalnEOYCFX9aa+OMZ88m+WJpsr06Osf/1MYNUkiUV55Awy0pvszdL2NQh
vlC3ZYMgol0SXlKTcZsp2c4Vum086jS3tVtU0hQTVFsa8FetgVnNBaOxy0eHtZ7COtDLgnCCLeeg
Z3K8jKgOdJU2TKXTkA0EAuYcd35c+cFAnKIrzHL0MBbA3NVpBsf+xiIsc4a0xc4glDALjpNjeJbT
WjDiPPORjunaBYLEyYDbPcLyJXn8Y44pzyMOtcAY/q/o/VhvQv5zqiVInezBuIBE5gIwXbpgs1yu
8nNyr4dq/9BZwNTX5vGiQ8Eb9JlLHC3QQxxfSylVX2/aluhBQZpugOOxw7j30Zgea0jYu9w2i7Nq
vgOFJmsYNKzYqZWNFFK3pw464cBawipdMnYs2+semX8txl0ezfED6MfyXVtfBdbqPkQhzCljAhcg
NnwIl8s17GHxGt4jBGLpI3DDz02cGG4TrkVlLAXqb69/x/fmrA6Js8dZJfE0Z1d2LGOf7rJPnntl
dXvDjNgpb8deaqu2VlNCKau+6BMFMHSvavMsFGLGZEFOJT8yWkJq007ypgWO/BQSe3sbGp4MWRQd
/1+NW4Z8qr16Y0ij7Y/XL5FprUbEGEySG6pNgEnBCvqeDU/tagr6tepbGTiOvAO3uTTquv2SDAWu
lhOX5+6k0ygmrB8T4uy8Yw/Kx+7g4SNeArS9wes/aJQmt4uOjnUCvWiwB6DYcTM9fuiK6dZuFW9r
39wYq8XDCg7KafcBkElg8JROmqtp9pwUS9fE8TLz92YLHpHwjqRF1f6GMHhMx/o0Z6t9yjl5cJvY
PERjkFrGISBzj/Q+O8O/EYkg4jLHGftYqIAfyrmgfywvDP5wqOVMsHEQNjq5LEV2a8RoTZW8cKOm
B/4iOoQukLEqiJ7i3Pl+hXI+KJqMLRfiXlB/iXqcBVL2i9PbDGg9BpMhumxLmF0w4C1U3Vsm3Maa
QB9qlfeLt2gpRIvWG33yzjnhMIEEczn+yk2J+ne9ONWgXRiaXP1d/zOBv2NCp9lcBxG/M0TSaO5w
D/y2sOzcGy/VE0BvCgLoGwBp4cnZgBf4o6vXoVacmASSzrgg17lO7fGI1X6HkUsDPdkVx2p0F7tu
/kCABHLTEofiFVzZIJlYoIJU5FYO+LGuF1BM331haftNT30f0EycRJsmUgpA/V0knpmnu0ak02ZR
dT3Ik3h6plvaLX3dUvmMwHHaiiqwGv6lJX1d0GWu/u/em/U1iV7LUEGmrnjCi9stSO16/PjtUOXo
CKBrc60qF68poie7dwyqeFUkb8fBtAsYGZ4ix/OT2s0xEau43O8h60LpViLYTofhGyhIuBGmwQcl
wLFFK89uyaMr1JZ5YC5TxFQEMJz2RwvEEtJqe2xEvBcwO/v775im3zSWcdiiydOuqrUofqnVkyQo
egwIpKHQGJv7EQKYDvCwTF2lkin+C0q0omAAmllrQZf/fMePWjDkkBTJlWeoE82ZdjpgLVbd/BbZ
nQK0XSFPkNjiAlnK9lnRRZAPokLO4BdKmVjxfMufsUxJnXA0qjLSAqanlym1SMvl+P1nUzwNrp+P
3AKF8rNbmU4+qochMe4KhySNJ7XQSH96jBwutllGuIkSZADQSL01Rq3/3bxjNJQ4VchjyzVzAIbg
cMMhVIl3QVQtreo1FEOf1Fd34/Fu9cAuu+Ia2GxVuJli+fglqssUdydR16jgIcjsZ/d+NowhNAW3
Zaxqk0LQsoDvviGlP3inOw53HJ7QKU7pVbI+GYzfgjSABbwZAK7hr45u3KXTFhC9qLGe20yOTOhU
tRi21c8DMjIcMr2Yks0jBjCrPw7lBjsStJtSzE5Y+AJiyhFP+Q+zWzV1IR9q6r6dT9PingANCdE8
kVcKL6WDo9Bfzv0Gy4fnUdXHa3Zk3U86JTzdfOQvlOwHb3XFhe1YVvKR3IEy7LTDzhragGYVdHjm
woiP+BUPJ/j0SQxUPiYfk3Qki/au+FjPrsAI5958rRNKl7OIZkryTZsyKMsqoqEeBJB5nffv97uo
E/O+1SmQBFOBY4IlryD6tCVvwMgOtmSAgO1UneZwal8UCKlGC3e3mE6vVYoDk7NOweVWddGpIvrb
Vupge+w63E5TojaTRUPgzVYt7n05gkUD2Swv8T4hM8EZb3UEpNhXFIpgGZKAg47fKJgHKRug9zWq
HKLouwv3hYBACt4Xxxhk+S6cnlpSBuKD04y/Sn4PXtbfU6WVmVBNXmv2dCXNdePxZyln3ZPcpWO9
tPTFUd5WIPbYO3HsfFgvbAkIv5jDX8hyCJWcqe7lJiNbgB4LWn5xUjQhxuwNp2sW+ensq6+W+RRw
bM9hbz+x2ltDpX1MCA34LZEsVnEOZvOarDPtKnU/tFmXefvnCSR4c/nZiKntz1nOE8DNqvBz85cF
17EZa6ad0JCFK5NzjRRhtEtppKxUXFFsAPdUR2gBL3ZVQsdTPaS79G2Z/GoglXjpqQuawm6pYLOw
xlsX5veVkYr8itQDgHIPGJ59Sp04Db5Ip9mS1qZ5esipW4w8Z1VfXZ2CUzCHquQXRpA1rTEJYw4/
D8SNQ1BNESRTA2i50cubDI57EOlJgnVZVPjoxPcXe/qxso2zf1tWc2w0ohaXdzdzuk+9s9PwKfsk
LwPnjp5MC/5RN0ZXZN/ZfEbdVAQsGK2tyqzGQbS71+utKHqL2YmWFUYDGOqUw3Mv7gKGXV5WhzMe
/eV6mMVaj+LwMzR5ouDeu1dRwNWoWweUBbdGwvWZhIYpW7qaJEVqQ754p4JyyZ8Zwk7thx9cnpGb
lgoVW/ZFivK7LYf8sltSwYDXHge+lW7R2vXvqo84mk7Y11M46Ney8Nwph6+L2PqSIJk1SWHmshC5
yWWiBAVTnCH9cOPZj/QmlPJSE7v/3FdKy3OaQ6SqjqnSkb50LOdyeSNYAkRdU5MUNOIL63QDpmcF
NCZwH4ivgwNZ3j0Tvde/8GpWzOwtLLbE+/bRDogfzwzAZHQFj6Jp9x2bVQZtsLP4X16CKlayTbwP
3ijO8MbhjlB+tbnAblIvVAw1RLDvndnX/UdUkOfxjnGcRxw70bUbPD4Zfi0zfshSyKfM+aB1qE7P
VyrEgHPr3PeBYacwcap5ZQRYqEmPNVrvw/3sP0qqMSpnOXNXTCQi2LK0Q97zplUBqQ44p07OMhY3
Zi32ub73dsTjIec7smlAxHbiwzLaoQ5LH6nIg0Y9MCSzQpr3cZ3n8yuaBf/S50mPFTMDP3ftYctX
KZ7xD8SxMftlkmHGQHeNCn//IMTWtSOcmUk01Adfpr4sAmtS12Hw0hF2DcoFpHsYdfPcim8ObKEj
MiBHRXk6dQS0MFb+tYUMz4qIgqvQTHi8JXKUZq0Vyb8V93ecamiyMytoYTPgy4v5zWCEopwu0YZz
mPgFPEGXCVmVCBL56uDWd8D5Nlv+Eqr5n2lQZrVyfDG8cKZiF+dLXCiRcdyCvNIsudtilWzDxtdP
lqLvV1WaUEBuiQuVbGWhoCbr2unlJb4wV/tv07PXbFDeEC9/qXKOsM7P6PdluJ9++x0w3LgrM7j5
vhzdruLHUPnBIWi8hjv5hvy2EIwbHSbieMU5B9WR+7i7nW2lUnEcqGLp/C7b2a5Yw7M8czZ7woSV
gxUHcyA1ockzgMoj1rQK1//uP+04XT1BR8Bn9M06oKvcekO3PjGS1WqsLcSPVUEVxLn+JlTAhMyL
fl/agt92fV1tNC9XeC5JqQNhDm6JcZ3HfGeXdF1fM8G5HxyxsEmt9UoKp/wV1ySD+l7ZChKC40Q1
1jPLNE8R6HLL7lkuh+5KMu0l30AGLmJo6xYX8Ed1hjCegZTfwGnpNuNsNLTb3iK5oP6zs2Ye+6jS
V+xucMm16FZr34Zg5dFkttts0YUiAZwBwXIHdIIOOJs8aX95Xa0eLCM0C9htnFVFcRNzJ+Bn1/z4
bznUaLt5gIkFFhOHXtqe1rzv8s84XwmC445vZTwo09s8nTzyXXcvgqXAik2/ulWfU7GZEGlApx12
jaagwsV6MKpPnFFfo+O2ZqjTEHz+bb9+fpiphCbFitciYtm5ZKE0+mqCauCv5vL0X8+OyXLr1nhS
4OAtmK1iQw+RQ7xGasfQrSIt2OgeZESecD2AaM4nBL6uU+OeuiweWh7CLrB+Wzj5dfW6iN1ngu/c
/si+iSZVSvxSwvcyhh0DSJR+i+B3MSTRfgWPBXpTxWKU1z5xpK9oTq6jTK1SXRqFTvWB02eNCd1k
BJQKqCVmBrFY5LJGUtkxMtqNDiZwfi7BWCi2GtV3sr5z5KXfxelFHKYVX1yMZbCttL4y3Ks20PgK
0nf3y/8HWwuRVHVrXceOSjFMjbgoNI2s2VynERvDNKYzgyQTDnHFzz3l8N4khTGHVOkmcBtqlSvb
3BRp/Rfd83LEYuFrZ0fXFiq67BfnIfGA/HAh5duTL+wV33DY7T7j074zHYgt/S7ZreLpf2edDAtw
RufxEq/YKuC/leixiwCrmQmWXHqoY0s1A3LmxEcuyiqFRFCUr4mSbF/M2STkq1kMZ6wc49PWcj/v
tnZr8Cnf4xDxrd6lHlqjEU6GZc30q92xIjzb8moRiaYb1l281bgmb9dyWU01nJ+KAzyksriFLQA1
riDo2iZ3pdJxJ2XPrf/hv/+H005Vdf5Q3ha08T192bHx2IViw272SnfEZ9D8zHGDLAbX/rYLGpa+
lhMMTzgNd0lluS30YWhdWU6IszRSE+Y9MNqrkqKkSM7ENu0z4DMJWW/9qdxfpV4L+LafQN7pEhsC
DJO2BESk6qVIeCqYBRfqgbXkikL/FtBKDWDxbd+gle4iTYZ44bDxrkinOYW2f7Xz1QnjSdlgS4sl
kYeYC+2gGcpRZ/+YgTdPVr53GgxJQtPZvWSpnxoj4dfUla31sCSelJx6UuTdTeo3UXoYFOxmA8WE
7zNqXvCfCHXbPu+NPTz6r7Fp3GH2pq7NhYVTl2cBVbjEzscRtbu2kVEJakDR/detsmWIKahFGFLv
LiJvbVwTdS0UfHCcaYM9yQvVt1O2Kbu9/YSTsw/CS6f+UjR+69HdOvadBsGN6g2cL+qnyok3wsQC
c3kHBBe8O+sc8Q8jEQh0WlUQV4rvmMdq/CUPSFOycwgd7fpSDR6uetIZ76EmVQjm4t/F/YTEqUT2
nlYK4OssJS1MEqusDK+6SRkxVdD2oUzHnPqrvNKHOYPthlDKP9+xTfsop9Sa/vUpHkQNEfSU0RFS
guCisa8whXM0a4+ZkrkchYOZivWRltFLAOsEIfczlsWGcjfFXNN6eHgjMChMiPMtco+4FH/SzXpm
1Qfpq1MLLzZOK6BQ3iLBlfP0lR2aMxzk/5y8mDVfLVsj9L2LgKeWYFhBFlXFRJA98D7rp0aS87nU
Z90NwG7Sah2/o+RenTBDoa1cvWwKwXaOQvJ474wMt2vD0R+vlpjAyD6yqYm/eDl9R60a4N7yvEBE
RYSV0w/bbYeaJCCd42AQdWI1lVlBm1a15YzQoQYjCZndUSZqL4WTvivp+NelY7t9Z6sixpOl/QyH
Bri7LoMc0gH6NiolE0NimdQ9y1tuCISMZsGNm9DILN34pmhgfoF1hEC9WQb93s/oIivwM6pt5/WH
11s9U7E87ti8F4YrLp6gVSer0+zbPWsNm8u6axwATJzFGFGcC9Y8rjblrn4f0zIzNyECpl/fsOs2
syUMxOaH2KVWgRtuZZ5G1s/CA5p1ac4+mAShFIw87zQgKNBOA8Ab3uALrnXtETJJvPa+BGQIXZNv
tsipNyP0TIoW4ZcopEmfCRF/HChyB9uIlfZrcRW/A9ANa/T6J1HLKW9oz8YdIR2lM2hN3gciL+4Q
cJerq0HfNXW4hcF6bJ0j8zM9f3Thd7OZugfMwuQv7XZsPJR6trEaGNI+nsVSBM2SjQ2akSt7CFWR
6feZZnP60LA2MMV7Fs2gdWl6DM/2eTgscdn/FmA6TEtjaN6pKs69D5iKVgNeMX5Ak+nJWeoHH1cz
xkJXjeXlsZ9jxCQDsnMCBI3TXAkppKcc+B5bFjsxKTQ4F7v5qFxwRYXdIPZZ6ov8TYqUGNjgM1p3
b2IJfd51GUdDu/2+e568pxOHP6l6inkrbvarp+5r3P29EOTg04HaF7q0NwbJRL2D6kjddW9d0DuI
A/DNl4Dr/DQGllndzYwW2q9IiycCX2EXz6f6C2BDkNVrxJX5ct+06bdTEMmmk7Dy5Znf/C/Dev+W
tybD9bLeZO3i0iLqTcS+06j2xKsz78B3utVw8y2ObIwKtwQtfVnMuIThpfWGGe0H10Hl3zhnUZD+
6e5STK6UriepsUzC8+9G6K7UljPdXhFqTmDLXZmCoW5jSInpaophG88XZYVTm2m3jem83yeoU9mC
iv6pH8CfAJhKu/jtL/WRx8iOaetRXEcR1aQoyQXByfjI+g9EPyi3vyJ9mbsXkVA8O0PDZrq4Khvy
8puZDnncSToP6Xoz0R+sEtFq0uxlxKuvll2HxOcuIgLHadg7CsUjg5zLJzHfMxFfXVq3bs0Aoexf
5gm9ljYi75zG+oMt/aLEtllIBgV+EAFgBAhuS7fQRpBGw15okh3wiOs0jbCpsihhRkpn84cBFfB6
Jl3Zccmxr7vEaJ8SBNIHdL5Biq7KRMtLhN/UkKZL1BCtUz8NV9iOVz3UdbBvdGewcgmBNFUUc+AS
2RtUeNYGblr3TwSFrIOC094uhWzVu0hi8rJPb3NJtOyOywDuTfdikCjQ3aVDOWnS+ajf9WecJG0C
ZnQ8luaxxG7s8CvpfQ9eF/eONDS9SM/WLc5zPUxy9+xJB3zhT8ofLVZ0OjuYMcHfUlG8Zud7xZni
JrfC1ufNPc357R9Hi+074Hbw/zKb2Yq2f8++FmNFlA2OvBWOY8mTooLwcUO+zIwQ/lCijGcDMk/a
f/CQYAbxt0E+aGalBmB3L7wjxXcq+Xsa/BfuJL7Tt7aEuZoqANg6Z2ojSeNGRar5/T9lXIe0Ulk5
rmx6Miz315CUvg72Ts9D8R3dOq2tvLeDV0wstlsIryijGgyKftkt4xgcY8YgRVxRUXt8L/zrGzAl
RDGL1XCGoPC3/pjdDtUdGuqnzy9Zrg4mMuKgV96N41EuP23XKgujN3oK4RBhPpGAqTvBk7vnXFoL
h8r3PaZSUyMGHz1Nk2G3wFvvFcP8QnDBSxXT7S8QLM0HASjW7em44whghwnNsiIhgCfMxRZ0Me2K
X0z6nwZ7GOeAwSNhr17FJ85p66vOU0D4Qsj0inQYTpW8Pi4kbqGWr8iQ3yDPOXa6B4Dehm8K+NuJ
i5BeEnFM6e+TtT1cKljS1JiKZE4YWPGaokZPLWypInmT5/ndrM8OxlU6NLk9ofaaOaOgYHK1wZEE
ot++tFLJUsFdN81/uN73T//uXvKTCkIs4iL55qMf0VwC7DwE4V8/X0h71f19eW8WD+h+GMWWdUUq
XzjNTlFwVLTaq44QvJ8U2mLzFsX+plvuf6hf1NsASoZeUIGJKc9B7jRP4BCz7QIpL6ugM/++nTGC
VLwMJ7TbzR4TWnVdehohyYm0g1avOUEiUeTVar1OkmqUtmTw3w2MSKVAn1Y1CSBjizcRfL0jJ1WL
Kv+9XE1ZE3/s8dHQocubgIrO6u/OiGTFnbDnWQBsqfbs7Omn17amxyMWXvUPY7DUaAsQMAAdYtYX
vLE34OCFvEU+VGRcJ/5Q4lIJEsFdTcS5yyYqILbi9EOhV5WoSbInkde04OcbwU2aS9Kcqd+7kUXU
7INV5wxbH3GxrcX2ioWDlNp5mXY6QlM1fhb+qCLKVQ+R7CqM0fMUNfguNgxAasz4hWZjzEXoE8gs
XfmHkvdh5OXNyvkxjrG35DqbyfCRVa9VzHArU+PqqmM7U3OQpc050BcMGUzjSqG2xr2nYFBrE5pI
2K4CO41oxPRLPh9NUakqaqX4+tyaadvnFXvYVdaLPivm8Sl6GtoLsS2oYxNsNu0KGmIOeuOJFs49
JnLMGiAggHoTDZXR6lYOk2/3Pf2+ZF4ASp6o6bb326FIpknxZYi4yhZJjmY9biXfopEqA8rryn8F
fHzla6NYDrvQ5EjL/Jg6DLZ0ivLhyGGQBFWQ/JPrxitvdgTlozqez2u2tCipZHLJBvHTvr1rEXrP
r7MHwXdFydZhXqsde3DjFSW5j7lyNt+QfQMDQJKwFpIo5VsAsbO9pull6Wztok8dPg/MQ19qBaJ8
4HZPVqVT+klk+M1W1U9p4T9987uE4HFwuE57h7KirhRsDcUSY7Enk6QEKkuP6A3Ta08Vs6+Bx/24
VY/60EulBlsaaprORJqRkQ4nZmqfp3tKvmQjpr5KuGwLRDOQbGE+GQhxmPslFtfkeDLRT5YL0PNh
j66A3IEyk5+mbGLiLMZKlX76v+58qsn2nFDvbfMdeRUyXS0lJho4cVXBlcHSdRh3VSruPxCXuUS7
TWsAs6og993RrxVSrm+9hnatSKCQHaLSEmaXFBYJ1m/c4lcJbO6Lm4fRQROESVoMgBYbEQwk9YMg
+aCkdctN2ZsRKWohv3B/WDCjTXwCu7QyoiZSsoatkDy+Src2dhuAB01KJIGMBdgArOQJUe7gbVe2
V4JsHFgC0UAEWK26+PvptySjtBtzFEuQHpL5XOj4GdcypF5liEOq3FCKQk0uiiMY7H+RaxhBJAvJ
a8oHLEz+gnHeeG7hm342XF91uuiGkgMrC1ISzithxjow4GBbJmElhLa44+cT3YUngSg9GfZBV4Ab
jNEJi1BtNDOFqhv58QSCOHc4b/rkrnatZJa6XvTZocwTaDZabTqyKo4/RQTCAVDnTazmMDO6GXrc
IFflOe8VwbTOGlXOI1qLpViBta9UPHShrR8sglGytD9yQxqKtK3i5e0rWZkTnsnsdUcRgVEwCDs+
A4mAE86fuJPJMFD8IiTT3wJvAV+t4a9081o7NigRBUzZQRXbCmcZ1NuG4JrIZkDYVsJXlH1Oq+B5
KDf9km9xI5iZa8BbY5jlnKuxcIVOmQX66DXrEcBVa8Ei9xllv6zd/pmOe/npm9nQG6DNaKKHy5Aw
axPly0gkIrRb9S+cLq3bzYeMghXeX4ALi4hjRVK61m8R5uCHkkgUN+of6z1h3DGmssk4C0BotnKN
BbxRmRkMfEURo//uqBBv/R/ugFCcy4zRihNZ6o8nrHO8Wq67lyyqKUKOXi98E/AG5EYb2VPqHBc2
byUYS+e6gFejImsKhzCJ4mYZOLhSvc/2zgSMk2Wr1XcSdc1MxNJTCeEuSeOVYaJ1ybltZEjck/YH
WuV9jTZ6Us7VMXLj7YlsokcKLjOCCAcZsfJXObVdQcO5h1lzLzqDiQB0hQRAGYtUpFmDk7rEyLox
zuWN0KjBiNcvwqVOq4AabTVCIMu3S36dNyghkkBgtphCwQvj6A9V9OmawfQs9hYaxis82+dhpmmg
zPqHkcuyAObHUOJo6tm8OEpAs3yYgHzT5Zr2nBx9aE5WjrdEJTvsFvdTQxmjvzekNsbmLCoVsVNr
+X9JFXYFM1BiiQB4/Qb2tS4IsLYXn9Ci7MrN/YO8pnbT8sSpPHlci7o2w5GnzlSxCvbtMVBzPxfW
p5szUfUYqBVcEQ/IYnwY2QWoFl+XWbhi4chvZvKogI7xiXWiSyfbR+dlIfIMqP1VFZ1YbFpS1ZUd
iZQYR7P0Wr3lymxyEfZnIHzjZ8hh45pNgMUBfVosQ2+Ur2WkgdaJVDwQdtNksknActb/fvs53czt
6VZEwGIJ/SSqWGyOZ+e94J0/9pHsShKVJT3L+AzFJhyNk6rkf8/vc2X0OLYI5BuGCrYI+D7RcqA1
Lc9L9L6UCJ3l48PvVc+19nNfs9p5hU6uyeM+rf21NhnIBanh6TvThGHq11cgoIOOoVX/zo4rAb2e
Akn4YLe0WlmlWeeD1WErWWWbtwTKjO5t2vzpuC6rVNTG4WNfEAtoAnVpB0svFpmR+PQ81BFUf1BA
nWbFxPqX9KK1ffpnrg4gD/P7mKB7drNqqw6o8gYCJiLsBDtCbQNCuh3s4PzNd/5s5o3s4NNO5/4/
oXxRdpRgtYzNRrZEch5Sv7VgtkYc/D02pGlraKCYFWgseeOeuD4Q35dbd7yvf76gjZdKt8u3FhMC
lFL5HBoiQ0WXkx0Mtanb5q+afgTlfJzrnjlnJJpF995WeSdG6YFH7QbKdXxKbzJHHCJzwBEQVXwP
VWB8R3W/D4njA2FsKQeKbmhNKMeoswjSuB/cW7zoakI8DCmf2vDcHvMDTwnGl2VFKpHDlp2Hgp5S
AnjEw1eJiyvFclW1dwvd8VsQKiB/qJNfobvkEF3/WT+rWUw0lI9qQy8UIa291oVHaPVcM3cJnM9w
Y7PrIEimLoQu9PLoMPuZ9Nv8MUog+Y2k7+OUa6fsFdqOHNGymozX6kPx/W8qzh4OlOVWWU5uGJ08
pPeRGiD9SIyetoAg39KJ5N2fTYsTGRldoGkIEEceivzFKKKAAiZN5qzTfevOd87gB3gryuMFUhPr
SaLHrCt1rQoZG453ipmJZEDAJIHIdHp1WWWm0HLn76MNvv/9gn/1vUWLWUwkcDWXqOTQu2p/TO8t
9R4qoW1ddZ1mY/RSgG/upv7kg7ZW5av2n/5brBYk1uvKmX6Rtl/F6Lm9e1WDB6NvjJ5u6agHEIxT
1CLbKn/haQztXz9ZNVw8P9UhkS3Ex5jcFsXXnGikw1yILWAvSrDfdS7mkZkkmzl6JBhKKCkXeMb/
V5PwfRnJAwrqvY/jljFVSxHjnVTL8A7mt+DxVAnp+6Nt+JrLHd+GhxQKKtbJn5Kim0yHqhUVfm1M
s2g8mO01pYafNek4b6ww+qxuX745tSg/QkYwRuXOWsvgghBLzNgcLEuD9cFW5NpmsttqTRkIDb83
Xz0EDdEJteZQcAOR6HEnfS3ZXmkdn+khOW7loPhvpmBhVhWxD1NqAwLYpW7+H5J6Z/fTwiiWaD84
TFqpReRKHKR/jI+dpgxMgk4+I6KPWnJfK5Dlju7XSVpg9oAKfTWSN05d6OiqAwId1kb5gyYMZck2
SM8PWzKg9GP3IZCsSFrGnbHpQbiJhEONYVsTLQrDQJAte///BJzXoDfUTH9wbHh5Jt57Hz30sv/G
id1c4jzJyIxUv2UBeLlmRn8laSX8L1CJwjneWj7f73MBHS+rj7L9xVYIJo6RWSa0Mp25JDAbgzEx
l2UmGKqMA0qaYP57MUBddFkyaLQ2mnAQA4mTuETdBUdlyYPuwd0VpcvQScsltkkFB7HXLCBL5JRg
6xQitBgmdUBtiGWZT2pPSap8aUDl4B5mmm/V4JJqtfMnI0hmF234x9H/vHH3Thydje/rl0WQFRoB
LCckjdSNB3xoqjnZIjo55qYG2ePvM7Tc4osM2TR3uxWVtN/GgSUdCB6Io5dzL9tgiF6cNauwo+6/
R1wTdIrlxY0dA++C3PRLA8m+HAXULOd72CVgfs/D9Yos2akUyzOtqWPWV76p1eYqYbqHQi6sOhb6
AIKyDaJvfiCfNOv27YtzVyLRKFmt7nsMXsUv6tWKSYcK+lmQY6dtJqXjKHY0a+HJ81kQqbLtoAoy
yJ/cA4roLNHbUCKzGnyUL3xh+fGjGOqxVchlj6Mf/tE8hSckwPDirDFWk1VPpMNMIK91SW/wlFkq
OYAlBHPpus7IraY2jGWRaCjQbX6rmyl99emLoU/uj2FpsHJWF/HREoc4soOhLKhm3zYv7mU+iV93
uXl/5XgHLsDoPl/iOKO92BBsDLBjqBJHbu3+R87V9a9N+3IG8ZX9sf6N2t7CxUX5cAOErCi2Cqfx
tumeSPN6gxgFdHhTddBCSGIqtoogJiJJX5auTKpOi3P+R8qskQ47LxRmVhpup6NEgxjJmhdnYi+G
+YTXohKxtOafgd9rEvGWBlctygWfYb7T+C9vT6t7Y+vFNo+w1Y5/VIM92qPispHkPCDkzcavKPgV
zpuzKl4rsLr94y06uiQS7XIY+MZOoyKqBXs3F84bnm1chI2OYuUQPzkyb/U97skCys2bDquoPkm3
hADPMFPMNpHn5edHjRryIzhQo3GTaUBqJq7IkxaCSY8L5br1hNSm1ttQyEiM7a1s7rZpM0Xeuy0l
ydOUkpwMscrVpAPxb+3G2BXGJ7f1haU5DE8/2UVhTwUaT6WYMiJui0oItEdA77dFf9jgG5kkKD57
/M/8p8nBXDJ+kRBNmqZXpGs1UFIU/JrDCxn8jbDRovPEfighKRNqBDrExooUe4nUVYwCnAWOIC79
bRZRgiGZEzpd2J15qe89LTB5SzFq9w02OrsWM7OgLW0P/bkNPZ+A/iMkeebIrPdbXNxtALKomARQ
m/u8yvbbCfc4XDeAqWw7AIbsaM68gZYU+VP8lms/+hxoPf0Y6S0Isthr/7fc9Qwwe3KhM994k3Uu
m3qhJ1IOQYWZSzIasyXaFdd4sSSZTpW5+2JzXDcb0eiOlVPk2GKhF3XgA6nW5G3plvdEVlU2nAjz
2xtVM5DLjH3dNvtbgA3YdP89coAb7PMsFkRjmvvQiqmRNXnLJ23dqzTu1tLj2JN2qpmjWZzIIreI
EZ8As3Clu+5SMJzCcdk2oRy1OlDFbRAHuHb1p5zd4y69zm5+pwRFZT/Rgu0RH/g3PIm1F7vsEvEH
9H72lBVYxHZrVbqvG4gvrBfOQA75pkUMnOiJXDUAZ82Wb3/eG23g5dgefw94Qa5rY6x30R/ND8LJ
pdYeyxIMbMUvDG0aV9VTtB8TdVz/ZF7VRDneyFdYxV9ajzocg0+Qm1uU5Xml/Wkts1hbnW7UFoQH
diGImwaTdj5YdHvxRytAoUxxz7owbt73UlKVT39zjj4yu7w6JEALss08h0IhiBRpWQCpipZ/tVfo
R7OJBpMfm+ePxcPqwNJ5/FC/sMvzf+MsC22vWOjSBO35NbbzFwBmA9JNVtPJwfuIXiArt30qcuu9
vb+CSO1qpGt2U29Jft02hXAPSUZ83R80ifxhhRMTSFkEApOdnWd6Tzd0NtenvE77SfGYuv5z0sfT
+21gvZ/ckbQIZtqaeEsqP0FIXkA+MkWv+Lxhw9apdb/x21kPUkrzOMJib1b/KBdus2MDMFUeziiM
PjXZlHm98r5hOQKIYNu/3GtxO656JIkcXIe+kTbZImaCQttq42lf5PfUCLCgE40BxQ7c0Lz9cQGH
yvHEo4uDJmFUutjUix0w8+YUg3Mv4H1u4SFcIh7YdO+IrJS5cRIJWCKE9Bc+WK6zD6V/Bspyf6Aq
Ps5FCyGayY0kwr7avDEhRQA804g30IyQgnOh/RYHLTWGMxda4nJEFarjn6nfJsi5z1Q/97kvDNyX
a5GBHTZ7hASR7HNif6EXnIYRO9Wjyxc1WTmzXDX7sCPeBnfx8w0DoFNDE9r0GYYU89zubvL1K0/J
oomT2zSBGDEQHvJP5drRupQSod4w4+z73xHqyI0Y+xvgHb8G6mbsvhYdizULTRXOfCoOmxlyIntJ
s+NAnu6wqwqzGOARE76ta2tdzJ+Ons+LqdHmHYKC7zbkhw8s51BkhTeLQhqcpyjdWeQMESdIs+CZ
cl3KSYXi5NWg/4s3/u9CZKG4jRg7Uxmx4lUQqLvVIISDORy92AGbRdTJJcw+3lXCuyjvfzghl6tM
q/hJVczwhDADsjPHxjpK9Kz9pnjRkaHf2oZ2Fttjnv6bxew2d7x01yLr6+1AKuk13KEAUScedQmr
Mp9ELx863axUgxyxjHVqcMI/RjbjmSDrmMrYRXc9YLeBhoFyBZsBLnLrq9wWYcicmYUVF1U72V/2
ejmANqCjTYauAIRcBXE+ld4eJihY1EAL9C94GKmk2icNwd7Ucwm3bsgiaEwWZw8QEdQ98m952Td4
cBt0G+8y0YnpvAiX/F3h4B96M3T3KhrmcuIhxm2X4QPanFZPVZNoWH6Q6LKirU35BQ9/UglUufBv
owzQc9xh0Wtr5W3wcisfl5r4MsW9Mgc8RGJvSPPOOszNPpfaSnmf3VMXVvXUWXia6QOxdBU3axsq
NEBQM8EAoAzEXwXc5FNW8ihZm17g4GRLmd+vxOFr9f0DseB0S7om/Dx0LkrVfqcFWSHsAAG2SSTm
8jiMrYAvRx0lBwc1OJrKzht21HTs8bgYTMkend2Zx5QADhfTjLehRl12lFRdZ+UOMUHkgVVD/ROT
/S7XGjY8BJ+tkth12OPRMXjuXiqLuZrcS7V/glQpbiBDmsz3N9vVy9nWg4vXPoqvlCbNDDTD5+9i
f3FZJmPre3FXU64cgznmY8NxH0A8aNeIUnwzX6VQdhtuq9RdWWwb1s4vc2KUkwjOyY8VyNdivQhy
Jyk6mFMYit27MVtm042MDiOTIqu1d9fFjMT+8DjiJfBUbBgNZLRZ5RXU5efm+xgqVZT/C1mrc/jO
QKTTHY0nbW7IJ7VYny/6SGU1EMYoebiNe3GWAs7teBShQUlCdhfuy5lr+jAHjm9g7IbXSNUseO+s
Xj7psCM+jG2eiUldlqrD0rTYUCUryn4h+qYbBJKGurks8Yk7hwMmcZiAhPYygAEM/BfVfj2TdsD2
Tz2t3NygWpmO3Dl8ifz8TFy3rUNL6PAoP56mHnMPFpOhmlSHAdpCKGGumJX03DL3JRQFKqFANmMt
jlNg3dl0ELr/bpW9Vv4fm7LWcoV4QTk89pfkCBNB0SFAUnKd50j4HEF/jGqoqgkSlXHnAp+w4ucO
6IbX+Sel08aoX/+dOhIRhCOcz1FWfwrqZepTFQT37gl+ZKrL4mcFy74TDmg2b4fhum1PLokJsqNT
iOyEoff09evuwX8Lyo/+hrgDbDoPBq8cpc07zngfZkoctq84Tu0dLu1sH5fPTrj3Wam3jwNZwsWG
u3D4OCkpBt7BK5chGQOAOFrNJX5e/KQR97zG2S0ZgpQx0FndkU6l//IscE+V7oSTHPPsWYxaw2Zb
JTFmP38ptpLGVvYVLSWW1zzP2VYKxTO4JZ1wfYzIyco+EYwbEGEh7FVAYNbSlIck9ZseLCAyffiT
AenW95heuY5b90Oq4Kxps4W0DwssQm2CAIIC9kJG+JVgSxVz60RAFE3xG7e8ozR/GDY65IlJ22Xe
7rvRV2QUHNjqUzJtdcb+CrAvSN6L9WHWTtN1bUnrFwzuBBS7KwhZl/KA4vUsCgOfiD+NyaM4zyVs
8T4iuAMDh01MxBmTnip4IomjJiP/j0aBcvIPizH5096NawnmdjcS1nJhHPNvZHbMprMWCcpTM1Vb
1vX3wbSSDYzaFD7/vPYk48l05RYALGSBJ8nwdS8eO3pz8bSRAmi/L3o6UTq/2J6aT55QP/Ypwss8
ibyONQ5syoLaQPYPGkpY1K8O5JOTcPN1Mzg6t3EOvfPyeJs7odAC658DoJprOwKl9tDpSvemjCZb
PrCCLMOqbIrE/C1PaIVeZq1YEFOYNLpU53A2Qr13kLH5AunN3LFqEyP3KyNTf/FgS5ye9dCPcyqf
IcytffDhKAfvi4cJeyWFjCilV5uFwob+3eIFUUVFYXxFEv/gZZGqgo4290L7dqbss15/n3KTQzb+
xqbeTJYd3bIWJmlqAX/XxW2UDiTIMO57smWmPP8C67e72UxCKnK+eHpK5UDDugJx/mPwvql540DY
ImlydCU0882GmX0A5RRGPdAYW0D38uW54qQ9aMHUyCilI3BoCg5Rb36koiczcvOJXVk/X+L1318V
niOxoH6odW8mGRArODs7+ZCZ1d/CLWpYnwxAkfBD2cTwq6kS9dP+Fr85h+rbT6meLH3lDUzYE0Z1
cjYJE/36gEYLrv5IBZvjTyeSnMwhcMfrRSSK9Mk5p1ExvUgFVmVPvJCu7nF8NuTlufX0RwJLVkgK
4eJQriVhFwXEwNJ4mzq0k16dwKzJndYeSyCb3GLmJspqtwE1ov805jx60A4rqapTlXx1hi5wNJKv
eBNTlERoiMisQ0UH7o8jEVUaM/KXRLkkoXz4BfzdlCT5feyu48kjgjG9dOaSVmesM80PtPBQQ8dV
K/zyks0p4IXcdJLxE4m8q+wu4bU5tduqvbpcucRR4rFyG7PTqCiVwhPD1GCjwrJ6LWf7VG63MRhg
WDvjQEpN8CWubk8/MX/TDktDLAhgACYKr0wLwNASRoX/OjN2Jh4aDIUPxY8pzGtEUX0pUV1ZWDdC
T3Plv7H5rWk9BW2J1K1oFy/GGP/jHU2hJIc+k2HfMx0+0OPbseFp35/v1jkGz0QvoVVj29Ox/vAB
fNiesr81q+dUh+TzMV/LNsHLcYvo0ZrzQd+HkeN7ja9FMLpexkkSIXL0zUjp/Xdo5tJZnhHR0vvV
jHJsVwMkiRP/+n7N6VtZEMNDC7ds0YKxOjCw3cSBwwT+uk2DamrbVWvFZHtNpewDYo1TxZd7sz2v
ENtJ9ThrBsLkX84VBP8VjAUojb+knfwCg9T5YxV64X4SN+LBUdY21Awyq2Lux60uJNUFYT+MGupT
yxUXUQL6/df+F8WVVYgp2COQlF/Qdp8TpMU0glBc4qEjAhVNHmCk7xW+8revBIkp+GO4SYmfxuTx
Qx4yrwGIrvgioGtI+xSATLW69YSLlBzDyUkxn5i0EuQPqqLRaAu0OaKbGgztGwBKfx10fHyupPYF
jmuoZSRdfUp1WTjiF4RZ9zgD2rGq6cQIupdvo6sXHudbkSd1jWAZK+jBfZOjakNss2qZwQ/8hPIG
j7ry0K5cX1W2JBV5FJB1wDgUEDiujrRqsHfmHFzIeRkPQZcsvJBxGs2ncUsO5wGCO1gftGvr/0py
559RKxPUUyJNLG8yBAFMb85UJieUk3eqLWjbvidXnD3+7w/Gzi+asj99OUbtpzA4mPdk4H2lRFN7
Pc5cT6a/w5H42x3S8Vq1waDguEoJ3EgGc54H5C5/NWebUgl2k5cxTHBgwZp9HiTKgaO/InhDTBdk
lxqx+tmJ2hZrycoOPXIAhAiVWfqRlvoFQOtyryh8jTGfY6psu62SNjAq10d4DeLdxhAFJlnP5b28
5NbkzjviqUZK+wXMqTi1mupYZSQHC+SKvLSVhljwTPbX7NM8vtP52nxW+upJZQvz8i8w4stbc3VO
iccAglw7Yy3pvVH/M+XmzcsJdA/JrC3+YrxWEuZvE1G72DpllXGllJJz0Klibmu99YufF8Z5Yicx
cnLP/blLk92+G+9+xcDzK7UXmIhmUAWqOoQOwFrcfRrPITI8cnuJ4oSvE0i/cUa8np1CW7YBTD/7
Xh3g9hWcrjBlxzpPH/k5Z9FVIBhkaQqDZNjjQVcX6HTX3XkulUi6ndjtlECjPmQKSj9wGO63VLf+
5brsAiLZz9i9yGtL4Qo1Z8NNHDje4X8/VgGKOv04zfqx6Bn3HmyQXUoCIrTzhNI+fp/Qm4O3mQS/
RwK1HuIKXw105Icj9vCTxRu0ljJpdE4urhy4MBk80k1n9bZgR2KG3O/il9Gt055rYqTPIWOdCKgw
Qu32MW1iBZIVOY633rJ3w7bwirN4Zb12ojbUkzQNxw3HhACJ+R+Dtx8+RPQyA8jyAxRiBrm3xKOr
SgAYGekCNxGW/hovVBSjZVXSNoU6QOTUsD8l5+oH8NsAAMGpSbfQx5GkAJteFMZlnz82kjuSyAM7
1SNR4VIrwNUoGqp6xBBcet3xrCFGWnoBq2GxjJ1F7c9/adz2Fni4pVy2TcuqNwbUJtrOGOgjmpvQ
reXLJwRe+77V4DYEqxHNiietEtxb3OJxucSmP5aiI2yGJBJRP44VpUSZUOgaGhwAE474gdDam1Yw
nInruYTVVP0naGz0V46sHrDVL1zTJ/9VzE0tIshEUznpFxgi8k/0/tQqbpeKRUiFIUI0lKk2yiCc
S3D7qobkViUpo5LA8fZv8ptuG/+GxwsPVcz6yxDX/bft0FU+IKDDImLHLo5Bxbs73KYnFdL2HbNw
ElIhoE074TKTJyygFeSwOFVLfPlsGd3f/umee/Jhl1Z2zbd8DB75+01jM5h6EuTB0ZEZcyWac6u1
obE204q18zsJaEiRXpxY74HUYDjYrDOctgiEeaFU9kjgRuXE1+0pwh7x34bDs1uR47DzfsJ3Xk5H
wR/X+clKIgFJ1J1NNucYM6Uq/qY6bYYyztntvsdlzX+72Astk0e/wKvnVppJaWtSBQfxmEKXSjC0
RFb+0g6yk9HSvsC917GqJUozlP5Qmp76OAQSnUCLyGzelFLJ8X+/r9XdhTAB5/nHSmNiLeA6v2X9
3QiMAQUftjQ9f8nrHYWcY2k5BOZPuSbk5UpHU2z5TGWLV3JhEzeGLNByFLqdvRcmLN9ZW7eV59ze
fCS5tCQw5HnWDZIc283JCRV2tM7tCY0bbhyfYnI2vL3LLn2I7iZbIqbD/gcjkm8PN/kx+teYd/o1
CzucsCE4EhM0eSUKLGLEF3CkY+ikb3exAYSll6j/1tx+Tgs7bgY+Gz/9qkhTZSKgx7tQv5GbByFc
/UQgk3gtzXwzUibSFKmqckTKpdFAVZkjbrz+//pyKUBKuahr7AC/cdPZVnjSEZYmv4XQMBFu4SCb
B4P3wzyEcCDoWJ4Vh5T3Wl4/k9rtGHpj8VerFvfelHnCcXCF1a0Qisa2jgt1GlaNO7/DgWbEOpBJ
j4ayoTe5jEpyd42SqqDtFiwIa1Tavd2Yt84AR/6W6S28evkq10AZSWH/gxaFRBY3vf1FNQrMI/qY
+6/7ZbWKSAS8FC/QRpsMPEH+Gn5ZINxAI2n+83tG1ZpkxxkNGsQUJuKNnBl4VsfVR9rY+jf07P/8
G0IfORNUwr464SKzDTw6CdTqJy2Ae/CMEy3iYmzs1u9zSU6ofER2a3JMGnOiueHliO/Y4XTzqFrZ
I9D9MW1j2MhEUxstnes7ko+98z2f4JpO26Jz2W/nzT2KOyqGZ0OoKWgJrs/YEd8TYo4FU8M6ac2c
9cPSQ7Yk3X3WXq4DerhENJfAT9S0mEFngyueno/EBpnCi7vXPtm7fPFUt+kb33p5VwzjyS0pUe4R
jtlQf7+oorwcB+/ri/YJ0YFtSfeklXhbKC7LEmfuLwnGqDmYnxM3jiTwZ/gV5xGlAoq8im7FvQrM
C89MbK0oeB3KT3skxm4KoX0tF2eFC90iY827LBIk9NqTFL4YRlmLskaNPVA3hGfl6/GNIA9EbnJw
vSrN3rDHJgXI9vUcqyWoB78LDu9c3M/MgH2KpHsJLxZZnTgMg4ia2F04FjWbABOAzVNlJy5evb8i
0aZiAbh2Cx6/pWiXsIvCozOndCnc+YP6YSxvJZLIctntwLGxPceUQxSM1ZDzZN9S4v4tNMA6yazY
tmX87lj4hJ62fGsHG9szmILdiA7OcqeEKg0xhGOsCJuE46vOPOjcZNbqQoRZKmhiO1Y+l9FKRSoo
3QgAcxyOXmn1TUB1m30J2hEaaSAGQ3o3EHUKPHvZhVfh54tR/5AsO4/1dPMwMcxZvR40Pd68OPHw
fN/Yh3gPuY18WSzR0UAlOwNOHM69UztAlZEwNBfCzk1mBSIllITCJgdGUdMvdFcxJClNTd+I7Wg2
aVwBikOesG+pzSf2uxxMZtmD/sMoQiYcXJOuzrInrr4U3GIl8t3Fu3vdaLKjHJ/Hb/rkdtOuPzAf
GV2dHWYwbuc46Z+gN8jB6AOUmKONaydOajFRYtC8G6fxHjs9I4NGZvmk7jeC45FXNlicJMNhYuQI
BtuVvIobasJk4BaBPa7FZ5cwDW+eEY3qmnBPpD7Cjn/nDk1a/jhnrcUrzJ4AnrIPN+3FTg4jNfLS
ZvBx23Q/2CSYL0pfULlWYUeXjDB0+msoYaCEiiyTcR5fmA4xz9+UCKM+IIIEhq366T6KmQTerz5U
8z/n+v3aJfxU/d+V/kEtFgd4+zLRWOidDIUxxI0C+0TTMwCqJlWhAyZm9QVcyEq5svGb6RblY9dc
ugMh0GLJboJwOUZbVEV/AuLmymGvr3vwRRgykb4p/QCWicdMiiVafOppsqCh/M7UthgSDBKBtIdJ
D6B3UvIkSBjS/sN5j/ufnJ8/0Mn2xNOK7sR1hYvNpDVVqJorEvdIq1uPX89yYQd+5C4KAC2vH1gM
7jB57oseG01o8HgWbx/h/0TtFPYf/eOhPAMTQbp5feJC4q0ZE9Q5a7ZbRQtLrogs67lTOMe+KcGv
tl2nonVlt1od7NwRZSJGcCrxmEFFCZH2gIg5N9BqezUltYbEhrOkCQn4QZ+cgWv+aNUp8g3VM+jM
8on3ULnV7+r/L+KFnfzNEFtE2tBkK9xojmUmLRYbAZCF16YXSnyHlr45YjAx1Dz5HzP82re5HVc6
oNX0zLiqWPcuGxNzGLtVSstlwdVBSedHcBtuyZIQGSxf6cQJDYW7wv1Zr5oq7E7NditgfbW8Fm/y
Mgvcb+8+TSaWxgskSi1PGEJU/PXjriZnVQJxxU/1YAmkMbRpIx/sNTeoneFR0qddIklhGcZIeA/x
rka5OG5wISne4HJH3KpjqhzHxpMPFaVuw+C/nzypnA8SIa0ypKX5aqSaEx+ryk5FbRWsKbTKLO8Z
5SigE35qbicCWrX87jIOl1yG8VYOyIGxL5srMbZy3fyc/4wcS1fhoBM4wFBiTVy+QbaEkgets1Q0
PYJbSbUKnJWfvRmh9p9kvkjmvIfIsMYTZ0+n4iB2k/Jx6Up4tcUCXlv3jthtQBmjgYnm9g9i3e7b
K+X6B6quYNsfvb3Y6rxUPthbj3GyW71vHqxvNExEj28rfOZDKifvDpQivKhkWFd2sdK+ZbDuzmvU
W9JsYwtQshAwIGwunRx0Tlt0Z0Zhh1fqISVefpeuOBDbKCPXwQYs5vkQXQbKz07JzE6/qVRgWYi/
XlYiOlnYU57M6bTVewGiY2It1EFAi0hoT6/THJyUQIe02MRtPG0WFRozqDWox+vvgcNpJA8Xygwb
GUSmtzo4g5px+ASpyqOy+75kwknDeZ0tZN/ILTi4KDECfsSMorIvPfAidLmAffceqbM5ZdQKCMUJ
JtY+AJ3hzsXA59qGM7Fork6HLKo4NpM7TL5RhnxC32aUZpivprbGYnZyd2gmmiLWW7Gzs8YmQVY6
NjKflhe7sI0oUX+2yuHZcNki3sZ496aqdjkrfrVas5ELLmx2QSaHziMVWTVvdhFzYxBNwd6kgO3i
NTrN5SaAy7q0fwyNtCLh108yppdZ1nF0uJNLJSPaprRgG8GqqAY3GMMb/nJZw5xZMDKXS9k9WN7r
h6QnG4oHf1DyBBgtdCT1c74EHMt3aPJH7gRGJ4VMubloZ4HxpuqvO93WGCeLr2Ah+jI/ihScIpMD
WOOaB8TxxloY8r3xLzGj1z8fWd4xp9hlf2vYI3EZnV3MwAIIz+QQ6ndrs8tDEXS0sauuXEwWKKbk
apKB+4Pubz8IYwwA7d2wwsSgyOyLalMyoKkrOyIfu1KkayGuOhT1gOZdJaWs9YhbgpJT/wrEF8tb
I1602J2PbeLBkHaR8HUL2bVrE3x+Z78oza8/oDp/Hu2/88j0xwXIlI+/QY0CNa7ZI73+tHRC0PaB
PPUfGVck/FZkL1PwYbQiXX7+o/j027UU3mZULtR+xZBvneKl+43qmRTZsDpeKS06DlptEqC3QQvX
/HUf0R7L8GRnABfuvmOYSFLIa+Tsw2nczZVVmJkBniGFjTZku4u/6haUfR8q4Ee1iVclwG+/WaLp
xfA2egEnGmmzvzwZuYHy9qZravRY8oHnZu2+p6JtUZR2/4h/BQjbchYAN/Zpa7O3KltyiH+Ln5ah
uqRi8wOMb2PJrQngvbXspqu2SZtoFH5mHRqUHgapg7c0XRo420P7mmR6w4DxO0oJEM/n5DaqVpWd
PyvKPUl+xexYfR6Cb7LgMkSJAc/SbUQ30AWUhveNwgpIus6iJIYnzyuEHMF3Kv445p6Mk7UypNN+
aIS3p67xz2D4noceGiiamymajous+di7tBvnvOcrqHyQH0btsS62egyi55rHhB8ep1nmaCD+7yzD
4WAvfz5bRRDd/Fz6/Ap5HboGyvCR3/zfUA+t7G/FjL1EuiZQmAJLriGQWOyhrCFX8Zt0oL142S45
IvkwawGR5PoKtw05esz/5PMrWlLNCiWuCehlhO6bPZsaf/R1phmb7KgS3Wng2xAIMemOefOpwh1N
G0QXZ9I3vK0DXeRn1m++glMgc2ndoInMkmA4CerO2Lt43N6ywOM81u2v3RWJx8M7q+phOR9Y0/oa
L/ieOq7LbnbBeZ2ac8X8u/WsmoywyTaO8YZu/qi+dMsZh8CJR+OONp5hl/rVQEQqGxqu8mJ3phzk
6hZlCJrQ1FUYsXG81swGCIPJ9q9cddm/iC+DJ+iMQsyTY3Zfmv+OQf9J6x0/Gdui92AgGl5bu68g
IpJM7YZ4FsNawI3jjn2eXSfb0g/gecwjHz8mUq9j/0wtjvmOb0tVS/B1fx9BC6lhR/a8gDYCaP3x
bPTThfq5e4NBiB0TL+RrooVZtSJD3uHPiFLBZsJYvCYvhbCqATmv74VtSrIwUMfvDGZCDA4vLD8i
IF43Ckqah9eR9rsWxJmDbDYyILxKgvxrx+JTzBlH8a1H4Vpaa13wWkWs7kVQYQSgkheX3nm3JngH
SG5AAWskb781RWDza7cnOEDrx6Z0029RNJT1Dx4v4jiqzCUS5Wl9bScE45cKnLRJpGibdUaoUosO
p/liTXw9UhaM3pBSKm7jyhoZPebir455EkKBd3riAuKFnKdtW6NIvKVKInVjYnTjSMihPCA8pfqA
dJ5c2hP8DpD3brjllnAboOSXh8TGX1kP0M0xY8QAKYG6weKOjt5xVLaLuxIjgYupStkasl9Z1u9C
yu1ell/aaybXEsNdbV3LwiAnrlYCD7kRzfs7qWhEpmWukzvLgNkuKgJ+vEJZqXWQYGr0NhxIilP6
wLQqt95ZRcYobIuM4iPQ4f8F58y84fM+R54FEtVJNAu6vGJRSId15c8RKM1i0UQnT/lhbs+r1v1K
/SL4cp6w4RYhLQKvCxIcFLdpm3S64jqlMNzT2R8LC/mX7aK1bekl7FNRFBMbbA9d8Jd/0CZjE/q5
oeyqaICgf8KmK5KAU8OeVI3aF8gumAp+XK1aVHvKnfzihcbQBJ+jnQ9UGylWIv1AreVz0sQDcEfc
rQdvtyDH8jafB1jeY+62rlP/PIn/UcKxm6IU0RqjOluhFUvr5jTbY82gdChy8Dq6mGRek+Q6OYw9
s3EEfwjE4liJTzIDHZT7oid7iqAO+73ZEMRJF1MGypYXXFr5Qr6h+t3qMz20kCLgBPDNElsphoCZ
bUUpcvrtVp+32/q1qgAEtdNRHMZJnj0qHXi/ajdeG1h0pu1dy60KWlHDh9Inzg8D+1nrTibzH9wu
a4m47nLnkGLQktU+RhDgyiRwnQutFKw43wupMj3CFmVvM4nVo8Mczu9T07SUcN23joc8cwOSITM0
ty94qUsdIgmqDAMG2qyGpZA7GSQE6U/tOQ2GmbbLWUQW14LGtFT2+g18n80Xoc8SB0Rvn0iALGTp
z+7+R0n0yJEZ0CK6sDWLOeWLV+Wu9NbPq1X3ZVnCrcX/e2/hJmRX6J7S9Tk1BebT18v8FISO8zgp
A9TToNovWRnw8ZE0/4WZ06TxMRKR/zpJmNFEhwqapjp+uaYxF/PiKAgVS/NnvTMd13HqJtzH7ZlS
aIN6nTtyEVZv+mUEKS9ZE5TynmUsyaIoGQ0e0r9N12boGGWovLhp9ZFpuKimo6Zg4rZ6o6kWUEbg
W7odW4ZdpMTwFsTZGqpIFNvi1f4RdCoRs8sMiwFLAfkNhasjXbc+VJq1jSVhJt7VNDKKdQLKLQMO
ehQ/G4VnQflG7AS6kU2pIxq4LJABrJ/pbodpDyzkF884Xwf0rGtz5kQ4jJYR4Dih9YRTUVE52EMQ
EDpLxekef3SwCntMTQmJ9mnYWzUb5eChorNLquZWYH595SC14IF0o+NcSTnoUN227p8jxe1TCkI0
4QEoDI8btbE5kKgFFRfE1e+h4UBSXEugXZDKHvEiHo7YXNOD9KvKnPVX+pAsRVwA5l0WJJIzxogh
H+FYEylP1husyMah/lFsRo6VKS7DEIHPmUtx/3jMWW2mrkhMnSgbvSFukgs3LKRuvQS4a6YtiLcX
EeasEGVtOpx0H4TeQsk9Cz3umZb5doHBNlExuC46dfWa/om/o7gdzgV+xGLPgaAdiLsYLko95Jaz
Fboe427/0RdGrNl7WB0Lhor1iYbMYY8nFd+ebiCMp8DOz4rNJ4Y63weg/DaUVTC1nTz8DfqjQ7SK
h3Oc98bfJug9sUFXtDYImTlpTrRPi4Nw3CCvu2MFTJZUKz/qIIn+nvaV3yFlJoa/BGFiJWod/tZd
WUutSjA/dtKD61TIfMeL/boZiv6nSIfnvUshq38sRCW3yMppud+hQs/r57oQdAOZo3Ex5umAdztV
qggK2jiLJIM9HMhMeWPu32VJNO+j2mA7k3YAPmGk8q9+lV3plWxPZ+D1QFfaMlKxcQFK89KZAsPy
IzZIvdUsQUpLm30aVjti2kZwqUw58UiWzhihUf9VhCoBk3JsMlVVuyYRpOUiyTJT+/85cm28gPzQ
1vb2NjkM+UYe2yYZmm3MWwjGl0LLx5RCp3pXGQyUB+FBBeSa4LfzXaEcguzQGbcuVsujUrgf811J
n/OjxMknhfODfMopf00mZiciKtfs7wApT2fJSIfjPg+4iD64VNacCjgM+4Gze9zXI7HLeWO1t0fM
6uJqmdCJZ2NcNRrjYPO1YzzpYA4lxqPBqV6b7mo6eBVb3YCgAE/0IeL8qgoiADMyRx+GV8lI06aF
VKt0R5mS5tAwJCC7ZiYw8vCZNHCRY5MY7OA/XVEUDzPPD7Kl8/s4cQ3MROF1y4UZosw3cdn1eg/7
wtJSspyFjckmwKsM6IthN087YxeVIrRjNyUUG0yuM/7DVOSJ7a/NPZYqfYqDU7t4GaFjGleCHXYO
ghIB3D0XS/jDhpRfd8rqq9ItQ4vdCiFHN6hgcirdPEdqJAYJoCkZGohINin4QWH31kxzvVhL7YJH
1nfYsB6f6WFTa88b3BKvOy9hmKbg4VgufqzvIqK8/LmthywOXeeu+scaaj6U0bkeLPUHVjh6bUQG
2hZYSzxdhyR1dEia/LMGZcFZi7X5CXWcJ2XdcR7UDJFdWrjXs/2PSNv3pPgJqBJUG5BVf3vVyjYl
V7Iv5fMOzv+iQUrTniTEf2SYHfcsZJG3PdxEP9s1anyPc3ELL/kb+VIVot1whQuOBHEcgasYJDY4
w4t48k+EMy3m5Rj9QqF7ZonHcNxeuKHyRtfI4EDyiCaTzCldYDk6EdWkcJeE76E+D/KoQrTdh9YY
pa0xFGutSuWA9W5ImQ+uOqK0vyeeVUhQ3G1OB1R4K8VIq4LTrRNRaQ9yTDIH5ASY/OUYIHRIBKcP
ZkxUxUEKnLLmR+DTDpknpKbu5pueIJCzuC08N8AeYfgNXB2Vy0/+b584X23xluMLIlPBZkgrm/Es
mt5hMEdWQ2lJuiB991+EKCo97Xkxj/6cAdYo1V/362q6Qqsjhuyo80ifFv0OqqmZQal6Jc0Lj52y
7R13HmlOa7Epm0+kOkYTFsfdsHVuqTM0Qtkz0M+aLOTYTEjV7t8ruaGIV3xP6Zp9qOIGg6AV2jgd
+XRmi2GEuYDLLOEyUgT+Pf48irYuK1JnkI3E4RV2YNjzzaww1IZaMS4T7E3t1m/CxK94+N/tj+bY
39jrywrjty5gk7xvsCuUHO59QyagW41RcNSX/1Rzgv//7ICeOI87SnsAVOq45r8MLQGSe8bHasRp
jQAiGDMMoINGuS9Pt4mIi/DWrQTS8JimOOBl2eY+Ir7mNmUkTKBP8QPZU8ddZm9jK52wBTQ46nqp
hWELwsAC4d3xKBnfVdWhlemrDVsUadNouZm2gIp+egDHkGSeO4WIn1pNGPcjYLbwn0lnob7cPgQh
y9Sas+FYDz+YYaSfXY5tkrwr5pci7Qcyt3EF2e3exV8d7SQPDOhpn3KK9E3PH8F9lvV14dKYz0Vh
LohczXosjyXweu7aaLoRfHrdEPc8swZh3YcFJuFdYaD1C/LFdwWe1612jAR1gf/dlBjZqbT3uc6q
gVSHJz3vxXMrdlrUF/6k3uoINdyEZw3FoCROkwLcr/lTIMAzrephR5JpCm4uwaU0fmiiPKLsJK1C
O7RKZz8vHceki2G57HgG2KuNFqDHpJjIi4Sfcc/fgdy54qX1jsCZlpIajytumbi7Two+7qUrh8Hq
8XnzYVdwLSt3F7D91riBDdidvz9gm/LmGyKOFmebOPlYArY8IcAplWEK4sUp5Lcg6tuJOFyHuS++
aFbOzpILkhR76QQ3bidJ77oQ2ltLEz4Jm1K83z+9CXFg2N/aly9wraz8xtVAMFEsIjqHLhP0xEQs
4GJj0Is5BqQTADUTOzWfZRCnYmsemvCk3yAsk5eKJTGDuDHzfZe75IdIapr8EWSGheFYcjBD86Ra
+aSKuKCUezAwwvzph0V4LF52/A6QfDx6sTILlRhyR3g/2FtAEUDLii5jAvzkRNApZu+gPGc5qsBf
5BOSoomiJYSNC92S4xU3nsnZbjrsZngtkqfFw7x2QN2Ko5/Sutpu9MAv5YVGT0aBE8AGfXf5KgiQ
XPA1t1+Mh2hqUy8g6Q5DDEgi5l5izKQsppn/ztH5eKFKAUFOTXrgycpDZf2gbyJhGUZasqcetJV9
pKCm+XxGZj1UamRcDBo1HTiEbsDYho26KupyPr0l6fb+xU54Jcsa3AxFbzNKgQFt+zpOftnkbZe/
ZYiC8lNtm/r5bnKriSWQls2ccbvwEwMmAOuxj8CBYs7nF9B2qsbgoa2sVFt91F73JwaB/PAJ+2HJ
2LfqWQ4r4IOVoQlvrwg0Cxs7215kQ9kX7GqlVxgS9X9Vpmf79E2n3Hr8KlecxORVpKR08/bmvxNz
72EL+y9ErnxJezuwuY3j7QcvWdv9Xa7dH1+hfKoQ9hW+zzNJqYVZIytT5Q3rXgrfiGYztJU9WrxY
trYmHNuSGvB46wajAB+tNIDGLNcI43x/Fs8yP2BdWsv2Ufnz3QxXYFzluHhT6ZpXHLzAS/Z8m2On
ZusH+Z2mrtBQznXtkAsIraCZ5UTyt6ETCM+w/0JzWDiMkAEDno0/dSAOMgrSPzrFeoaDSLssC/g2
o0K/KY4mGK6N/QBo4O0q9+dlun0fuXc21wvjyH1VfjfHiWhXbt2Fr0tWzbRgq/3rCfTHvZzBsKLV
AyyRG/0Nz00ifnKlYvLQI4zCcQtSWVRggqRwLxSvuHZ51O26zxo6xL8WWLn7yIhtyD9M5d3obNTj
q77yASa/nXOq11yjR/dzqb0lHLEpeXq0tn2V8W5TEIi7kX+hWJK9370yPeJJfijPPjEZ6GzrakY0
XQO7VkoC45xpO+B2eLgwsDKa+r9IHWeTnwoK39C4ZVVRtwci1+Fmw27WXQ6C30MswL+DK6sg9EVr
Y5YaQ0w68bi4HeGi2Q4m+rB06Y8NxuwjBVBl/SPivjzZKnLjSpiCiG8L/FIv5i728Ca9Gedk6hXm
LTJtMrFuUIG9vwQS5E4yTyQ2TwicSAG2nxmjn7tVRHj4GfdANg9LWHDOcSNLFMia2QRS8j2+TdeU
/4IEZZxmBfo/8OjwBRW5OrZAO5iZYlTablcEqWxF3icgQVTyF8p4I6acYri3XB/uvst3kAmZlf4G
4q79HVgFjxMVsf1vmKp7ECCAlyqOQ/CU53paKsKpdWN7GgipqX9g5+DejR257KDcCnNuVmjdb57P
h9tfq1S3ocQ8XL2JWmSJSU1Ntyw3nvI9eeSze7KCNy+jGJPSRV6wUVbdOFow/jLAPHxrDbvItE8G
33RymLv+HbsKuMZAod8GGigvsKrHbsqoHiyT165bgb/u3lyynh1rbRH0wxw4QxUCSFKh2LHxW92H
nUUinNG3tUA+CJuQEogyj5ZT/xbnPHKbYJbdHN4Qoi3+tcumjHJJFdwW/l8YyYO+QFnWZGWg3JAD
RETHl4ETyLqO/cr8/zzL2mwfsPZ3Is9BucceKaTioqV7Me2MO1WxoCdXf1flqHoUdVLNyvTRX3+X
GZ9SdZghJQ1Nt5gbmzkp3nZHHhb/v8xGr70VqKBTH4IFVWOXsd5JqsH2TvBZC/q6kDFiuOyKk7s/
W4lScCG1ZjlRWYYvJHie9ff2ZxpUkGf8e31Lm5wrLmMpbpI8ysz0sHR4Lms72oWyWCDXTKrEIibN
JYAAGX3NQbGKIow+BOix4pGs+bl3JsRGKmj58rWob5r73Ha12zN8+QyNYJWTIsFRXuflRn3mPXBf
zQXUhVAz0T5LwjtRK8eBVvVvXlPrazSpsOBx6euFsPoB0osm3JMY7C4aWKKr0xTuBnCiOSVto3Ot
d7N293x8qIJa6OUUmh8nkrmE4iYRTivFQdzsI8uoVPa1ySHyfPYKko4nMSs7m3A+D+xiZI7YHGWm
UZlH0ncV6xpgEFWwOwTJYdr7SHtcPw9HGS1XhqaNsWzFN6jb8rhUYixHsKhz1z68dLmuIyG0RObi
WkbPS8k7IZlVoa0psVjvI3i+l3AS2ajmqoypgy1vV9l9VSNG2Ja/0OPpK1P45WqLmMj9Ew+i3keo
4eDTyk6dU362+cXMi3TamtDHHQh2XZU4bR/rbI0pE6oKXnNN0wU7rjC0IybMPQxElOjqKkuCLYLa
taKm1+i8A2e9fqxqy11hiGEKkjsSlDDaMxl7i/ORioQ4n/yYbvPwE7qp9YJdAmgZ7LagiZnxenea
Bv6MzLGMscqAeqIbr93pi284egskXygokOP7Z/DGE0m1eQ7CTViGOO8G9RJ+i/e8axtRmfkMikPm
BUqMT8K0cNmfZKmwm07nkMD4SWvhRxbvx0fsTc79VTJhmx7s8QdJg7AmNJ1cdp7fLRwS/5xbUzVE
Q4PKywFNw0W+C2AIPLwU/6OWdVckGJwMwFOE35PZ/uFdSI21qnJ5D13bI+qKRt5JhNF6/QEZpZjL
uWcRxEtfzSq1CGlT8C+9+vta6TufqyoyiWDs4L/76WEdy6HryonJRn2ebELPPk0Z13Mqj7cATz6h
T+yeG026EJ24ixUBvp1IcDavMEageejiehbH7vcxSd38N+5LXGXpRTuJF7FJw/p7Gq3cdLO+2wuu
GN7LCgJjpwsKPvj+58VAj52ReFvIWtNrbMnO/e92SWS/IrKwWyzjFCJMDWvFZibtGxzX7Fcnnb9D
/dxVieqP0cpiQ0sW6VhZ/sCQ+DYdObZWojjuLqjsLsyf5IztXUvB0nF9H92fpjqAIVwFEtcddqfH
yWmTmepBzjBaIXptufx04m4R2tYZmBaHRqBGPLufyWPXJ687mEmrrAPLEAMgC+gIvCccjQiGfP4m
9YqeqMGwzOXQC5BorTlhOVSebYMuNuKgVRjCNXfLqNHI4d5uU4IoFKPjpe30w/GbMMnKWIV0cwxo
IxWvwzEC/0n6argqQnoEDgXoJskboT2LIaX+kggcJYbUPE7OQkAiM6G+K6p7l/qSf6HsjwPNmJsx
8cedUe2USeXEgmld/yrPedofKksP1oYQ9/CKuBoHUprFZwAXDimQNEJRdIx2yKE50hZtTckvy8rs
8rVNFsuJ1DQlDF8fI+J515yNvYbmrjJJmLzzJ2N5DXI9/A0oFyN+YPmTcjT5ABxWVzTbWlod18NV
WQZc3Ojoce9F4n9XW3ZY8d4NiZ+XpEJ6e9klfum/rqVDzrcEXL115fyiwr3Bb/TuzX+T0pNXm0iv
YR4N9OcD0cqWndU6ysxSTPY//s5rB7QTzd1y0fD6Er8shLCwvOpafPnWqGtXoMWaU7Ta1Eovk2Sg
aEnN/ZWVqGOepy4GQ3XQ0K6g8u/G1LFDw5hvE3xzCBfmwXDrWO6eYYfhr7C3u6ZuQkTapML/302N
tvoJwq67n+j0BM9g6YNWd2WzmBz4+9Is797U/OiPKuXTM2hAOncjakCxmTHiys+asWoXtEl63xcm
Lul+7xbMBqUB9SoQvbnlN7C5oQ1vDc1rOQWMeceYzCQC75+9dXHlD6zdglEY00ubd9xvwvvh5NYo
K3bk/5iBTcaciwulsNoPA4WcLtV6b0JxGO+PhHtXBF3l9l2Ts24s6qDBuRYkFx4C/7EJ3dXrzBz6
ugETmx/8OWo1OaUjyiwh6i1G/nyrTr0dU/fPtw11csVuk9bRrAWVDqdmxLVMEzA52YlRRXWsQvsh
O2PxKUuzpKgyWgC2pTG2HW9J+XEiP4OL8fpNSznJ4dAEfBDkCm9FmLBhxStcg2JlCj/KOqY2WwLr
zfiEqB6qzOZRt8zJoAwQY4cmOgtHIyifKQsbeQbeoER2eqIMyRNaFiFCBrZRbNtvRkVw0DCu3jg/
oQ2Q99VIUAsQhgnfran/mXIMwq01TDRH0XW26OKXQuySQNDotsJ53/4YY4YV40z9n1knvG49aMHH
TOGVGTXl7PhNPh5rcfSeCRs9jku7GRztK6OoeVSMF0jYM01oPFagtUeEEWayiGX++bLJ0MviDe3Q
QBy4HbomFo3V+xf7XdTwf+TuUF6oqw6mcMv3Es1rjfgtlfYzC27UTs3He3fak2d2FIBqYuuS4IvD
iMM7GaGqsbL9N/dGylPEcyEes4g9/IS6/Xrchzdhxr68J5S6RZxFdzStf7MNX3N0eQaZpEQPIXoj
mt9rlP058fFDZx9gxpJ3S676Pmx2zkf+fLe5ItQkxbykJi7OvxETXzV0DvTXdoWZ7Bf33H2FKIWz
VJ46VZaNRK/QQ/LQXJgL2iQJcotrzs2RYNKilrerefyjz/zL1qwGutAKE72ECF/8Km85tfyG9vwL
WxAyMHAmy8Dp84XdmZbWPdwAXEGKmiMSVYDo0Ey8u+Jn145FrEC2KS7nrTpjZ83x06Yi3gxo0PWO
ucpEMuxnYlHfbthi5PkZVd6jWUqxwNSQ3NPTJW4TNkuFz8oTwc4XqRvpitCbJRqABVHG9IS8qfcB
XAspIAtSWF/NNQuCPuvICsmEWaOfZY1Yi927RNhg0A2PTf9/ZC2q8s05/a9y02QK1TaXao+QkMmq
LMaQhiTjJOVbdkAe4yeWwWVI5i2syN9weaFrLF3IzIDaGfqKEMpoYTkLS568B1aoClzC3KznrDkl
CCMc1aQEV9EknbhcJc6rVGtgiPOhszXFow9rtU0d/shLs3taVNwuLHE9byDZvCBGAGvypnhy6jXr
ynkdPWVTiZuqheK6acxamDqbBdNRdoQuE62AxaraqAIrCsG5Sco5K4YpPv6XspJO+bvOzbHkz0Yn
2j2b/Qjnz1kttBjhTR9p5/14MdWK7uHl27f38gKjCu6IFjYOD2SAJJzkArHwzuLp2nBh7hM6lwko
ybaeju0TtmIb5zTwNMM/9LcB6Mth3t6cKFKBWkXKm4Yaoh192JQgDraDSc5530IStK2gEPb95QgC
QUXQ/rA3QhMMnYlcNWVpkUs2O7rXaZakoYKCb2gz8UIhFgR/3jn6El0as0cEj/iU13TSi3s5GcJf
TNMUsiYUN4EvLvtrx+y9gFH1UM+Uk37g2wFxSr2L3I6+jRIg9vfXn9fhisZ8kI7KnEy77ff8NZZG
Yle2l8LS6v88n2On89AA0ljnAUWEknMHzsefHFmfJw6e286bJpxoBo1E8WwJ+5bqOwO96Thkq9Hj
vZ5n+xPUspazXYroMAk53Jj3k5x8R9T7fVxDl3VLpqnfvmfGsDa6o+ybhK6qv9f1NqiUk8lREZ4M
cocmNQWcPhG6KLg5r0XiLUZDCUNmmFZ8odcr7zQO0OZ1E7J97D4udV/WN/P8gFenf2p1T4B9Qpf9
isYGhFfsHcLVmjHyAWXmfeBIPCLYEORgxC2tYjR/bxFAXlpf1zdwMjWQgJitG1uxYjbza+aOmdpP
EC74p+SGQW9ZN15jPacMqDr9KQ7a8M5lSjV8+tTiTSdnCozKQKHPUGmafRP8eKLFTamO6QtnS0gc
Boikh6NSuDWs00bGtwsammpORqM7dC4022wsXP9epAEC62nES8BITDOc9KLasMRroRcnM1vEOikL
UrCVfAXP9F7C4Cklmh/UZpsL1X2s/kIHWbZ+lpJ6AdSLzS3398V52eS/ekaYyNjlcVcV0e/B4pK/
pPxhFovaaU7/zcxF85LsW5ni8jYcA41gGOioqlWQtDikmM9MJAeU9wod15OsWKGOgX2/gfk2lsB4
4PHV/SN3gdDVV6KmR2cJ1v5RfU5Yq7ulRmH5N5mly3yRgdfKLgdJP3UDjo0V/wQNrE5PHDL9JT+S
rrnhx4YUZL3/lGQHmRL7Quaz1brXpKFjqQJVjckNhD2VJMOHQeSd8iICxi4UyiyXi1/fKqhHbWza
DshLqofeLQsGpNYqrfUL37+amhZoIKeKnq2JnwtRU8OWI6HrqKkrwWLHaGdXNBLvaDayMZgoyI50
HIqRVuVvPwzz/1LAGWb0h0RiaD/WDIqwFOvNR4N1AYrWwknacNGO8lczUi1hU0WgwnJCCFhRCYtq
2hRNloM3fr5pKRiPY9Qr3QhGYHikYKi63f1miZpYo+fxPafvYYCN+XWsGfXtXPY0rkcGly0U9ouZ
uhfDhS8b80lB55ci1A0x5MHrdXHE0cpW5/94BBAqPTqF91Mjm7UbZUXwQOGD2OJSZiNNAnxJRXL7
kBLcqKhtWM+Ew3lB6vD29IZZkgCSe/x1EsaMeehM+oYfHSabTav/JW6iMROMDtm1HMLDJQmGsIFS
zGvCMPjtVT8jQKt3a4iTUSGhEKfY/JpEyZQnCnb0gsxSVSpkA2qC7F38IV3ZtlCYZtk+DJGiIOmC
k+1AzA6/M03YYn14vkdipHB1g1/fs4t0mHuSUOALr+UOBwV4tr8EsbCrYBjPNwUjKr4Ye99x4Jza
tFnDeiMwnvBE/R69O40ayQZd5ckZfud8KWlfw09AnMXu9LLeYtzyNj7TGJPFIVDYB7M3h0XdakHy
R608QucZB6G73dprvaiPqmejs9zReypJaWz0u12TQ7NCTyxm01rS/ckzFMzOKNCMFukRKgzWswwl
4K9Rzk9n38OH7Dn6RqDPBcv90lJJkXrS0r7ww/sdEG2YkGIpUHcoT6ek+pUhycXKADX/dtcoB+id
wcabG6oBQiCuEHVJKyr6Ea8U+sREMpaa0bBbf5ogfHX94brIj3OL14hNySuAnfr9F9aKsxwWECV4
kvBiliharYC65yeIwc0t1xUe+D+swMoQVAPk9qPD1Qr0mQIecFTXcqchXcUxq67YvVaDzVEbf8Su
IYDOmb6sQKZs/u/4Y7nBKX+bQKs4dIX/WBKIFdVB5OHXypBx1m4OCMljYY/LjQJP+nBCRlAMUN3p
61YnlgyVgdFooe+R5ARzJ7rx4V8OeeEiN2U76dvs+rRIZ/JQPk/PCEbZnX1v/gOuoxE/69hBkXwB
567vTYVZ0wRUxJQXde6klkEogd9D5mPVlzi0CXpgHHBp1XKtByJO47SZ6mPmSgluTE/SC+bFS4J1
z3k3pTkZ8hX0hoUBrWCngrSAjRhv17I7RKw/fh9Ue0xaWdXQxKpYqXnK7rH5Wwyg/p1C1BIapFqK
VAIiIqk6czXboOONAicP4j0iHgDYfry37E+ZdY4BfaGZPbbZ0ejztI0QSlNFctfcMQLXV4T6mMOP
dES7x5xO1BC1P8InCPZN3X9wPuib8nou5TfB3kZcMu/PU97qh7kyalk8Lki6FTk11ff4r6gKJcRe
PVL5c1Ap5NNH8RqTEO4BKV/2te4n2hNXpKYp/8CCbT9rrlwjfmShdHw0tKyWk0mpK/jFWv1s/FbD
Fhb7mXGVK/HQjqgTIHbvbiF6/0NwE1YazNSdrXJJXc9MpsLV4f34JE/bCBl6eiVgmJ3+H2sKh+bK
j/wgGSeZTOdQx2K1BVDJvEDNtcxQSHJ4HQ4Guw9JP+UBSnR8E5hToiOYfC4uRqg0r1zGO7qpy81S
F5lfY2u0X00rWS9XmzbL6Z9xvntLOFXyGKdPOQKvaJ6hGKxp+JNDb2GNpFLNgFEIFxUaBZp0/Gxu
WnKZrcfBEzi152c4utA6iqZBlZX0Rsij2sw5UmVgRuXpM5FORk3lQitf8gtVuVYjXKxa/XTWtuja
EyIfwv5v/RvO2Q7uDIQu9PVq6ahE12CrPS9N82LfXk+KHut0qqDYli/jJNBEOIFsBudPJuU2o1tR
I3s3lxSYZWtQLBeMs2UhVgqBySMxTKWs7I34spCGmTDIsVwpaNbU3ii681CPUuZUL7BYyL5nwmen
sR8RVBik9gg8BPuLOhEuVV0R5FH3xsboKKX1zwKGgKEskBiktv0hXfODHKpt06F1/R2LYemg5/vV
lZqyT3dAgKgyg2foLtJpbEkey5rlTWtDz8aWbuWpW7tcY5TeamSB1bWWGBrMYNLy+iYq+S6PQ96Y
CeFMwYvyg8as48OLswrMO+pZVOLV5TCaeRA3WyOkUPYmF+3EJq+lvsdb5MTr1OnQHFSuF4occ9oB
SpV7S8bNXNSw1v6XRdikvBPMpdWcdQ9/I+ChAjEoB1LXGiui3VYmljTPpqoDCpp8zjutj11nc9OP
MSOlRTHpK3rHUIpdgofEaUqGll6cwsiALCymg7D/WRclPe/qOjc6nUad1FZyOnByYwwd2em/SIKr
hE/4b9HLFLMcaTHWvoOp0EkxKrDRD+QOvzVynX+KsnnDraekGht8YQsllVjTbWr6nkbibPlE5lwY
0GrgRuNXyS5LFF+BHInuAI3OY9nR540CcYchkjQVUX+58u5wZIkngjbchtZLOXt8tEPcgmU3TOGi
Jd++sEn0KtD0xJMjOtwDDMK+RKJc/nGGEX6ZzMbgiTljdc0Ljg5+VXum30jWDhvK+CqB+lVhcYR4
lRNWFGwKkjYTgZWaxN5zreCCNR02v8piGNf+/m/FJV1U3MViEqYtIVf56YAclalwO5gqCneW4k4u
ykNkt9jOhORBQ0QPcQ1hG5ha7+UIQMv6GGAAgr5zRk6eSBNZeVy4/CKmGzHvZ4lJm760b7WknVHj
/BjX4jPkeAxSvUl70Gsk8vU7INfMBR3AoPRk6SXWLtpo0wNd+psKQg92CWsW0QVhVzyRUWooN3Pb
n1R7LyD82bgDrJ4r3l6ak8fAdXVdxV7CH9tx9UhXeDFcWg4xyqLXqPq8BCb1aQEyKXPQPdkRb6Th
K1llCICHTPciRlk3DqCCB94yVVtVXqNVKyjq0zDsoWvcv55NiHsoVXZp3G3UxFtg3gj7zh1zE+U1
nTBb7tm1MdsllFnR9dnjFJL4r8uJ0JpX7UxaLzh7DFximotkU8wy+6VSCEXGOaH4dNmtQfzYI6Hu
kwhtKY2oTFPf8rlMMSyVUNpcvug1n110ResMFrIVF83G3dMyWKCFK7s1Ksm2Crk7NPjlVAjONlhk
7XYyDyMyRc2CiW1hWNW7bQd8jIA/wr6BRbgaxCC/Uivs6hGrr6XvLtLe7F6R4mKQeUW1D4K0DsLa
9RmPHliAjKlhDCZcn+HcE6TpPWUPE+eMX+0Hw5GwQVbfyo7OpBI2gcl6jkE/K/iAWOYHFNVY7NKR
TCR9ywqWvY3w/K8uXB6eIH92HR3DplkS/4S8lrqI5ouQilallbgexur8NJ9xgUgla3fnf4x/zgQT
sTZJJsrTsJhr3ddKcZccRjFdKYunjV3iN654hsKXEihKaXQs34YH0ejA8SW6FFovwBgX7j795Yl8
xeEY/szRm/ulmdul6WT38YDjY1BH3YXwnNvAOwhQkjvpkyQi1lHeOCOUCu7nms5xOC2EncbFWsnD
dImOLrFE6R7rJyX+AbHAjpRz3ZXsMQtMNZIyewcab4XdY7cWxPTlcpHoUIbQcVldQyHoxDAYgKcm
Hl7WbwbE+SZczF/+fT7ecgcuKuRvu5YYLk97GMWI/wUj/yxmZSr9Vrr46qhy539WxeJtdgYnt2Eg
tKl7HVuGiawFRYA6ozI4pljEC2DQkbbAsgI3nK4q1vl0Jeiapm/OgCSJUEsI1S0lwGliv/YbHgCl
UAEEZM5SNDsN25nzeV5A72GoWQqOtC7NUlX9LJQIwxYF4dEEIiBApMobtM2K1S40ddIwrfkJKyFI
rOG9oL3WvQRlXb7lBnT86tCItO2tdI5F5RcVd08nWAKJ6j8UQPo5ziHP7MGcD2vIZMoc82CavNyT
FYw0ARUPSr3JZ/2GvXnqkNx+5qvaOpkJFqBtkitoa75EhBDehu0hzcb1o4krfejuTfFGh6ce2hd+
GV0q/ozlGVwJWlOkXcLhBFbgjl76iU+Dg+zJzzSICUNzUjpwE1nnPXVwtSjUKZxoWcDvertiXjai
zyAmewDhVMSQm+4exLHkrr42CDq1lRBNpssvJmTZORguzWyVFfJ34Ld9iEfDbCz57j6eR/7VdxG6
9SLHkeebTdNWY6eKtVc8R8s/TDqqxDwbD0jn5XoMTQ51bbRe0OFQ+oCw2VLNF3YqTGSwd5h1zBcX
teubhBSGk0ea9b1/C/GnLMdrGLfUQBex2e6uXWZcbxqWvsHjVFW7YZTKLKNQK8OavW4YrZeWaVbz
eAx7d1RWTgRyBSndK6TTgpGX8Sman1X0jWwl5BK5eHxhxdj3nTbcrNV2sZQ8jNf8BxWNm3M+gKjk
4wafVBFRYMiZsyGl/vg8Sj7cGxxjjHqIOroUkFGHg16K86y8E8PiHcc5R4kvZnnpxq9Y3o9Ok4Pm
sRuCvr+Cf2K4xuG3HnlQFytkUVxyBg5BCz26DwX5zYRCT4YDTi9BwKlCf1CyK6BCFZfOCotDZmUM
beJ11dpayNvhxYqe5h6aqARmuzeCQbdZknpesDsZW+F5xOolkt9WctJ+GVzn9yaLr/BXSesYhQCZ
z8Hz4WTaVE7/FrGmoEFWEeX/Ic1dcE314fz3AZS9l4XshPYIrHV8vhtK60o5eKzWbPeFFbhVK6OO
SZo6uioVrqNcn2TWB8h6STsWdYZpRnSJKS2cSZyj8NYCMl6ogx5e2YUZUeaZQBs0k21AZ5U1Ylmn
+XP8ZOLGW25rbWUMNfB8fRq8p+a92NXAKSUnZbczdF6tZve6MPHRR6/LpLf5ldEACw2ibQuQmiSi
OCTEP6mr+RXoV14Vo1PktDgPlnV4dMt+X7v2bgovsXE07RZIL3ZvJXx5dUqRhThSsa13ebyP0vnP
YiVdjSgBVPRB5SI/7ZTBu1eAfbcXxkRKc65ozeG1BvT3CEoSZtgv/P9Eb6j37gJ9NvnQVuuv9QE0
DlEcgytvj+76xKFbcUzqMvzumMKb+3UE5mXVX8YNDO77hnMSE2oWz4mSuXrbYoN/zUDsnHAze66C
3n0Y9153LvU2JnSVOqRO1eMEfXR0234s1l0+dUfDg3Y4eamJ5Cl9mT4PrT4pRIjpRog27L5yDtty
l9tWPlPFjW5eYqiGH/U6zBLlIlizArPyWGnAUcd6SE6+wqZzqholtFZvwWm/JFz9/pYiXIlWJ4py
i4GfeQ0mmDFFBM87GfTU5IH7NkPTFgErn/caW0ESdBJ5KsKpzeYg7iutYauGvGaXm80+1UX34jl4
zWMJFX/w7uEy2GBQg69oyXL/n6O9emtV9qFQFH5QMgvwjDpu2x7s5X2BMHDBS9dPAIqZYb5G30Uv
WTV9fzOyeVUWD6rCy0zm5uHafrge+QSnQlnOY2j1RQH6yBd5rwMlmoB35iv/RYe2w5Kt8N0UtPUT
FMJN4C6WBPS+qdHf1Yd9DPzml9qwQtWInT95ajhe8PXASCDfTyTRsLo/MP+jTfzzxLDGk/av+k6a
lRs/UpgwZrKso0zUmoJ8hX7ofnnLke3EGm7NLhJsBQvxyIm7+BW0mrmDS7ok6idWD86/r0u+MtrI
pUepS3jiClxT42Qh4mExnBa3p1cxewZ/glvPMRD2YSboIPiDpWu3wlGjiL+/BfPX0i3XKuNxKDhN
sQ4b8nIevL63ZLIDvlctRVby9NHocy7jEXZJ/SYH+P2UdnHx+jJk/G2gqM/DuR25V7c94EPbRq6t
aagI4rqOn6XeMce8C5M+6hoUFctZxCU5HdzJiuqOoKZAGyO5TNQJ5frahO3q/MBtnqKlBoPlX58D
Nc3WTxkiPU0v22S07R6E15HSUV7IpN/NnaMtYbaFNNbDqp4zhlJW1lQrl+xg/TZLE2Xj2MUZaRNm
vxqsYbk0o+n53SOdqccgbhMZMm2uGvkt2XmdZdSI2WxRJ15OwY2hKNGxFLKJsIUB0ct7bag0IzOc
wxLN82Q8+nwEqnrEdc7Y8+bUXIK070VeR+eQMMzrJGIDbRils3bysrE6vbzrPO9HicM3HQcuVBPy
1LIXpf7NqMczI7oawOTvKUOVPSIgimVdgCbFiKa0YGEn6lO4cZWX8etZxQJ8BKQ1WAKQl2G+czJn
A5nyFvqOt+sMB3/nWOhscJrz/bI4z3CXiqCOmRdE6JMVoXrg19uOJ8xV23kixssKylT7ueI1OxKZ
VZOxhnvkSXi5DP0x7FW0kV+AeFQwBykJ+rm0+sgyvuUkqAk0nCwbHA88u3/Cf2ecsoMgnE4HMB9U
3WALnw1HgdFo1b/FMyJAAh5sPmqir1dkYn7kOfySNyICo7X5T6rSRcvQmHXHsxrqZ9SU8OsMpeY9
Fr2xHaWcBZdje/KS3t234dJx0Zh508AIhqAnnPJvMyTpXg4gFbAhmMP+yAGioMN8uJCEZxIkPe/T
EXz+PEO2e+u4j4fZ6voudXC2DZ4VD4eQ94CIfHCybrSjbVuuwyNiE3CeQEGfRyr9GKajuoIILcnZ
1+yseiswMGxqs1K4F4jyulQO0dY9vt4ID7fbroM2Wt9y6tqTXhuy9Setuyx0gz8EpQ8m2mlbZhr2
mi2rWwItNoWhmBcI8P2SY+N7PzrM61JSgXRyNN94RWZT6ocd0yOQL06ForwIlGfXKZaLuifjolwZ
AMbtqDZ3nfAOYGH3nC9SXlHhjhUrsi/1wwhCE/lsWyNSil2o91J1hSg//BLL3iswGXx5Oy4poHyy
Y7oGGXayp4nDBjYsvu8epe4szNuV2hMrlRLxHlaJFaLHuyEhOeHns2C1Oyqo3bldkcl/nq0rhvr7
P1gurNZ2TWYx6tIlpEOcdRLbgKB4+aFzHs9oJs/24KqhAgO3eMEdZ0ihyEjRlXUIsnPjg7UbBWzf
HIb+FkmtovjUES6WQkYPTcGulEJFIsOymCCYQ7JxKc1QbQDh4zGKf9tONwer6Q+jWu2VFV6nvhWM
kRx8rrHQ7SrNi38A+xe0izOXGvO35Et6CNEcHZJ4yOkOYeVaRwswI5rFvSZD1Usye3ta6/EKcTrs
r0pEa1bHOsfeMHEEcYWYMBnhOFQG2HUfPZ53JVhecru8LwqpxWhHZLpL6NmeH+E7CPSVeqJdcBu2
pyCu98eWoJv0+/SnXLymZMRHNNsZUXfRZj30PJMAqCTgcArhONwrvmNxLclcbWlDiNHjGGH58YyL
qirVVPi+wj3TEh0Oo/tw+KTA4rw5cFIDQVRQl0GYETQuTIwuRNaEWrIvGj0mDs92bL/9vsL8i+/a
gpSSqXC8aQDkbIKmuP9dyelsdx9flUDWpCUdtj2wUpNHEZjQkmpIGfUXQ6OF9JEQvmk+t+mpWRKu
Jch424KR7J78m/sv4rWteOfg3rstIkOlLiL7IUqK6hb2PezgEQfTA2ZTE6oGCFnJxLy62bXNNif0
TCW83ZNXvUiWcrxs0XYHEg4p3M6zfuhARl99D+7/QmlQt9oATWO2WWLDrBMZ6iorLEiNFoROQb81
17J86461mjB9/PFuul6mUIw533rB7qZWSVbavbxwVL/rXRr0FgoBAZuGv7sNusuK/M4lDapu5ZzT
V5rEZUae8KVxJLxa7AebUZo13Y9X50ZwXURzn0RrhnFSMwv2EswuRDL46emy4Wvj3qDDS9jh3sE3
laQn66GV/eJFl9rSOVefKNaHZD+IqhMNqySru1D0xezOrREChua8WPleszbz31KKfH9QSNXRGQC5
U/vd6eOATPrSj9dpwcYbrlF7e+chxkz5RXyaC4OerciKHu8msp9rds8DLcZ3GPjLlAx773F3ExAc
sXjh0SEkWLmiJHa+vnROnHZ3RXQx3bgV8EwMgUwdpJeWkWM4EbaKfj7Qokj88RTKUy26FoGZjkK0
MeIN6mU69JcR8AP7vSgu6PhuSJLkWOzncOdmajyz4RBpQl9bnfd9lY7k8BS/tE4GCAfKY0KehvaS
m1q1Qx3w1bDocnKelaQF2KE9M/PXb1lvGo2G6WA90MCN3l3akWpzU05yud1pDvF6qHwpAi5FcGFn
/Prb1RAXokIV5aHfegFcJG/SlAlJydQxuupeD+iY0Z8QSjzqtQ4Ipdo3qDOnzw6Lm4FVPW/y5xzz
q6kRKfNZANVNWpP1QhM2xE0CMJhOQJp/8Xeq9nB/kijOSpu2hkAI2Hw5CBDqvicPPWyyegIt47s4
ouVU/lxTT03+jnQclWUTqlwqw2I+BIXUk/hIFOI/YtPlIkgjryMxZcbvrdj2OHfBiyEodENmbUKc
vgmPyUDrMhyMrYe/j+Pbna7yDKxyhtYSEFskDrk81rUIYGuZRoF5ypT+nlvtJJ7XsTsR9YO2NzVi
fWgYHclZq7Uhbz/vP4Xf14NNSRGeRTeNjh+RzBjlrU6Ba0vBJTEF4CjuylIF6JRHY8cTwepHDkDQ
nUI7ZGkAdIBsGWGy0LPx+IEjNcrrddEBeJkG2fP97j/4uvxspM0z4IgKceYDSJlX3FWTwdJGx8Sk
FdNOv+P/38QCks8Xizw/UdUc11uEA1H12MYPLNgaZ8eGcuvUe5FU5Hctk+5nZ5QAgIeXUxyMsS37
CFOzJ37mAUIapnihiYwAFnPIGKBhu6HyStwrot9bZDdc0S6xZEQ1s4mKDTWTyyyiVQaET0tHSRtg
cllv4bjLk+kmYFLql9dvA5/tY2dGN0TZguK3AjkGpqUsm8izgy2xhkZSm/0w+blkESg1DXZVF96u
m5xoW9ecZy5LaddrsANxyr0AM0OkZDcvzAa6F9sy0mxzeDE0GVURW0b7Lkct0LTaezYuL3NC/X3q
gdFanl4ZoP8HK3/tVo+Z12mUMMZNr0trIPpIBcea9V7mi8wA6gn75lAZsASb0nDCVPc3uedCykLe
vcjpVs6d8qUj0rPmtT+ijgz/FMnaXngS0Xwz7v3XtyCh0QhZIHGi4FRP7kMgONaW4ZxWF/B67irl
IMWD2o4udSE3kh+1+GCj3e8m16GoHJuHSEiLYjYD0uO+MIOEKqqwkGAdLcvrtjd1/siiy24HY/nu
vKvliHPeLM1EIof26JdZVMhiVQtWI1IyBbn93Vez2AVhaEf6EOJDvJ2zuPi/0y/Tejbapcz3o1b1
sDyZb6s7CUAF9sUXoYWwGs+Lu36hogFzp9SNNLruZaLwKZwamJuPHcC86lueIbJgYJnFbFYXsBBB
DruY5GiQIodwkRZeuj6PCWIor4rgEVJpn9oUvNUZ4QS3YdKHpqapYiJDLNIDJ1gQtuNc/wtv+wKg
ozlj0cZela768hFPBh4G8w19v7u2pbD8vaxprexu+B/Ptxg/K0N0uW2GF48csQaK8Os+nOCYRjBU
FvlUPt5Y6wnOR2XFKAoo0Yc1oSSAzNvIkOTeKkJN4qEOSRuh2qFcfXGMXZlsczgP4CoBZR/pULSz
Jt+Z3/AQ6AaEvRXAoMInsvZVY+LKDtkZFobeIyX6yG9DoYHy+F+rN+zz73ElE3vQb3dXLP87tqCY
0cR8kc6Q/gowYbpG39wSs+2LQWNHgA+oate5HcetdALuKqFApaYI4zJbzIh1VDxm4pG1gBvoE9Ez
6xYUdvgkiRqUhY8QvmAFXtVS+4gIhcv557LsBlhLdvP2Nx5ZIGEMnEYZD72RoLOXb3lPtt9ExOa8
i5uqG2SYho4a7xbbUsr9eOOpgxGi0/IdzV4H3Q+Ga4YlaaQlpzAJ5BlNZxofpXiambsptWDvgs6A
L/i1/DLVPJpzhVMeacp8uekNBOv98djEPhGr0zzYl2k22/yqJOY3XR5Q84411rLrON+rjDCRtqlG
3uw4xPW2Asen1uS6rjhF306tWqB+F3C8i60cQhlXFm2fhmBN/ux/CAHAirKSY4BEnV1wjYiX5buc
+80sl6fPPgrK+waQIumFT9jinYIZkgYrjEQx1ZiS9Z992gusNH/0ANsx9K9CJPCJS4PJUj73UrKv
Z5cD2SyocTXUAzPNsNsud4g6m6LVC2K9Xj6OHq4h64HMOdB5LIBhcAytUNenMEj1zeLOmZp5QHkO
eKgU9bVkTvRmP09haMjlKJ7HFCjtN9A5etKrrTgiRuDMl9bxkUnSqvyPmLgHzpLqWAEEnoAkaXlf
T0cfEa9esjcmfTQaVD5jiyOVYTgIRn22HYIUPGyAajd8/tivBnuQHLFAfGgMncv82bW6ZJ2mC8wa
pb+Zkk/+sW+kFTIIh2PTfsTrsb87tdn/BYmin3a9yA1PrmmMlupdycjnk77qCVP4DzygqxvyIr0/
Ws3TrC57PcFyfLbn/BG/mokzVXdNc9DUklfrxWvrXOoMWvKM84HQRdZcP9ITW7BqjrTh7+oYbbxy
BlXRJrywX2O7oxWN15KnyWV2h7HXTDlODPkpc6S+LIu6kPfZ0wpf+E/h06Rna8HOTwowarD7cdFn
UhogwCLjmEo+bEikDOUfYQteQuB2l7+nGYhCGOYGLHfoUxeJxa/IhDZb3S7NgUntlN2MBRq/3EX7
l/ZuhhgmD/a83RGbpLO6C5prCU2QnR8sLfJr7U7lxL/S6DpONQ95++j3ls7FVLP9Xg/sfUNwiXYE
nSlQBrw/NABj6+LPIeySGKQVHz1ux11d9ZYA5SJIpRXe10rnXaMaK4wvqlipivHg+fysFexJGbSL
1/BKQvtRl58S12sI7JEOBMTBPrB1LXFWVJ6tOzQ1IVH3ynpFlgYTYW6NrUdtSgUCejvnMUL2LYQX
bAcMv+CgYWXtjJPyNZyKmq1cAKE0POIQg/kB1G/R8cQVBpWseARoUEDYCjUpfvF8eO/48G8Uis+t
WIkfIp4PPZXOCvr265NBcRnDd4krfLyODqI3G2/TXeWr18S2WRg1gd9oAYvVd58F+wrAMV20Fcy5
a4DVvYiS623zQcQGmZHEaSr0svatcWjSepEVJWPW8+Rw9VMQhFUDDFIQMxoBfaHGtZTKM2ZSlOw7
UOFSmnqO7WGyb7acVytJYhK6Us6sXRzSrTEXv0aHZsCelxcLN6PsBCQnn+teGS4tvuqcswGoZFZ2
8BrQEhcRJBBrMsU+irTA6Ccx9W9E44lr395aa6JYPCl36blq6tsx9T2p1ZjstQbsDc8Fq0EhC9GE
3gw0QDZMlGrY8O01vRUXrLiKTyIKMK7rQ3LgrqY6jiwTjzV//cIGDpLVy7GmJ0EqzS+H1QXcOUPh
9dgFiCyfO37q0C0OWlI6tBC+utfnGNikaM0hUSJTlhPjVzPOwTKl31LDP36+sRK/CXvtzTAkVXyB
khJe7pzpzo/A5etPQsajHkX1qssZYPPvUtgi0jEScT12+/HHKiOcZJSF1cwi5lKKkoojh33YcfVJ
SjdTkiI7ZeA4ZinHw8zqWRLDSZaRKojdsqj7CTbZtk2n+eNydPtGfbJutusr/uAvQWAcHAQ/UKX5
ni49OfRw/ORxHpoJHVv1A2OAgBpkjyu9GbjD9IM+E1b8xhXPfHA3lCoQTRbX6kTd51ZPIRrDfDZs
tsDaGpMM6a5Kha2uinVggeoB9S67gQyLxoGCVHr9SPQDjhjK5U/twhgMDc19zBgtgiNG9QSMqp0p
JczC2sYuxeuqKOB7s071f2APWqrWb86b9aSAZxGQgAPolb8golvEamXQsBtX+Uey+m74i22fKVHl
39IK0aqtg7FjWaIGfboxV0GLR+mtuDO6IMfNPHhT+kuht1A+yAfhJvJ0fVKRnaZMjESQ2BQMX0TB
xROe4CrirYwL080f9w8tvbb2PahE7EEegkmmwlpaq4gOEMqXAd462ijooek2WljhmFymlkGoVZf4
l1rUbHCj2LxeRvFrjhuOXF4KkHwxPhrUJM3iSopDHshuXvEmqan0EL1+aaFQg+AvO8yB82MwZKkt
fBr6eL7rjhZQnh+oF/qjq1wK0aHA9nyiuO3WbZyBUfQdt2u3+/4EST7gFUkre3x4UU3oaZivWwHK
ZnzjQaFM1qyN73h4tQUslju6VQWXI06RHXs01bpl7xKVlY7YJ/ZpbXVhOybNBljj0sMc4vnj1LvU
1hYCR50X7BTF9EieZ3+xfY2BwBcMloyKH4aLc8HA93B1udQIsgSXByJs7aQ261dh2c4+7l6EKZOv
7p4Zr7fI9fzulN/Hphx2QIL0HgcKIrPb4BfXK6h9yHqF9LW0N2iUcfNtBkYRoMmd1Boj2jqfRkvP
a3UFLjMFmbwNAdIiWvZKhYlLJ8ha4zgsOSbHHEVRmpZzDHR9WBGYBf+77FviJYltfteE3gsJ09hB
/Nk46YDNx6DNc30IwiNsouX36I/Cgvw0S0ScXdNfMAAwBcX/jcUUjryY0KDy7zn7yGRdSH3eTkmo
eHveyIzwydzNaAjS/vra7NO4bmccXPRmzS5J8XGiiiuRDX0fLtUDG2ArV4pCQT4MwLGC5GvsuH7u
EoNK0IJ0ogGoot8+/2BXE+SouKwwIoRke5/7OWXps23/X7i6CFTZI95EFQ0OQdM0vWzasqs4UXfr
9IMs+qp9qkbq3s/FeBr1Oc65eZZz4a4pNVcMZI9z97jd0X7/amNZCWYY+vujFicZH83mgUK7zI+N
DrY+j9ip6op/+slWxjMjFtJW4UswgcwxkQj1Xv03yvxBKXjdbMNrF27Xx5o+em50cHNn0oA5Ajy6
kTMe1AnF09hoH1QfXt+LsPx1pN9mO/oCdes7Lm3sicjQt/yESzxgFOKNiq2OdtUNljMJ1lEtv3f2
OYnhaKRmX8qDYzjvCL2E1wkOM4llsPNUHzzUN7cOnAo8D0fzhOtSmExIXfetvz20Am9Ms5BcXGjX
vMO6OPnqv488xOVJsdKcWVd/WDGEsL/Ues7Mlykz7WUl3wn8TdBUhWqHX0POTwd+AU2kOVe2x2XA
iPURwmWjhmtOQ46ud6Xdo1PFhAFcPV30lU1yxXdbrRAtqG/ggO9afZLYfmv5DELBAziZArRkz63Y
KNeq9OG5jWCEcenJ2ZneLuQSktIliUzZiq0Q0SyZ3LXMAjH+TovHvAWTxutcGJ5ga+uTM0HfvMbw
Ns+jaQk1mhQQaxha/xyVKKz3nqGrolnRozUP+Y/e9l1PD2r/zR5kxhftlVTELci8WXjl7JGm8Efb
CuG+ZyfL30e3TdKdtNKS2Z42goV22z+Zzz1wQmj4/+gXEwgjaxLpOeYSbMjj5a9TwtzpYH0ER00i
Q3mf6L9pYeMbIw14tgqLHnNROtvD/Y4ng+VAhPxW5wPVIUfcseCFtCOGjeAHbNrxUsh7XBmbmLfA
gmOI/nhJtATRjOm8B2NxdTrz2i3/CGpihGuxyQd2+F2SCR+jlESQtPMJLLtUySZN1dRakHzWvs1C
5G47UHt20bjrRIAyv0iPEBI9QgpUGO5Vtm5MvGb8LRlGR7LAPvgby16A5C4IeKvRdPFbxEmIM7rj
a30wiffHmbNs+tLumUaAclHmUMgaUFtvTs9nK9GZiAafgaFMa1Urz9QrXOx07qx/cu0azxPREAE+
M26aP3ZnI9py5x5nasoWxYcQNPFoBFzyFcLK4iQv04mn8ozobjcRU9jksjBRrQeG+3IFIpjDn3nI
oGQvbkvYRWN/21Y/GxMzXH3UHZSimN9njYnfnmzxGqkV7KOHN6IGh+e0TVRdv7CuFhc5Zo25fCHd
3Rd3ZJSBcAwXHhHTc621T+50l3IJ23x7Bsa/9dKfVVqxUknUOu+bWPAdnDOx63EsTcOJs2p8CSXY
suP1nrjk6Ais5M8jY3W0W34RYMfox69uqMSrSWoad4FoibFBz2YTtJeV/l49A6xwF7mzsXcmWx56
QJuFpuL5egCA8W26o9Y0fixra5o52LDba6XOb7eARhfEJo4G8x/G/TXes1NdG7lO/jOPmHMMzJW1
r3PEeGDDa6LeFJtG0KB/gtv8MjO7Z4y/doDgp2rz/Eu4zwmnoum1oAiYtqlDVTsiMmSJD7+EiCyd
k5Mzz7APZMWOqEeH0qjO+1sPggfKxblCrkCu4MKJVnlL0Hf5E/ku2uyKx7J85KLSHoi17yTNOVYA
50m1lat7T312/bO3KvIIesT+pvScCBVB7LAmgZWo0bXTVFsqBU5Gg539XTj1vPOSYVZJcpiDrW9N
0+sx4L+CRmSEQcECMKJ5uGuUTolYBJrsAFdh03ipvHbVv5u/zHIpchhq5CtNX0n7/rEfKZNHaMdn
ZzaKzhSPIzjLNJZJtZTooCqWYIXUT/A+iDWNCT5MESdVgkDNi10RL6WyK7o/HZvBf8t+BZFkuZYC
+F4RcedHMacklxYFWstnI+gBmznCOzMEZtt5kBidPNcv69QF+vtVt/sjJTUJOkXpVOF8ukQZgpOr
wCxQYGbcYgVulqzK9Lu4YJYvuQKLQ6PLGJM+1T2xLL85Lqo64WsGCk4wAqXnVGg9QKmr+KZf2Gvx
RztGPVNAdozBmEPTeEVnYJ3ul3QNpuQTmdU9HGixHVgshxsXkCajMGvdKT73dj2ezzts3ExW/wyu
LYUIpQDKOqDB6mnrZ11fZTuARkFCOqZFPAUKdTMa/QoCMV4AR1fa45akldEpSVFljtsWOtcYE2bJ
oSp2BXd+/cgglyigqUYvEeliUrbAdvFC9iAsPoC7UkUGhbqWS5qg+L3xP7zOpfFN72jdMwuDeJob
xVR58S01tQm92tCB0Y7sA08lxlizRkUqhPcdLfU9/YSeE7LtynmOdiGA47n8A8Q0Y0hDxsEorJJF
7US1DIplG6gpM1O8+hw4vQ7SzNzzi+wnD4YNvBLW+tcPZFMHMWoXzvdEcuNfSZVdAgAqftmCBTwR
5yNWCCVRa8uZftQsMrcRqgvY0G1Zv9XmdJJG5XvY/+X9gkFPIZzFisO6j5SuS0iv998gpUBlgo3B
U5b9FSF5SG2rRRAwzUc75aV/Vf+Sjivqtfud+kXy4hw/17zV0Ko/wt19yJHPSD0NmswSUENVxTMR
/FKXh51d8h94BtjgoUB9jFeIOi4zv91xzn8Nmpu9/S0PqzxgpGB85n9Gj65QNGxhOwT/IG4S668J
7ShXKix6dIRWQP3bSi5+W4YhDEFQTEPkUIJZgNhcqfQAZdC6KT6RnaDvpkivR4jBUGqyZj/9H34P
57RkqsN1SUtmjyBlFuxruUP4bWoPZM0UbAOHMfhLuD8u5U8Ko6pGtlUqSMiHjGAKFHRMXgvKwS5I
MzK9R5WyrlQk/bmrDfyoXW57LWkt0o9TtmpV+ZJmYbsGRgDcx05alO/mU5dlJFa6LyPCmtiQccGY
2epPFPq77RdOLGxJ3kpTNMT7uJCyGADhTiZDdfMZHFlx09zVDAK97Fu9saTaqV6CocrW7GLpT33p
aCHX23MA+UoBk8v4XM8mh7n8vRyFmUY8M4iWGAe0Rf7QuvyYamIyP4nC+9C88hzDRLMAwvwAIi9S
0DUVH8q37mH7BP1atbde5Wuga4OdInpug3aclMlXjSAUhneqzJGnbhimYDo/G4Jv2FmJ1a5NazbY
txz6t00Z02WPF2skRj+9/gF6QnkKrbUKObEuQs+/gcQE9QAJlkwWtFSLIMSiN09OnoDS0jrbVQxq
xdRK+xJpMMJGO26Gr4rC+myQ3NP891FVMi3Ees+Yk5v4ZP5LT2b5cr7P9ti0QIkGFgW+Hj2ni2JB
YORRsQlrInNzE0kw6sVn9zENzsK34BTXbXOKkdRThhq5E0uijAEh7xum8Fejawr1o5NIWdgefe0y
jOQDCLOQFbP7RfP8f88v9StGAD0rF54LXAvcIQvlaPR99I9XYNlGQ8AU+nQxOYF53I6wkMpd/JdQ
rWzzJ6GD5OKv4IszkazEBAUGoQmaL91MwhrWwKMzVBKih/7z5UfIQpH+7Bx50JYiREfoyvtjBs99
x9UQ1mZyen84J0O6w4bY6Lj3+PZagPVNTqaCYkit+XUNjH8S/uETtBJXmHCufzdr6uM2l8SVCYo+
0Kduqj2+mTn6jf62BZadriPk2aCUe10qgJHQ9l6qhP2hQ6prOInh7d1igIpRtb0oFv0Xo7Vu1StQ
fi5Tf1SM2EGFNlJ3oqt7Sa1MPwS7nlqzKeV9xVuDHpFfcQo5ERbmJHnB+ZPfHoMB0fSQInNgtXn+
AtyqzMKmAhZfaLwyDkshhERMG/HI3vU5DQZoDJIbEdYzNEchNlWF0T14YDZJteZu2iMEPKcP8b7k
P1JpL3qs5WdXuuwsTRBBfHCsbv8o5hYK2d4Z76HBcn6p9kDPatnfOUan+JYhypnWkSsS4KRJNwde
MDTI04SjTQrm6uqLJOfimE4G5Y4uQQaoEMfInqXb9FgjGlyvZMO/dShvszMCklO+KhiaZFMhMdoM
DJIrkAXNrA5akCelUMnGuRMIeVfD8foxOi/5tkn3bS4ed2CS43IPFABMrpui8kzseRa2fnTSZxcb
mQ3lRJqVMUnF/oavIDX+/983tJ7CH+QQTizKrKgOqX4rpFAKiJ9tSMZqtbwY/lpaccc9v8vowHW+
0BEyfeRDh9OCblEsPR7WWVxrpvK9UouaJk2P3RdSIdOKLbM5cyYrqpbcdNWVHggwAmukCaq2uclX
Rm+q1bxyIdXjqWemx3BZ4uFqNjMZHZvpCQEhxaXB894toeIbeZdXBf+v0/fphrm6t3Y8Jdw01U9+
52HWvls5B4+K4d1HTLZmjrFfLUOolmAanPymzuGM4eLhTkp67iYmsJUwOMclkYJtbs445sSJfOaA
x5RNaqMgPebO0CQSiHcteinFDND/XUUOF+HzPmfvtuIa1lWV6yx4okcn16zaMDKjfSD3ek7BoTNP
aFNzMDNKZoWuEI7ZC6CmI1ZDeZ2ZPrTgIe8owNLjc5Kmsu59U9lQMklFUQe0mIvXFtF4wYxr4sg+
rfyittTv43jRRU3/a1lwYYz0kOjR+XvejdgZ+kJTkeuD7gSxR4B4GLTC6oNyvP/taY0thwmdpW0T
LKNJof/w9QSsZo1toyPCsEClceF8WcQ6n+a4Ncd4BDKMLhvOm3JC7d1IKHLxGiMNx28dfKYlTc5E
tk+tC00HZIE2KyIeF09i29hxE2Z4s6teskguqxVUnclLOSL+Qex0ulFLUUXrL3NeqgxP7sEQQzLf
FkUP924ASH983Ip757NqOy+Gxl6GYWY4QWxs0did+FbLVczOfOMz6GKlnACbQp8pNunieB+APt49
GLKoedgtr/TsFdJEJxcjjkcu/ilvmKlp3E8Ndaik+I3N4wSzyujZxtfANS6EOwm+RXBtWmep+5xm
JDK//SyI6gnm2Vh2FCmZrNDbPP/dYQXH5RiL5yJfgwXGtp53wZ1TnYUq/EF1lXeafLuLEUrofuti
69p9Tt90CEx+bAemaoZIGQ8sissIyx2dTWg470rUv/avQXtHEQFfq/JepmZR4Ko/4ddF0r5xFPCO
+IeD8bLqKThAheg8AJs3A5qZ6phApCcDK7EUEZNfeRKMheFNnjHdDqCcAbvwFw9Lb4bhhPqV8xqK
0SGaTtYkEpkh9uIaHYol4rRd9P/TxA33E5ipQGPDWPxuoW3R3BOUWxAoGdOl7bnbAd/yWC+W3Ll0
Jlw8YjDJiXnSZ9u1aiUAZaKSVWn6jEZZOMKCFxMI2CThMr27u4ulaBR+cRMdKMaDoPA7A/phNRX2
lyBnvR2H/ZcUBa3BshFfe7lQiiTov9XxSQmrF8toMdJfa/47hZ83IepRdXpdJr733KSo0b8g/vLY
Q2THUU3UjYmZaUVa68Hhq6EsZyYwBAndooih+JV21NmvIO8ogqQUi1AOYk7E9lkZvTKdUXV5+YIP
6c9Ji2qy/2gNYPCi++L9h5nAT6EYi8mke+KMSAJW4WTNc/DD+UX8rzffug7sw8k852GoB+D1vHLM
wnJq+tP6sSY6zaipAZtXCd2MP4vUZw/VoUDjoZznnh7yOPe49Cznz/H8sYrNG/uq9vxiXi8E6bwT
nZ413vUemp/5l6kZmkh4+PxYZKjROFIGfxmDFHTpSRO7qe9nSJvXlEPKwkWQDYSjWrMQkJgpAy2Y
Ys9tAeyuhL4dE925wY3KCZwzi24bDKHVtUTRC0rpCRPTOFSYMHUTlS6aOF5TqJya4XOpOqXuYA6E
I2w9e1OCLC5xxpLzVdonQ5xAms+upq9K6HI+xOHgT24VhTlOYH01yyuQpKM6zDIAWEYHqBjdHCOz
w396pNsjN0YDPbFoO1Ey2OLVVG06Dkx3WNs/DJ0A9cv+W4ZQ56lx8kS0cIdkg7sCSU7RqU3ILo9Q
no4lsjyyUqIEEKyijxvaoCGF8Jxp+Xm6NI7rSaK9LJNVvcGojxTNeAZ80IYIKY4frivTFC242jV/
9sdInz1AeEnKeAMU/Xk1WlRYTqKhPnOqlT6fN2S7Ym9Ejr7gOwqN8S9nV4EPD9PyBq7jpqpSMVBy
BZpJab/7/6RCnfBtiMf4lUcvVGvulUfK0X5WuBz9x/S4NVy4LFX8W4Oi9SYum+4n42WHR9bjgGZ+
ll0ZUr93l2dTN71A7WuZ8prPacljvJVB6gX7di98xNeI/jywC5cxYfkwhGfJjdahLejP/4fJxRLu
aNx17nhMr0yiAYBWhDKL0z2fbpzcnF2q2dWvW+FTcMjaXTa/EpF6Re+an6DxRDQbMiDGmKCr2FH3
DixT7YxdiMzy+wNfaLlkDcwgKK17utfAbQKRQv1l0BUjxgvQUyyI2Mlmy0fep+JulbRPJIeYVzbG
l2gr4TBFuMO7OZCggD0H/UiEt4+bXjnEqIm649b/bllwyB9U4HXQaf54mq8iLacxSOsXH0uf7O2P
v5R0tuWB1sQH1Zpuxe/bLZTmTPl/r+XvsF21uErYxm796r9fRHdT3jnIDvgEDjbAt+g0HZm7ymlL
Go4DTbBt7N6ZS3s9pM70cytNN5ttmDxmqHgKRL2R2vq6HsuqOBJcVdU1ViIwRcaevWBENwABTj+N
FB8lZ3TThmHcw43GWguYQmPldKhlbfcjG2o1oghY1f48Ofrkm6qfeW0NxpLXMvsoarajap1PiDA6
JSK266/EpkGsaFhL8hSer3ingshJYMVvhlB0OZ1cxHYuqOkDlO58m0vblqha8GOALFOftxXV+y60
hwl7BCdogeMC3YjHOg0G9/d9Xjs1Vcl04tUusCwZuQo+xPnpWMaKTbAnmc3OgMsgFCGGWTDr4F1d
lQHYQCXGIaAmcOYTNMDFbdvnAOh1TqVmD1xD86jIb3dV2if+nUNP/KkCREWloG9kIGov4RLEwOpC
lFp5X7+PTDaAmCRpYT+ohuX1c9WWr3kBJcDX0dM9NMQrBKDvuYIwEBIeHzr7JbBmxJ7oGiBdIZbW
vPmX16F8Cy24EfJWsimCHPBEIoJaIQ/qABUnOh7x/NXz143M3ZMg4ylfQytAFalCK2RtPL3c+t0v
7P6SocN45kI7JO46I4gfMmFjiiYGGuP5q7cz7RgWTaokVvbTGK3+v0lAkPGNNk5VXA7ZfBlm6QIS
J6zgMJ5FovYLibJFpWisdMNGT90tUC43lzumBuBflzD/vZp3Q6Zk0YK2sqANj4et2o7TdH+sQEtc
162fYM4F6dcpOg/Y6/ZtmX2omanxe5uhFnngWs0HknV6yC6I0k/75NQaTC0UgilcFYcxYfDVKUvM
H9GgxCwTanPE8qJHYhQAfCx4EQ97XEvIThl4uruFa6p9HL1woayoL16uNqbvQ+u23ncovbHXVkwo
8O3UDkbdaUZ/ufiTfjhaTrMOYlQ9zy0tBSlKsZhxwLxJ8WZXxo3ZZoFYOI7Jz/Avau0DGiflKxKa
4XTUUqAhoA7QmKf2NguKEWvLIt1dz/5OFRUhC6td5gKOnYluOh78sPK4Y0mkX7CwATSp6vmP2xW2
60hiy3079Kbkzj4b/epHDowPOLyo5OBT/Y0AbAetf8Nz7PbpxOZtbDYtkGXlSCmKvlR7u637OIiT
w2/ATGsFfD2ALw5qcPa94/IqfBOnBZQtXIwnhkUvq9Dtr81YyaonRvCa1HRSb5V6t8lgEumsgDLx
rO/DMFPn2FvVfufPx2v0Hnj3UM8UnLmr8naxh4yW652AYpYJDLlPQmyBhAU5DLbh8oAwZY8yukYj
fGzxqietWLy5lgCIB8SILivaVxcm5q93E/OnKcxGhvl9dc5Qaati9iT452GknbZf1K9E6h3S3uEA
UkNqdWXd6nGvdgyTjcuqh5MxLY+gZxZCb2RlFwJNjCn2MXgqsq6tLH4GwlM1Vgc8jw1EPWPRWDWd
RvHHCjvEzxSDpt79/Ap0QVpGhwBMXl53N5HPR6hIQ1m8ERAnjFmEL0K5HpUCQU3ODamAU4QNacm5
8jWVLCXc50zUd8R5gFJE2zDw+P9u8Ys2R4A+NbG4g5jZ1raNp/2oY+sEIoIthHt2g2QNpDSCBksj
J3qIqCKhpKzr9vQ/e/DgUrm9IS+DTKgRsnJyEkeTUQmIeFNbnwAcraY3HXlJQ+gR6vH0tX5e7JIm
Y05f/u9CIdKhvUV3DFLmxy4hmylrK5NGpa2sGR8w5XQfDkl1o8p0E7APl16hlnKCrfllFCOoefLK
PgX1gsbCLAwCnhmzLx2RRdD6eqPvkXGMpdO6D8xolNxqGYuo4jcxoUkMMAK64CMK8m71+A/OOk/4
HU0/8ea246efh8/nOtjJQX2bEjZgysOuRdEwEGz0F+zZ/WHMTxYgbfCMaK+frtqHSPrfTNljBB9W
pnTHNQwXziwDcdL0soh6glR3NWiuKt8Y6x/5/ARYIHxSkXrZCvx4VqlEDgIwmKPMlEMJ6zsf2V2u
x6HAzgeq5/dAcy8R9L2yQnnRltajZueSaOOahT1r5is8NsH4qtyQxNyCGkg4O0oYuHohRCXN/VEU
o2PrXbE/MvrDSFnQLWByO7tv0NNeVD0BxArs+A/H0DkE3hlzcDzqq2GriSFX07e4hENmPQ3Dk1M8
m+it4/6Y3ldX3zX1peAV/3bd1Px26lNdYUnGEK1FkEAe47KNdqADO2eTrcG22p/3rHxeyf8XTx0I
P/gkc1CIJIzCwDJeS7fQqJISaI7dKMyIBhAUTEysiKZ1/FIIenXrjNrFT7FuO2hXm0lLxc9FiBDM
ncj2Fs/RmVOuonnwyWrwV8XTs9sXme3KieQD8qDVQGZsFJ2oey9rKeTrdLmTsO9flLICTJJym+k3
atSKK6GJjc4HrZ1Rs9pRgRdCLyAN0/IfcxTua5dsu7wcjx/tLMf9rNhnc6sOYcHSCEhaMmlCYJds
LoD6wTcDXcpmNk2KO6MpGm+LnGUG1xwIupde+cnygpTKkVbxtWMATxtGXaAcay13Ig1De+UxAu+I
BRPQrmSuPGPozYYOQQVtiBLZvcejV+8mTquRIw+h+3yjHwrvKkrw7vn1D81/1GwxBnni8JxnkMt3
Kd0rQL4nCJd7UTcSXphLSo7RHVzZS81oNNZAlwjwhkGXHl+AfrdawUqHDLQEn4knxd5Fwh7TozGY
uKdlaa9mwe9SY+H3BJwM0qD5S7zGSlAGTOGhntqHtpxBVu3JEZbt12OjkDVwA/NSLbMn3xfgVYit
7juO+utAluAb5R8BfxwSxwctZJgBnJC6+OTXO44renWQymi65z/+ONVgwzzsS7Y1zd/xPLhmLEfP
HXFOmaycANPAKBCbLivroZh6eMLCB7kApeqkabggyl0avpAqAeg9X+/cB5naDwxnDGwjwmOubwUN
mDUKIw9O9vS+DUG9pYYHST056TNjzBbuk+ApM/b1c2QmYHPKDWm1SSYEPJYSqwXomLG5QpibAhpm
QZWir7gwMjvm+4bppM4L88YyQrLiN/YzUPotboujqmPfP7Xzg2LcZ9PeCTxKsZfjTK76WDF/xbl7
p3B4Hb4uAQOhl8cn+5SjP490s5UAS7RDCZ2/6t6lhdrXjRwMl01uolhinpi0vve8vF7XQMyVe3Wy
NAP8KTD5sMiGQ0NUUlevUh1fPf0AUAcHMjRmFLWki0a96yAK6xgaCVqjP/KB1xJOvNgHRWmCvxEr
gmLsDh+I8cNY4ryT+Qgn8yJRbjuc1pDrm+MfiYA03TOJxNSPjOZU7xpSojGN2XsVr4EXx5T4dDbq
vSUVeCljUhb0XitNDOeDYXrowSffRujBATsI7giK1/EPOG8kOCLRapL9ECsuvhv1I+TAaFFUK3KD
29CKJVfTSJ5Dqhy84zaBGwf1KJq+m/AqKS0yikuGObp5RoWqfdcdwegskl1e67opFmoaeP426st9
NGJ/VVey6CNFsIy4OvQW07sFXCErPq0sPBLHEhfglmfCG0bM6FjeOg/LB4/Ax2LC9kn2FCRkJZKz
cqp+ZtK0FnvztdJaSTjOh6GYlKPkQt1DpaPv/+ZgQ3uET5zSeVEiKmxkfG6d4VZzog1uzkNw54CT
Op1MeZNMmZ+iu4LNh09/VY+0SVc8sv2KvUQAluJuRbLd2IIzamnVIPY/6EaR0Ebrl7VXHphHQWqn
fKttGGraIhZ3fiYOntXwdHIX0oKBAhjHzhl4lWFHDZeWRE+5nhtxwk1Q60p9uOS42+nJY1GfS+es
rAKFBKXXo9PS+9T/wDBm4bsE2bFYn/PBwdKiu2GU8jS8lAfNH+xoKfyZyb7THV9n1Gku65tKsSht
ZLuoBDKOWisMhhpo/NYvbzydSjVWEC5a+ndsSphN3WVW4XKdPIvpE/71TMnrayX73+nJ5nGl/tXl
xyvYyo0sP1mC6EYc6QndghcDuGh5M6gL0OH7HEl7IH40+CTcu6Yzr5OUOfsbyFiQ8xrOpB5B7co3
fwpmrrNxi1FiX3IgPz2cmzYQpuhxav+QrFdSrjTmuOuzww2lIYju5a9hN4lFCmYAUP0bkwUttIYJ
XN0CsHFkPVMNVl/HB72ME1zTr2OzinfCgR69PmFeFwhCrB3/bZ3hLizyPjwHeGMDvfG9PAqqyh/I
ueOA6BCCeINXSXS8n++dTJ5//tk9FGQuO8q9t4rIlyWgLChERO5Gyx2yq29+ju6zHS/jyZYHnB78
r3LzS1Xn6ZNdzjCerTBWnxRjRvT8wy/cZuI77HIPsIXN0IE+fkVBXDK9NWtxEmLE826NMp6gzFp5
cngaNNo0u0sgVb1aCkL09NYWU2tTXIaAm31UZHSaNYxXBxZpxwYdIfYak3x0EwkJRI5MSun39rjg
3AWo7ayaTDEt69bhzYgKQBTcXPLgEdTVOGmkqlyW8CYgdvrhQWvQiAUYJnp8t9qDAqsrLsnKDvCC
KQZ8k7WNJheoE5r4+FFogEvSpD2y+5xawO1N4sjrU7V8XCT4hg8r4WAls96xhHHQWrOluo8PXIhV
w9N6iTqF8Ijltg1/9zJsXQTGPFRHbMmVF0vYn7EUp0gHWkjb5nJ6BT0nC5bxtGZgiIBCtYt+UY4I
ljXWRNxcZIMAORaGNZSYqAYUetm8MB8O3n/edjzP3y2Oogy97cH5Xdbl4VnlH/HbpuosI+JGUC/P
ZgaXq4N7djVm0josRKtGt545Jr81KzAzsdhykT8hx6NKcpMpJ9GDTFUGbt8aEp/vNTDyKci/wzwO
MKRhxR/9to1dgCidgCcckDngUl6e2cKQbwBlcsnwiBKsSvdNp3b1nS8z0/tPrRLpSjeJHcNvJQMI
oNyxo6YJEkmOKHoSQvvMnU4FAVLjLbOs3KTRl9ctEKGr2jSe1ey8OdoXOgLRkyeM8tpePxmrDOhW
J+wm7g/M4Nd88yviKuzKXY5m7/zgTxN96XlHPKnurD/YI80azDAzDIlZjCRL8A/88XTpQKRIU2/e
hV9+RbajJPRLNKnU8a7H1XRuGb1CmGaZeFTSh0EwQ5D9bZ1LMDX1Ggbmqn0Vf0JK0+xQH8rDKqX9
ok1KKa4uzdG4dwL2urSQUxa6n1hWmAuoomvfM68Qb3FRmfCTOcxpbzh/6HpoAN7Zl0bRF9eb4SY0
pHJOVa6tqlfxZ2og8FwiNZbRtdSe7ikJ4b9wl80L46DhimyJZYbmCDzpR4nG8KEGXCehOxKXI4b8
sQmfm9A24UvBgIC9EmbdK44PFtQ0Xt+p0Es6+hnlOEorF1iXoklW4I4o3xN7+w6KnEFbAbq9LJq6
g1nBlMXD5ZLKLbWpgFgTVp85mVYBv/OiROIWQvjzelnWbyKaEOCYjX4FaoSmhx3CHHXvP6g4ni0Q
Mfyapb3w2uq/9Gq7V8hGonNjpjLN7MhVWKn3fiym7tkTqdoRPHp79hVN7PjqqstvXJbqhspzsqbn
4gI7tVaRpakVch8mLnSPWBBPFsAaNlr9LWLo/hBRKhV4zs+VzZwn8Dk5b6qi+tAshe3p9mndVS0H
LUs/3LV9YvrGSrQhnJgEGxAkWc6kAVldqjpamD5OnHsL6JilvBRRZCYBQe35JGz1/vTijtXxaOiB
aZSDlyX8o3AYaevxmzQFUAQKRQxHFU6OfRWGbT1GJzIXBDejuZIYosB4Z9320gBWF8KKFyc6fJh0
RSmxG+k3dfJcHho621f1KZtBMLAx+53iwl+4S5Mj+kkOmZc9fCSeMT9ZzenNig48oHsHZ2S5UhQh
5WVWxhV2/dEnBaSbpyvRGpr1nyhvbWL6qqNUsmWTiUTOdXeCeUZvK2twDcfhOWw8rNmwOKrPCkuH
PXU3pJ1CjwDuJGdCrOj1oE0JwmGbMHdf6znUOzrMqI5coyx0Ihx9+ok1Ni9eOF0PFpKzzj5FhyCZ
pjbJwFEBRdZ59pZR26NFlh7Na5fDandJTQVLy3HBdnGEuVMHmTZWYT3kOf8esKPHIwG9TTKaMN5G
jOoCasQprz/RRedLcO1maBcV15popfWtHTf5K2rLfHNyxPpn/VbvxKZ70nJKuKfebSPRDrwxAB/r
oK9N9WA49qUOdVnmaHR+kLO7Hr/7G57NxuvXWaRKIrqtU74wwT/PPdRSaE4kXi4dfsv6NqS0Ube/
cKbShSHxsAkYoNC9oyEJL4q43W0cja/Teqy+BtRLh9B66QGmFIqnD791QtPiMJtec4GJEDdhuFjQ
HuemKthKzh2KzXGQLXJP6MhD/68zXQRWRKeb+z45nN7AJHkSdZNFB4Kiv0nkVxdvrXC+jlyLJpj3
s2q4TFM3VMwDzHe+TB2zogul76RhhpitMTbitYdRZVPsEK/4EcvP8XtEvUrP4M7TwDKa8zy9IDos
9hzxcjAqs84IxZZrx7EVVscISoOg5k7Ql121m6qX+h1K/+59ssRV13Z9f0AwZMNhtP0ZYWQoEKXG
n/tXYd6xONyJW0GoOTDsoGss2yRNL4zVPPvn5rxmjAZBcUfrroXQKfZJcTCMbpSkmN1HFHxhMmA2
cYg/iYgonKNyp5hHhM0V90mntSgt4mYNdbC6BzxNFewpXn6hitLSZrUJUq3ThYpR+igYhYBtW4Yw
QpKKsd4D6j/Zp8SvLBO5klytpwEm/KLoPb8hDFE8LQ3Op5L6pGnQWXGKW9jCZldMLOE8L5Gzfghd
EcAvw0gMADPmnY8gontutDbsA6Y6cY38FqdfOGO60q/6TT6/2anh130ml8GKbU9JqLOr2wctXxTs
rY9tCCWZZi2Q7MtVwFHqDkiyQs5M8VCi1IJ3brtdAlEtivYXpcZ5NdTDqqBAFx2lWeBeNYYu7T25
GvQN+UgQ5IhJJFk246R5asj6p1sxPiC1RQqNQB9JVk2zvOAOKprv5KGas2abxscaTqWkEFlETe9g
nOSRJmiJSt+1slBYfSND89yYeDf6397hRhMI4OyIH09v3oultMPOtqUzBOFnkSe3tjHEzGROvJrk
mPU2L9zq3E087ZLaZZFVc7siPPwSttdzDeXzYI42Fj88g6lwbF5zTBm8uJDAYR3RYVLlk/K2Kfts
8S4ZESzwfLSjeFd8baUUBFAtUFsDt4pBlLtXzTShcIv2/0x3vee2x2QgTiur5ZDTqeBGoGKgW3gX
oqGN3luvYVUAu4KpKyV66nWH16meN6eoeq3GGxdrpKvL+5c4sXMFePpwxflUNU3zAADNg9Wqoxoh
Xh8TKPZ4qIULnW3Yq6GeEeqKSLV4AUYL2wmbwfxqovO58Hq2UYE99IUUsTAQDRYtveQdwPQ6SU42
ey3n6CCcCQV1TEY58iheemhA15xZujibMqbOpHrZDvdjDRg7DA/R9QrGhRjid91Dc7KVbgV/Qs/R
KmmEMjR/YfzEqtnMOc53l+GmT1nHdHHS+4OXA91xBexW0JGhC9mWpE2G0gMyC0I4mv7ywt90aUAb
En4obmofU/jkAHA2OMPCS8UdGApHoJ+rz1LnZ94CMIvqqy7ClKKTHb0yKM/rMKeWfHor2UNHgYbg
/B3T5+t6LC08RcFyMSvJNxoCzn6rFPiThCAUkSKm6R0i+17qg2Q9ctQ0o/bG9wtYaAwMSq00aH7S
wHDKyt0svkF6nr2W7IecsEuA1S665v8ojjveNtqqkN3agfH4ChdirKLUwP2WKsQ4uX0M5oy8JY0g
mU2v9nk+2Xr+hhvPNxhfgehh4tfRhb9MFnTHN6l+nkqHBho87eY1XOjxIonAD9Xwv/9Dud0zow6Y
dqtBuZKSRIGPFfuU4Iehdrz6x0+FDNWi4Kea7DFdqI+F3iYc3+oaq0z7pTQ8GF0Ju7Tre/m+q8Hx
2lc6O4FzTenQ1uGbxddUS0QnJOCuV6hKuoxQ7oCU/wkawB3fG88RW+NNOmneq6F2AcAgCd6upPEl
bB78/boqSXzLgBg0O+wHF0H5fimxMIZjrYCLDWmFmKlAVWV36C5uGY59vBrxiuZKGUVpozYeJgXv
QZuWsAg1ftJ/4wqR+J5X0UW3srTk307KtagjMPf7QrbEVS7yBwgHp80KVdxF/BTkgMw+ij4YKX0Z
qGr0XOaabj+iDTfmqa6d0zfHHZm22cz73AUIGvc1nQawnQVDUOO3vSavhvFcUYQXWci6/BgOga8N
Bsq5MFg5M6BxY378rtWT2bEkC0SvdRqoOBgXa8Xvl5kVGK9UBrH9dROmnbjfmHeeeiFA63Bgzm7x
zO9zNlZmd5d2Ld4JBff4spSn2t7Oa7Xef0NhKjkvv2uxq9XujUpYg6MxOXNkvd7Su6e4VVCEK6Xe
f6Lq6MdIU4Udw9RiF1oe4pYUFiUzutJdNm/ITMyYDKyz7TNKGCiZZ+2CKhrA656nax4GnrfBXdTB
WG2Tp1pkrY5baqu1GFJ0lbdXJvEAZ9PVdOFlxyhW3iQ0QIxAxAymfMnZCdgz25RYBkpoTcRmjq8H
1hHI6Lk1GCgopp9S8ztEgnBTwbpvE0NHibZgz+ujM7/vZd8qGaz7plq+PYlRvNtOFad/589bTAiE
HVsJKiTPgkkjSIaET9xYGyqSHXV74TQY/ReC5+HqHvVZg5w4MYeUV0Sy5yvgXHVTqBh/8fJoimA5
zc3mumaQD91gFSfWl35TgTiLVhsqB+d/xD+fruET7lk7DMpPEEMmxQVhrppUafmYd/sr+09Ev6I6
ElPJzFcWKQOiM/wxXSICxXFLA/Zhr3iGNx4fFmNc/LP2Dr/aNzc166ucYedBIpnhjObeEqE3ikUZ
oNohZ6m5W17DnAmTaE3hJ54mErVmMLrfHY2JCCWeQVeOOPRgySSIBvPAiSylb65JwoQ+ENbnk0ud
56b29eQkzibDebFoELPAtZylYK1Lsndrcf/rdfOfVwy3CCzSV3VBItk9IXvelUIe3TlSQjf5WLVb
CPODVzIkKObVLRiQSMaN27+XRp5GJQKtgQ18R1gsFUvXPmDuh7ebnQIwT7b4XID+4h4XRUkb/i6o
ADoskZNVgGRos430OqZmjjfA6cCVk90rre++hbWTVqEFKIwu2gCmp18f31FMwzOy7OKXmVK4QGSc
y3t2giwUjHC7mE5HFsOKmK5ealtMo0mNLrSlU8C+eB1qiig9iKKxgX/s/lyP3gkxSWSkoKqtNSiq
armS+QBA3oLn3vTjNwLIm8ws4q1G3DN2rQRRNQz5mjv2wQRyrKDZGr0ayU/Uo4d6DZh4O0mswGik
l+mJWO9t9ash4iaHlo4BIKOg3wBdnsg1Ur3MtN0k3w+0czTGQy1zzU/p4oEi1GkRkRWso5UCvQmN
QtnignJ7F5oOK5YoiRNxFZynbMzNrn/d2wunbtFYKSdCog8PIzGRX+WBfXGk+aaduihO7SbvX4Y9
MOW9GrJT42MYcoj1ADDcHcQ0vB5OFhvOSuK4eATE8xcFyVBcCI6JdLP9Tv5rLY4TKBz8Wk6JKPvg
N9ecFb6L+dTBH/pfbERU6g1Ixb/aq4JXmcKitVGjBYWapnOp3Bj+b7LXFAuT3JhWDVMOu0uDAFxW
ZKe4M4kvdfTzINzMoRmFTirDHqLaVIOdT/KGy0AD4KCXL/0PMYitNx8lmdkYpGesDm1X2qrXT8wO
mhj5t0XBSOG0aI++fzuO5FSFYDtI3EfQ5TUN1BZXKC7FwnJC6/6GlnUCkP9oQTdGflNs6cGe5dVV
XHd4hkS3RI+2p8aBNS12DIP55oUPhGJn0OJRRntYZjiWYN1LYZbg7n9zSubXUBaiNd6cUlDwwYPl
aRLIMZQVDFhmBKNt8FstP9ff5iCw+oWkh8aatbxvHem7ZlDarPWr1ead3iIdQI/CdcWZM4RB7ZCj
Zzha5pdk01SPTwRia3IXt/ZgcaCsLH7mnUmHtCFpRcYJNK3Z50J622+5+6mJv25kFkxGOCUJBg0Z
AAL6krzxP3Ia8RkY1QSkvufjgKCVSyyvV0SC7TvVZK8cOOvDRXfr2u5jFHmcDGv6HUZxeRXCF5GB
TrfswwvDO2qIXrXxOreLgF0GvrOLK9XXsaVL5EuWlHshE1C+KbdLR0hyNf+7H3jzbC5E1Dwv7l3Z
hEO3vECpE1J/TZJ0MJx0D8r806Qhu9CmspEJcmbGTG1tHv5jEOFMLTgUUOjNVlLMDB9d7aIMW+W4
qJ4uWZVjSB/5vG86iq2MXZHkHPUN8Iu9oeyUozrV+Q5ZU3zp3nIQ1VaUvt+TMdnu416zkq/TPV/y
MrZoS1sKtTP+JIadM9EwARsnnWFLA63/TCEUJYiBJByMlb1eS91kn9g7NxSbBeysvchyTtXaorO7
orZjAuQaFzYZmQEeTCh6KEC7UrDo82lpgy23+/lfwnbhaisgKYJG/aDagskxLyvucRyuxz4N38RQ
tyF2bxnG38tB7bGc5/ofdYPbxreu7tWPFWVN+TeBHcGUksqG7I5vyz8z8+V956JMPcaedqOiW9j5
bTODxmTD2BUjJjoWfXxhDlumhKGNyQvAJbiIDlESF6N3gqCGXC7wVP8ZXGPTtIvA0tcVA9PG3px4
PI+tltyFZtz4PuJl3KgIo5XJEetbnXV9fU1hF0aEr4vyYxoecOqH4LcAHn7HKncMfOKXiGhW8csg
q5nAYcl6mFXhCci+R18OO9Dhy3WYcp1UqIJzLOlsfhRJCtNge5aO8klHSEs6qPrIS1uownJCXc0b
q8ZCZbk5YbVzE+HEco+kMuEEaMyuQp06seQRt2cqKI1L8bAWlTcCsFVCrjN1rY24MjMS9Xb5kyip
JeAzWMdHBVDmSdJX97o17INxLlZ+0p1kIf6IEOSfVQZLFd32gPm3S2igsbtXYwccAwQrPN9VUCiH
bm/SghI+79Xe7jft7rUi07LyauI65B7k5U0Y+0Ivjm0/WGvoeWnqKIt+ah41dXo3toO83adHlMhO
ymK91Fz9eqbA5oAGrNqYnhDYxIgvDqSunbZtXYNhE/wM1EnUDC9vdIjoyDZRy4UXveOXnBsQhK2h
B1If1BwYq7Wuf+Rh8hsFvaLkC/b9hD1DcxlDpE4xbGrkZXLctkrp837/g7Jk9SpxGD5986BQHbw4
4trfG1JdgM9Oylhfs97kq8sOityX6wkdU/tXRaJM5NwhM5ddkyrtnSLovC745lTHFZGCpj2oVp4n
uswI/2fvOdQCdiN1qpSl67Lf5PriqhFCw0sCQuTqxt2XI1ddcKkhnPFxDiRQu4UsJCwBYA49/jiC
HAMQopLllMHtey0V4bVyafQjUQu3/qZ/HY6f8R3f0sharmcI8C3ngrHN/z6NToQVyqfoMDgjrsZA
gQygXXu8oQ7GWghrMR9P9JCihwG1nyY5bHi/rHWWeNUc7kzPjbNhIyg8l0+5PcymUz/vqM3YIcXr
wf4X4Xmnto+EaE7dpuCGNFrHF/TZu+N5/DRFW07K9ThZJ5aoo7bVinqyhm4u3E/D6pXSUj67nRXS
Zg+UuoeKX5QfPomndm3YrfMm5aFwImOtrQjpb/R2SmA0rzpn4xgo0TCamYmyVdu1Nj70P5b6VdX/
J2fdyK0p0UI/7gl61GPKlAkKXu3Ey4yo8jclnI59IkplIL7VZQ6TJhZzdZ4708DMnmIcah7KSu4e
/DcaANPMC8DhIgtAJaSAaLCydjsEoBzFSa5Lpol9GVWCRWxQV8THqoyKRkCk8FlmgjqYLApyX6+k
2HN39nAVz0J3AGvxTAGElAl5mEsbwwkkT2iIZDw8BVSDpesIFQV1R8FiCu2wcFRu8+f6Wr1ZLkEz
1fd+EFNBDLrOHo0A3F+ATs/vnp8ojTzIzx03zgrLEG9Fj2baU5XWMssrRL26h4q+UZZ/zEyYAQvl
CBRfGsgUQPPQpC0eLJHplBxATShfpbSLQZ0ji495fxP8i+Int6iW0qNJZkRzdhUlHur57UyjCNld
rSQZlTluW2gGG06qjOF4AS0tlJfIlj95ssXdTnxKngG6wHfntAYuK7bnBFh75Fbl+KyQl3z/cI0D
APrbTz7E4027Pwx1Iujt6GEaL1h8ARFMLIcVm5t8Ldi75LlMFJD39QRvK0Bdgaq9LeI61ESAUItj
0eQhPsNOnFWc//auykldlLj6iJiQKKdF5L37ciXHym7jRWvc196PgPYmGbIozqnnaRVODjrfkV+m
mMrOAgCTP5SnDAQqDA74kXqrOSZ+wAy6g1rd4IQanXhh3oYtQ7utzLmPPfavbl3chla2gbFkhAjX
RPs05wp7iPx4f6dohz6IuZg1dIdcNoj47/qCytjQCKx4+62TGGcSoHm41czruEct0XY9qyHub1lF
nCpLF7zOhwQIQw5vS5TD9qEB1tMhUlsoxEmwZCFeIRCv+r8jR5/5bqKZZtuoVK16UkviTqG0obaA
1kJEywOD/MzmF5ld+n53NdQaTUtU5u0LzOlp+6D/jXi8Ro6Js6987d/K6LwhavcXHpFGssY3Vdfl
57vtDIGjblA2ko6fBj9nYqUc8/oZvYKSUdGP4d/DlMT/3Y3TrqlK7CsuOXiqg020ZC4EGQwDkrdj
OZE/yiDWU0dSEAh8xBab1q5r50vP81N1O/qOjQhzC1AafHw9MDYsPSFKT6DNjgOnz78S8kRf2Srg
g/wqGcrtT8zZ0lhnMR0L3No0tASWZO60sjyM/CuzJkR8L2S+XuIoNsV8L0aTCF4zv6va6U0ygQ/B
pWpLbauOXgqVakg1B2huqm2nDbTaOcHTLoiRRSDBmZ1HZot5w3h6hN2s4GcVUPh4d3tJd5EXttKc
9NUx8gibbp301zfPIA/d5V0ZJalFVVtHhRQQ4LpIlX6ssy6xWihAststEAZDzYT5sfsVLRW1k5Ln
FgCHJQ37acy1qH8xKBYxR1X4Qo63vi9pK/vbfEk7kJbHbDQV+yz8qLsYNsksSjtCnrxYjoqn3SSw
qRCjaiTpIbhhCTOfEx4IJVGcbpP4EtpTKPxeXcQ2GKbf+/Ww/eQsLmGLYqD7hY2kbNA+G+eluQ73
JWzIgAOHsbkq865BlgT7Ilsqc2H1r/ADKKC0+01wj+jPg4wG2UfpFo2MDRXm06X+/CuK3Yv4j28a
1QdnqdUp/J6LxfHYivqTyQaPE7RFbQM7bWwmMhyEA4mj32hTx7av+JUUQyopB7CiyP6TM1Z6LddT
wThZiHwX1YvaPA0/Dn5nQxMkzn3frcahfDBg4DxE3EI4XZBWoRNpiIIdYo5XVtKUoDUELmPb/WhX
oaDovV3WKrPCf/ya7jHnWcjckRcRrnIzYjgTHCE+LPBvbdldtl440SUHEc6HZEr7roI9xf0YMFW8
j6wow79lYWN4zh0M+i0glkz0F4+LvFbNI6fgLktMKrbXzL8uhbLQ5oMZdJiDNFtwOdU6x7Olx+UB
/00TsuBNLQ8fBa3dPi4W4gM4jfmEmyuB8WU7pByOz2uYCwMBlUVe5YKa4O5ZKXEgIFAAwoZQ4Mwg
G5SInTED+MoNSVt4LLPJv3Mx1To2DOVIK6RAsuahw/gnCI2JeQN8mTBOeAtKp2TvIJUQBzCzyviM
1GT+jzuKm8swGgzNLZumh5Hep7tNhQOGqTghQxn3nA/xL16bHHvmQbTyUPVTeJbCM+aWTOfJ78y2
7c+R07QAddFgGX1ePSWT9X6k5wFZTi4ZcM53R6Mij8ebdsJdbnubxqGQdRoSv/G/MLvO/SNPzbw2
0qfl/+wFDsUxV1cCUMaQ9M/TmOkNL+UgBYffQQfDBbeVw3ix16T8S7bZgLJO804vfx7JKus/sjTr
lF/m+RyUOX5A9lDGaXFmnr7Kk41xzySuAbWij2Ce8+lxAzGQdlhRL0M6p2txi2HKFZnGMfn0UDdo
+WpaX2ZxKHjKh8RbUBkadb7kSpsL259bH2Kkvg+Ou1nVJA8nExyUdq3LUlhlomp0ELvwiZYAErxG
5+U6yNDnHgyJaHfQFON/Rf4bIfNgF0ly+vB/i6riROjqosQ4QVu2zvcmvWLlCk7ULI/nX9jrLVHN
dNkir55WcoDF6RG+rkgMfd5QlRKEd//1CYEE8bkxMjrrt+APdC0tXXzgbhCPE7EwVCVib1g+t1Xn
bK0AGw7Hmq+kyramUgiiYoZ0jgOLHYa2HT8Mgsy3D1sC5VmEDRnqyGFc/N3IRO5LgldLJn9fyBcr
Woa+7GCkLY4mwUpMIn2Ymyq5Tr9LknW9FrRzSpDonMkGXMjB6vj8JlmeoWE8FCbERLBOcT39ephY
C8txS0vtsvn+pQTp8gURMRPfkrRdK4uD6Mlax6SI4ltizuI17+TYfVaI250VenhKsk1Y/kmJTRl1
Iplw2l5FKzkvD81l/Nql5SA0I8b/UaOcgLBkVUSvqICyymh3knkI3k+0HRDUPRt6KyUjIgO0nqrF
cxur9gT1yrKqtBQTRXWeSgDYdBNQUF4BG3eyCAt+IrZcpi2t6hIWkFWIvXUZ0hgxETSgGUvhSpIO
7+oqe01WRPSwqOa9BD7em1mYIGBwUum22Pu2I1n/OV93NRmMnv7hvcTiy17hzsCt7lvdDa9K9AA3
y7M63DcFjsXY4EUo9nW4gGsvTYf0zEksGrLGW68ZhbsTZ26VyVRVGkelYuzqMEXPHahdDHjz5OCA
NmJ97qIXM/gQyjIbhh3Lh/qkOm+IHuTvzBNlGR6D/r8aG2ThDL8XjU0jHry/JFa4KSCk89BDgEyi
7VQglZ3iUp3hJjl5o78aOCSZU8HWNOmUkQdHbRn7GMPp9AaJQ7VnLRxm9pMkWyAM6yLCp5wZ0th5
ceKSLlq/So9Vbo+hdAbnMhd60ZkWeAEpWs0cSeEVeLPxty1ZR+wsDIXhruvhH388vt9qeLH0Q54E
DP0NuEGbBDbElPcOshDQrWt9n00MesEGkjegTCVgxly3HdH+7MNF9FLabh64XtdJmD9ksc/UXiAy
1wT1f3rAwNcr6ePMNIrNVWp3WzA685fudXQbSznYzTMM2uHbUX2S+F6VCfwWkAmtkWEaPsRpCJjA
IlKi0wDZB5aLybOqgD1tVXMzy/npcXYaxHIK4Qw4MnMmAWXVNKxx227Zu7VszknhQKmHyS6CRunR
x3axZen+eyJd/o1k7y5MjLtTnYyVSjhFOUx4ltd3Ca3TkTMsSbgfV10NVkBrMRWRfh1ZGJHSPA1m
HLpiw3iP41/St1XoWM70sYLPh/XAlho/Ly/qPR3rLgX5WuyGf7pChUAxpBkL0QgpinQ7CtJS1r37
duLbL6Mks5m58XGjzjkeJPP6KGVkzic3NXDjas/vjL2zYFUFz+NBNUsR+VehL9htiH5Wp99vo8Tx
7dbIYWiRzQRVhUpy2WxQOvev7qMmtxcQBse9oy7BWaIemTLWTEvb4QdUVGEMhEUx1bz/8QxuGsqu
pVd1iIPe3cECctTKTELbuXmg6jL0yANHefkcb2mqcOV3O0IxZygWOtJgqTt4BPVoiaH7jIbMla6W
5pUZx/+iiBzhKhg5SVGeVBFTT2drsY9Aua7n6TEu+X8bfyLxJrwNIx7ByRRpe+l6FQpHvRaMy3+8
XusbTC6/CrNrH+0VpwXMXH8xbI/KdeOQEOun7JZmaN2PphH1A+IgemJ9m5PdMSYrkkUspY761Wwb
/7rjbvNTomWB3yLq0jYn10kWfoxM7GO35TAmxhu8A/3yK+P/WP3uOLYmpqFNdYMimo4S4a2G097N
6QYoHG860mg+sdDvFphFClLkrZ5GGbViy0PVP0/TPU/sPtpxeSFzi4b1KMpl3Ov3zYK3ca83V6+q
zG/HCh07UI+7GhdIBybgpny8mFaekqagNITt4VyHVqnzftT1Dtmp61myIxb5IwQXJ2GsuJ30D9er
BiBtlTf7RoE4PtgOa7KpMSyu33nTBk2MzIpfwma/uWQQPJ1lK6ydgDEtjiUzOuDmp7hD6f+GQddw
g7gy2AFI+YVEUq4HtkRRlsblx0BVj/HmQO6CVe1kqMmcBj8GYj4aKQ6euoGfMqqxueetmMpI/31T
vFz0+YuVCkj0PjK7gdehBXHOkG8hYLt9cPMfeYQxMeaj4kr8fa5vsF7+1Rwk9UUvN3vE5jkAsbn2
nmlUu00Q6TcY0eKpv9lce1z+UFqa6fzyIwdqNoegIWECYXF2NtDyhUlmFcvjM0PhK/hYuh6VtSNo
+vlx3gvIC1zs0tkpky4gumd96UGoFvhlnRVJi5MuEr4f+YqWK1hmI6DytVPjg+mPYciaRDBsTTlF
11VkyU2v7NP6X18PxgjCxNHRmzIgbE0rzGPejTvS9MfPk68yoFl7uSbb2Dzc/U7OUVKqzcZIk4rW
jFCSBGq9PmiJufrAa2OUmXxIAyIkb0ixuQRjIN4S+JnTqEsif6rPaFjWDUqix6gjVIr2QzfoAYYS
RibgGnss1eWFz7oaQJ7TfzSng9R2yRBARBGh3cGeFW83RdQ5XJLlgfgJy9LT9JqsBQMbn9udhVhF
/Sjuyi64pbmxfZWZqyHyB5GWZsrithYbtMV8JZb6NUrWd1t/pWIsT83yPpl1TFz8+u0epROmfj3O
h4HSUYv7lec9T0YRoB/S/+vGp42M1D+szspKaJRglqvR3gTM38lVm4O/Z0lrlaRArAHJkz4PXoAL
vAAmh1DpCfN8hEqq3m4z6V5WfPkuhNJ3BViaUbITCDMQH7RIGSkCN+l7rMdGoYU9HMCJStqXMTvl
JAd6OGCiS+PLX78sBUITPNmMxir5OWWgc7RBacu5zrF33O69IiQKy5HoPxnkv/dN2AC35JLk53d2
vKh0M95HOG6dIxMqDNp3vpwBczCWJKtuHsZPSw4MhMuAw+MbqZXKisfoNi4mzqX686AiUVVh/5Vg
jyc4sdbTUZXZRSTG/EgIX0DAfzqd7f0Ct3RO7CNgyDA1LaBWVy8Hpy8bjYU3vJj7LElE9Lo2gFZK
KuDfCal0cH22GhPBT7aT4gvfFb2uLX8NRkX5sLHs6piatY8/Cw596WQd60yM8rVvaKRKwTvtYqWM
bkGjHGzVg8kY6cH3pq5tzKfYm+Sj07tZ9twInioQxaLqfjyrgxLjwJFO9Iqx2GHAYckGLk74IP9D
5mACoUHFeF3PnuKIhGKbvYWmijVP6wj+nv5ynhiHz4Cs/p6JLIIxQU8VugkX6Y6VuWQdK151Np2f
TQbLAW3AqWuzbE4zy7f4p8uGxpicURVpo+Ex4pqSd+9I6QcHqYZizY2o9ioii9IRKB8J+I0xY12b
cIs/Q/HOTmMBV3eQyemTPc9r6JCfUCP2psEFdqLY8s0OKxhUbntSczE9ekvFYBU+Z0siRst47kqs
GL0UkcQoIYe+hwXfrm8tZ6g/r4LwbYFbDlobLsPUzuaBHMxOVQFqETzVpNXGYcs7xd8S3F6x2kvT
Y2CRKh2LIQr2Ub9KpLYmQbURbyc1A5Kwzt+5bRC2rwtZvilhguVIhDGCtYm7AjFPHxW2lrHKnH+J
4f1beKYC6GCGCF5vGkmWlfsxMG9x8X9WKmXR5W95D6xFRmNKFc5XfxD3UZrvXQEnmjVDtorKFzTU
fkLyZKGo/RvXFloro6hDlCGmyD8lPL0G3yBfWyW/zu8SGtsFUh7RbrZYJ3+88ysC1Qm0HjcgQrN4
1N2N4atwzkc5mDFZ8xaE3v3q3CaYnogJIclyOVxrvKWNM4Xxx9GniK5jMhGblK33Z0fp5/H7Bkqn
vb7xUw9sjL6GDuOuZiqcKMpNG5GrWxb4TmUk2TzZ+8xh0TVXjNuQrxFA7KcW4b96cSDITpzLEQ6+
RmbGPHP45dijcg/cqUi/FoVCe90a9RodfwEPpofrHyTwhfiCO49KpRsKmN1x7Im4w2Bku1yMWXP8
7CqA+HVc5U0N7IWe2FI+Oe1fGHxKmNLtJoFv1MY2ErUHMJZKtElGyZvb/8VLjBZ84+6nmlMH3pkl
LTvMbIN6uj0V8aqhWMwkUH1izVqPNez/p8DpaJ+3EvEWmFIVBI2H3/TCkB4kaCWLAn5yeyL9lyco
Vp/jTslcq0MeCZscVsAvgHa1qa+/Tt5xtQvAMltzuFiRnX3FUvFPzbuQb88HGNBa7ifFNuXUnJ35
7Qfac6p2oKmMwxTOaqHM5RNHRZpZanXjpUFnA19wDUZHLzGGn0Y1I7O4YKTODJkBLnOcOMQxWQyZ
dVRBv89Nt40YxBSdZxCKBPH+FAmrsu0sjlEXy1hOZPQ4g4MglQ5ngCssoZcR+ZLxTo0Mgsf3y1sY
6fqhpbeZTHVRPBsvMDuzlXjAOxiSq2rO7ojfPYjWdj7shkZYeLHfrsR7WPrBqPdzSoFJ/uyRDjbo
wvRMzwwkot+6SIYXdHY5lGcfZE2u0wIEwSNWUDE9rkQdDq3eWqT3geLcnIcFV7HZKbkwkOa64YUX
B2ynIS9tSeMsfydYuAYhBXAC3kU7lyqRFvAJAHtpB4m6a6mqb0lZbTVvw+RNPhUsmNpl6xOLRvTq
3bMWZtRpVE/oMS7OMY+xOLy9cXgOUrxShAiYQGOzjN+nWKMV4cNWp4afyqLJdZBEjigZjxL1hK+D
qo4DJ6a11PY263LBug0OShoP5V93GzYR1iC5VUvgBgn9DhiB4eFw3/AGJ/i7f+4doSdYgYPs0/P8
oY3tZIEumBthpyo6VIa8NKqW7JxZYZLuGJUpLWWklvZxHt4+8b4kF9emE5SboqKyBTf3gj0Se3G0
RyWgQ0GzM3Gy6DEnn64KwV5ICr0MNUlug4LcGTzA0q7ZKH7KzFPjPOTGLBRGbgiqsg8r8FJuhi1H
bVZHdvZ7UPj8As4DzcoT9ZO5oRuhBpfAwVdDBQq3D26ZuVzoZsL1fBNTZbmr162xExKTwUSv4aOm
rUgwUhEYZFb/NywNc83MZgrXh9iWgOCoSNxvMsDS0SNUgtYWHImkh3jgROwZImNbFI2O1ZryPoGc
KbsKTDTI02WIG+v84Wnv0RSDmkSEakF1rCr0Rw+D3Lzzi+vp9UR5VzbSHrKvbgMneI1QaLWzrAPL
ZGfzaLDvsOmAry/MyJMbfP6mgbrrGr8qNmjwQBWI3GXYAx7hakXLdlQra+R4ypR/mEuJbAch7WEP
3zZfH1WiXUw6MIYSrQKvqErNI/1MeBRuCI4j3DwQrlo9K5JHdDdWxlLWRLU/lCaPs4YfpMvU+R+o
P4uyvgf9eYfFTlw/W6F6RFglZAAyPhCvAZ78XbkOPQS8IZu6OwlOQpk96WEkQXQN2KMuqKmrwSb+
j9bwVFLctpDfQQW15vS/VY+CVLKLXfrmkgY61Jaf3ml58fWWBS1NTbpAhqkXFDBgB4mRfpXHxT9e
BMQzVzJ0nGB28hTP3qX9hjBxK+Nbih60/Q==
`protect end_protected
