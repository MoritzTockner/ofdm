-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
W8YO3p+K4MGqAi8V1bkdPvmtTZwjpz1YPfyAIpcoBiAC1l29viOhCuh5hK0TaZmfY1OjK91YNXkp
PM6j7ekaEvhlmqrz+jQyFqMJqRHjD+IKjUN2AyJQjRt2YSyl3YSGqkyRZ80Uwz/m/CPSt6eZdgnE
vO4R6lvmkAfZcdxEPVCrz4dN2VLWtHV8v3Z2HbIeV4RY8C6eVGAlG2+q9QqvuhdmvuGC6dziPWaR
A1Y7UCWpQwQjAtDFWaz2QW+pB5eX+YAmoD6FnSCFLM+WBlBdpAc3SUSrYox3z/tIP+bBZL/Nbf7X
JjsP2cmKZw/JFYqvr6pLdWK3egndSxYgOYCX3Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
fT17FVfjOnChq4a8QJHVouGdyMyn5d5QhSLRWVIefNC2EUb6yQ8dyt+CtHOMNUY7Nrhf3VzDVKzU
8+MZo24UFs5H/ls/CAP3xl3VYwJpMIYWkeKNaG4Z6dRl2KIFOYlzqRDH1N/O3/MzkQQY1RQfcHke
syxwfQY5kv6XdBa9+5JWM1iHPGrFB+Gt8VHYJa00j1K01RPWydPjNy1wzWOm3KlP+uGi9ranQOll
+fEtWKp/QXWT4n7YHRvQEVjb/dKf9SRiRY0JiIHRrh9u1l6ss3n2eQjRhGWik3hrstuLOGdctrRu
71YWbVegNI3vgzUh07DAA1NDOwc3Tt81PJRXaM0zDjD1WjKDJvwPYzkBMbNjB6BhTEWR8NmGA8ws
3w6WWhutrNNFKHJMv1cd5ndkbgKK+MUE1YhNkeZ5jMRNzrZpulzHyrm9SYD4jLqcdkWErqMbnrLF
yVQeJWLYH2sJxzd2MKVek97qkxeSrB9o5UMV4RaH7446VIwWQisVCA7rwnb7kX4GPdA8y2n3Ko6Y
bcxcc0192NwydJ96cMdVfTZREcUiA/dC3t600mHOG5NRp0uVKSK0vqIxIiUjTKzmULB3eF3ccb1L
47KQ8LBrwPtLI5/3YZFKeyRMZ8KVQ6d3ekGcAENln3fxdq2pl5NBARWhB/MavUiqL55adsGnWA7b
In6AAAht2/obaKpYcBfLZgyc1yMSy86PjHyNWWct3O6IL/UsV22zvaKOi5TmrKvlnX5+X0Gi15rJ
B92KbQRYFNtnXr1sB7Ta8sWIPAqR2DX70W4W1J8GIQuT29O4dVJQfgL2EOflTZNuPAxe9ZP6OLGS
rGMU+G/8oJfXcg2ff22YO/dQnq55pbpifmh7K8HLPdZQEwWruqik1wa7QhxwLhkFDkFr8lfkH7S/
hvMoyZXDGOnyB2qq7eypixAZ1fR6ES27RY7ZU6qPw2A5w6gj4uutYQImEStwItVMBElb75xhzHmy
AiqX0P+ioZOFYjNqWufYeJwh4NlAisvxx11b6YgdKmBfeiZXYas2XYRFvHJyijw6x0LnthEv2qpj
1rdqv41H6ME9y+KKvC0tNK70201K4jetJdzwOEXzNYfHSB7M9DjAMDkfbC6dyD33n0sHOoW2Zua4
GXBnJp8n22OL0pi4jmqfsLSgb3kG8/Fl6pykyPWc4QV3Au6ybiDZjvW+/QVmDWMoFjQa8PCckg5t
IMgoP/9EQbWe4BpTUhM8fakLUEhz1nj6c+kiUSZ1wxVgUAUqortXfPlsRCIWYyhVELBxiIoC1L0B
CDpo7Vk/uk4nKX+SRh5qGSvqX57Xjg4iUdSFxgAYQRGt6D1IQLlkL7Vado0El4lXSlNBQ46F7YFE
WCb0mqK04Rz8xY4ECP0MLS8wrGZ0ic1C6WEqoHjaPDLh8tdK/nJQE59/STjHlxLOqnv/MZv2sgxz
e8TyyFrG0gviI8y2OcmZu1EyHK4FCXKtMj2tveac8Y3nKDZIUUvoyUjs+jtwlvMF0/tvd3S5U+bL
RCrYcMMa/s8aFxyZaZOJ2NfYM5bxPXmnVhYm9L034IPEd9kN3flVf9y5no16d4ZydOr8Yl8pJf0d
APuzCRWxI9pIhhYNhSAC1WnjVwy2U8VP2uyQdTvlt4ScjqSFR2esw3y3BLVM/SZrjOaeg+jZb6CI
M+H492Mu04FnWvb1jdaTVLZQNh7eHiskNm1JppUDVSczAIv3ZcPpWbBMX+O71pGiQrLKlMs2rI1k
GwlqonOw1tZBKb7XTSVZFVDSOGryEVVtLcuMjeOPv603EjkdGF308SZuAV8uDEWWt3oQ4FHP39bg
Kab45MHKlLyY/ZtKx753srZ14l5Fwn61tsrnavG7F86lnPimqIglwhFl/l3zuJWRk9kboG9S+DdZ
wppQsRkLLFb/FF/w22ZJ2mjutAtP9QzsHU54fDTrl6Q1ECv/3vrk68l8y4h2g6YJBusTFwF+hz9j
LvBs0NetGwwyeT8Ny7L43Hf8/8yJuR/j3VqSG+dc9AUclRW+miogq0qEN/E47jm5JqFwkOXCq8y/
bK0KD92GPGurTDUbrtTJJodcqFWiq7YIq6toBqUvjfWvSHIuN64tqhWJXSN0NWrHJEV21K6OyyxS
GBjUspVCC4Iy8dBOF8GzGNRN4vJECEHGP+qLQqShj2ORvLnhutB7SGLYOLo7N4C2USAyuePvEDSF
EYxN3JwDM+7zL2AKZ8uLk6EMh6X8nBxf9tQDNAyEUmLAiCYDyIUk7Pymzi4zY3ZOq2/rERXxrhXV
tJ70Y6wNExmYsuLx2U7KB9/RDLozbBPm2zyvOeSb26RBDQ+1Fud6CKfddCEManWdXrwUA5mQGFBp
Q9dSURZN38vx1p/24VNm7u/W564FlBfEClW2nGhXyR89NZZQhkeEL4rAqEca7zwSG7pH73JpF6O5
ZRwsgokOYH1WkwhztA969hC2227XbSi6RC0kV0yqnw0HNjid3mYbWCp/ptBPgpOcWrYBHcm3pOtY
5v12Vmy8MzkDUxJ0g2pb8kcwZzXtKb75N8IalqBKajj222F44lwtrp9HOw756K8ctH9x52BbnFjt
EtOonvKfVsyhLWXzx8TpHTa+pEHfDIIrn4zzPD6Cj/+fVbS5tsOU3wiaNK/VVcbqTO0XFHBUONEt
A8TbYXk2Crxo3h8RvK2b2CBSsgr7hhMvOP5HY8XCKwGBuWFkvJIrz8Wmqa4DN+K6S8kBTzFYV0df
hOUziJrEnuUdN4FVlg60m/OyVuhH+Rog5pKXXa6fS1og4LM0Uey0hW4uefdKEwH+nFyXIBlmqd7D
Fnn9pDYqslUfJMWKeinJBCCc3pG0YNrFAqape6pH8gPj8yEk5vNtj9Uo4VkvLnualu5N4lPYc2dk
FqJByjkyijI8YFdknegCiMv7o6s6slGNlzahZIJvAJVs+L0k0tYJL4ZgAMWYR3NMP+K95wPXODnc
sRJSeHus8Zg+fE1/uX7zJzN7sARLVw4eHwF1e3KQFvhzR9NHDKXCYRiykW6+UqF7xpHiCIhhJCG+
/AgytD3XD8tb5Hbl1igF8SfwwVi9G/ThVa7LkFj9YJKF3wcGEJDEOE4c4efYv0SqY5Rf1lA07lB5
LXA7/ebir6jn5hVGipeoVIVHeX/6De/JYvQcu1hkHjmAFzZ2pEKTsmLm2HpfbxatTpv+B0XcSBlm
zi50n0mW7BKohgM+03xSxTPoT+w8NoYd22CS/yikdUe9zDbp0jkTXdeATRBZIOqcPek9pD9GU+Vn
c+OPRQwcY8GwqIIsIVim54/vlgBe3pBO2W4jPmZWJeU53dMDiGaqeurxaRJMw8hekto9NCZo7rsJ
DwqJC4pThgXJOS1BDFNMWs6gwr88FWEEvp5myzI4qB+KInfdftxtBu6H7LCWroIACqLsiqhYhevs
qXp88LfeM/DrorsUilpCNeiqvq3p2GEhtNxdex5n0f6F1PpNeIRWtm8G1Y9/iiVQs2PYqB0Et8rx
3/19eyYg2evbC2ewXgV1B4ERnXvZxieANOvUrlunuM56RiXHYJPo6r0Vz7dheW10vzdQ+NUEaJ/v
XifC5qxJTrCtL9D9KDvHoZDgV9Hs8mI0tAJBEupHN3W66qvIudgCLzNVzx1Sp9UIAAQZMl45uJIy
DcV6kzzF0JCfKZy4e+XgJGuFKn1HveDcNrue62xJVvuIt9RPmR021D6CuFKeuTYGkr8cV6aF/xtR
qEqBaKIBPGybRve8rrXTlcSE3Wf8KYMkXelBwObB1PAJxktyh7+HvgXqbr3NG/txZ3uXkIucCfyH
bir0WA9L6a1ALUsKiKm8gK98uBDcFQDI7wBmTC5JMC97vU+zL9CKBP8kWkEDGge0m7N55L95ekrD
2WtiCn1ut1Np2MLPfDCC02x5dkPMDtGf+u9wI+uFtjhsYtuUk/XvFl7U8A5Li0jc0GqF/RjZUJS4
BOz7ebmDCxAhYoRurSkv4TEi5Fv7P5HWCelphjz2jAe7jB02SPkQaS49axhA2Wsz9MYDT5lof4Ve
ypAVEeSo5DUrsNgIqoagGsI8TFpD5lMeDkWkxej5NVL9ktZ6PHKCyecqW/odW2UGEVGGKJvXMe7B
igevcjsfuExTW+9PF9JPss2mgEAcpUIgNikOOPNrFNq02Aw1yrxR89V1GWh9II5zbYaZ30yXEOAA
lkt+B+t2epCvVWbpyzQ5ZpGZeyaLqwi24MCGIlXLRenNy5RS2YYkIbrfGc741yZSHQ3nBBK8HQ7+
46FG29NEzr5Rg4mr0YHTRbOHU76KYZWvAS31upPgxVSP2Ic1pI06YValyLGIjfw9PWm4RHpjEuga
g9wuxCUvgo3CNn5zxmr7662mmi56mqvzLSg/X3CxvclwwFM9J3FLoRAy8yjSEgc8d0wzYO5jiYAQ
fPCW2pXgrNm4C9CVIb2+wneQwvPKhxZzEgryq/oP6PRZBbD0+SjEEIKISbhBCGsn3ZLjmwusoXdy
RmXAZ83Up5Gj/GmEUEVIb+pOjj7DvrPWr0VopWXsp056vdDXTiV8A76HS/81PUWLCZrv3wTYPzmh
VgXyh8yxGlMtrSkmy6f9SXFOllM5GCWLJPEyFzAr7QgGEcNryh5dKOzpH1n9V/uhbNywbABJlXRI
RXqOP93yVZ67ttLT1jILnFZOZ2aPFQRuMhmr0U45h7//zIuUaQzwtRtS/XYJQ8En4oCNANcYU/xT
EWWgJzu6Yb0Yp0k5E7RADN7107ESMVdrLK6vql0eqGPi1I9ttHPKd7Qxf7m/g66GQ3InpQvx/R5P
UaOrO8DL8ujet4Ed4s34teZWY9OjKoP2nmvhSH4t+b3Eug0LWojICssAwPYYtTou5q5q+OVK1gSJ
5d9NtZGDJ6q1qDs34wG27i5+XnEY6FOGghRDz4WWUtzbCDAQzg+o9eLHcK9biJgkGKw6ZZGubDO+
jjzY7ixfu8402IdVT2eKACDmm/OyDgzB94kubYRwfj91C1VenYKfcNj+/TWTQbzJRj5DPAY0WsVo
C7ySC58HUE9Jc/P4WzthRZ0/2jGfON+ODBUueGaagEbSPY20g+OLdQxNBrkw1ZddcVY/pgmFHFV+
YpyiLIN/2SGfevRQE07eBgUDNlSdODEFx2jjIcm7d3vdQM07ctRTSWh7aErFZh41zSp2qt/IGMIJ
/3s+H8cNh74L13FwQa+PpB12LV5un4Sv4QP3lHjPecToPBsYpK5Y8RW3LQaKcAsHO/WUyNoxfa9P
o9lM1jwZeGRqefuYgMeFYRMjfE76eZJIP2Yusey5u5QhrU1KEy49uUHN5RigHUtXXEw+w+mtIIbk
c1IWro/99XqYyx2Ca6HFYVIkavpwpX5G76G79B/1XABEUnBhx7kUwm982i+UoKbEsLthPniQgIEP
cs2CU+7W6Sn9JRyTeTfSK+BJoPLU8huTnQdNHODnYVuGW+ajbWBkhDGmlyB2yJ8dkEji1WuHiNsi
/INnAtI+dywR0CYsFF19dTB3t9hRAlO7M5OwktxnWm3gO0XoVL4it/FxQerqap/ZkByhrB/57+gS
ksjPILEMlIepNJxmFBxU4kqQWGH+HBTqJQT+ewqBJUMymIzLCV25f6FJlIPJoC35F5TlKGyd+COr
38MXCVhDcS/cf/h6fW6IepEGn+eVqrin+HVU0SFEQyQgVYSDzjE0FbP+qi1xBF5+n+YADUV0Hwg2
uzuT3u0aCxGfsIRv2vxknrKZGoNxAu1LvZ6p1Pa+m1o7BjFj9ypeJU6+FxqZpkRC6ts/aOzRwwyn
EoMIgT7aQU2mWQSvwjI+vBGJx0/Q09OcmjLL+z81YGCo3oCVSntdg6GLisRSHkPjeibK53tWx50j
5WpfE5+OkDHvva8wsbSXQ/9kR+b7th+fJtj0qOzLkbyDPAvLu0KWc5/GrCX6gK7RrWPbWfRoo8HC
8kor2xXJp9nUSP7kudhq8X0nHcVuZRxBgA3eQ9594n1VuNfcOh8KPGCeQpXkDx7w7qDfPo40yeoK
iU85aWRz+6zjlumCntgrRIE2FU04cdhhsPcYRT82BMVLjGHb84uNCsRm0ytJKrTB5I5yDPBsTwM1
2HvDul+shUdE0VqP7OAyTgbI1NcwmQcUeij92BM/W/SPK0Pv7QwkpCUYMPuXcgn93lG7bv9ag7SU
bLBwc29ZtFI6RuB94ey1mZ875MkmzYAtufAFZOncM7pf14cP5dgWSW7492DBiEkr4nGAdhj+E7kO
oqklasvl0HsVj71WGOSdREvS1PnUL+F76di4u0eRTr7NzWKPR54trzVAIq6YQ0q4U/WJI/40Wa9M
2+vUkm0QlNK3QdSEmOL+taV+kGu/bh7hdu62cG/k8xnFzCTuEyvpyOQxJgIysD5WmFckJxeMjaaV
TxFtYCOW8mFgjptEsyonu1BnS93c7TnMl4IS/3+eM5wr58cjCZHvc4FwdKL1zhjePFINW78dRsJw
y69wi3WamG8No1eYrkIIEzeyF0AUpnY/CEdCdQEAtGn0nWtFUPy1SZ4ADJkzt7Lcah6pjYSS2yvK
QlLR0Xnk1WJlqwZnhYxAOinmH3GQKnA5vbani9FrTxCNP+XG+J/2Hl+rxDZwYTWL+KD0LaU8BGiZ
DlG9wVSBFAjV0Qo8iYtJ9dc0HHzBG1+BdC0/EXYd+FJ1iveJ3MUKc0AsiQeOPbbNYUTFGosQtCeM
LlHEQgC0WXrd3NjbjsLKYnAMq1TPGFRW22pc4YWIQe8Mq0yHDQJUSaY4q0GaYmOjE9kAyySGt3UZ
IZ3OPlPUOExN+0M/sDMRZKUOssqD4SDfKckfFyyxdI0KECPZ6OAwiTIiavnDTnGcVBt5wOZRRA3P
oCEbbm3kgCBwFZaJqIf8u7G6jwxKlsHoRRn6bKP3DIr6+/qpUAdK3BM2lfGOOf1U1sCB1qDIIiiN
bxgyMrE8r9H0ORG4NcFZdkJBTorslcul8dp7MiJlXQkbr1k2n414u/f0O+F2BkEpOhPlkdadLwI0
1NjBkqo0GEOk/ks5iPW0D/PxWgHReGvArOh85fA6ooQmtCBs32NxHyb7x9GsTw30iCNMm9ov5AXR
pd9AZx9wDsNtoZV2tj6FC9cnHraupJLhOTO/mMgngya+vF21d5DFqDYKie94ShQCXUxDi9HfgCRz
dXMORqKII63P2DymNcpQFFD7tKIxtw1oRypfbBFaKj3/oyZGG3HyYx6PrZHRFZpGwcqPGlww4ygG
nnlVPTXie9uXHl0PBJH7f/eTWivP/esxAICRn4hrm4puyx6W7CDGtQRGCvQfi7Tw/nADPThLSWox
dvWclws5Doauyv8Q4iHCZPxS0U+I6ybPZf/izED3zNevOjnOoYulyg6a860fRg6/7CEFhWMdUWCZ
R8GC795frB8y/PEiVQOeCcJaf6MesEjlY9Mf/3Oel8Ihd8TG7lVXd3D8mcq5ozxmEJ//Jztl6RAW
ZQnpYpAYDP+IYRPm9tPN8w+A8vSU/fgqPc2ZJChofHw7aS4rkqgPrf1/WbP+RiEzx7S+7NuBvoS3
LoAUOgChZyrhYTCksN17r+kDKHlCyZA7tdwlFbE8qRKX/HIYDIURrPYtdTDSGhITGD+vh0uBeEtO
Xb3ussR73pWhnXdnma1cw2P1rN37qxUBUXFB82VUG+0DObdURri+AK5+ubDFdsrcdsQ2SRCL1rS3
SHJtb7tXb+tpZSwf3x9An5JhVrzm3V1YJzlawQl5S3CAzZ0crSjuYFjvnMgYo1nLqhe7wdxjzrmW
32gDLm2c38qoX0K3gobeG+/2X8ntXKL/+EQ9EXASfXL9HiQ+JB87Hx7VMpDBBf7/O1V+MUlfddQz
JF33iaKYncY0S/i+U6NtbgueUq50cAmgVyiDhqCiwmySauvs25uXUJ+wA9OF1qkvMAUxeT9NEzQe
lJk4mmu5jvixQEz/WZLp/LD+QFZ9uZhcGwqbitSSogDS6evnjCHhlsHYJQa/glo4aBmonqRNnAaR
62yonJs75hZx1jk/XP3HxcAUAT4ww8zsL3SfOxDd7MPnTt0hHizhM6LN16Z87dj6P5GS2H5pjDN7
uNwxok6/jhsjTJKN9nFzomFmO1222TgFwTQ9vfO2f3gL+fCQi0DqJ6rMYxihduc+6fzDCVxqnCyU
SU+KshV8bt4oPLFV+m0NESjZWsXiZhkUxmhuqSRRYzjYP62fxk2m5RLTq0NrfTBKVmJGqEvgjEA8
N/Jz5tTjdq5qoCCb9QIVTOv2nqPPiWYE13HyfkLchK2oM3dZVoI3H5rn1KmMzARg0jvXakqAv3jE
P9w/IlqjvX9ZKOop0avW9Pt9I+p5gQOvnsJ2XuzOQN9b4ClILCRO2mD1KWWqZFuLVB3d0oj8ndg/
7UMcm9h5MeCDNNW0GsGptydGLXR9UI23M2MBqcwtERbWJTQtcMVkzrPVVP8RkJcxowl/cTcQc8sn
cx1Srwdg4JbKMOCNGKjvDzG0ebxL5b+kY3lcsFWuTGuoJCHFctaXRE0HZcobGpowZ4ZUrG4quy57
w+p+3IEIB0C3cz7P2Wev56Ryifm5gOZMtkLkG27t4fSGYly9TJC0x/Hc+dqFXphvsu81a5eoxXBJ
Kf9eHevyIEYFkqchKy0411itM8Lyhvq5IGP5wcJ6nQ8IItfuPuKtGeQPBY8beLpdXEhnqcWRzcaK
FgSwcvgvmxhUrVGXCZz6NqfOQCuA1aBE2NZYFjDh/Vol7QK0gefxIzXquDyFUOtEtxdyFYek1Gub
XZ0LqPd1fpd9yKc6eoq/zJ6i3Knb94Gb4srAWJ5VzsecV/yAtGHRZ9AkiMqLpxSDHdrAcR8kQFYa
K17aVnsr55Sl3/RmP3WLGQeqYfWXc7iR9/ZJl4tNaolBiffqd09wL6hg9d3urMI39WkpcH7ny82x
yCkIOPzh4q1XF8Z4Yxsy4A0PLqPeUGOYFLZMYJfj9A5dFWJrybZXtrNIk9TM83UCP0xQzZZ9zaRP
YABTCirK+aM3sszEqqhegv/LgezzxrA6ZgglAY7o7PFTVrwFri8r2Nzyb+xj36+bCpWnMQtHiK8P
5cgjt6ScBvlnL8M3ROFuUVL+WfyKrGYh/SVlJ5jGJzonUYGO7lUxQMoD3IOqrLlK2G8vgPm8FY12
dTtz5F1PRMU8A6+Yu5WXI0rGiWBwWg1ezEMRKwQoyg9IEu4X/LEBSfbtBYLGQky4yti/pb+7QeWw
Sa+m5SvDyd8JVEibv5T4FV6PobAXFacIeJNVRkBL3ed0kX3pJRgxAyN6IX8PCJzpqcnO2X4OhxI2
LuN3zrKJqpBjZYzoshcn+G3xOCYikYxZUSmV3LagLwqApnM2Ktdq/FsXqujOLvNCUMaSFDXl2zC8
erXTCengEpcAlEQkEZExKWRRrJLXTGmRHxtU9Fcfj0ez4TDexmgqgnWw6rrc/p++ctAImOH9RXHA
PMbZYVmzyHu2QMCmjNi0y63WYAK1l5dsEofGmf4MdmI4/ya22UJnrhqYQ8NABVlbkpwuQC7Us+8p
5V5cHVmmip9VSYNXoHdREXiUVfh9XfAStJS+9BrFz4KCSyhX+NaA8tE/0UnFtzv/69r9jXkWZa1J
PrEltbBdSe+1WGZV8qRCWIHvUtsaFtBgoyMnJnLPuzi4Ljtu/haz/YP5i6ENy3ziQ6hz9bfjAPb6
6Pzf60ozQYNi8xgvmdUi+Sfq6c8L2bpsSXjjMbOWDgFRHmxa/0HJMZDaMAYeMSDinBRchB8mss3+
XKpoTvRf3oZ8di3ITksKulSAlDuvvAn1F5an/O7i/Ogh4JV/VYswgEqooRfyhj1zGbKw4XIKoPmO
xF0bjnzOOr3ps1wugRcDoSPc+YPQV3rVZ1nC8KoNxTmmORhYYdiyJZNyQZGhRGHxl5LnH9mEZ/bv
U1LsXCs1kBN2+wUNbqK9I3H59R6+GLV7+7KQVFDJqRp3lyygnnCob2dJ+63BmsHyjsfL9C1oFSLz
iqlDsfvjKoCOr2JoGakp8hcI4L3Whptsc9G/IIs7Jp6TfQuLnZZGMYIS+8MrkOYX+eflqCxzRX1M
VEoDFW4s4y82t8Nxt1ZnXi0GI5e6n+u1+3gcL2/57LNkBQW3aJVvHVjjJKQF8+0MxL0BZ0dck+IO
R2mdUTCIMtH8PrRwGkXs/bxD43tfwlFfJgdrvXePrxS0KQmScD2ldZXXuFZf2AvW1nwoN82o8YwY
n4NZcdheWn+ci3OEscGF/lRWj6gmWWRuS6xaHAYdwKafBQRsGbGnJZLsbLNgF0362a6uf7/CyLEG
CznviAq1xM9fqfQLQJUQzAkw1mGiLicv+4bWjVvpIGKhC71nRIFugzcXO0aVvWVqaZu2pwO2sFih
3FOSLK1WRI8fuOUFGFHRg+5PRSRQVH1sTiES8DHkiwja1g+bNoUBCba8NunvpedgKB6Xuhxmr+pj
8cKB3AH2aXk6DrRG17/hlrKpOzvb3RJECngEcQQMWR/88X7TOFoDMcwFkNfyysrhkTm1A09cFV1y
GAuyI5Jx58GjbDtD8T/3QeQg3rq7nEdFxeYbVY6vxXNCwSpzlxRCkuWccZkQRcQZHtXxXanOII07
ODPp2XKK0bK/prZQ9YD2zcU/PimLNWGTiQFOcBnwq0CCCzh/0aGW/UHoaeSEVY5I8ZMHZRfisoZx
qj5fmh7tdTl6vd6m8SY9/r1S/Gu1IFGDE2/A6GGuxqtL05uIg7yyY1sCnsq2jCdsrzHwnXojMeRH
2lVbLx2ZQSPtkPMZVn9PvhUG0cMD7opCiNCRzxDB98szPy32xXBtrbd9fDb7Dzx7/7zBNPwOKb0C
hT9Rd1Pgz+Xc8yZHKKFtj4nhvjGzehBKn3HBd6p1E914Ux+T3J7kvpafHC6mnURoPUjiGl0xdO1N
E6lV7/tqT3rQBVdMSwlJCpHcOrIF+q+jPoAY3D3/N1WCD+OaK/9XFBIfzCX1kJLmok1G4qdW8FGz
v14KiCv+PZblh5UPY4Wy2WHV4KQSk8YTuwDBH3axvg2nuAAHdh7cY7WCmne1HhyBBc+p8GBuZ3Ap
DCinPG9z30I8NpfspubEs+/GpSoMX6+UTZ5dNAtR6PJLkUwJEQXL4HW369wuXKehprUJEvp8k0Uy
lU6opHf/nsZ1Cq+RZkpt4F5ueTXkmSt0ojieq2F+sssSN1qMBgtew1Y7bGKJzDx/fR2e3g/8OCYM
gnap4EHRO2yiNCyB1I8MOjxftUfYkHsrQZzQKyKQv/qm5wbQK3iP0HpnfdiWYyY5279l59hLSTG8
/I5aXfSG/74NnnBVrbJAMwtS9uYlb3618bBTL9djipsuTXnqMtnbN8WRjxt4kSt1f8ywjZZExcbC
ewp3DMsAVEUAL5/l1oe7UQ/h2+XokCCXG8ZHBUK7t7iUGDJqyrsEtql4OhbOKq/w6rjY
`protect end_protected
