-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rD9upzKph16UsqtDqvcCWZvHW1bLuMXi9RB1XZPv4tkIre9ZOmNqGSfLx6tfAgCcGndE6u3dpJxx
wimHzwtpsPSPLZV+0WQ2kuyBnjLaweXs3lWFiu+6164IMjK8wjrVYa/YB3lZny2XmWsxhGzJSNUC
32fq2bLBbO1/Ysj9Q6w2MWOg+Q40u7c6Ertu7pjBYg0+mJ0mLMvivTaGlFfU22hP7hHeWePEZHlc
bcZaEjqSn9ZEUj63rNeUHZdIT4XgEqgTPQM1f4d92XC3h+0RPq5WQfoMSWb2y1WfDefznVSUp569
rF2OM4COdzHROBwd5C1MvOhyUi+z35MHYUruKQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
kKiYeMRBFrybrk+Eu388+9+wcH52+1lAM3nIVC2zGYtEF1HdigZTLlQgziIMuvnLR1BI6U1/NO4l
xO0jj0kshiR27vzZEWVTFTa37K7LkJUnYHhSnFmNdiclVOzY8V8in1mDVrAr3084SeXRGeyEwtez
k/Kh752FkwfYji6feZQbXq7376TqhweODKrB8MaEd64MfLSWcndDMmR8aFOpYm59Cov9qj5vVqEt
/58pqfIrYmP2pS58fTFnSI1qLEWNmGDUljm1dKB1QvBaJ6O+3R/bhleca9irCrZ5RRfJBExMplOA
GZTVa2w1vuo65z7aXn2fnAkvzsSYslQOlzyrN7bzMAWgjkI/HCRfp5izjtS8zik4Y6aG5KULUF7q
6tRgR2owg0WmdLyCVMmTbyanjzM4Tdl1tOxaLMLwVhS2d/NPf/4lhCJVYOtwG9Qe9gGmUrOb/tQa
lR+n9cud19y6JivhancKq8QQy55/1ZEFYeHK1NOHyMEmb+D/5DfmsDKYZECD0JgjouIb3qZkA8Aw
/n+RRKngZxyKC3r1KcXHWzpZjgGTOVpu07A/a/qg+hlBK3AADJeVoMA6YlfqBYHOEIxPaxhwb2Y5
QP4EI7a2MaiHLFwIfuylgCY6ct+1/oKh0gubTMG5z7QtoNjap/XMDN5zmzTJD88BGcYzleeQQ5+d
nzYYb4uqPY6IWgCzFXPeLrP27EvKo/7cyhdMvjuHBmlYqHHAldokZiVqFBnLtzbOLXPJF3NlOQzu
w++Ib/4VcJDTpbiNSpBFI5TSsiljgx1YWHZbvMZ2mToBr4EBgg5zEHSTIaRHHnKEXJZZvD6xj9MF
ttyW6h/mWlGIljP78F8SnH0R4XHkGU/9SzUIfdrLQzuQ+tzK7wx8DsFHLK/69SV7kP/eY5eSI2/f
V9qAb5PyHu9eIDP3j16VjB6Qpj7EOgUGcS5lKuNgjQlHgJQ0cl2qSVSwE+J1q8dsy5Rml7GgyWPP
+KME2y6k7N1RPFJ6zn0A4qwBJOGbFn+YG+xumNOtS9rvOBakTGnWxa/AaXZSn5BEytLUlZGOjoJD
xOwgpN7j/lhYCaXcy6fwL/XymOlO68VZhc1u9wd3QaUK/X3NrsB2quab23nGgMlVE4TIi7od20KQ
Mz5BfN1Bv9Kd5b+60ePLOT/87sL7kTDBMcfMndZBDOp1dXPLy4cJCruiJhInkT1lQgV4YCdQUznX
RnbzJNc/WgqhvMyqCziqspNqBLhVzpQs6wVAtiNa+4aD1NMZIfzZ+Uh7RHTT6jPT1gpeZNS8WD+i
fCQxUcqf/pewgLVPe6aflkJr7UuTBGKDdn9r6kkJbCSYHpX6gfxnc6JIFjm0SobiML6xdRACSAoC
1QUZ5t833FWFh3l4C99o4GtajRFdBN3Hm33xK0K022hGr2bE7HjqV2KdzXwjgB+9H1tHmTY5oZTq
rjYWvDVyixpOLh6Zv3o6gRom0DnyeIEB037aNe/qzlP0aaQoyqW751OYO5OskscDb8+kiCRDKzTg
mIt8Fdup8DgAqpQmz0KxKN7oxXYsHGdjprsQBO3AIqG2ygUiZOEEmivGqWfGQbQZHMwMrdJPDPRS
Boc7iCo+IhncnodxFJcOZ9YxdvfhWJB3A5MtKO8SXx0brnchDJmzREoPTN5nfBywJKH4o8Gt6JT6
Rt+9ELCjTs57jfBXWw/Wb01GiE//7JPxpyaUQLqrWi31zBMHSBNw97Hujz7dz9uu0IOeyQicyozg
ZGObojoYY01quElpeoZD2J2flX2r7HlHszSwEoiwNyCYV2aai7D9znz/hvadH8I81PesZagTCSwc
UEfqQJuyl4E/EVwnrbr7BwcFVudpsQLWGJKGjtdHuVkhpxpSEGUoKvkO+gJFWihZE7E8DqBSXodc
gaglXJBVanrBH8BvH0qYGYKJWkGkbxeuVFkz1CY1XAQ1L5wQ1FmGd7/PI2AV02wOBsMhF9nk9RGQ
sYLi4poKlXA8ASqtPz5T0UxTpBadWWo8C6K9CKXGLKdc81SM5ClTSprbeD7QxXZ8GaCtzhZGK9Yh
JK7Sg1Pkpq5UHup9n1LQLF4J/pASZGMzpWjcyLRNdqLviR6ZoD+YsjZ+sieFXExNQwWzmsP6apAh
YtJH6WDNO2lULz8y78ftwifJpk9YHj8FsAJ8F4QrCVBxtB0bpKR4wZgAsfN/du4XIYk5Rj+vrt+C
liwEYGZxyWKty04A+YMeinD+MbJ9CwgGBrKYfH/3MxdzUH0m6U4oedBNXonzO2NNEbsxDt+AU+SX
iKMf3j7O6OUIGHGPl5V6Bu59jz+P1ycFn5dp8dN/KLmNmayEUP318fECbxBNVTG7E8JGTr79Af5U
RDgNrEq3E1dTqHsrETL1GdSWdZHDGfQpPGLThz5u77MBXeZPiHrvsdTtgbCzicgjDqoUbPKcSRle
HPxIUmpRKsz4+RLgdzVIvsTxrNjnQ7cDOmJh00B6AW/g2MCmL0XXVUUSVarQDKxkwW9Y3TTUzZPS
V7BD9laoXWocY9ml8vagQzgl4O/aJCOpIK4JcBnZomBmAlrWj/joqzd53kNCdeJxc7vnKE3D1Vgr
S44Wx6M6nF+bHB67L+/Zf7gS6dlrIulmKmb7QoHJW/P3gtpbPLs6QGz/3lHRX+Wiv0U6yFpmLZqN
0jTpCmxxg94+izd7myyYc7syU7mqPhLD54+BC8PkcQnoTqq9NdbeEV1i7Gw2zrxlU1brUEEiMtAO
kfYqXvmGv9XgQ/Wluc6GebbWjpiUQBr6okDh/3cwA30TFSkvth5WbT+vnfnE6SDo61sx4bzbPMRd
1yDIU3wIJo8uE06dXaeLOSDavQvOSb05pA877t6rvwY6MSdONWWPpGrpGfTlpIRM8s/F6HJW01SX
Qsj9kniznG2MbKEBveBAcF1vJerkw/Q7+pn3hcmeG0zLbUcwy7n/n2OE1Gm09V+xRm+TFEa5GDPl
VKZEaETyZ7AYI8LpBYKjtA4eiWJtz1QgwtW0IM9LDnK3Cr1J4RpEBbmpJnjzXVCIuzDPoSGlAjbZ
NacZVNGK4zY+LQlO7kQuB3tHKAe/mShqhj74nSsSQFq21dRs9S4mtQHmz6qnJbd4md7UCiDtZTP1
dpY7TxBg3ifDuRpK0PPtqZdnsxfbZ7DnpDQc290P7tIjhgkskRcjt71mApKFi9pDHI03sXjeTNV4
vFMelL35yFnXCMukVeJ9W/Qe+vHHfLIDVl0Y3RGhN65yxIcM1Ksjs8Q/K+Zgtvx2LBMQanotkEfQ
d/9aKDs15inXMZcvgR315sYC/mK53S4GalEYalXu3a46N02EBlxj6dx1zLOVQOiF1LdJ6C+ES6o/
g4ba/Lm2cMMeM+0fdHaQGsLgqKrAPwoIepNAcoJa9yoXCtXuIAm5TrKqBl1PasN8MsIwmCeo2gXD
F0nVaxB9T4Hj6t+UvsjpNhk4LUxPoc56YW8agXcVeW4mU/3/uyjlXXHWWcyjWLGOcQjoDtp2SdKT
0yhZTQzYx9xGi4dpM9GhIvGtNsvEhS34B6P/ISn4K/pO5pZxhgeb4TmKAmAST0o1gEAP1AVMTtuC
8rTtbMRI1jEb1BdfJPVGuD6Fhk5RbiAWcjZH++2DrokHw5Qc+SheW/bcKgZ5zqKfSmX8iIvO6aeZ
iZPJSNLKE6oLyOx8DrsiBlzb66qzVto3kX1Rf5nYOGnstltLAC7HdbNzJ8ayXJAgAAq1/ToT0psg
oHe16Pxr+vyQITeT7PzSTy9LyCrvRJZDVH0Ix2JSu4GlcM/nHgZv5JLiRPQgeUMPjd0ErrZAotTi
BsqKh16+l+i3t/Y55CDBPd2t8+ORMmHry6F/CIIqhgiSbzyNemQG5vHzf/MzIUEw85TZCNry+Al4
7Cox2jmicoq1wyYQv9ExsnkH4LPzIpdvruNGM7WNRBD5VWi1Qg9VWSRVcuQnJgD6KMoa1nzmdcqe
URhASUaVp8KurgMscYyhobSS8udH6gRxZY2xUEvdua/nSlMnoI0V9t81JvD5MllCABlHyovLakIB
oD/Un0qsUB++D1ZXEPoP1X4u3C7Ko/xmLB7DS7lflZGxAGjSFsvVLtz9zReuL2t3vGBvSgdLQqgy
lhKl06Y/I0Q2cHkSZi3GwlCcFereIaD8HlGBEpxAjyC9yW2uU8zolmfZApTyEvypZMmQvfen/dIm
Gz+yM8p2m2V+M9CdOTzX3jsYJYHqDY9TgOs43QHaz+R0UOzhJsw9U41XBwLdOVtaKtbtCzoFiRC3
hotqY61+IuikCT7Mg7w0AyTiBA1UOuOhVbTcw4R/pSS8HuWUSTzMom8STkKHOQyBGZdmRsvou8po
uY6XWzp4vYWY5b4CbTABJ2H5gPgeuhdarFeg2kXy5/3s4UfYlp2lu2i5aXcCxKLWxwT6mxLgOcwR
OBlfGnCdVgRstrHs0Q7iWuiOW9NvDkzag80TAUyno0Q9/GxpDIDyjyJhRf1uD9Y0uaXG0yMnGFMN
HCKVeY5jsB4BnI+4dRcGGZif9IHQ947UVeGR8xWGUH1qv82GNafrZcdZKrRiaIEkMMbA1jCrnx2+
E4aRMw/8lcKSw3W7QWJs4LXcauO7B/HX4DpL1hbcz/zJCLqEsu8LABdP80WMlw/lCRMR64tn4bfX
GorG/JKNEs+TyP2h0UxLaaAp+hyD9z7qcy9F6ewlYatthvCnjNn+kg30zjHZCD5Q9NHSzBtAqy/K
MsNjYuYu25+RJOlxL0A/brD6f1IZrmCbGNnNy8qU/ugXKYJ8LXfOdoqA7i84kmP8ZGOlljJfTDAI
SKv1hJUJ9+LpISXibH1EmAMKRT79dLpWewKQNqTWY5+jSMTzxXk1sd2BIReY/uveEwIsChhmQY0r
hHh/UtKQFIM8njE/wM5AP1NW41tJHyWH0E5TB6YAV5gJV8fXOaGJ/OQtl/FXaHOY9RKsOb162Zl7
EVX0iJAKZfgoJg4Sy5A5NBX8LvO6FI2sF9CDiFZ5c1VeGNloRvX5Si7jHFKV4rRkxHBvrnAhjp90
cVZHC0RW1MDdSZu0+9hy7MNeUxxGqWHbh3s8r2cSM2w+dDMlNay8KfVh4GhO1UjtYDKwjT/wuqC9
aZ0c8OxLCGdqnyLkZA/dld/0diduvh8Va5Cn4IZRdd4N7GgERADVhZ8Z9WWtBYV8SrrfqPiNNqfy
fjN2nYRNujNEW/3eRhxjBKcaW7RVGsCelkIhz+Rz4xgffAQrroJ/O89tspLTKtGCqcOr+QMZlhGp
IdHqoQQ37d1aTCxcIW+PyncGlWzTUjQrIcjgngxS8TIXx7XcMBT7v9ui/TEZ94JLJmjIWvtVGWC8
E7KGHqPTcrWu+zNN766MfbGBSalqwX/bifADa0GEhTTqfqXzllRcBoD1kOvUEeMlIctL5rqvpjMg
7uZOfG1V4FZ6xlctX2Kznb7TEwJmPUIp1wUvkU8uOfehw6N940t4s9orSGVCfvfrvgqL/cOZZnKd
uG+IL05EMEaP1TAKfOLJ/oA62qO9Mno/qaym0UlgXJTnjAcNY7Z5nF8TIhwi6TsFYBZhd67rDgRR
r5vDoD4HeLgPmxcwJGZRlfjjHip2BXr+CpBWhCcQA5XprP+ttUazSWyKDGkLlt1pB6M6cRrRm/Ra
PsD6rScfiPnr54aUo4mhWRoduRzjE4jEeIhy+4OsBL6qZn0D6HNx2AfEgPJYcAyiAULNXdWTPbJE
Xq4/YVLWttr6R59SNBoDnbfh6yhcorZVKN+403+dIXpDOS1J2MGDbQxb8jKThMiIV/pQR6UL0DZh
eIKdMaYvDxpmrNySAVGaIkZ3YTCjE+AJDJhTldi0mw4R4I8Cjhc0sXZ7XPtwNlaAxopL6y5AG2UF
nGgIfKqQFK5UZs5JWt6ESJbXRVhoQGB0srUw2BiFkG0x2ln8e+TdNA0D7yPjNWn6fYSkliAVe1EP
353qVhNG7KkRbOOaDYUoH4W7o5dWUhsH63DVT836ubdU6C5aYWDUHqY8An2FFmWAhtQ6qPzrjxBK
ynPJ2kAu4k0tcdcm4wxiNDtNYBxIk4DzrBwc+LBxgE6WXOqs3NBOKWDoTVRkzZ8he/J+VcoYfyfw
ojZgSY+zi/A8cokDQr1FCh8E3eOFQs6/IVE/959c1/FFzoaGuGb/CNdD0gsfKhPM2/hTkCPDgDiK
+3FKyehZA0k4Xqz/brO/ls5SeHAA8/32M+drDskAwtzPHfIrBVzBUlvQZiyvhh68y6xR0gtWVw==
`protect end_protected
