-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uDHNMoWpLcHyLFCZPXH4O8OoCU9bUgkoYyY2+pVr83KL4CGfD9OmgTwjw/VtAsRDGxPjEHmkhyS3
YrWO5Y0WU2Zu6h7hotHMQy7qzgyBXFrEs+f2va4XLq5oOymgbKImmDzStVT9r4dLgPKoBmXgXKXr
zuYX5xfbSCKCzOQkLFxRKsW5X7nqoWGlgFeuNhoEVenHw4ML57dqgiaCr3LcDYt8zI2VfntQpfCm
24WfKW2dG/pVAfOc18rnmySi1AD3hoC8XxIRtsppakesLJ6qvB2YD7zipU12rmsEyD62c68w12nj
fAudZ/gCZTZbm1cX7Ef1zZshUdmJenpiw3uGdA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
6ozodpgvPbbHudVNWgPWHDGhNB9Rq5QuGmGhu/GKxKt1xp3sFtpeOaVlMcinvpXm0/CXA1XypqRY
BfwdlMQ8i+pOBgrIi/82SKtYgM17foQnCV9yudQZwNkjf6mkLMjFhL6HL1vZAtfmp4y9NIC+4+nT
/+nJkE+bpuhGXGBQ8vWeWANpkbYPQP9KuRy3kSxATqq3YnkNo35RmBO/gZ7Gw5ZcQsyq/eLRnVGw
85Hpae/wQGD+lvtSDVO49VcYf1KMh33JJ+mh3ARI3LlD6rJuC9RSzDZAT4JyLmcthcG4SJKf7ME8
atnJscEcNS1ziN3+dGxK3F8BDV0yZImh31vhihI0Xt2eywY/z/Q4lDdPUZwl/aeyS64TmCYidlWO
z3ZSs2OmjC3xk0AIrFvhiTJQy4eqACv10wzN25AswDiuPraaMQusV8+MoUWMSoxh2NJAnxwgYl5l
rkaIRyqtOpPL3/5JHyfuQnMwrIohXAyrjxmmu7Q0Wnd6PUGqdN04qE3Qp+AfiHZAZRIuMs4OQXNT
8E4TAn5aOzj203axzXN1pZ/Y9hwDLNlAxmJVr4B+2Jql8Lpb8Jo8P9AsHUi97v5SYj0d51LitcFA
sy8PZ2mxvwmCezcOD7aQ8jFl3qSeYhF11N0Ah27ql+Ww1Wnt3Z28shGOfkEmoh7TvmmemPJP0Xle
1mpLmtaIQuDeKLUCMhNtV1Y6DqiVhU/IS1V9S21gUasljUs1nt+/O34cApTf7zKhkHi9wM7NQGHg
sgriEKBseNxm2dggWdryfjAgWEm5hSHHM3jg1QdRVtUNU8dIFriibNqY56E8MioCkFfP5q9U1fGQ
A+UjsntIeiqMaARBa4l3prIuJ21KUTShHHkbpgf+LO4ejzosGKURbMuKY5q7lZitdtluVkQE7SzF
lWwCSwnkX53hhCdHB+W/+wG/5O8XGJ22Vg14C5ikkkpr4qzBUs9YHiULDrJ4DLq/1LH7mK/KHPBm
Gl6+N2lTog4fuY77dfDjSi4pT4GvbhtBFREqz7BxeASHvAuUvv5RO5iHXZMiKs7pNxd61rmxyz+Z
2WVVA+W+S0qc2sV3BaDeRjPDvNPhOSfwUNLEDOFs+uY93GlMif0no7zHibJpn0/DPWbxdCic9/fy
ES0S4ysm6q4v6UVJaQHQforOadkVATwZrKhzAlfiJI9T+TYvxkuvDeoRAjTMiPMFo40A8YC+o0Yq
c/Z2h5FTFRgCXqnQlwoyDOxDZ92b7b2Dg1A+ofgIT3v0e+ZvF4rtRXSyZw9GBJH2B5E+tk2sQNVM
6ljHUjIYf05LwvoI5ensDlcsol0QVwmQS5B9GYe3RVJwGmD/x/O8Vxs9o+n8e1BoNAkpkaxYfRP1
qWCNAFoNnnLN3JMC3agj7ziEcu16nyq/ZLpkXKmnKlBvoYxEwdYFAHyeQmORunXXsQQiKL0kVUlg
HCeV11mf9y0vL4zduW4Pvywpi+S/ErjDwiGRMYZOr0TwiVanh7yvqKUdPEXFV6qIlY7CJXM/Xc1B
woypDusVicoroVQfL31dIx+geSKeFHWjmjdnxXAEEwnMkPTg/B4OJQp/Ey7NiGNcgkd0hsdwghDk
3y0JOLTrtYfC9kGXyhZYs3BLvSMeimW8gtwoN7oDL1CyOyo8a98BzCvC59ZlNsFZb7+q5LCSjMh/
iAutPnKNKL6y7Efs/rLCW2cWoearHoYKVt7ZZwpDLvpYa3BaiprQXq7VfZh/HRxanHmw3NxyOM0x
7Jh8m65aPpQWZAupq/bry/XIE22JIhq1Sx0GW6zKbPRrt24I22J8qPYKqzUPn4osBpCLYxzuM88/
KBPVFAGUemwFmuG4B5pb1yYUXcokg0fy/S13rWl0X0FwP9DI5bC3u25FMyEs/GVK8JcbLatbat3j
RvJItY1sGABAcMyPGyO/fEgwrS8X5xkEauEDlwPaFvzF6j5frqldaIDIA2WyPk+QDZRmhc7f8NQt
7HYiBEwpWe9iowtDnWijNp/W0m8amGwvsWdug83fI6nwNw7/lsw50uFWd8DIK70f/YaFNArVr/7/
3/nfsY0jxAPLz5PLEjNp4CPCmjSZDvI5A8buXHUTuz2tCnUquwxK37gJumU7vqwIrboungVJRghL
TBs2jZkvJEcLWc4i4MQKb7AVhwoKq6eMoGLlQNE0yRnp1NM+jwsaXulCpxuJPo83g7oNXbYp4/iZ
hdGtK5K7d3z77pRMLEad2nsG7WvJ+b24SCg0Q0JQDwBY5L7tNScnEVrjXfrBXSLqZqT8EJaszYA0
MUJNoa+XMSJhCk8A4+nSwfhDOn/aeevYe3wdxsa1Itd3MwywASSCLDzMIGDV8QiwGvkmIegLdMMr
fTjrv86upts4YyMvkvSOBPe8VF4l34tLVFyAU0XsPE8/wFuWHYeelRP78PnCrqtbte3vea4ThIff
naCIY3Oc4qpE4HdFWvxyRLolT4a91khcHizWvFsz5+x8IC0OsdeDMI8N9UdQa5o7qBOf3z4UUi53
bWyEf44jpgbvolKdXHEVle44XoNzjvMLGYUXsIzZe1RTnxDJm8cMRv42FKyqVq/bs1+6WGoIpD4u
4ko33s8d98EG2DDbtobFf2biQbxUenkZNL4tmPNhxGoNyKXPimfZIJaWm0rlpJXkwjhvoD3dN5jv
yPNkLLQEF0L+RN11Z7TUCK+h67BqFpQ88oLWfwjsSc8qmj3amkjMsHYmS5yR41oKjzlPsnr7DcJb
6NuMtT/q5iPYm7HhPTUIX09mYimp8sHmvRYjsToZXX+kuMkK7Pc9onOCT03DsZS7zHLABGMshC2p
xFt/19Qv0gz9v5x7KxTItm705g2ymOnDqmSvyMVxxsFRYD/rNXM7GiJ7foe3PIz/IuWo4/ze43jK
WWA3e1FhFAQtzcqZCxkBW+7S8Lc59+9AwQReCuBiwTijmAxrmwpH5I2DG/xZKMF1c7Cu+LHDwmJZ
WH6RUyvDtTg/MdYK4Owsy//yvtLB9zP4jRpWd4NeGHSfIvDGDUbXzGfVlmn1jWFtBIvTqBcTznd1
XCjwHtOP379zHqbUCLuu+KdQuIiNNcVqjPn2oKkWBkZNwFf/nERlVvBnSp5qOloc7NyUqntqZ/OH
VLWu+lyUjJ0y+SDA6DNl8nq0wZPAa0Ko7IG1TLecymINxFEVQLBqOJQ65cRiXcRTpmFTsPsn0qbL
jCJZnBqbyPKUAsQqeRps3ajKfxm6TxmClnaTEc57HLjSB//65q9YlkYh1LaUpphzrQuRtdHkQ79Y
fRmP92oVhPJkR/SEwLux9syogrqBxIl7oJYX8O+LGrvaNRyoR1m67BbZobRyKP2H5ifupCCZVVCA
SELV2JpmoW1oM4R2HC/jk17voOYLJKI+NfI6jAinQ4fPsaLi6R8U10h0bVfj6Y6sNkC7IWDyPG5Q
C9UGOL1U4z/7OXxc52PPaLjZB3AhGfIIs284YNtHxtjznmI0kS43Dxsxll3clMQo+4fsheMC7BEg
IjDnPH65MtVW7Mm70RT/Z4Fo89N6jRz6GPc6Ed1NPe4PnwVNj1nS/BT1Q44cRJ8kV9M7W0b7i9gs
nlvlqGn7UjW2sPn1UEuBC83ERi9Vu60ZYkA3/cTEKb9xu0a/o9fGpvCw/REFhY8BejL0y2+CdzBx
+GrCxWY4lT2525+oS0+fYD4OuXjXHz6VonulFAZiUAQiSOZbAh//YFGVdFjtMhkv2xBWdDXqkNlK
eStoC4TdE0ERWVH51nZFWhOGu5pF/ZyqRhG4iTIKpodusE3OhCJ34IW7lXaoec18DlPGvDPKVv8i
nPc03G3bLlCb95gwdLIzarTN2D+gkpLWz8feaJkr8fijw3BkLYaMy3dxGhkB8VbMrqA3vrRjSDzf
ok6G7cd/R8iSwRqbtwrJzLosxjGlb/7YFaF2eJ4BEfbgeIdTWIxYxLHiNIchUtkvcz9Bo/xZompC
DcJwArg3BH5xiBi6EkoHJlOc20k4xt/pr5weQwtkmSFibjQBp8fs8ukHTrdc2eIQupcGUS4M3QQD
38MsuP75mxX1ahX6Y4Xg3iDfZ7BvYamoFcmYU8FRxJLjViep/y2fTeuYS7OatHkPlYtvKLgiopsd
swJyzPW//JEgaKr1HnvFl0+gRWFxNQ5MhAhPsuTk1Gdsz0AjriO0LvsHPxOfDHoL284H7sWHA+Iu
jLmRj6EXLLjlrde8hORC6FZIqqGpnTxuIZmpTzQ7KsgKQyKkE7FsGw94bny/Om4yYo901vYItjzk
5pIzqdASqBwnz70pWTU1CVhXPWYOAdO1ajGjrTZyfH8lbnBqZH9OJNtd9g7bJUMOnGTE5kqsY4KR
IMNkItGvB4QAKWqleikJDe4J3ja7/jgFHiQEFI4yIjGe1wv8aA62fZ/PlRoEPC/JytLykzwGg7K2
Vz1AYF+CB3BlebfsMFjczxVC3eKhj7oEGimrGNFuMCw7kKSEXvqZruAd0B+VmyCkVkImAy/n8GWw
ju3ri6QOaIBylgjcZIcdNyJzmJfHPQ0Wtw3iAJ2byCcetvW6o2LQbH+uoWMWjsD7zl3CJ7FaOuYZ
z2dsXmUAjOJsK99u6VZoPwcRREmMYNkSh9x+9sIcbXm5/9NFuSEEq1bcUp/fGK1b7yaYlAnYC6wq
m5gcOgkD2LS7hBUL9q5TlgJzhw4Yv9zgsIzUyKfAZLZjRhjd0scbc3HOnJdb/av8hEcdnH01Qg0k
Z+JiQZfQR1Hd8gyq0bvbLsmyMZV84Rx+KNy4Tsu0pbeOd0UeLLl+PAYAT/UthJbfEUB7baOr2N5t
AX3h1p/0RHgy3wohjz3HsZsC7GiR2zs4YPYDqcSFTF1G1EK92GfY8NpyPAh5gbrJRnRv4V1NYUxa
ALXqK0fiWRjFUPNsTfaxUZEDF4NBhPAnWJM0rLW72o2Zj/7IQlgEoZp5mI4q02QRwElZ7D077caz
W9ZR8VM6PxvHionK0YZOYCSHanldfgKcQd5PZPTJ5vLY39Rrb07F1ok4Pr7WOAXJIrJAKYud6Es6
1JMWnb1rmyK8M/8SKivhde2TaZGwzRkwabI0KUK4DNyKxZeG5T4UTi8KsG04ra401+iHbHx5TJJH
jhB/qni72WRnEG8yANKanGN3ykGamAHlnaRhG4x+pwl21UCbe4BXTUxkQS6pV0XA0FpJUfOjSuHh
+MMwntWKeLnrI3+DZw7Rq9gL02xBkqoxIELBuvi08+lDw0dnoAb08XRVNv05lBo9U4d6HlitokEE
0AYGOsfMKKEdrSAHu24+BZCcrf8jFy3SFsR4g2lkBhAna+rKSmta6rzUVdSnrj6zro2FsmyZ8Kr1
QB7B3odMssOCnK51rcjl2Kos8RBI0QDDe9JlSzlqZuFBxAVak1VfNAlKOTimQzGXRcyieXUZiP0Y
Oc2RRbg6gepoT0zmmcfeq5DP0kbQXsNhxUQgDkRaVA93ybGEAy3c6NNnLH8Zgng1OVMw+XOb7fIE
AO2DmGLAza/AyyeSDx3MrHyCLG6qNhlx545fptwVzavSwn//SbTBIIGij+5NskAulHgZDOYzHPgE
ui8YRbxFbkG5aaHN8iIn3C6W33I2spCA1R+OavtBqOwQYrxqf/uq89a9zyIV+NUEjmMmfQUNdNMn
tBFdb97Y+pO2mgFagVmrzTUjmGXziH+MKGyz/S50e2NgJGhAr4VegtXJYH9xzx2Eg1bKsgnn6ncl
TFluY1JLwXYTipfMNSpxwbKq9zE2CZrDMVu3ACjrDhQjRiflEw5Xokz9yj+XW9cPvwOQda4rqsHo
wqd1aecqCv/Et46l8N8n0D3mNta/VZESmm03mQr2WPhEUjE0MQ+d8qDOWMcGHUem1U4lgtON51S3
qU3FB0tDPY6LFTrN5BLYkrqs71Z07xrsaN+tcM0Qzu01FnUNldl1rrZl/rX7ss3PXAErufq5ZC+E
xRwH/vOT8FP+gmMWrQk1h5Cf/PXcQfY3fnQXwq7qb3ziEt7SZMwZE7j2Z1jghQnO/pl8vlx9NXjR
R/GtflRZswyNmwy4gwfeW1J54owwsJNArQ==
`protect end_protected
