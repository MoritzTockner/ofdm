-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ppJTlGuc855unsr9DIOgnfxT6B6M1+7FslzN2cFT9qUOXLU0Ms8rhagblDYSJHh0hENfIMv1gS0e
6F80zDJgKqnu10rgf7PBVCFCDgYUBk5a6vTtPNszev9w6ud4vDmd9DU+6WIhOunOUzxxirt3ojrw
mepRp1C/JkrDwurKPVGAhcxnlpBUDNHASckGAElBfIs4hdaG2Wbb/bTVP8zXsvDVVyBiCFp1fd2X
YwYpL+vU7L/4tkhZVqcXS6gktPmCFixhMqPhu3+gvhMFUisXdxSgQ5iczTXDKGL7YPy8s+7z+oaM
y3ZD+xRoXu7yQx3e0LjByMzSa6H8fV6Hm1iaLQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
lYf7//ZApDoL3G5HW1Dr8RrUkNmWYpX3zwS60C7H9DKtvl79vWoSyxLwfXQWSYvd4uVftmP0W7sa
4titzx6r1Tmm31s7meBb1NLt7kbrv8+AiVbdpesV8w0Xp4Drm4lvxS8b71fue7nwY0gmec0ecyRg
yAoj2SNbb40qw8KWTnDg7S/NJoANpezC+BUAjpPDKv+jG73uc0x7VXLccLcPWrZZAGhv/dOZvaaG
Vwm0wSmxXtBKrjS10Ec+iQ6pUJ9rnY31EaEqLK1KQpJpD7pHvCm7riNpBcTNTr/bXcTcQYDHAObH
HfCtLegTXA20YySLZUD/eAcQB8y6zRKTFQdlYOHKX5Iny0BoP8sTv9ZBT2ZhofL1u3YDO4C63Bi4
XBU8h/juCP+YZqR7+La6eb4bmsd8Yoam1OQvGFAMPUyclwwlCMtfObvRz0Dp+CwTVyaVkHrK1GwT
tHxGqSQO3qB37Wf7guu0G9mjd/vVGq2DsF7z8QBHE2zB7ibVh03A2ALZN7QsTSzw8F92ogi1eoLv
rg8kOokgAyhvuT9rstZcsOXjM+jA/9F4CzSSLUhYcBt8TygMUla24IGfwoz8GGb7bIWv1X2Vca6J
FjHw5tOxuZIXxvPLfV3VWhq961gFkh+5ZdT+0YRwVb9T2LLxIhaR+7egr3GWT3jetpoCEnh2V7V/
nmqvZzhICfHX8k3J1P1wq7xdTnRiKitg/ACpPgHO/YGH1KfzvNGNaswshXjVcVH1PIwXKiK0D2nx
AcwLKzbHC2Zo2mlpJJ8Vy1akm1GWtxpz8KHw1OmlH03Hrc6wcojCBNCluA2Ga1Emj7D3MfkFqg8+
kP9y51v+Ki6fTCdf/ySsPSbKZxCKJPWR/IUNunGahH7SVLPFr+dBriL8+0ApfYhoKiJyr6LM3Jxn
IyfExjfWWx1FWvT5OwWSrPI3QAYOGK9rmn0ZxY2LvDZelaz+CJ1DNCbzKGVuF0Jhud6nbdSqIL5A
rF6zVcOfFbMiaZieC71tw+aVgJFkeU9vb+YhTekicYfn7z0EvG6LuoNcU+VkY/7ZgcmPoXlhWD7U
POwsPgHAx0myGz/GAaayqMLAxZBJT3Pu04JTKyIG9rjt/EsLEE8H0vicsTplg8RBvg4vXr719v+g
EmORJkTo5Cf+D9FDZ3DYgmO84zQ5yp1X5xHNlSXfB3FNQKnvmChd2161eqgGB4FruexNlOXg0HNM
sMghMQHRS8gZM9epimz8XAM6GIXBDbeNdyVexxl6lOb/zCXeEYLuXioYVsq679Tb/VZRoavSa0JQ
3++B9ReZj9Xsw01B/n1/zb/A2K5d1d/V+kZsujy9mQEyxjTlDxSGvn/UdXmyuVNVzRG+Fv3GANQ6
DPWoNweRAYOYKNsIA2/EbpzykV+A4sugczcisAmLTOXh/dnU2yRGG7gwrCdrEoGZQ0YOQIUeIvkh
s7dbRFDBZXs+8WQVWGPTR/PASNkQEaALtCzyc6oIaMjQToJyib+O5D1vI60TZaBA0zqo67PEct9A
QYSbQWslj3r8ffUIp98uxJ6WqOT3QTcugAahCN3KgKDdHhsd42dr1nZwF/GO7XAK9MXGLhVtzyGg
PvN0va26sT/8JiwGu3504p41YWMRkpUSxu1Bcpy4//Q3LXw9CG6O/7u/9+B2y13PLLRwEPBchUOp
EaGu8+JHooDEVgINnm8NYKoS3J6WM3XawngyP3FdXYgEXbNJ8Ly2p0De5flzbI+Hz4HPJ9/qKzFO
fhBMYhR+s0p5mQeqMzgW31Dhd91dXpe23oW6tgr39LFbJ+FN3/qkP3GP3fiH6yJBkzhzYT2Qxm3H
t2a3fEfXTSDTT5hRKIGLMx3CsfSmPJZ93UuUJuvncP0AtjRtczEpBlC59M0odaG25dClodlG9gzQ
E4OkgZTIhoRCRCW9atUwR+1I+4RnacVK8uLXeeO5dbLZR6eRjtTs4MyfFBLzEXxdXOH6NV1Enrg6
voYZeJNJsayEz+Z78ZFno31gfaOVaE9Vi87OZFVpahZ/LEaIArKPcuowksvc8XYrFVWrGnnILqCC
erfhN5wpfPBKtJhU2ePl7kyT/E2sjaZN0IZh/NButP5NjhfLR6zDAm6Xn4F6i5LtnyJMMwr90kzm
MjSGz0vQMKeLvVauYef8XWMSkiKyraNR9E5Y8AZeiTw32lq1+jom1oizT42QTqAM7QVZWc+pBPB7
NUOBG0+ClFh3fKdDWuTmKuWERALGi6pw3N+aUix6EqwEsOrFRQ0AAVKB51ye/bG8PkQsTYPrg3iU
YVYLnVBJ6KOMpyJXsLTxcOBfVV3cgAT8GkYdAuib4A72QuBRzluuB4Z8jsUnorZk30h8TsoOxDA0
MehgYbzfdKpzNVDpCBxCHpB4H2IPDxXPT66MQMFv3Bvf1pUI6JzS4DLatQG15xyH5zpSmNALVbeu
87WgqqY3joj/xpmf4ZlrF4/nj/5M+6NLoa/YFtJJXcUdll1BtEGQsYTF0GnwHY4spIt7bZzD+KAS
mNhZL3jm5/jsAvMBvb/8SLd73eUM7HJ5twejuNuYCml5rKJD3Mkkg1BBWrrz+u15lPCDqaK4nkLI
I5/7HeK2egwOOJYAuaDCp8aswM5i3yNJ8n4PWu+ZDJchpNm5fwZ+8NPMNMom0/m8sCyFDAV56Um1
1CtynxOrbzBAAVEWwEpHYKsq0UNhZPoeE3eplG4OxFFqIq+62th/QBO/6/tBsMBG4VrCQfuMpXyd
TZqmqQJUXLa4fBYazExTK+FPkvRb1vdRqcw9d8CanbQgQ4TxIJ/Otvv4JwJTPXtiozM3N+BdI6Au
FCG0lttmTmaKYs8VcordPsP0cS97hdmCRTTPpL6y5R1VxthR8BAAosJAEy0BJjmAi7g2Jk9mFl2X
i/p6TxMQfFp8/bR4CSvggaJ+iGwXp3lv0VCLAkFpz4kU9l0pqR29GQSYFNonuz/uj5hT/4pARRpn
Qo4ryrjSpDLHLd9Q9tox9XiHOlF9mmCAIvoeMgrskLWFgifvAf1lGklDrJ2NMb5zwKr/hdSfULWX
RzrRwmqwYqtRBt1Imaa76gJo9DtE0pW1crKcpz329Q02eq18d27AVGADEK0oA7+2+FHlRT1sd0o5
cfDWp2Umrn0d8KyB5KB3Yob9fOBcsOFDnmd8aadhC6zbbiNqGMTLOwCGDBpLHSdUu4QbJmSr0RwH
6uTQajMF8WXdDbBsoFcjHWyO2ufBxqv5HrtmVXem1HLL2CEDMIh8ol/OHFl1BTbF6cv08TDCdW9/
peV/6/kl9SxSrggzslcN8eVDTz6NYfVPNvzXd49JsCEmJtf36yQ964Kq1PYxsXEbqJ4gBcswNuve
BdVtTrUREBora/GeJn68Yh5n+i5ucOsirWip/0vd641rAZo5cd6tLMpOMmyJl2yxom00d4B/cXMn
nLzZ7OYQwsqJW1a29hio0nKh7OkLwQK/R8l4/XvG59kU0QSYPUhbxsec12AxZMj6op0Rff1ayodd
K86BaQWHgFX5Zoqon69Oq/w+tm6EBMKzjjMlrT2v6iVs+0btKQCch5lgyLoxtyxn9RXFhUquXO9C
V7dxSL5617w9Q7coPfwKYD5+R2UbIsskJiLSmdvAfU/7qJRJGCTIM9JRukxFeeO4TtgV2oQiWSIi
JNVNItupSQyqnoos18WccdtHtCE/TRMV7XC1dXNNUofG0V+Vyfb9wlucZNBQyl4vIDTNf/oPNJ2Y
xQsAWORITqjiN70TxuaWcQgzv/9Ol3r2w8P4mop1zDBGV/kwhMzTfV+5dkMjnE0MVLRLigCPky3o
USif1lmQkNRqMmN3OxB9fiILlyvlr+lTVFWuZfWfw9WBvGFdo6U+6j9o+Aaju9cmEPCfmnu6Jba2
ehlzu80zoa87I7q2erz1VeiUz/iPj2ob6KluY7/ZKYIAqRbQ0WlN3eUqkr7EnyOOqBdkr8axDcU0
TZsmMcQulMQB0hf21R6ETiXNDbUiCgwvSqig5tJDqDW6nndPgBXueeIeysHWuRB0GCmkyOwR3eQw
c0cZ+L9fDSnAC7pJxIpSbHOqa/6PB6cYU/3NP4MD/CxUBnS+Cj+H7y2G1vjY1wbnKZ3UNgGi0TAx
fnNHFFLK5SwgOg/6fBWx6pJMSng9JFq/0xoXuX3AoMUSFsyEUQ8mkDViOcW4v655gAvXAlBmFcpl
GxURfIYj4PiQFwol8WhuEBWQA65OVuJzpzC28wNJCv0a0xt8lwZZZDCSwguh4OD1oCOqGdvV+cIk
ydTbWqAVvXX1soLRWAL3NDFyw0wLG9p1Lih6R4wWe+fX3lxO+XVnUP8YxHukHPhS8jLemj8Gg34F
yo52ME92RHBxDt+vNpogpURBBKIST4ynGfhoSew5rmoWsWj0FEiUpFDUuN6PU5t+KS+Kja5Jw/J6
ecYddoWCuOtcdBcQylcFxdtg1QhO3RGXoLvWP4rkYpefq5sItYK6Ys8NVKQXu3xwgupXu9t66e3L
xhytJyo6ucWpyfCcrQJB93kwWqYFnnxXzno8oEKI27MmL/BxZoxQ3lL6G0nFyXHjxN/j/tNHr4xk
RnxXlg4mPsXXP2uuu3kSCYddJj2UCbpO3341d0gcoMTIHVCsrtQ8TY1o4xjPJbx0F1mfBns+6lRt
iPZRt8swxcColHvUSs+xQpV63P/DgiAoJx03kcHkU76U3/3hTdjmOjbwRukWG1+gsT12/PHuwExH
tu1R2TAzx/6ABzZinDqL664z8youoK2CdFIRz7sEckMirQEJOLPeYqnT5+z6XD3mtmxnwA6adBBT
sRhZaV7H/oMeRiI1xYskk8502wAlaeM7gtQBCMBoYjgXt3Zlhs4den3P3Mgb5Kk9Uj550Q89A8ip
k6lcBjatU2sEYJZqPz9WDcsq3fvUYmALjvW7CUQw1Ok2+fep/RnYSHCoxidVlrWYLQ3+BmitK/g6
nKTr+cKsBlQ/4fihGJbkDPPA4uBOBEVWlrxVqGkPoN8b3JnXT1nM6YWO7Qj8u9awWa9SwFzK3IR2
zML+BIopJn8ZIJjUwFqYaaps/9HL8h902JGCR3sPvQQD/fZmHqGg0+64/OoFWmoUFuL4rQxo51Om
fPErc7ptETTP0wnVDirVH/MfHwwG9KSl1z5G+sX3msjbtf0K+dDjHKKvlcJX3CDcxqsl/p3ADTEv
PC9v9gqRsPEJLZ4bCo1gu8AdtCdZ932GMcjYpPFcWObZwHEaa/OZLGrcvDu9JJq9UxUsi4B34O8d
vsek9v0qdzbvtTDhKyPqGm0EVp3KKjD5pvYYswNpHizavdb29rldyIu1dkb8c2jwCqsEULf7fyu+
NUjnK+BydY9f7OJ1znvwNdZud8dyej7TG6uG8USPHf9FBC1GVlS9h9ucY2qee2C2ullMHbmzntjm
TTBWWvLiHZ6/BrS7r7eBApVJSVzrCzngUzgvxCgF69bdio9z3ibcqGosNHzn04hxxjg4EE5bFbI7
YYM1Oy98KF9GooMKm3iFf8pzxTxWa67wigku4y2Inob91CAkzPj34Yuac3ay3dY6Vyp3wzRfpkgG
UorP18gZdpFOIfOlXmGBMB7TrQB6ohRwA/MZIg+PFJRwfFsiQ8RP/jeTS3g+wqjKXm5YipIrGLUD
VjHwOvUqyV2+NLggCuFcWJFkEmX5yjoKcYXInZSVgS2gJO5n4cJrQgOiqDxQC2MDDPHz+fk8r2eS
dnYBwTWeiHjb6MwJgCfK6vIHiVdEgt1e4BFrVIGxrmkjiKPtejKofNgw1YYVauExEyVTjRKl7Llr
OBMmIxRh5j1pE+AQvYc9X7qxdnYasm8hgB5o6lxa3+rZHdwi4Ln4eGjuC3BE40q92RrHM/YJw/+o
bMilY+4WISmHiHDiOuSj2chzN4cYQ4gpVptMzcCyp3ZPS8Y4iE+P6KVwTX9P5C1aTntER0oBMlSO
2G1fcyagHQdQkU8EturUdDBQO/NQlbBIVX4AtOLxz9AsUuTFquQyGTytAY6SDxjahTo1C71s9USt
6F3OGxwO7kPjT7RSEvKCJvFv5qnlIFfEti7c8uPbZdS+ygkt6GR+MpSbHvevc+c/KtuATH3n0FTf
RYKQC+Os+ejlYeKYP+TNsymX9NclL7q9IAe/XloZZdtPCtgQBR1pG5i2SgGkha5IoAiFXOrItNSG
UEZzNRuKcaDk0FG33JkQGjjXLdvnbIVz9TDBnOb1zabpMpRx6QtoQrMSMOxOjoWW/iKq0lxUld7k
iCig4m1VHhiIWcJjib4jx0MRsZsUDd7H3YhIZeGcpB8u3pBqwtd9froQdPg+9yJcuiInnKWqSpU3
RgjzWYRPGjcOJJxuxiURzxssCqdCukZiGuBRzHnNJdRuDG6rxxwNivQiG1r58aehj1pacHi2od3v
kjo5eFNDF7cngygMnoILlcQzqA3fVihB3qjJth3DhYkNwWl1Cc7recQhDOXtQdil3hLIu7MRh02P
6sMcZHznrEU8/YEDlkWT0h9pEUZY7ynbh1wu1bpEvI6zB/fGgzlhLq3LBpylpPcv3uTqz1FE7ror
UNercszmQD5aTsaNKBg+0YHzx6vBPaS3gCE0BafxJ7oXKUwn10jP2yfR5Bp4zu2PgUl14IKhZqDl
1yiVSwl7krn3B1g09YdNzLPVT+zh2A2V9FyrgotXL0vDYOIAJ7CBm/GEmFJVgZp5h2hysHC1AI7a
87Afnof9sZ3hUNiSYsyG1hsAiKrrT3FBICPvlK8+9BflSkrQx7q70fUAC4yUMOJhivEE4DkupS7C
Sdr7rjCE6x/jvfxcOV9mfWLuUX9q90FcsQxVaoroajp1mgnn4+Gpu9TLFWCvvoh9Yi8Juv5ZK0NU
rRuDZ0GxduoYp9kXP2gkitEF8tfhiEZ5qMfQYAtsqBsD3EiOhlVisIda74n2nYoM//DYDBivKxyR
fXX9tI6HlpRqkQKb5f8vcW1JjmGiCd5A88BEKpJyuQnwg0FlAL2H30pzG8T9/ZvBhnyslWb6p+po
OMxGMf0iOMVaBwNxcC7erGJf0mHA/zGgsQd9csOfLD6pZAAB56/IXFOx5LeV9IOZRc0PWyVaMZHN
ef4EWRLbJvVYGdDp3cgm9rongC59U5QOqfnoZdEFf4PX7rNWdLrLoXtT9mjksHhO1ucdnO5uc5C8
3s6Kw9/BDAt9fNN7VkaLVL0A/1+foZYuhK5ts6M1OiUtLaS6LMA1wMMO3sHcsUcw3l69RHPfLGxq
NWQitGSPFJTcnyWDvTGOoDhsI4r4o2591qxfyTzA6GtS/lY9yWGePgJpJ3RspeUOvj7csZcB2H8W
wuHKWekkpivEN8UvwWpXC5GklORLIPWPi9RCdltWSjSgfowBaqNayYVLKGvBp6O7IDn6/ZYzemuq
UB0/J+bO+KBT/8NWEk1hO+eAcu68BCcqqx7tn3mQdyQvULby04cjsg8LbSVuSU826NZeBo0NpxfT
Yno1Z4BXFWqJvEqPUxcjmL4xnqC0o+oDfDlnFvJWh6S2L3U/+7ufgNpy0ktBXdZ7G20aKPSBDgtD
iqLawB83B9DtG1UdUaEzcU+m0gZONetCJ35OjSeyQfn9mZFVky/0mcWjXNzl4vNezD/oDrhtv0F+
twsLoqtdCMM/Ruqm1LMqhqtRMpTezJg8SIwiFup+99um36/RZih1GTtty2pfrEb3tWdKe9s3bS8f
2PLEDiA02xfVLpJowyEhlDUuYB6Ti8os9Lf8ffAUBUEBMQLIjQW9e0RzTbP4d7528ptCgJnkUnpe
DF93o6y68Ks30DDmYlgbcbD+291zUBlhKFGPx+2HrkVA1MrvGHDBvUiVEG1WObyEk4bX7OKrRNYu
vUZVFcAUa5VCtrkODxvWTqmmllilFdhgsRS/Wgp8zVq07G+66aNVUY0QOxrGpYZw/8LA+KvyaLh2
mg59nSVWgPeJgo0fWEMz9bofL/naltdLJTk4DgFKUtBJ4r3FkOD8AZpTWzJC5d49rdPJA45iWvdx
cNhAyfKVzHKaLIgXWvghV5o4cB1LmKB1i+GWhfPpSfp2Oeg7FdkzT6DRiS7XYoVXlAKJ5a1AYeHV
p3sd9fsajpVe8C4OKUbwJ8GGzO/f4z6DJUR7pSILk8k/xyQRuAQ8LnwPJquKBlwF8a6LvpUEvD2u
XtHQiEnSnukwwehM9+6yx9J2xHEQY2Ea6tasLOkRyxAhMIMA9Nj3iA/4mHjFPAlLBhXbN4pCC7Ta
k7DwEiFb16XNPxp0sbll0ImOl1fQz0xAFSuMEqPHL/xTxK9SgUxgkhdoWNx8dOdwGv0GEFp93gHq
sY1ij6CvXxHYL8tjNlWv1+046q1G9cTY6y1RTauP/etKKhQM0PDNSZ/WAbz9gb3jqN+ABdFU2XOu
ozb2LsnhtnAXkMRoiATfg8vsJTkTPXtMj0nWAcBliRyAKQLyJ3C/f8pSl9iL6CKYtfkL22n78GdR
4lebXVZWOqUpOoddFJf//ZrJAkXzkYt6ee+if55QC865h52BOLowgUOdTUxiggsIlc3Zzu9mO3NE
IzsffsCuOlGCtT+0qWF+XTOxhs2BW+zqJcl4zdHc1Wf/Jc//g+6EtwZsQ+h0oc9GhQ9Kg4r3SUok
viWO6SkFAIjaEeNCGaRSDyYrmRk+z6dXRmsa1Dv4uq/6iWdB69MhcvDAI0ZGNF98JW+4KPTQVDly
QZkkpDoANmcaoXvBQL+oPOlXfmwDZ1yqM7zO4yJ5IW+WkHol8YB3zzV7vB9D0hEsQO2pwP6+vmdl
XNlB8+uHj1s9hycvWc2zDW0JaNEDtHiRwZDWU9HCEZf4JBdRDAuVqFWpBvSDx5Fs05wUiOuxt/d1
3caHDeR8zfgTAprxFns+N54H/OykDoje6i9QCkSx0BTYbgFiyCE2yz1kzB0zxmSa3+rFsBZZ7u4V
spRdDKgGjGx7J5O6UPYk3JMS7+Tke0v06qeVvzQbeKdTyvApNbBrCzSecSkKSoM9ZDILxwdNULvp
UsM1djocdkRSs6KV4mAfDSu0TBiGfI27JvDuSX6TfZkZ1n9adh6Myb1H2fSnIBkobZmTNPFzlkFH
GWRf9frc16W/NOWSt2yawCYm53zAIxFtWU08DNmGGXiGZad+LUfhjNzSae9nmA1NJyLj1KNzJcpI
L9cT8uaghuCW7NhbbmXoro/YR3zSFCyAvHE4xPrLwbEIBqA5ejcVQjY5LaSc4XPReRB2ECVRC4JH
2um2cpG1Qj+yKFyobBquGZw19st7ym8VNwTDWO7+jeuC03WHVGaZmsuORMpsqUhcevY4ymfan3Ez
FuYqQHYqiMqIpk9Axf/nPEc/AYqPC/wTRhaIxkESOxT5nYNZQ66NqmNde3QpQ6PPaRtRDsqYL2+n
DvHI99YTq8GrgBkm75Dn+9KGi2ushdVz5EWDcmu76JXX6WBicJghofWkDjO9dsCSVuO5agsoOgdN
6Pokq/UW9cYaUzTwYOs8wWMoHwv8FRD+z/mX7QlKvTfSdh6ELeqizbPfxHBvhT3V3dHpbzeLoxAN
Goo0WEnxxR9tBlTsGnn2mMGlszkwlMCAQ3kmCLsvevHB6Ry4ABc/wkSsPtmXGF7Xe1notkE0eRSd
Fub/TbylbZDCXWEmstGh4SPKUIf37GTa4bbipZeFhI0uRE7UFY70KjbsPagVTODVi5sRUUQG6VlC
/6jrObCf4TerYCL8S6O5KmDWDCG8neYcBZc0kACrH2oXRYWvCupzwekmanThqjBXBvZ3gvre2qRk
098RT6HTSf5a+KIUUCEQlqfOAzaT07a9k6QNX6B3XtMIjQeqmWsqPvyqbpxyF0iD1DD6T7KAxoZh
//V7zn74jY8+xl0W7Ey3+7ATPLYxY0Vj+jHjkbLLMslSAq5efTEXesgYXbef/MKGoLI6YBaZM1oY
J51oPjggx35sxTx5+PUPCKb4GwvnflhvcYDlMnqSHoNFSFJeGwM1D7j6QO/wf8o3Dev/sgWQTS1T
d7RZNWOLGWZowFX6bNCfXtkPNfx8fCqGGMZ6ZyW+/pRML2tkys/i+DMGHmXjoih4KRW3L1Gdbgin
BzdttnjW68I3VE/o19jsnSVTIgrkVVqeiYc8t+RLu5cojKrM83qvQnZDPdQxLuMywzwAy4Io2ceo
5a5/Eu7+4eANjJXogRcshWC3P5qfDi6xEm24fDFQMzEMNhosc+XJHpmeRjem8EohjXBp2iKbksG0
rKlJYyDjOMR+CGFcllyUL1eJ30VFz/GMlsbTXMQFWcgTncgwQa0TDll/d4IsHcYB1AJeDBa9iYQd
ja26ltEzQAq4z1C7YHBeR+YsiMXTPhIrJRQ0oADSJrgXaD09LJxjTn2SuqTD3YS3PiQcGJ8Aqzre
o5kEt5tcSrb4zWHu1LKhhrnCkchtDvvUB1NHDwizeEAiidbFQ88FFmQsYHsxQB6ExHgaO8oRE4F5
dL3zTZRYKrQhNtd3PGynfKSf6GRrCtclUKOEvIbQ90okdH/9F50XPjteduMLKnMubqDixR4LIYk+
JkpASNKnzvkhkGaxUjXAJmalqt4MTUd8G/MNw2ChYTMgKTgaVyfBE3BS28r5HaBK7Wx5M9EbrmGn
8zWkvm/RULpWf7ehuyk+3gyMytmfO6HqxGA8ANb+nRlXWsGtT5MPf1h+mlxEe2t3SlsnSc5ZcRQD
lz7CODwXIiP74U2oQ3pxw+XMA6jaKbx9PZL8o7nzrLJXRexh/dyd+AULD74qCI2kA+m12y5A4RZY
nkLKbiL6pAqgEU2xL/ixtu8TFDZJfQdTmr5EyfEoFZ8Hqa9aZ1XYyDysdOTUmuUhL4dLr+m6To3b
LDE5ZdWtg3PIuE1nhIHyN9Gmzhv63tnR6M9wzA1Zz3/6RIzT6GpU0zwCnS2G6nLEkln41g0WMe3V
WnX5zwuC3pJIjNLa/a+Yszc3IrQwz3Ou/eBpjAZvp5B9KYQJG7a7/DJ9WSM+E5SKXB0j5QpXWNno
GpmaZLGnwU3AzBpMQRDdCYNGebTdfSC78bUYzaw+6TZbEzWVlOH+wFmX771C9ijlHXNlQN/ONdvN
hhTbgH1fXty7PsPnHuTJ0Sp+Re7JwI+rplJRfRnu+QIqx6XKY1AeZyqVguf6C2zH9qfE2fQZwtZ3
fZhxzvPawB+A/Kzc+tLTnDh3P4oRHjX29XVFRBQDMMQC1tKp8gAjhIF4QBg4OKv4gJgaiqDbzEqH
9B6yub8aus23Zn4drl8ouUvhSfRWwc3AuRtI/sQG4fl+LzDMY9NFMlaj1yOFgxo2jSdDo7encB5S
8Dlk34VMJST6TQHuGwcDSeMjme9mAgBU5Ro8H1ZOGCVfsVX+CmkA85LpS0bFBNi6IuC9NCuZqaE1
fSOw/7pjEavTRdWoO3pOjNC1R9HBokrcItxVk7AMpuEh3C9VV5MJM03p+JBz8/viB9RTF5lSHems
GSJIoVCiryVDoLY2osXeSu1uD+PZ3/dWild+h+Nd721/hbFNow9iNywIcGbdr2xYnYf29+HEb+e1
pMHpITVEFlcvOc2pQuTOWbW/tabcBqM56hOqTZI+2IcGFKUZGVuul45p4zmp2ieXWqTitY9ZGe0Z
hZFDJYM1h25C5cscFBBFL3GyzwIG9DHJ0dn+m8vmi5T5tYDUQPPUlp5b1TWz1nogWtDMNBoMxb+k
ayBWjJ9RsBGkk4XGhz0PCKCbVgVn0w9owEiWQS2hb5onPgUrmNJdJ7f7ISj5+a1W4fcIEKNtKinK
uAljzXbojyZTW0PNFXXr9MYThtywWJoOSyqIl5/RDjW2WpkIT8tFSaYufaU9mBG78B5hYa1MCbcT
TE36U66blwy+EbvUsj9xOBKNnPHQ3NxPc2TWr6u+sCg5SNlnt28zl3Xmkbz/bbZzYTHdQEroy4EI
Bs3ZnX0bNOZDYchF3w+yvUTD8qw+nOO5GssYjr2sNzLQtPmvRudOEGOFtzyKG0aAN/rlEz/4T9Em
YMtmiGTR2q4TXGMdrtYs6zzdemQD5+yfMgfBglGl45RYCBQaPEkRH//yzwiSYNCiUlr1aadVAj+A
rOEecnoASGLkiKJQP8YoQp8iwWrGPr6tlo6XiJhgj6U6i4GFsCZar/HcGNfLSV5BwWHqYkNvyxaM
GNZ191dARAhNf+89bdHTL5jrp3dwbjOvnaxWd75IAxwPd//XfzIqqHsectZh4qKndnk7ASMwiJpg
1eWtbzCNNxWxYFFqeM6jbPAEJtWrYlcEyB+FmPg+4AOoR/MUHu1R+iVB8+iWwz+OtrxeUVzbas5A
rTtBA0nfGAkNlV/jpX/hUoYzcOPFjyME2O/JoephGuPNEltKBC0Om4BR3svy/3cR7tWdUgkEK6xR
/+cLGYvQpnBFJYLILgQiLqEYKrlDSV9KWaGcNuKjVL1oHYiF/R1UN/CozxBY2rKaVGDEs9SIQ6Nx
X57BaRu7wpF9kAre6YmeGcDC0anDMBffVox8Eo/Vg9rW1A04iY14KumZmrOmXty/bpajry35UvVN
p09iVqymG451b+/9wJ7cUuw3YiAGFnKJHhYPoa4wvno2S1PyHLNSpCdPhpD+NBI1Zg4fO4P9rf/N
X5crCkhYPM2t6vkT3LYfrwnqiAesMVtBJpEqdnOFHWEoESMUfg5yMLnOVSuqRj2j7Da+MeyStQfg
fKMmaOtjnFw9JhIyumYzi8sehkfTmmZJ3wX9K4fKatMu0y6SE5IXwMqdFVMEzKP5O/SKfdDVvHXX
oysI4ow3D1HvU13wGxA8R9SFsQQemESCY2tcGyOqiKlqwAqJtHr3nDsxeCKL9nW0MBKDZ74EpAc/
X5v5iez3f/lBpDOy0hhz1mirmIDglmLL2nJg3gpVhyMaELL9OV1UUsQyolCJgQm0wQ9mJmp4hnIz
oR3C0BTMHTLjddEuk10klZojj5vQ4d/FDn0pwhrB71/2DFGCGhNb08tbTmIsrvmExdG6aiOT342R
ohYpuymSbDn7CtE5+Eqflz6+b7kHEUPVjJvh2uNRpusP5MBG0CxPGv0rruli/qqE9M5WRvyKymF9
3CQDWKIPegcS/4e8Ag8Z5Z+WF3FzTPeWQyYXaujErDoFWLOkW2Ns9XSS2z35lCifZB+EYHLNj0Pa
l8YIYPj1HCan+ldGT3M/eZQdOZFCnQ75F9P3A3puK0j8n0F3gTBOXSCSkmdH/0mCnYkggr1yKRkX
JAwJZrO2I7bVBn4EEO2+xGcR0PCimMt/z2+Y5tiMZO9fJdJey7Z+SrwOkC8iNsvIVgYg/kGdjgbs
BKAxgm2GfsJiDPzSiBYhIow/BMjZUzcjwfXRC6hA3HSuwa769k6IRbi+Ms6syD4VpaiNbW45C5BX
/qPsxZE5TGiotGDf35j3Cc6P0nAr+L/IiX296kq4YgxBtRqQMlYxo9B9fQ3odSotz7TG9TXe2yom
EDxOaIVIKq0IVXR5tUOsv1QWz4sAmSREnn4o6Oo/Fa75tRcFtlLk848XoWsF3RkOdQ2Pe70vCt/p
FVUmXM7vaVkxPoYLK0ePwHEJN8ldx79mQgMewBCyCmGH/tFQrTNAhYWEeyinhNLykZmgDa9hFLxs
/rHk0gcsCxmeRd99SeFlMZp/TaSqhkHT9O2loCmy5Kci9CrC1hB1v6rkq3BOxeZk9OqV23ORnSYv
DYkCZgN+mE2UNFNYyxy0hpN6A4ESdGfjhWh95huPhVzn8sQrVt8+UX3RDCz/cXzIuT0FcojasZQL
Wb3Gfcy0H1zDbeeRYrL73Uq86H9tIN0pHx7qgJxhsYUbxGgeBLr6SU3sEztpfLi6aAl88DHN3cE2
A/j+fTOHClGpj7KOl3ibsiBH6HsqmyzDRBACeO/t/4FqPEy8NMhtZaveLI5Hys2ZMGA4nyvoJGNN
8jWYN1eyLRwtbvLjfHvXxkHQRyZ1AoZWBv8VirGUChGFKLfwgMil7IX6pDtj1fy3iYhdgsINPV9D
i97F2RdyoM7HhJAKEgDhIOVACh6I78qlYkivqPnZAkYrIZdFNkzn5hwX/A7amTPiIYWH1IwQPdQF
JEXqdb3k5i+pQlijhPgcCIm7Yet6LS1l866V7lYXHod1cPo0Ofrq3hHrz3rLCrPXMyhdK3xSJaWB
VbpqVR9R4H7Ij726hMEOu3aIQC+lwSKKtL4+9Yv4QLYwQf8nqBFlQugc/ZlPxJlFEU2a05rBOeT+
W/6VgUHIgdqza0aKjV2WBGCS++GoPXeui8g9S/pieZGG9ME2OdtL+bRkqqviwVBbLgMltVhUMdCO
8k4norRqTwpTk/2GzZATZy/dpwTgNyoO1+s9rIRHJOcaeM5Ts9dwwruwLuw60tcb0i0f9ixsaAhV
AtU8nFiinCR7EhwJH2275kpJmw4MvAk2kbBuf6bN1j7ghnKBkWev99lO+fztlq6jKrZ0xY0pF0aF
QGxtlDFLCeAkWq+aS3lazT0OEfF3l64O4B6QY1csi4AojOgfAPpPSRkHehpmhj2ZsfQ7irfAMN9y
7nPkOCWOvmpzYG/Vlis9R4T0MPK83NomIALTtaDl53ilMi+Uer+xlXY+qmFJHp6EVyDrVNZCRIrl
kk+ViHO5biq66hVkqyf1r9bo9OJJmWYBRkcGqz5i07iTSWWjzDUj76uj9NzNwDcfmNvARB3VohZy
gkbDoDBLycOHUwUBXMAEph6wFdboJErzejqMJixmjRyVbkPs3QvgcTJIkiQaRaDzs8yPkEKGrtdN
BG7Rd2fo/p5lpWb9gy20pY/xnvxIJ/PjqmJZ7P5OIjVRVNxTK1ELu74hXg+B2rw/w2YaOdGz6Jbb
mY2zoWz8AR9JJv5yKRVQTZS9XsQLeDWoXt9ZhOq8z1QBKCW8/af/lq4+Il0zuwjGrdBflhtm3aTg
g3Qc6OQ5xHCUgsuNZ8QLLLDTmwAhsZM1YHMGnzpXMx/Sj9LKqk4n9kYqwSJLivzUlatlrhKcMYWS
PFG7bx+DTSHH2ArSzgpVUJtfU9AMY7xznsubF2d8+JOzNg9LfxFFFX7qkHmPq/efxbKB4oaciGVK
qDBCxkTDMsdr4a+cMQVW54GPm4Jj+xuPGI8vI2O9XVMIV9hazEYPQe6q8buXj/R9eE0dnKmIlItM
9RGN27l/LRxDjmDJdqrwnzhLikfQT/X0Qxd6kWCXvHxYZMyrnxXEwzXXoO7PV4Qc2oFgvQubyz41
Ep1vHGkvP5+y27QOE3ERF1GlkBuX6fFnGQL8fKu1cqfEVIhlKAhdlRz5gcVtee0ooCZUBe4RPF76
SXIz55z7PPPQpyVitZEF1ezM5qUKqVsRkdJHnVzKMcCMsM9frztl3rtX2Rfq8QJTAipSGQLRsnOw
z808rLaY4n6Ud3oWbVxyzar8h0lifoH4Z/pf7UtaXfauEkJW0EgHfassNzS5/coM0o33zg6NLXIr
3vAAxSQRYvDS/mR7I1dgRBUeWSH4hDPkUUo2pmKb98T9Hn2CO4CkBzOzvb4b+WoBFitdCD4LogZH
dF322LKC817pqCy+/hLM8xpmTwoafNi1WBPs0qrybOFXymyUTEjLWGK/GNN25bMObsfGzhXCXta6
cgyEcu7RGARE/jVub5yyS9DoI0ptvAB/BSF6y4ohrJiTjSmTuvJN6KGX0ric4ydyAPLYmlHH1ANp
8Vtv8gBALplp5uv8UAHzKEl5mIidqCOB/DWEAJWv14MLcvJH19XKAUZu3WoPUT4mNtoprSb4x7CK
AyhomhOOZ5FjWZBqJ83n1PskXLFnPNZdMo8ySCv2os5fp+hJ+6uW0aJt1x6Kp31QxPdR95bg3L9F
35PNNMdaQmdWti+bA2q7GCNrW6JNZG0BdvaReoFLNHRplodlJt6yMtsWSMET1HDpvXad8ufnfkQQ
3SDGZcPNX2J9Xi7mJeWtLUVwvDSjgmePiKVdZ+jxout++TGx5DRbC6dMkga3EMyLqY6KWSjl7Pzx
01FPduffwIT/zms9PcvxuECVhTse5nwpSWKBH0nUW6cEMnw4plloTeXswf6iYEoCPRLfu+581sZU
QAbXw6xuFNilgtBxpKSG0T9BpFUP8ZRljVpLJky9AmCXDKVsQXOECBAXTCpgJU2aHgRlNmQihF8T
UUr65UkGmbuD+mw0atGY5OHfZwc8zmlrKze+o4qDlLGxgh1oyT2Wju+ADQOyx7dZWrLT0NK9nxbF
RpF2oYvdfkjSMEMeHiwVXhaW2Qct0jXOgofK0rxX74mblB62Hmrti4uDd0qV/HFDT2rGhY/lk7fw
O5cAdccdf6d8N4Nh6U4srpuZiDudfnfYB7xnNP7mH9qrDaZGFr8dGQaBxFCJjCmbK0h14PYjAQB7
M1a/wwrqyQNWC4H5+DIFx40uhUZXNN+RFvee27QWJfN63YZGwuvfvi2L7mcQ5Tg4sL1vCIbTobNw
FMxr5cVwSLT79clBmKg954ThGkXd9S5qurhRZx8svgCqExNTeZkMKEJaY6CGjyOcGn6s6NOVmYW1
s6eqZ5MhCfaKGstKN0G1xXKnXX+aG468FTP3q+evjB8LFQskzniL2UctzJ53wDouwaiMwXO4QX4F
BSCpdEXtHzoaRdTDoQwK9Kjti+jMv5wALibwzz3ckmvSHi6ATxTwl+pFDS62DYFSc8R+NgBzdgek
gRKNyFcGohryPG5Gh53mYU7ISoUpHKrZO2sDSyhv4fzqMfoHzravQ6w30evSeZDF2uzLYRiWBS7E
b3YVHkf38H+Zx3Sle9LL/DiIQiYrwCmvqwcztcVLnZ4xzmzDEiReg0MF638fo7HHWnpQbL1dgMz3
zhUhMJDanrfAEMcmffi1NNpsya4vnX2SdE1V6HZ64OcxEI4YSONk7HbCn6yvviisPkWNZCUt34V5
74Na94mq16iEumEUwlAYuozZuhnJni1gnh5FTu7A0/UbWLPrgqyfBkLX3L7l0SGNA1q7sEcOHurT
O/KDOwk0tF4VXxIKPxLDVM8GdgmNzQEkNznxeavUtMJV45oNWHGz61OCMHKV4oEFndxvt90/tSZh
DIbj4Ndi+LJyfgK1y54+LHUdS3ox+lVZn3CimYjhlm5N5SplVhzL0CV2Ec59tITW9l+qN7OyNTeN
zXirXiW3AUKRxvU7YzAgzSAvZlkTntcp53SQelkgEECuNhdh70cUslCO6UyvM4ywZP2HCvSXJMtN
/kHI03wTBoNGS0RHpxalYbt0reZDAqUz7JI3ZhlTPyK2dVc8GbIl+TkjNUWHLUuHrqdivMXkEHMG
smNStRdySYUiCPVoQRy/zixRjAQLqp2Pp7OqQUxW2CKwf9vOt7QQMlONGa3NnBTf7V6EiaUxKOZD
x7/4eDZ7KMMVWIuiQpfHz2u/py5xKMQmv6Y30k2EPRMcXOkkqh6qTWNhhTaRtvCzuKREROivO+01
f9GgMR60YnA1ZcVjXPBhKVTgtZfPuIFI1RSPc0wnVyT2yx4MXsIFWAnFd9Mp0sL6WsGndzGKM7cp
0gfloBzgLptZZw3L+twyNGlW7EmtvmOg4b1ImU9zt5+Fa9P7jiQmWqVyxdf5mkCJpyULECEqMjnj
h/QXXS1GdYkYxKsbAOmSLOIU6pO+jiS0A8SiHjA+DJozHx2v2ybo3WgXlfeGaA56nQDNRpRwEV/O
QSy5MPHy6+WYRe07OQMwQB+QNhh+z2ej8ZZhR0iNRX8uJv2fjvIv/Tkh2H+wiO4His1k5wum51XA
lJnPadDI1a0TTWTYhP1VS5DQ51Rk7KFHrvnxtqnTBiV+HSu8f6eA1lUAY+Sh/P9O8SKIi7urTh9k
LgfYV3I2BPdh5uLn2Sb8DzK5bUUWeGqEyEn5bgwtR/6dDlJpEZFespu54dMyfKyCOuft8FmfN+m1
ABMF9QiHhFLIecsGjYw85M8qhLZczIhKkSxJaIEZZh7zI10Ey/tNPxv2uLzrdHiP6ZRo+HQL/2mq
UPL+3Q+cJ6xS+uPwARd14rk8LPY1pwPOPp94TYo+gXyaXYgM0LNtRpOwQm4LTu9epd+TuEAffrfO
SXc9nJeGYDobsA7UfaoKGxBBFRWdR6XmBJpg5aMxReW6I/HZgm+qe7K2aeOoJavrT/8AqzMwQvrK
WJ5DUWlaXQQiIjk1YK211PP/bCr+++9lLbubBSnAtcOh0mzouor89Xnfc+beGOVpZOrp3Jr+m0MH
D04GHJmz8IJtqevOzktFGHLTVrpDNcHqdhpMj1mLth4/jYRVTepBuRNnX7TxkqF1Wgd0pCHoaTsy
I2jSWQMNV4J2XN2xDYnEt2lqX2ugIfJxiRb9jtDU5gaqN06/lH4TUbtFmkpU7kEkzlxFDODkbtLq
wh973yS0qulomtwo66jXhvKE2Mk91lIMKx1KLeZQzZtM/14eH6HDKVsQkuBTHwKlJ2vU93vTpgjf
CEAG8M6WFDh9mYs+VEq4qTUoYiOMEXlP8+y/JTXjt4AJhYyK2WMe8IriegQaLB5g7YDjVsBUzcQB
eaFbAZyl4NwcuB3qJ+GjZh5zW1sFY6bUUmX/esyZ6GcyhFlg2O4CUDo6lZx47YnSG/vcNtJZQHOJ
5wgHVRm7naGE3fLaAC/+OwCw2jh4oyw31pnAKdzUzAsJpTsCoLwb+JMUwyGjX8lFtPN2SJKqZL6A
GwJWc3u2JRCa358X0MNFQSQFwYdwYvajhdAS0Co0MsHXehaMdtGUgM5whFs7kvpZQj0e4N2GjWAX
hCecenhfDXQPamPDQElQw5lnHQshtda9kUmB67nIp2OvH7fNf7B+EjN+RnukKdvzRUTs1LSj3zJ8
QpgBX4WEY4DllQFsRpZqBQe1S/e6uZMRDC+6+K3fm0riPa93Xd9cS6+uitkfSK2CWlRiUKORP4IJ
LQEHfAcrrXTox9KNuQaPYMaUHTlu3tFQBkEZkMyWCKIGAl5a6OMFxjBIclRBn31ipHPOyRBCGQoY
6urxGhq8lxYWqSbl+DmJ6hj51g83dQJGF4IoZgP2COOTMQsne0OvfMV8Zc8ghj78akKtIRApqYCU
+WLYxOQTL4nY6Bc4GHQ4EXv4GsRnhuI4Ge94ZRuPI2kz2WlV8QDpd23qVwYzTqjNXkfIdq4qfxHO
yRr9he9clOaaxSBMDQ2mewWHwo8+7VhmHlqt6otv9WiuWuHKEb7pUcjxJZ5oyNie89ZDz6npmffh
EJO52tuq/Y8yCQMotHXHhUTE7XiFZQW/iODnFtnYD0keIhOv46oSOvXA9A8HgkDs5eQsJl6Dc2s6
w67ZrrxbGBPwA1hyCgLUbEYlZkmfBwccM37+uvDE25j0Q00GJkZDkzBqHDWl60kbtWaveQ5SH5wA
N13NCSXHPsHT8Np6CN1Jajjg3A3kdcWnxGe3U2rRZJ9BuT7CZ3+ADi3biOIlIAR5E/gC67ZIorS5
k9GDH4KTWLr+CEeE5qAa5lw0a/bHWe3wOHxrlUgbPoHBeOo2VtFlvVw2Np/wDDqAtldXYcGgC9xM
Ai8KeFt1RGGk6pGrRYTxekRfqR0eLO0qGuYNN9UeJS0ZFWgwhDl6qquugKqs7qk/NwHcMu+ZXQj2
k7JkpVgzKTqUF7x0IqM5X8Y6/SVur7LHIZbht0tQ/qgXtNE4ApJ0FS284q3DvsW4DEB1C6fJ2I5Y
SPf4q9YkZaE9T0orHnsSziYG6tHiGf7KHe+2Qe//f38dfsKGeNhvNPFZY3PbWOHikrRm8NGwQL+1
70jaGYKgG0XwFg3Df2SmRAL1Atl5Ma2tkHhgBVx71tLzB1vvpcXYDoFXxKVvlAjc0dDlkkz6miDe
Lvs2j6mbOpx5OBuSTYIybbuNdslxSX+1zVcFO4uWcX7LQnkuupLLG8D+nWnbTYtrHCX3775OH6Mk
HPctw/TtXD5GUyjxDMfSAOfuuFa3TZGdokNwAY97bMR4vCA0tHIM4NiSxnp6gX4NHoFdplH43Kp0
Hq5akSfXMMl9FdJA1vDd2VsKh5v6Gu6KGdzvwzPHLdOKbxKETQEulnSImzHE8Pkow1gjuq3Dg9wE
LBDeJDU7YYmIOx3lA4sRmJYP1nQS6AIXD+1b2s/Fusus/RP7VpLK5G6sYrD0YCswQAJMdYNb3HIs
W9c2TjrVysqdnhqpa6B7xVNEhQQwPB+s13yKHeY0FGHC7dtDjTpCK8dOy4hocSer5JvBryg13fQ9
GtoeUQdhQfeuqGDpSBhnckeU6t4DDEIlowS0v/6Anu+9RdRuSH8Zb29rVljePmHq4z8A6r2TdJ3g
vRfv60LZSpq3g2DRAluT814dNpZAVa/BHTQU8wBgCXKieA47JKxQQREDa79JyMsasi6tU1gWO7Me
nMiuTUcCc2z+2VDkSqdE0U1Gta8UG8pfcjzXwUyE9d4vTwQDm5gsB06BGPmpDHemX8rdta+XG0K6
fAdVmT2Ego/lkvJQom4LIVCVQR/ztoc0Kh/Jzbmlygb2GvaZYU3N7+y9M8a7uwA5q0NvoInyXlbP
ziCRrgCpZg3fDsUAf56wXSf9ldYBlpGpPs8nyG5s1eCas3yaTf9R+gWwOQYn6QKPc16YP5z2J361
mXC3IcSwq/RZBmIAu980KRf4Vs2Y0ngQWNEDpxKAeTgHv3dq21uYpcUSUOagFfuQvm2nw+Y8dB0p
oY03TJo89SNor9MVqp+uV48a417wDYA13zBiaeBVCn9t4dlh1TMC00jfmFzx7NTJRkKEJ/Ymqla/
09c8JqSgiaRLOehXbkpI9BpeYC2MprzbhLzBza/y00zPpRXlZzRKDbIjgJZiCifnxxPV/5mB0CVF
Ux4a3ySlOGQfBK/mRBlxGF+azmmmgaRL6uXHqvpXGolIyRku4BIlY0qtZgRAs4QbUBDhPe2CUxIS
51XI3azjJ+45PuSHoeah6tc9JlxXgg9eCPmjBSJU0olw4cHoh2AwQ2tnqXgMzu4WHird++ytnplf
eB/rQTfOO7oV4//dN33PBPxIzpzfW5XuQebWMNE3+YLlBS850/3gdSgJigw18kULhrD3Obe57NAi
C6XC3G5yFZxTIq0Xcf8vVmHtVXReblHTassEBbDbsqVqsjEWf7el24SPHEc0gHbek70QEzgxaO3W
/6+vj7RMrvC0D4Z/qQRU3tcgQe1YP0A7hXk4MKuqTz1A0P+rc0OHfP1LnBLyTBYcT/ze24GqrT8Q
1A6CVAItTDBE6Z8xLlhJelpEyW9YTgkHQ69la3ua02wHXdAePJ5ruRyCnLGSc9M2tQK6jhSshcNJ
mb/y+nzUyRUQ41jYvTiAxno0uYidTA+gVp9VqGWUxoWTOnF3VgDVCYIo+QKMQ+Gl0DfK7LvMcQHx
C2Tv367cEB/SJK8l1wtquFGLtrh98t87OUo9+GTY+s3FWpZNfZlJcYHheopJvU4aaQijdhx6mtVL
CjMtFO25YVBbNnrWN7aDi2oe0nw0YOAlcfsGPEnQBBufh7UiTrFraxjNihU5dSiKpWzhSYUblJs9
qoK+/OIHtzb1PXQ4QvbnPHfdm3XfXuzJ/qxe2jZUvmp/lrhCH40B0K0vAQvs6DYsEsqgM+mLxcLT
5NybzRVCAUGp0yMQqO/SpE8B1dTPnEW2av4Uvb3F3XDXhWqlvC/7UeAjdL9kNuJqsKL/FP41FGAG
LjaMrKDDucAkhMo6s1h3QC5vdFfl++MXLhe7oqaQA1hiW9ET94G/7GJoPUuXDhYJdsWcNdRQPCrc
9eVOCFNIoKNme8f6ybX+MlOltEPwkfRiFML0APOaEwLsOsiq7PmIsDklYGDqd6RTRfl4IKwpoyvf
TxW2E8wRK8GLvNF48yPlVg0uEtgxvByjrsmjjBFI4Km95nkwhZqAl1BhL6x6KsX+cJJQAn7jwS4Z
iy7A0sP020lB/h189iBXtGFddiCffF5ndMyD+Kynvf3sWYJCatcHT08HYE5y0jQ2K1rZncbFXs5A
rnVCsCTd+ZHRP2gfA+rcG3YeATGzHYDVs2+KrVhI+EPv77N3PE9arvwxhnoiucY3sB5iopky+xpd
xR/fCt1hIxfbMHb4Xrq3mK7Nq4VGZoNJU/ROCnWvv/xrR++NBkq0v+0WWVnDL1ilrbM6EDdCGiwV
jeAg+3MPrRihG/ReHHpSIvs7hCk6drM4X1+7ghiySiZ9b4WQK49+bVQaNbIVOjCgWDbYccd6V7Rq
dbOqVKhFFG3bcwN3Ren9QlIf/4AGULi/7GDefHvdZyxq8em12mi/3+0EUuebtJHk5/b++In0v5yd
AjYPX3Cn1l/NAL1ETs9C1EcogVcUQTZaZRtF5kP/TeBoLlJkA5G4WAk3S3CUnnKdYnaGBMkdfT2T
esXRatAUFbN3qkywu7ZOCYYkbTZ0W8FuobjHMkj/YdVDG7KUC6AyWBZdphQWvzvcp+cSmZjCoATB
8U0pJckRliDyoI+CKqDUjCXWeBgYqNTNyjhFCJxAX5nAEyjesk9ZF62kTFxj359DP2oe2sAeXEM0
IAPbtxPSxqID3IqtgK1lG6/RIMBIkAMSTZ5vnSaEp+Xoxcz5RFMeefqumrYBmW9HD4y7aqEYkn38
enSLXSjHceuuWxBjycE94CWSS1ZRrfsO818+PGp55Ygr4fWDpgsFhYnx6vBk5mo+lJIbBKyz50k/
IVF1MzwM1sMdJEi/l0NljSwFbxEhHBealAfzp0c8tB7FcFESDnYbxZAPVcKRinDQbFT9rArXpJ1p
RuzCoX9HJb45yHEVIN5xf1GpV3mc69aDmIOD+hIRJPhzUYwFT010wFfvykzEnhNbTIZMhVWcuCHq
Zh/p1ooUseVoeFsDDdE7EazoFHEgaaN0MEOhcTpeVuWWyKX5pTFp56sWDTaEUgNkphietK1zH7xY
Egqege4ZIVU+NM2BMnvgWNtwH5L8qN3TVcwrymfw2juOr4qT9/Ti6OolUisWhYEmILxp0mdyHw1i
4k1SV1YHSga2ZPf4QPwov4refTOwBvbE8e2F4cUqBAZjWq62k5arE4nWh9dmJeC/cMPvBFaNkFuD
XnUIfLP7M95DEflYQp2z7/ylJxnE7EjggSZEHMVCO3b0tWwU2xkyDaSmCDKCPo+ruL5/rw016rQy
bywgESSJft0ou90InnpbX6/tWzLD4jnChrE6aXIi/ntVauYSUdTb1wy+Z5PohUNdtXxIPHkGYRns
nLOoyrBbtrn+tki73VGrEARlL/5FfdSynI+GqgEQwYWg5X+1Fdqt0SqoItZNZsJYAlW2+bJUNzxS
XpcNkGbKBUbW4WTbgfcrPqm5f6qwdXVEEf79p8/Yss4PxoTgDRXQcFxlU06EDOH8VBTqG6un84KT
t/i0Hu/V0uJ0b435WToQIGZrRjROdogoCrm8I9eFC6bR8j1Szn1RHhSDFwpv12u8wNsr48AhfeX6
GHhFgVFeyiBEiKNXcm2WD9xhKNOc3rHvOSwuyXOavkPI4BbIk9inW14PyaWzTmGW3jtX4O7uoHjJ
6pWH3pxEPzZAx55dKdWGU6gi5lPPDu+alMLE+a3hODss3xzqd3TNqXV10r7JiZ52fNNy8spiBhkj
pgTSqm+JimBydDEMl+in/M/AZDxfKHZNRTWxoPjBR+css/12MShx9qi6uQezGJUYCQx8txo3SVcZ
ujbSxrWuBFeh4XOIpvLpz4FCCpqI9+4/l3K5A5WinL1KKakfzNBsrcUZNQnl+FVkJBB/qDGdP6vd
ph3OYXbHgcth8azImo6AjpLaHEj6BVlC3FX7crkBEGiiAvzoeSEYQiVPPmYg700ZKJdb4nN8Ad2T
Hu2GgJdyiy02oIEKL5goigTGnfqJhtVhu45kY4YYivowTp5Vp8KaqJ/XKrBNPZr76w6sx0sK1b35
kMg8M/H7GGLQr4s5KB7uyhw1RntPBZz5a+KNo6AtNMVa3ZYsgyDpBN2bDPQ3dUsTvg0XKSPjp2Cy
5TLCq/VfiUqQbKQ3c/b429wyjkJ3fsexQGCzNq+c0xJV8l1lbrksWjOxdbwMvfDQf4bngKv6JsyI
ft10b8MP+O1Ha18t0P4yN+eXLUVWZT0NAvPfQOBA6XnSnEkbi31mOPpTrE8WmrfLQFWpNoPbNl3O
xtGhnXbWg6+vj9iM8S6WRHK73t9oOiPTQa+dXQiswpcfuNJyIohiBdln/fUOFS0YDtaygzbHMbMD
gFOdx9yfym+m0Mfnh0hOTinZY4XYU6VpBoBZ+PRoSLKLaBSG8QtAPqZas/q/XKKgsHHYFQ2MY5Yt
iIFHJD0HleSSVOXs8NyyvO0PQFCSvMlmXSbQX4b0k63w4ZFOl4KQNR7TuHYPKydZOHIhEFLWh2Yw
zvC5gRJBU2TLjgx4sehlRtNj+E6yCnuLuqCHJdqhzOrvc46jDK88YF4ery4c9C0mGLqZwU1wugR6
lC+vJplieXaPZczXfegr1wQUJJo1P3517JIkMnvhFlu0as0CQFvz4Ai64dh9EUWWtkJZdkci3QLQ
9hMEpt8sYe1wdu7WQArlv0SPrM2ZF7WXM300Gn5b8v+bqy4z6nu7AgrfG9oaJ6WsUqxs32jdTst7
ofeCe86ZL0WqGwsCm72M8TI2gUbD+D56D+AM1Xl/qtncLhui7MjSCh8GxjvHbdKTw3TFqeQfPOfZ
RlzxdO4yU2IVPRVK0Xk+H6N+7+bZmKrRXblrWkLkEbpGdl8ZXLCi3JCSZK0GIxDJ+Z+ZxkdY3gDh
OQBmUfvm7XOrwWligmOLczVi3qOC98k20GwTrRdUjeLelotDV3faV2ZDOhOx4O4jnQy79yhJ7o+Z
/dnZ4apaTiKmHHU0i6c9nKL/98iWON+vzAfmI3BhqLfxbPf8jqxcskm6tBMNjbP3gLHkZhz18NAg
c36FigevK3LKQgAThmOHvvswn/b6WTbfE008MANOqPCSp5gc+k3UzF+gMp1SXdZvtBqZQ2c+T1iG
QEGS1f7FO5ZEPt1akpoEhwnm+PlUU8qA1NlEAPJQn3rPSexLJQF1uz+V44a5PZMd43lRZ6+uxP3e
hqWCDcvd8ryWIILrlpA25b0V+LNft9V5AALSpr6Uq2VUDaXrn7mTezyP04gVoSh5QEQeXFuA1QTd
YRywUMKmdGEA1RQEYrBeUS6e4exnfHVl7OKa5yGwRMFi3wGemFtgWfRi4ppIW7H9sc3UvG8B+4j5
60xrc9VRw9cR+eImZeBZLqM7pnZ0qoJ07YpcLgDCx2rKhEtjdC9wcsuzv+61PYKvxRs9BzXXnHBx
BPmENcqrxVwhGFqt/5qua6IgQNaokHWtj15rdbfi/mtdbpgDtxLOFWVWiKebdIZkwpPg+ipxOh80
bFkzes2zdXQe/ihU3qMNCKPZz+e4drfMUY7nXyTMWfOB3+6mZb1TCUCHOvF8Pj8Fn7hg9IZ6YBTH
E3O8qvN0k7jrSkvX9z3RJ5zdg5TrQvuNdpKVBco1+k1spcjGKr3ETgdXsSa1QYR3ObXE5Z8T6ggV
vaeUCqB0jMB7JipwJGiFBSuRlDbVenNu45G0Syh32sbjxC8ZEunmyoDOJl+Oy32zQDj7HESoRQo0
AxALLN7L/qUP+euzCE/+DNW9xYtAyi82YDojalKhXVfp/hbrDoZhAx0e+mDAb2cQXKYMp6mITBFi
AxUbE24l+EFhc6r3Wl/UmvtiUF/JrXt99iDl21k5E+p8a5AudaZ9SeVAWWrfHV9+UnViroOhvymT
2760Po7qUJrl+6tDtgO4wXvkTW5dyo5OvLr/oepJIYiHGHHJNNVeHhVe0eBsMp2zGwQTxPaBx4DA
Hpq6LRg0aCTPpCgRLxKZelJbNe9+zTcG0GZHuX9Xm2ToNsL+iST+bM8aBCCG7nNjBDcXAdYCr7Z/
RWPU7vLamlZAcIvi0jjPc9CmMROyyNzt60gZxCR/bP8QcxfLhnDIxw/h3EMIaFMSAzuvePDNZroh
CS2T7gSJCLFWTDZGmGZJPxriPM/dGs8/asD5UzE7r+ORmEXFwlRkoLPVL5BWZtKIDtrIsbj0KYne
HZfXQTnYwFTcKXm+SF1d44Uy3mhLb63D8iOwEAfGK9ZgBmFlrC1IhVOVo3tS0nE/idsPwWI9UJvg
MNm98Vc/lC+Rm84dtvubWSJ1wQ/QSeKqhLFRmLm2A3amAJsfkNQ7OwY9kY4HmIuZIWikAmZHoRZJ
Sc1u6kP11edyhkboh2NLLwvn7LG04L154V6ehAeeBQSNYtS4nvZ3REcaxMRnnbtXpGcV9ZWZy+Eo
KHAcqx50menckP+/05W7qqOBxvRfI6fLCjdPPAgUY3khhVlcztYadUpuWBSEEaaiafCjV454nHbK
newqQBJawIg91KC1PvuEjJwsOv/gSDXL8abI1u9mZKKBsXtCWjgzjqVa/xPSujJ+QUOXPMXx4oTk
QJPXip0ISlkJhCOiDZ174ZIM1kpdYAZU9091o9IDPtpUQKbYYD15GzNIhpP1047KV4EkMnwSmPAa
PhRVxgSOfkFMOoBjLZdhwC9j/IdUabxXEpZweZUEvRvclaLBwfTNOVi+FxD83jnoj4TnyzGR5rys
t0iidZ3iHfz21jGCoacrkMvsQliQd1UZvW0yRzp4ocsWF7ohC5g7VEzh2YTRrCGZLxk71DGGsW0A
FdvryNqxbTBc1BFLP6xWOt/juhYbp0ORu6Y/oo93nnzRglhRXhQZnVTC2wTqPOAIbC1Twn75RLRG
/8NnKWQCsUl50K1xR2lkoqCxunZzP4v2cVbvpCyR9fl4vdyQXpTyuwBzqo0tFzUl8GcgKwsfVCgZ
0bhOPLgrvNIPP20of+/PNwOXAcqlekzO2PObDOrAn23gY7MituhrPmwu+MsyLUshUR5WO593rjk7
J1eDGbh8sy5oC/dQpxYsAGqUMd5xvD6SDZX0S0O2BiwkaxrNv0LxDuGavBlk9UIZBOPThv1YoHt0
nGrZmaur3ucBc96AD0s5Tnra1hy0bWL+F/eQ82jMid7Za+DXKAEtt+x4FbEaxjrTorUPjPe9ZmKN
yeRrJvjzeGKwjitnc+RscgJ4qj7i+GNUWrCVnY9rBcX5uXKNCHT83R8cX42Krs3um/nG9sZSwY7V
uGbJZvTy91ngIgrW+xJI85w18ZEG4egE8HdXQEuV322bPwjWHJxSOy73agkqxG/wc4XzHeWF7s1F
JqSE0CWyxe+1M4gP8ni8FK7mW2nJrNFtXRYr3Di14giHLhYFRylXrhgJQLYf4P/n/e/8ka1ZKoqw
SOXEgMMQjZ3B5CnUTkngtmNwcxNdX6cU15M5r5iqmprRcl86hh01YBawI2JH+kjPh/b1LNNvhb3w
GFIkPmlmkpaMmQbTuJk//0obiW1Lb2Vv7L2cirrAHLx7i37+h6DLjspqndcl0pUkrrOZxf32DBJk
cZllW0eCeq8zuQyAmTZ7TwhfxikqXTGxrm7r1br/lPWHxXAKOFByKga5Kh21viTbuOv9Of6CgXMJ
Ek0vnUaShtvS7pDAQs1Jy25QC1eog1Ib2VNOInCaX0eK8Z6aMqf7xmnRnXfxRxh6IGIpqqCu27mU
5uHShjM3TtgO3YSb/z7bUIzH/bEKH+0c1qgBWRMNbkZqTJrKT1BcbJrcequuDceN8WjthhEpEPyO
79uwmCLIHcls7VBhie+phoExcZqbz5fOzDiWqpAx82k4h/s2vfIbjXVn7gkVHw1GUm8aea+cLZA+
iRPyWQKua6daWvvvifDpdrg0yXc4EI+ChtCAv37RvF8gVAGs0aPDSUxovyY4Zqiq+A9ZBCF8yrsm
oHt9UpFZFS3at/RR3aRF0qLWbYqOLckpBy74+lm0X64LtiNiZPAPnzU00YT9hEy96suDiZZ7umAj
Le1h4DI2T0MXgWWjBuTpUTWKWcVq+yNqgsoe2+YQuBhkAP3xuG3KWaw0bzjunOSj5ssUAp25zgym
JDfQFLiMlFXHiVqiABB3dilJ6D3uEi9vPlEPnLS7COAoQiuLpL917byptn7e5kPfVmK1Qjbx90UG
QxgLbJsWzZ/IJ20ufB/vZ7GOijISbexa0WQTdGMKX1FerjKIZNSaS11hCw9KfOOgGgxse6hLR40T
uA8+bczCR9t1iU0acUZsHSk51LLa1IyCO3VzVwqLRkgEJVaca5DPU5Ixm74PIWRILRsNvAturB6F
8mwn+r7IL9qT5fPiw2TmLfiBqZvLftmpcur7FiH10ClNGVzXQAvah9d3jsNYhqXMddW3ZW5D8yTc
+lsRo8/2jmWjb4tEy8VQLqD2feoUHhwfSe80utpSxM/c/z/vh+vScGy5oGlCgsfy8/t6AOMSXfPW
+im76TvZU4zBlAkL2RyyOw6NcFE0PkA8v1+/JUmy/w+ZOYKYe+b3CbhSO6xOrO5oT39HE90H4q9T
S3+4W8hNidtP847Ms9qZmNAcoYPEKp2vuHvAikvdqIckOaq2Eb4Lo+sIIQpK789TOVesu24wYjMg
EKSG7z0/vju7kSof40NRHRh4hfioU+2yHkV2bO4pP9OUri3erenlOlUF2UZjdp+78A0quZJqnvlk
RETOmrIYNVNs86zT8a2mCQL/i5NGLILVJYyhMFcgR1ziou83rykmOXHd8HE49vuEO5vswtN5a1Hi
CE2s94miyRG4eAzSVA5PNWwS0MS3lOP3NDJYamGmfXYNW5AsQ+g7YPNobykRKr+6xx05nYlSs7qk
7XNzIQvL7nj3fnowwAudYDGgdmfhpTcm4VmRfTS138kgRyQLbzB5cK+MIpB3I3tRcWnrW2CRYZmm
iBMmwS5Qk3PHbfwYK+1kO8xs8n6/NXNLxz8L0ZsZB2dIXQIKRK/Rxmx/VwQfGDl0Q6Y+WLFfy0Oe
oTsdnUoWIgHnMGomIGnjt+fYKmrgg7bx1q1mQatLK9M4kKmFxzSOt/0ZWhnCp6Accs/BQTDDlDQ7
Vqnh3qv/GrtMZJeqKH1dY4z5GKFnYABGioHTtH/86qAbreavhuVMuUEcD3M2jbPtc+QDiZIXg+9s
6cOXMY2Qi/ugnd6F2E/qpzHvNp3MKU2JO6106rR4BJYYP1xCEXggBj6wjbhnYE43DFplNsr+0Yo1
VIR2cdIUzGRnBd6uV/8QbyrzQj03QucJP6iRaiy4TEeyjwHC6YuwwDleJnSKiAuO/bxKP7FoBWwS
M7lXRJbi/J1kNwFBWVAp5+t+5cM3+A6S4hsacdyvurZE0UjgKDeZV4zZz4egHFsyf8NFGSiZ3FKu
Qe1uHX9hi/8gp96ZCoUuTh2ofpxoyzR+6AT6NuScaRDA4ICpoAt6LS3sSFHFAOHr8pHbxDUfH1Bd
OXp6YYR6GvwmLp1yz0fMNwqY7ofpf37e4QWYhuqYrEW6Fk2ml414jQIHR7juB5ri4RzM1kNVftWz
1DnDxsemn6jYfY2O+OCE7ZGTOTH52yJZJCqtecQGiFPfekoj5e/WIjtjbaNLgmq92BpaFHDbqUZN
0Ams0XjyqtLCyDapijmpBBCHV1x55uNJAkdYpbF5na6CwvzCj4+MtWZxfokeLREhBR84QmSpQ0rY
dBq2ng91q5I3pmA+GApQzATXwoDU56PAKUtaCGRssHk+Ky936ulwzBNF+qGlZnNQlRjr+im2/dyF
jGEMutGXu7IbD37nHQUCTSd6lOtbv5Sr2d86qT+nLmP/ND1OIYf/aNCC1NYpAwK0EsInAHDEAI0k
7jTBBqBSLuCKoUvSt3fHYhAO0VD/EZDIRCXRnKVYqEc//8kFzk+C2n4aaqpZ4iuddOWRuWz5KEei
dm0b/GAkLCF5afr2dVeoqC84S3qZY+YsS/SjORKmwZqQ8cGz7ryzDWObBuLLas6uPgYQ9BU29Ppr
FIY4NO3z0l02fMvnntfSh/Q+/jk9XWAwv+jEBQ+8yaKfk4eaHehFKOT/TjhydMNdaGGG+FwPJ2Tg
SS8lxXate7LWsFhkTCTFaf+fgxAdv2iqxcetLJ5ndy6VgQaZBaGIlGl5BhJM3h2VK9dbxKU+vLtA
qpUczMIHYJoi22OedoVowjXfcTeSzgupSIDWP7TWYEDW8ALZdONPBVzQ70wtf2tvgypqMB2XRUsw
kTTqn5sFIA9sIx1pEGNEvaDt+N26V7BHuApFoPK9mgw8B7K8fWqbCTzQUtxNhAoIXETp6pBIjram
1jDoLIuLm0uZz5aC2PgQsVSWB0VSyUhpMRXrIHjtyskOo7Q0zp3Ob6pU0tiVW02STQBlGeUbEIkM
ZU+VH1vyhvw5l9BUP3BnGKYcmkNEluliOcQdwqfvIzXPVHUy+CnShFNcKLUDUdOiiAZFY7adrnyR
jcqIabQsLML9nQ6XsZGdktUGirLjnJkoxJYPIm1M5r+3yx9hcQUVybEhuHeD0TLqFEcVUfr1WMFg
IspDADGPWXEAEsXFaLc0ZCxZQZK1PWwA8iPBxwrNAvi9olyuhqyMn2dCOsqJU5vE5t6Ss4bXxw83
odknIePA+fhpOeuDRRN2UUV0pDq8MHJ0BHYb/SoSzcNZkIZ8sMOubru2hzRKT+OhbjSPGYvg9S6a
lcVofniqJuvX8XLbeydUUkX4Wpg2gfwsxtGB9lVAJCCp1mlcURxv91AHhjP3Mqgn9zj4fT0fDMJy
81mZHPzD77qm2rHcf5S3lWiHN571v0IRAkoV7Drm3z5XrBvhEj/LtNyZPHK0GkzGbqMOZx3DDe1W
MsjYx4MLyP/xEZzytomCYviJBst7XAC4Ll5wXiHg37CGox4t/kTiKUzRsLUULIDV9miDyiAvS0ZJ
497DywME7j93VNI6Ocg2n7RxhQTWylACO193aL7n1UTZPWlhO4olorXEa2jvVzTB/mgTCxsj6J4+
ZBkXtbed9UZOM2c8lok+qfgbOAZflsQwcUsK2k/brVER/LwTeiAD8oKR9UaTqMvLqBf7tv26XuyV
2xT9s1rJ0c1AJsWDy0cNDjo+shCgDmQNF5DJtKFKP/im7GlRvuUr2jQ5gCDRQwQUOboL7Qv629R7
9jUuMbY0RhAWFEqoT6yl5KL45YWUDu5eUHY1SU8SSeU/T4c0sutHib3a+afRz3CJRfGnTVLX563R
GiGtcGiadf4cfnBuZ+vzVaSM2TmTfanirwF05RFSua1Xf8MViIxhf2Z/KhxrdFSzwWcfk1MHEUZ6
35t8nyAxuHrQzmf2Q5SBGzZoLqTxYcGSXymVN+daXiwqMETM2AszZef+i53NlGTv/KknW3MW2v17
8s3hapDFXgB/qL9V6UBasD4lX90ndURHplnN5YnJFez1Gw7i4ydQbcoKcduh/owtyBAv8ceSVkp+
5OCdUXrPLSWYMPk4+6uUx5Ucqi1cUeptURbsgDtIURZEg4drw7HjksyRKD9CSAdGK3p8I73qdBRe
OrXhs/pQ+TAZyX8K5AtpF/FfoJBe7FU9FdDYaRClmj2XUN0kK6a91oHx9FgHeQ5fTq1U85ozEb91
KUTeycWvRYban36TCPveineExmzLLQrTh/zownoCvFUHS7b7NDVUZbs7ALnp42ZAAH4ahJII5XFg
EIgz97TuT1K3SPYkebx72+GBAoyKW7ETJloT7omAnqxSby13mnO1AkQNhSbMAfHrNgLY2ooYcydi
/fPJY3PSin83F6WeIYRQZdeYn6sTX38N1+q1XUCpe3QihT8q5XC6uSk1ojiys+7gLFbbIGgsagkd
LXvywcfgKodTXqDwE7aZI4lSISeh6dIEShd/LHnea0SJy9muELMEvM6KeFY2eMDZA1za9oAyWn83
aPBowT7qVf+592N05yH/KDCT7e/CWW7L1jNhySDYsKBUpIGk/1P9zIBGI7oCPv0RNrhSLk1HOZqL
nM05GVkZU8LWTJD1hFyNIaRoQ9UD4HLjJASOndXmJck985ql4ug+QeD2S0JU3ur+lGrKd/Kx8YFF
tnCcwpvGqFznbt6jRHzpcBWjL3FNLYRDAXs1cRPayuaWFIZK5qJdaYM7ZSzz3ulsv70VAu4Lihx/
NECntMJXbnM6/6ZeA/9Obz35JjsdNmId13Qg7kq21pB/rWTATF34UQYjBNXMNwq5Dh82RRCkMrGG
dk1357x38HXIxXMykLt+aBOnYhL0AIYQrLbRMGqDWq1z9B6R5oXzIQbCPLdBtfMcYdtcWo9x/U+5
/Xq/22TwSxUn7NgGcRPt5xCE/yvVf02MPIUHf4f1s2IU4yUd5b7wvs3lNk2Mkl7PIpqVb0nChDzQ
LRBwowiwFhiS+YY48VhxBCAAPISXYCtDiSjdjG3IS60PjUX2FS0QFsm64INpVj8bgJXjfFr7m7Ru
Sr7vPKtcqyDuXjir8copajFDu7aDKaDXppNlAyi2LM9UMgnLFb+yD0DpsWm8AU/On4KMMSCx7ZH9
rZHlFuJPXQz/Ko0qXnfiwVWDTBdpw/MsZf8uJgp71y1O76CeKXwLEYebFyTAMCXlQlA0KnQkdFdA
ylhuviEccwaw1hSAEb5cfl8TplgZoIAYQl7OwhavQMW5K95JidVZTkNCoEftc5L3SzCdcuTc+4ea
MOQWpN6ReVpg22X8XBxcrW6ReKKAJI8Iy+1F9jMLwWsr+mmj4c00fmfTMtxhBS5tt2sU3ZEf8S7Q
y0GYPL74Hgis47TbgM8aP+cqFvEL6bAaG/fG8wzXKSQjJhjKRUUvNbKpKfFj6bc1RQ3YHS3ENZdl
OLHCkfjMpMeL/sJPFcUzeU70CDwS7L1d5QLXUwZw3ZxrKrfhxsYM6/D1VHkeF69kLrYkh6bToxNs
qubm0YWVBTRQYzaIiNgVyExumxb7cwuQ4ry5dejYX0cWQ13URbmsDuShaxOVHej/nXGqW7KYGmBM
Lu8Z8rtdhWgHzi8LugA8xeRvfWqGezL+XMP2L6nGup6d9HW+fp/hyv7tnnMKSoahrAIxojITYPeX
Ft10y2ExWvxC+cKi4s4oKSp8pZPNCFCpeTOXFWWD9e1e+t/ko6TK9ed0fPieG5uu3S8LxQaNgMVI
CRCrbENFNPhyGpWyYETioYi6F//WhoflbFLGylLJm5VffGLF3ncHHr/Yj7eT5nIRnbotO3cp7OQL
ibNgZUYhu95qoXC7QHY8fiotDKmynxjt9dqlBJNDWmi7+7/4pMsmT2zxv7y4hS49FfJxU2r9EMKX
NeRSAgIXtVu/dPwT2LH1mN8rSVhW9Yx/nfzBM9uTVyz6dv/Ji/D8vofthrzfvlE+Ii/j623xsn7u
FwGgf/jypWJwRm5ttVHgj8Wl+axtnhz8Z0+z23+L/wl0vAmorGsOl9LUDrYFg6a2rfnJ0rU452Wf
0EkOADXUSXuS4Ny9MCAxME42QWIJe+oK48QrZhY0SlXY4f1jxut4g8bos0aNvvh6jPHnhuGtsiNq
eRfHspdkAb1GDwuOe4lPrKIonTPE+GoRLfGQ2LdE/GrYHuKXNk1vbg1DZB2+ffmh6r7pjVNFlqAT
jkjEgJxbA67STVdH+fN1kSd8EBMmUaHss2RWOUB+hSewf15UNIGkdfR5xnqE0cPLB1WgMATRtO3R
wngYYKfFORLjtD8AnOMKXme7XsA7bcZme+UOi+xg0PPWNR4pVsltQhxi5VRf7EE6e00zFj8nnP1d
vaaO2P9zPfzT4YU23Le9A28CnSFv6z/AodEZ+on0Z+MZLr38LaOh6vFoFzAeGrtbkux1AgywtR2c
xmzoWCFsdQto/QzkWJK+5qddVCB7MiM0OCRaQoJ+ob3D+QdyfIp68OlqFRuQtU48ZCS+jjJ/yLu2
2OYSNBZTMEpCnDZb2HZXzS8FYSxewz7NZjRkW9UfibjclEpgsFgfkFswG+gay+t93CvIAlpdMDAY
BriAYJLeZijTqG8Nm6FbdmTaOc/5QBtOOmmuXgKEnUEnww7Kz91jRTdHrwrAFrflKKQ8sdzSQHYt
6s0YWF1D9tQp5jbCMYJmq0FE4ejMa5DM2tKolqDpAVEvcDaUpohRKu4Oc95oYKUPK3iPukZW9Ufv
NRN8EQNEBD78TdksogpTgbkaGoQx7HDY9b91bQU5AIaOGvXI8cx0n4raQvhpV3x8Fx6IyZmDqJY5
HbJUnQ4mahSj1/sTbXqyT/QLzon9KqGU7OTPIeIZVS4Tkea6tJQ/fLm5dtbYZaP7hKV2wK6WR8NQ
SNXjkaunMOuuep83F3rWvs6qAovzDgwIWuBiHUY84QvTSZhctacslbUdTuE2bFuecCrgHPTSlgyM
4ADHQL+0ky265rTdYpRmgPfM2+Sn5fbAw1dZJoVM6DVki6csCBFOMMHJeHO1SVdJ6Dp1vQ5SEfbv
XKDWyRSJ8ifrOemLfdyY1HXQa13+KXMxxw/cdQ4q2r7S8trFC+6Hm7QADB2aUftVxjlyng3suxY/
QwbZgUCRKXYu4qzsUzSlFf7ndp5CvNjsJe7b64PG9mV6NGdp0jo5s2WMsMLV77AkG5vz7gdFJpto
K/wIG4fI38S4FSC+uY+WJaV/VEAlD+GgX1y4hq9Izk6bm1SqCZjRGuyu2I5uy0LC4LMovTYoi0Wk
oqhpU5ZFncO+Z+P9re906hLPfz3UrJHKEnhulvy2abwG6wuj5wD0+XwB/jkcOCE2S0MNj7MpTX1b
bANCaxK265vx+5qXywqykgvNcovgqYb+TLd9ZHVFGpNaX262XJu5QXh2D9vkcbNiWYY2/sCl5UdV
dIRNIF7Mud3QyGxf2gpaF4AkZwe8A3s0sPpkOXw9ckJCVFss2C35O1CLXaEABQVnop6KJk0uC9PC
kzL2A8gb/Ll95E8GtnD0uRxwjGA1px4EXfPj+aGZIBMCU8OKxNmyitDDam/WMZEvsfOXXlFI6jyV
iVe8DZxdK2k3ixUdR001NtkKiQ7l+ijwfC0acXdBH4HL2XGcL2sapZVDdZGQsQnS8427qv39M68u
iJmpnOfrqx30c2U0x695ERru0QqKNL020UYfdjDD/Ui+kpUMkMi2FbahxvqLCVosQ3TQmEtyKlIw
V3oT5XMhi2ivvftCeA5uTVn3vgRKKgzsueW9thAAh9ZFGmKsUzXyZawcOTl2kzPQHlm+euo3NGd7
1BNIDK4CuExMBrBaNcwK4FGQHZadRNQ+MRAkPuQPbW8xa8X48VCI/lZCTKQ23CJyIv6XISbIQphY
Fp1rfaRolMcB1Dr2LZzvQi7eY8VE42GbjhA2hhufcT7BKBSUMtc22s5XkVVOKcTAS0gst3DDD4g6
wxnLfDGG3+QnRyEtQkBfONESdCE/qG9IXsOof03ztkRg3e5p78HUwL4XbJ3DNlA9AMoCJ4gC9GEi
HDlDY1p7od0eEa66kF3mfE7CLoKo7L2kG6AbgBNOqV/sVnHCRbzFDQsNlLiLjhS00wUsbcMTo902
Le3G9QJqgQaxxI7IOSDZGWrz20aCEiu7Yo5HVRwJyuQ+2SjojSujjL5DBxgsDuWJc+tVvk1YKNKZ
qyUsZ4mdA9Iok1sLDamwOZKx14IYJNPmWLQGviO+FEE1ptka/SG+mQRHKyIAOaMhjVdTShGXOB4Z
CoeaUgj1QtBx37Dg6DLVr3pFNxWnMstYq/ZLecKoc1QIz4RfctseDIDR8bSPKpJ/gY3xl4KHmYdW
j/xrvO8KBrEzGhmJCIZnEYhRZ05VGBTJLRxBUxgUh7wPATJWJ+C+kAkPdPPEB1eeO5Amq8nAfUaI
UQdF23JI9MyE+ajfunCmfbrZbTWIfCq5p3k3aEETKePcxgKViCh/tmHLW7vJ1Hsy1y/1G7u7LIjA
wA3O/MAILmE7B6LTZmQYwlOT2X/mlZ41ilw1oaO6dtWVNaqwEoGD4rSwuM7uIE/9qM6igejYoRfM
n/OK6gIwr4pTGqR9vZtbSX65GSu/DzWei4fKKhVsBx8yXhZKh1Eua23lmuGslAcDZwAQh11EFZ+v
fJ3TouVnQ7RqZSs7gMWbwX4S7tmtsmRyKzRpZLVW53DYZgkiEIKNF5cmfAI1L3cF1hw7v4+EsORx
TUE/m95pt3hRVYpolcenLfZXHqa0m1PGeKCQtHpk/WhbhZg5FnUiqZqab0RGIrOUqxGJZeRuh5BQ
RcSIBgGJfj+omdASQnPzwXD7SqzV+e8qSDooIe9FQkKBazhDCHJJ+Kw1EN2gdm2hbS6dW78+yyoB
sQJUmlYzGVybfkYNiQ864/J0niXYvuyqmsAH62yfMII016ss8H56jr9Vv4nE3Dzq4U0Yx9HxzjQb
YDidGHFASWtwrTx3o4k5/ZtzPTsUOIS1w16N8Wt8XK68F4zcgpYLEVRwRBPqfA3/70sSwTmZXSeQ
xdbRLVWRuKxcr3++PPw5RN9HhYLWvpd2Ci1pzYgfhOWef3Cglo1QZyvofd864mrGNSkKUGdlJRnI
Y6U8n5A4cw4Jc/HpS7t77oHkW+Tn+/LZglP5EB8gAUVsDfPge53FC92kSDM5c+4wD+imwbLtoJ8B
2A1PbiRkprJ8dqSKnhERW30DV/Q42YQBUHK7vnkLC2NEAxbOu30tyumcPb50IHOpiC4TmJtkvC2Y
8P4vpHwJ4H2/eYPCfLGR6vU4vNy2f1K5iBnZ2EobD1TgbgiQcsSxnJ6R//opezpCSV6DtlJl3Z1x
FOjin2k9iz4tfogMONnSytXawZdnn7gAEc6RV3By88oldEegjLIUgo9uHIMHx3sOxqGR8n/CxjdZ
9ZZl1gAKj+nhMnlqRaQspvrffoiAYm1wwZYb9bfi4DcUPQNfaIVfXRHQ+jcXo39qZHOZvcdcpIoe
CFRBXlbb/es+3Iszblvv1BlTA9QvWx3eyNGeqN/pAWUGKihpXIuKWG2xKngogxFuL3ezgbg68CTj
TOSK0LlvruwdbSXGvmAUsN8PQ4qB4G+V/VA69TgBZ9GVo/MTpzC3bJ3H4G8VurDx5rMicC0eHqQK
QpxfWODSCl5nvymeIfpLqDQWpIGfGWYUv2b1SGEs1lNhmkqMNrbPMBDF/X5hjbbzQVbiIDSagZd+
oqz2deL+69iST14an67STZsuCiFXf266naGc8KXo4g/W9fBZ3fY/zqkQ8rE0HEeOfHnAAQ6Iaine
hfKADAXz8grA4R6ryYHu6cRuOWws43WwylDfkh1oSQ0AOmh3kXvP8xXPPunhgcYY+Li23QqQWjIC
DsYlTu7CZjBSt32tpkZRMZId/7V2LB0GAjVygubJa0PMaP424+41zz65DA5mwN8GX3USOJPZkXko
mnxJulnH2u93i5hIChIa11vj95Zp7Jwqay9RV+mQd7ww25CelzkWuY9PgI1NBWGVK06pmEKgrhTo
3P+A52jj3XfGARfQWVsU/Ut4VF/CdpaaQ6UHoz4J/MELnew8Uj9TAHs4KsWNnN7xplTlXh713iVV
sfL50A5WZJNPihBYofmvlWcmIwtV8eBjd9m8G02hajKDc/Vkh8ppQy560d5w0VvOusTf8rfghnMN
oPXhSEyj3nCC+R6ZHAZ33k3vMMJLG9b2Eka5QclK7IkrBM/GDxDPRmU1l5sNdhBUOjFigmFvm4Qs
Yq/4l/7rGmilCBqcUKiuJ0b2bOVLZ8DOxz1O9D6IuVbcKQa+ioYbG6d0zua83+51ORFrYF4B//GP
N3QFKpJMnMGE8qZZ2v/v8Ibj8UOOiX6fZTLSGEbruIzFBlgf1Cb9KUrgPDwCMw3vowuHBCND0sbX
MtHDEDx8Q98gMu0m21grmGOChgf9kVn+HrJrYIGiMH5mf544OPgbUsQ+ezWF23yu7w6R+M+aQETn
ihuHhS69NET0EHH0yNmGC4EQ7J2h+1ETXv1wpqdZjiWxsvgJTltrkNpYNPWGIM3S5lPSX4mROV4U
v+95fPRAHX/fi7oOdl3raP3+HhsBaGlkIUX/XEIgk/ta0H2h5LjuEFd8Re+md6NLXfSPINKOVo+s
ChMoAMrJp2yYwGvwBrGdrCPA810r5hQA+JUlI1+XQ5gTzgxYjHr/9OWisSsG6+1fbQFGikFrsLxN
Yenh9NAY3bUZZ+AUHYMDEAVrM6WDUIZurxTbTFRWHjDZHk3CW7Bf8+MX8k2gawE4CRTQF2MRK5ct
k5FJbxK3WAV9+YM9HY6IRgF+Hf6/MRhuZdifQ8IyFa3VbAZiB45EaAMcSFF0YrSd5lazWbkoTm0Y
A8pRs/kx5IxU53jwz31QpbTavbDRa+j4iX8cq1spyzDVzRYIP5tMPkkwfeLbuMrTiljJM3P3wp3n
zJxRCnKglR+V4A4MYkiOa0xadMfG4HM79Ghh9ZdONJtMXLqWE7mTngIX8cSjKhZ/a4yrKAeWmNVi
ufzDByXoViLYBilQjlP+8Tldxi9u+W6W9dVGVHMzAW+3HvIJDliv7BKtvvnL2B5ZjDmcJvZoGXg6
hNPa3Bt9KOvJaRlzdLc5wG/kVJGDvrOuU90kfMmhXd7jYRId3mO3MT4zpT/56cd5kKLuv2FnQtan
X63fnR1hZe+gsoIQaewIiuSnDEHCee8bxY4BCWDqyOp5xXs/ieNfNzAOPhMF4ze9UTAQchOhBflX
Wf3GnGB17hxjqR078PqQ/rffwdxsWuw9LGMQvnSptJgWQwnKzuGFds631sC418706gXeZHnVBTzm
+RWmd6wAGJCHqH6rJWq6xiWmN62lI5XQCtQOUUZKZVT/2s7cJYKFJ1ba+IJC8oe+3rTxMcYUAb2i
Pmc3LynLusp8pgn1BOpHA2Q5zP8zCPAWlzBH3QjtYRG1CgR+m6tuHosdfNEfYNsUxCV1Un0J/SdO
uYhh9kBzlF0Dv2HRDMAxVj3mGyhx7spvVyiUJtfuJJ2gmWt93grgy0v/rnVUQICRB4ivpgra2lKH
5DEYQRXM8o+tf4iCZImVCaZLG6SxEdphaxuqIzXl+5p+/v+DQ6fSVe5mhzIjFxRsys7BYCmW4qFk
/5qOTzmHXtsMHAgcpkbRP58bh9g1iLVfPXD0Aj5lScPup4TG0wHH6zj66gS5r+PVsgHuBbFCqv6Y
NQLqjZNX+DRYpfRNb86X4BhbUzH65KEJSk9X/+VV7Idx9kMxMEL09JMRXZ6haUj6RnDu8w192R9g
K4Vu6yNYJYBt1VgnEn9QXw9tgqWv2pDqcG7Lqnl13pZ7xgqGo+vdY9toyoJegMo/J790cwphfrQ2
zCg8Nr7rr5GsCp8oyA384aRwrQrXgDcqQhql5yoGUjc4iAstqD6tFT4vD1qNKemGSBfVoqS2B/xZ
tbhHxBdBDISH1rqOuFhL8M/SKk9CqLG/EUdkd4su2FdWwX4Uh8BGY8FeGuLgcQzmWcOUpWbdAevj
pQ4gXtmjqdVenRQuLVVLXmeibSCYhqeG/2ZogIgkRHk+rB6xha66zvX/w7MgAYtZKcB1miyDFpmD
+6Pn/vYt+Jos9z7eylTQ1D9g1D+bL7VqfJ7kCWHkbnWW7Jlua4pijhjZXboCEgsvbsJqhZhor/Ce
sRi/RlvP4xg+CHM+luoe3vl7ATFSbDoUOb+nOlkgmCxpXHAgFOSSQSKa3dMjSoWBwcIy8Bp6gzTX
frC0MsiT6k5fbmvjC9W22EwdnMnfHRJvRWuai8AdeX031pbaakHazdRDLpCG7vGZVE6vr8OBYxc4
3An3hnbfK5ZoSic2m5jwniTzokKvIfib3ajbuMHUrZhf9ndcsziDJZAYowq55v14Hnw4wggJsMiM
1NBYMaBzTGqq+qLA50+AJdgSsabY+EeI0ifAz5wpaZwsqxtItaq9+fMhWv9DZ7HjangwDb2kSvhY
3wdXlQTtXINd46cZm7m1TAYfIbn8wQqlL9tn+SHA/cDw0o1mGCkhzptRVLeA6RmDgM2MzOAPDSeM
yHIYC+NAD1hH8V9WN8cKFJbf5dNHY9O3qsnG5WoXWF5qUxc5S78F0UnpwJsTSjUJu2ozl0nVHT/w
yDBhpG6uTrpt95+W4n+1mks9Nr6OYwWxJJvRZMa6qlgWu6TArC8XjzQLtBrIPgkYQqYETgFtHZep
mzbeirC1HqnkXkopxz+Vg7TqWp7eZ1colAoFHSBtVQFKohkmzXgTUNNh7P2ZnyASTdIFZl4NDTKt
wTieHfKoTkTeBqRdM7OgMUWCCZBWOFXKeqwo4A3l/+iNxDCV5cPQ6ibsG3IlDhiSeaBTTaLudw2O
G/lYpG5G6oV4j6gePN2p2bWkWIldxXHYtkB/TUs/vTH+iRd8hM4uRuJPrH4169jAr5zmFOfF/uXM
emL9Rs6Dt9VpuMFw8uIIiGMuIG7SmeEnLgvtcEgTibCCVlnR8jXTq+2BL54f7qE1obmg4WSa3/Sx
GIzDla4u8KjeG5D33XgzxtXQ/MF0wiAVj53zoUwRYXP2fvXg0EseMk1lVonWkeCxYSOnLk4+gLph
23C4i+KhEy4vAhfjmCHdVXihApOAxneQIrvYf9oQ2d+ByloEFnyYo5JWjTF9mlPufQpOdmaQYeie
OFdiIO7z8nrenq88k5PBBvyDViQtSBVm0bMEiPTnS/N83ADSLXjlgztPyp4jUitjWIiiEsDhjgmT
mSE0U9ZXDC0Z/dlAaD6We0ciZTDg8YoeqLOzdX1W0J0t7mqnv4+ekHbAJZHYeLBFqLcU0OCZeGwv
Qo7WJXyb/lJjAFKsfqzFmw5xbLeOxZLdwJwgYwE5j4vGvF1sBkae7/qiz7xPFDWpzbdCe0qOWEUl
tJ1mBZGwDmUTmXAlcPNyYK1YU+JWlpTPB4oLckVYcDxSIZPKLd2TJV1DYDrxWZulON2e2iH49NpY
3Epxz2yTEl8QwEMaTnya7SA83zOFsaSyc0DdBygScrRoLak+lXKfPMGyIPcsyW2HpNiEJFfn9lzA
k3MgpP2/H3vyqcOdht4QKrC6G5Yzkn3Z7Wm4BRTnBfK/a+lgBi2NomfrdkttKRyY1FEEPeaCXGYe
ZBTmMkbPUPl/ZdAKgjrBbUYtEhmVJ3j0058/6VCqtx5e0AjxwfSLfEuUMms2SoCBVpaFRbQw9eCp
DjK/jsk952S7bJhHBnaTGxtwHJGEe9ChI3JxS66HZ7UySQg2xsuN/2XIyoGUxJE6pkywpk1e3Wh8
/m1rDw16azfg7m7fZ420mC8KmMgp/TFBg5tvqXV259TnASs8mDx7dFHZVRZARYOsHjFTL7ax/zXf
J3YFbd5ePYnc91YcUNAkXkbwLrpOwiKL9x4rfiuQOZdho4egDf5Ryg5omRbtx945OuSKXa3krRkx
t24eJmN8cW8hfeqf7bQsxxS1pgCLAIjN5veaXY3SS25Md6SbIvCBWJ0bniqPbk4MlHNM/s5KqoGU
vL0zKB9odoh3yEpiqzQU+1Dnbg6tHO25jKW0BqHMv+nDu6xeXiojMKA/g/LeysCRNbOO81LZEw7h
McSPuq3vTW98tcxcJqeGlZmGaixpaED0VBBc0CtGXZGDS1nhsnDvWR0JWA59U7Mf5rMI37yQANn7
23V25jY3c3nw2oDRhEvEjFvD16Bn+bNPt9MMvxUhU2DNyBRSU5RPocb+fkTJplUJ519vLeX/0PHF
hIXP9+U2nVom6qLLX7ecdtoGUdyXJc5gg/VjGDXsEQ/ukPYgLcU3Hp7tRlC7+Lhxy+vwX6Dz/ebl
aXah3Cwi3RXIafW0YjwhdakJLyhYc4JEWfX3VQ5HD5f7rN+PPWY5ttHyO8tvpeFQ7xXMJ5o3Ue8u
yF9D2pEvJhs0+z8kx9kvvAWBVp4icx5Y47lQtNKnucE2/W4Ti8aGkCqcIJAri8ycml6pNg9MsK/B
oI8gQvRdyb2NZTJ2RqCjGHgPqoOJLyHJAEOfTVssbnoKWcvpXRexPis0VsoPFA6bJ7YEKAzpe3xN
kGJtw0ZjtddZ0yj1MnBUvaed6oR2crOkc/bqzKv168dZV8rJ5OXOjzgab84nC5LNBiOFHzDDk9Wv
yKezlDLikV8UEVxwyhw7GWXpdtG9+NqoK39+1wIcQkEh8/wlG9gsd/tYaQib0Mfi7V9XlKvmpeXo
2Jk9zXHq3p0RkNFx68lRYQEngEJe8XjAERT3l+x21u9MW4rFQ9bDTnSs4Nwk/wWwBk1dNfNFRgv6
LrXGg/jUIQSlO06SdHg11RmVrKBZtWlyL0xEKR50pDMTtaWTIoVy1m886egJZ/kITnpr7r1Z2Zjt
BE0SrMjez8CS+XHRZ3He3QAv0yjtyg/K0isZ/tY7Ov/xp2KP1mKJ/4WYjASao90p6+YI0fGCqWMj
6D21JT0A4tXQSGHHOHCDQM56PGFIwsmw3AIsfBb4gLUrO8pKqk9OKsYZfK7w/DJalqLEyb/ctir+
sKYepkBPGklRB3o6OViSsDnu5NU3iwDAcCPvEyjRqgb4SJi5VZDShDTsszOUdn2NiKrY8wJY+rvX
lmnJEOb3xu/hyWy0A1ZrErx+Pph22PJqRu8ooExh3qD0He+Sqe0qkkvPmCEMp6janDf3jKv54/ax
vsfcPWb7pJHGYjvUHvNTEzNEwPGaHoDvCsBMgite0QTMrysD8lbaVZzXqiM6ILj17Sqa+0SN8dwY
xXc7/WcClAZvV/UUj678bOoxQ+IJrX1QDnAzh1TMVQamM4J+VnP4j3Vutf4Q07iU+xZn+00iRN5f
OJ7iubhGynJ2doGYO0cTQcVXCV6fiY+Q6/pQnySqCKxDRMnEJ0ZvcuYZN7EvRLEzCrfImE85vUIR
QNqU+QkXFBpDcd+E7KNw7AZgpnmQDLJbj7nnwEj61v7NmVlEhVRdD8FEm3MdKmUtjFwu9quFfuX3
ta3xIpbdlKoE8XiLtKm0BAsg6dd8ErN+EbqB/A2Cw8RDkQEftG/s3ayH4TdfAEDMpN+KFrV7yOO3
DFvINc2SQxSvl0zwRm0E2VZS3rjl8BQO0JziA/PcmGzk9XP1l7i3WhOSta/NU4dEoJAm6XQ9hg+c
uWbsSMfbKhwWYlmcPzE3ZCmBYK6Bsxu800UV929ZWC0gZFZnpO+uh80wKY69FrXDaON+pfT4vlUw
KbbtRWErXiE2O/afWJvKyOLUMygAPzQaw/hNWyIVr174109zysNmfs0A3HGh4iEXTpmFyYFvDkAr
NrgxOI1TOn6NY5AIZbol78vBcsxy+wR3U3iuM7D7r1XB4Oz5lxjZ+CjHxoJyqYFhG2rLLTUUqJq2
p5TOR//htQwW1O/4Zh6VuHxKm29m1FGeeI0Cv0x0Iakim/usML2wUEJev4TERptM1HgkqxLHwJUv
MpBiCReoM78CK6+N5EVbfMe9F5GLy9k9DE0xbGirJwziavPWKpQeV4CsgR1LKNk9X/HKvet2ZNUT
vq5FwvPch75RNzOchvfKnvT1sN01mc2um2FYQfP6fg9jc+0VX9wC/Rqamv5K1SJSVNBbjPl5dF/Q
Vn84/jXMFtt+3IgTAXbtzAOdDOQ6roL5/f0DnxJHC/ByJ6yCwv11mm3iZQO4M36xgC79J0+dttcL
kwfeLyKf1KXrcsDLk2h9EJMQ0qNFDo6nvU1Il6tPcPm8rlhKePhhfalPL1uqI6Scj8AkEp0riQ1G
6ubTjllgwwysERqXula4Ww7X6HSFgyGaiDneBzBjp0vbezL6ZlyYMAlES93If3YCAPMhMtDz3By3
BtINNcyEtpklZzdprngPH2UdCkQlnmMDGcZEzas0IgE2I+pMURrpPrbp0nxWbw5RXuZxy6bqo8l3
ByvAZ8rbv3oGP1SJaS4PjcHkTd0ECOvhrHyDuszcJe2dRcGFaerjXrBrBZq4rVn95YRGdd4DUcbw
dC8zT6+tK7bqI/2ZCstY6dvlcazpI1E38P1se5hEq47VNc1yC/RlRBd7vBg+c6cJfoKtS7CPFcfG
yz1a2Y59hPZMB9r2KLSigMgqEzyyVFN7VnFpTUiyRcCae/Ek2kM+0CIQE8/UrftEhJbzhyWQWCV7
mdRd2CPcc5HyzM/7PJHhi7ASRoGtfgK9I+2/bmAPWrWQvfs18AETBnONnokNUsNqQUVbOne3D5q8
HENddEijR14BSkhMJncsW5amCqun/3n8Ak/AXeNt/7QnhoY0h5I/POUCMqSP0L0fyQQ1ZXHaym6y
aw7I+bbs1Fvb2uPRgZNHapfOwoHVK2hmrsylJPlvuHgsO9b3RQyiSjDad5JWbpRgRNe+phady0Yp
jxXdQCOP47CZnD+fHjWQhgCyh/oHvYnwejB3I1KOpVopsOLrxHJqYjhDBlzWbcUvwgcePtYHoPP4
BzeW+h7plBEJrqCuv1Uj5UpyZDJA/ji5n6ZPwiU1aj1R+/Kx4g34tdNwDpOhU1H5aGSpZBN4hcST
EMVzrBO9ME4kOcVt7Rhq95o078w07ZUM9Sxwqr1T/17Ik8k2XFgCzo3ILERy9XuCNARargr02q92
FQQSC4Zw4URu2NToaOaybl5F14VYMaB010+qEQENfD2U7FaDoGbpAk7Km4Cel0ZhcnLqivjb5QxN
BkGYxUOB1AN7VlplNWRlb6gieymTf6kk1mQ191LnONe7UV/Xv+UGBKM9oPtQCVBvhqeeql2CV1q5
v95yEDvXfJklmRfA6fCr3ut53CoDauq/vXNQpBu6DVibJheoGu6x8HpB/Zc5z/L+Wx3g9nWRHQ9F
4CRaPesFWxfEQInWcf6MhudV06UQGsO204I8s7GpK7Ni/rbSDk5dq9eEXsR9ULWcIzeV5NmrduKA
7Ou2Hm1jQ92I1GxmZysWRaRURq3ewt5BUchnRa75W6DQaCnS0NplZW3FoleK1sDdKZXam3hjNv9a
reWQXffATMxP7XbXdc0IuSKRbfJy2+7rWphAHIP7azZw/Ro+JBozM1Qo5xBsE+pX9MXttZvce3Mo
kjygpUvYw3khhxD6mOK3evXZhAz04FNj2yO+WX8RT1Yy6y02mAjfw2JfzZcoQrYzWBRkNh5nM4UX
kg/2P0DY5yHlW9deiMHa63iGFgQKAg4owfkrko0S6fVMjJb6NIcw85mcOsxu4pTdDdiLVrXG/pIk
mYOoCBtkhOiCcF8OKBo8VIaZ6Li7ZebrauIhyTdQSsPzRGHsK6O376IyJBmrrkaM4Dx5Jr8rSlbi
wd82RHlAtcMcb9yy7L9MNqMoa+60Ka9eJ4iN7BclQcLjBYyZcXce3EVmt/tiyoOWLGYHOnrWC7oN
2p0AQRh9AxtXsry6wrtnpOVYrL3KOa8h4edh+4nvYLCF6ew8oANAwTmV+dTZIilD8KvJMMOhSsG2
VpmQ80UDWGnCi9B4HUhXJNfnuRUBjZRrsbrSKqSDJ26FwH9yhA8FfZD601/tq9kBMz1Z27hIi589
wMKcw07dUgm2TmnEEedn4crPtPeyBdS7UBIScRVxsUd726oWYa1dKbTmmpmxI80gidXmX9dNh+qi
xnEredW7wMKbgOL26ipafcduXW9m9Mic9E/diBPpPxAk3v94km9wiqkLAxCD/wb2MvyABI+lAYNt
DvE9LlnauZ+GuIzqEWcoflTMHMbi5bMObIZ2bxYtVXso2g2Okkdkx0QwiVOOYOiH6H4l2FcSLzaX
MVhJyEaStokUejJSgj7TtxnUxQCMb/bP1w2lD7KWusfqGLXNy3EIZ8sKILPgaIvzz3heVSvcbFqZ
M+r7O0bqUTD24NkWrzhS1KFMy9uyesYjccSniJaNhY+xVV0Waufr6fzUuWyGcgafc3FWFYH1zVeW
UQRxjRL4M3Zsg2EPIdKHF4AhhFn89urukspiKtC+FHsf3KVkFXjGn7/laNQ/+/wYQbj0SdzB+mUJ
5wmjpKJrqbupLc/CiTqqOlPl8fZ77lNcIeKEd6BxzuA1SB2rS5ekm/0a8s3MoGGQ85WNH2HtNMy+
9ry23TPGftReiVEQbtAieXDm+EUI9sGDE31k311fKn6y7cII9gnbUfmYPVpktZ56NI8WbnnqmCwa
3Pfqies8pK38kt6asVcjfq30Himk5Rn6JRPARY8vDG4qsYIKNBgCvVstutFbgEczQrN5Rk+kERua
clZokPE8sRt0EbP+YNhqLISgEbF9UJ5u3GvnF3XrmG8t8ypJOPp9W/swSX4TE6U1E6nK1ldORm/2
OROH3VVDdNf14MRHzFhu7wxLainCZMDoEX3aq8xOBWCbLf6xTzG6FC+DoysC4189E7cnONfsmnTO
PAGaM4pzLPAsWsm57nT2YFFbvPSlEu1ha4hNL8ME8btPGZJJZQUjtj5Kxmdy0Bxx1niVF0uD/U4B
2Gb4VPJ7oIq0KegwoehLPfCj2oM5UFIjrtmmyiv1u2/MOhWOuX8p1yoFkqY9PRNqiOomGXLRgOH7
ZwW3mEQF5hjSa0KpVMgVxtec2bR4j9iselSHcWn4t+V7x8e5cBYJYZXrGw71bUNSMBPCkhKhQNUK
L3bjJFq9YJyMBtS0hNdr0LFObFibmlQBG84hPBy1VqwjsS68H0Q8ofw4wbTaYPTGx70BwNqaEfFu
6g1qj1V7tBTMn5EJsGi7ZzX8377nn20MB7iUUtTDkW32okxIEGmp/XS0nkucnhYPUAQKvwTuGeye
ImXLZC2IudKhs0nBAl6NK5Ai5Pd47EYxQ59ub9EkVhIM4n3u8rscTzr/TpdOqNV0nCCT6tmxO0mW
YnequaG5o+Ljzw+yLh7USieJLVEJQB/0mOFCwNa5vtsVZbGqe0Oc9IqErnO2cIedVuFaS/FjBBVB
RRWLCvtRoohlLkD2VU9PVRP9ut6gIwAmWxiMoha1Y9X81C7vnYMqKX5jqMckMeY7h3kPqVmpmRSi
w8DaDu2ZIwLBO4OKNJ4yUlJ5MJ6DE7KISe5OJflCg8i6h9wbXzc6Bx+z5Jf5OumjOSIKYCXycOxb
yuYgExSqDkksi94V1KyDzGaeSwDlTPPYnZopSQEuwyrbj78tKjPQpZZPIS1ZbbRcngBcBy0ofeCn
xnmZhY8y7rs/Ex5vwc35SbJu32ZjtME6W/WlHT9+Yt6TLTCSPcJ6qapX66BXmujW6tGS51sjx01e
HpmLwYLpf584Q0JYaQVXzNUNRgZARsWndTAiSQiEZ3ISztAiLPMgAjcV6FFlnAyKndtoJymry+v5
sddj/OIwVNzRewjnRJkwlhabknoCBJ1hJlRcts8XlZARF3zAPyxZd0eGakRfXCdqimPhMhziPoL4
gjfXFXrWGZ8/W2c3wQotrj15YbcmFHjnxdmtvTorcnBA/Psnvw0xn17DFxUjiq9MMFRviIu6QFnH
H/kB84dftBq3KJn+hJ3N94p5S7sXUVofIRIhTZm2Qz6mfUMnepDeSJjgd4JewQ5B+xMvU2qfV+Vr
Dz76LlpNl/ZvCP4VSK9e0ilOq1xcH0rmL0M3adxvf1ouKPm2CF/fpK1cp+7oA7iOAqM/82M6WS/B
8flPdRSqO0Ej86WCgMVQ53G2wiLf0MyO9E69P0fpa5G9WrAStzFEbZRF50RsC1SJqM7CWdSraJ+f
LO/hnnVrhny+OPV0xyImMyzAshb0YIMMjQh2NXyJ6WwwM6fyVuoPqWVkN5RykZFh45dhUWAUpS/i
3kxYCI1xwbXLgRSmf7BWZYYxCEHsvIhhjwAbN9E3EkSgJ6NkQIkipZtrVf3PqS8JhDcSO6JPM2IV
RVzinEZP9lM/QQJx8AP+fbFJ2+1JDPCRhDA2USBDIV1aSPdGNxhZisFndF0N9BagVBgNe4wefnQ1
uO7eeUFpyqtcDRV009rQoNhAaT5+BzDjDWzSs46xtQl0DSDkIoWM/x1dc6p5doMdcW7D+S+ivg/2
r6l1XiPM1xhfjNQ1h1ildbao7XBCVw9Em5Bft25hRJPtFpcVm54EZ/MvkuIswKBwfoaV8k54bJ9j
IlgQKivZZ+nKGwY8+HAbVXL09afjtrShaN/A2+zndmvI9AhLa/nH/tvXvS8FVwppDtAKfASgyotU
G9k1TkzdBhru8mezoIMqgZBd3Z75ret9rl9dYfon/aAry+Z65PRFaer92rZmHCvtg+yOb2hr1BwS
A9hnOc5JyecDcr97ebfM8HuuYfJ4VthxkbA3MqA9QP89um3iG2q50HFQ0QlYRD5yVZtwGhIzOxmD
WHuSciJUJxw3JIP5fQ3IZRori/lrsgLo4FKROv7NudVnbQr2seOpwifqLXmcWCt63n870cvMM/0r
2lxLFwrBH9CIBfDwzUTKEpP3SIb1OBW1C4xqmmTpDymmEoRYVC/srVzhExZu8WSUFj3nfk9O+wVw
p2MpuiSKX6MUNlocdplxpbhJhrQlWE+zzVX8QgDpTVljnAekmJQ5bG0JTBUnM66T/yTmCP/jI9uR
PgY1U5i6HATEQBU6rpebqEQY3pyLAWYBBM3dbWKrntOwpZ6i2uMszOd4KueaMI78gXpv+zWRj0bg
BuFiiosP6Dx8y74gWTFQBZQ3ZSh/726tfbR7EliCBEYn6jGadIkh9KfMvYkkWpbicT1VuZPBjSAZ
b2YD/0dswFa3jxgXdJAH4ei+I3mrUhSdT2FhqmGxwP3xjIAa5QHeUbDJiUFu3ICs6gc+Qwi2tsXY
ulwJoAXrUm21k2de7ZJr4DvRQ/rocozoxXFtntKCcUNdYnG4We6l0D8SLqWoqP3wk9K7wB7Tme/P
9TSCkPSwuzFGSXGwNeFvkQ+LqvwbZCiW/MdbvNEOzfiGn17WMAm2QwcfgGuIoYHtp6ygyypZAxX3
RlEBhg4QcE+/B3/V4lVxHwtKqYBKGWk9rgKDhHnk1v6npuWVGzB0BZ6ofiT64J3RC3vrA9hSVMsc
XH7Ey0Tszg6wK5kTXQPyMw7R1oECI8vugBz1CF7sU1gjP3y9wcSyyx9xtsi07P8qC/IIUOl04R7m
yYcUWjltqIF0fe4TJlemEas8aWw6L2r0n2lMjZZoQ45MnPMqkbH+/uo9s3Dsl5aSmBApX6HYPmnZ
bz9R3A5j6Pym5SGSsRIfJ7u5gb50CQ9/bvvZPbT2MI4n8ov02NHIuDWhIEegCv0QQ9Gezex1A6lR
YVCmlwkubHnQA/NT13xIb1vRSJCZkrB5qizWNKIJ1k7oe2q26t5uOwOQIz2PbPZf4L+rZ7voPzdw
2qiezOJBuJUTF8brD8boos+HIUXdsYcO/R7Nya3rWsFUyrw7jPFLca4ANrIIV/ExQK1ZEJVjBf7R
t4CQ2xSVZinuWOo0A+ZUfwpcjwIekcX6oA48i6dfPm0iNHSUMAYHjWCz8V+t02drmGYWiY0MS5Gu
e1+I6GFG6tOjXq8dT79w0oYTNJ2/dK3Ehd/ISVqg56w3sgxpj5ies4u2djeq24OCo9RokC//uaE2
+9lZ3IKXqz8kW7d31yrNGxCB6PkYdKtQ59ZheNQm4b9HKlMnEAGIk5IvZi5MIAHciQ3ZNb1dNjGH
3NfrEjLoAgqZSm84iO70v8UISu1c9VQ3X/B1XvXft+1veGrAwCCL1LWo60LrFT5DLAC8no9rvMbE
H3eR0rk25Yv2iGgGu+3FD6pifCxCnb3kMpKONmsQr+o8/uRa+rykBRKBM2FKW0bplHm7K6h0/LbZ
NxBaqQwI5Dc60V9DYtWz016wkgcqQS/7HhuTNSojR/b/aRN4un9Ookrg3icxFXyosE4mO7mGET01
Xy8VIPXfFwrb0yaJCyHA1MezyoBK5bC3Cf7lXSxlsG6SUU3AiwXDH9KPu5WHcYpBLH1yT5I06WaD
CfYlO1hMuJDEb/vFqv9LFIfIcHmqoIFM6TLhyktXMm6KsbKlT9OfnzKVGfBOXRJ4G5xLmfAmlYRl
vvXie08ftpnXu0Uacj2eMN2WN8alMdaL5TCDnnAlQOGbozzbZJC9pvUyQyzEAAvXPJA9J9aUIIOm
eQoy3gDFjYXDvQRtbP4ss7BsiEz3XD8+rktfEjR4QfEx9pS1eG4k2YgGb7g2gjV2kn3+yrC4PKfk
4YehdP7ZLLlJJSyprQiMovlxMuPIZdZP28ypERmklVodk8G2aj5hf+wKm/dJzl0+ZNsgu6lXSxWe
OXLK/IVmc/hQ5dIyXLGJkjpVg9+DOmiwUAvtWmIR0Bv2HHmE32hMaKeE5XD1ZWL59dpyQAPiFHBL
Za+gEEe15M39puq07OkNVT3+ovKMFRJTW3r0y09W63F0vnmKrOHwZDZ6rt8nGKK3ql7D/NjKYNKT
4kpQ9WVuCAKb0oR7pp6ZiqKe0Uf+R49ou5mT5MTSs/6fiKliG2857giwDiIyiSmwDewtIZQxGoCp
YIjkHe/64XHbqbjsPuP62PU7/sNinmt3k9HMBd2jqFgLzrfNlP8zbLyfLB0rvXpehvSY7QtR3gex
UByqfZKJgOz2+7ofT2Uo02zhVt+zh0jPNS4c1C91lQ7DmIqh9RiuY7DrKvK3aCNWGn0lyXeMdZR7
Vt5IEvqdnbYqVuiL029P3dwwr2ssTHXZ27KnwD/W/p5IC2cpPgFYr0LNC7J9R8LZK7sGaoN/JyME
6LKeXgPcviMxlhGYdML5DhuJ3t07n2CQ+VoaEeVqcYeZJ2buGEjHuShLvOiwYkX+1gUG3tfyAfrt
FYdGOVjXMXuQuQhCCEzbu634NPasAhhKooAQUkkqANUzfkgVd2x07jo7l1LHTsw/MBqHrUpWdMF+
1xW1xiPExHAyI7LgyMJVuunQfEFgRQnvbnLe58X8MpKG+sBOzFplHnUXjntFxGdQbBTVvt35y+Ih
9+yprQnQsu/DofX9KLzVH/X4carHyh10710DvG+qLLY8+wT9VqzCcEMysXxrd+EOhvBC2PFIdk5U
wD58hxAAu0ykrpLNPRHzaUb2PzDmw+53wg53SPkSz2bd3m3b37dNHu8NSXFyxPhFRm5FiAsDQ4Tj
u/xW2cHfY6FU1c9A1aULiX/YoHSNb2N28K5KRhVJ05lgsn42hFCcgRubXRa6geA5FZJ9GQOETTu3
37uFU9G/qK+oT2fRsTgrdq7/+uJ5rDQKMAjOZsXSgtfP/LRthGJJlT2/oJ4Y1FTnb9r0YFT6e3Ah
gMrFg0vWfSjCJSo9LALBWQ75JH6ajqx8aDy0SsxObVBVqr0sZ80rUGcwM4ZS3peZRrRE2D+cU4Qg
ejFNklINWh4MR5ycgrgo83Qi4IuoJi2YpVsNLh8W7qNyaaW1guNJSpo45glxBiGui52wz0n8rlFM
Amvh4b9dZDJIYXdmwujd3D8P88kqZA1yVzBLzhfJgVxQcpg7qO8TgcmejcTYxjcONbQRhpBx0w+m
8fj/w4Y0Ruwyp1rNgLEblFCMtjIdqR6I5hXSyt8zhA73Xi9cdhD+cpY1D0NvYeDC2BkKP2XdBUpb
FvrhoywTygNKREFjCV9IqGDGdK7OU/GtVj0CYnUex87nz2/tnigey5C/rcir6gWw90Z9XHuiU8+X
qn8KmVFSA1Pv3b4J/RM/a86IuxV1EwHUnqq0XOLsx+KqWClKnyHJ1iCAE6zmjdzY9zrd+jSk0EvX
Mij5fM8meYTrJriOlzbftAUyhDef2IkehntboAlsAvX+PJsHRrLrSC4uNII/NMuyXY9AEakEaQ3K
yw8ZNhhA2kfpv6K3/tlqk3BBcDcpnvRajuNCZ+eFHVnlWPMEq+SRl63csVdgvBoZT4qvUqbuAPY+
9XG6oULCYL4T9FgyT86nvedXfok1IcXJO6gas1qhEEBjQdXf0QVyszDuFeMoVzBBkQw2MNTSTHc6
OmL4A3gysC9MhjiwNYv5her9DOC5O3xHChdTEii6yXNSb+7q0JPXdvXjSPllqUl87N6RrFFPb2Fq
hXpX06Ks2/l4G4C1sKjQ2kp374vixJREkCiibX6nmqMtSMZOjKw+hIE2P/2s+vKBZVS2+kSolK/H
+yHk3QMPXbeqqPMOyQztHQamDvUlEFEYgviH1NIIC3MHaIw/UxlseDy3+4TgrAVY4CI1IWzSFo0Y
XBuxhmoiXwFZHKheQrBvJq1JQAnypO20nAGIcTJw6b8sg3/H29Kdqo0857d71+kPXfkKXFIRAvLJ
UPw8y826sPl81HdDS/gJCPXIOTAuPHBCnyGvnX3+6xRZ+intOnvEZhwZV/jPch65+V6NeEDp9dYz
MR2oEX99HNzDiFppQcWRiT1whtDQylJv8Adz/xJNjn84f54lKlLYkdXqtB+8yqeX648eb5bn+tW/
QVkqIzIUH08k9WH6jgfcBdzIDa2z0NSqhIsnXQdnR45bVKIslwYf0V4kjMLhvPynwwZTQzqAzRxt
aO7b93TWE8ttX4wh+Vp2sh3X4BuIRcZ24gNPs5KQd4bmTNRVtguYBbUreLaI28yVMiVnUPjZztxn
ingWyw0nSoz4xZoTiSas60dsyOgfk0b4THCDvz9YSwe+yMZLtLGerXaGjsf3NDvJs+IygeT2uonj
VT3nlzmMYGM9cLjhwEQMfvOGlQraUkyBNY2XqnzZ1VVXkIHMHc6e5lyuHJD7U1UIity6eplxwvan
LP1FvCwBpXPeCLRtiIvOCE6F3HOgeEI0tpQJBq+/h+UysS0JeIxVii5V4HL1Fb5KTrvOpA8/riRv
fAbsktbpG7WhOeS6yeUdI20bw4v9Bex0XFz5zRpjHcD1wTNpaj1DLFgA5O2zNYndWAAnz0J039Iy
qV5NNs5g5booZO++pvftVJVQWlDAv+t/Y7Q4xDEPIbZ+oQ4ABGlBdQU5ZTl5vuDS9T0WQo2pFUrt
Iu3thHYCORrz2YCpQLph4N2yOxe6hiFfID3/WH/BD6f5MDDeNUniNO7Pda0tsow+1HUVNicaBHty
DT28NVBhnocQt79uCM+HMiENhW6b/fc+3bXJU9JclUZVxsB3wWSqP72JhDVRLl7lTm9L1ukXDB44
e+lC9eFYSKFyNnpijNE+VZGHXbRkeETpIXLRqxrNDpOPZ7sHt4qyNoYYgRqJ5SKvEK3IbcEZxgrL
WZfghJGyEl5wyq+xC4rW6Wh724XC1L94xDRGWs8dObqOJtjzumjg33ffeQ80ZRPAD1a8oL8LE/w9
stq9ddhZaDBxPSkRZEBEsUoHRq4f4DV6VkbHiSaY5BBQn7okCQx6Xu7PhF+4b0095+Ay2LfU/NZK
rXf9qIJgsmAY1R4CPefWlfSIo5dczYOKbT72SR+dZOEed4eBgb54S+pLgYJ3Rz447Px0lH//clP2
+kOBqRERq70TDMrgz74/4HDi6mBSV+n8Jzi8MzLHvTNKVhZHTu0t1NVoZMCJzq39fRwWI/kGlaYP
B595Y5Tur1JwiongKfZZU92FKECzNV1xtYZbhPMCb4SrMuByS6I6opogKcD8J9c+Cv6tDadrF4ai
Yk6ORMQYVgKDO7kUo0FKgc93+2KpwpKERlXJ++UM2WcoKAte+hBJkJP4OP1wcDgs9uixJGgkQ0ph
yIzOg7DdbW0TV2owYjB1uK/RvB7K4ivjYQrrszJ8kLKNZfxC9lSAK2Ml+Sna2G67UWnKvB2m/Neh
bWz0rNfb54IdcsuOcvvufwwARnz3/2K+D/ArL6RabvAmYjogw16OkPOsNIP7sXkX+nQkuxRQRH/e
KZrWg3U5GFmxW+NEvpJqWAYx0Vag6eTM7Y2wZNBsl574ZQ0pocoifWBq3+AL0belVP1D2IdLK6dS
tgg9dDOBVmcWiIiL14/YVwCHK4b6N5lQMEmLXQhZ6eicIzirAlBvf7UX7PY2ytX8oFzg0hshNwlQ
fyY9PVZuCN3/m4REEiJAv9PyMoNFxG6l8MsO2tLSRUWHHXi2odE1vYeVaS9qqKRGz+GNydlY87Ir
w8czi9OFt4WGge9b0RP9kgk0NhCZBasvRPpxyngmhLPHH4jKCXKePf7jyNNtxrSYISMGr3XFhy9t
BgQjoSi+1dRTIkNArzs3NbtrZVJvRQuFdHRfaPvuYEvfAxB2An+9d9D+KupzX/VjIWObw+5WZ+ow
rL57Kip0LgFU9JRHGK3PnoWel51/QiU7ioACtu4a3kn4L7MkUL7eu6hH46nOluuaWV/7sRhC9873
zW+CJMSrvsOIhT+z+PdW0WRKEB05rk3F4iLX26RcI9tSzZ3pOob/VDi6mv22++hiX2HrLWhYhLmF
SDwD0FsfRNdA7hIyVEestMQNAL/hX2rPLecqKCEIFv7nBn7XCpE6G+vfRhWQlcDl/Lw6zSwjQlhx
zItZ6wxkR1fTx95QB0aYq9isCCY4HW+ZEH7pzpoWPX2xxWp3JC7XLSfEDYrUVbrbnp1NgXW+YAYy
j8te2zG2quM6mGZa6vYqwQ9jwIN5PIK8Gmv4OmPSi6vhCzmy5fUcw9afqeRJOKlHrXOhdRh3n5I5
89ryFvW7SDNsfBU/ATyGiSZgf9GdoF5kW7bqEbMLQU1k8qAFVAyEgiXlJhtdyEEFW01zP+raGhvM
uWTySdmT/3ya9CA0Z3zeYGJagRIpViz3xy6WCjEjW/VkEePlbMNKH+OomIa65vF4WVpo41L2lT7A
WzJRM9tup16eHjbxkiFbhDW/laDJiGz0PBYbFeC92lszFZn3VHsyrOZVnLnYMqdBmyuXxTvkF/1U
sSwBfz4WLqywbqryV4k32Sxx4Nf/ymEW9jenoNR7rAUpp/DQqxivuKWjB0kjL3mnZOt0uE5kqbUJ
V9dgj3dqOf1y25IwZCtwOxJSnFW5UrYPVdi1+odM2caQ2w1npSpWHE0BZyaXPTQt+ApkhwiWzjEv
WcYELiHUd3eLX3CXTa276lAC3CW0Ykdi37l1nVr652+mk1PAjN1HSgHbmcv1K6O3gCIdWsto5HjO
bp+fCstMDXPxQP4cic4xjUWS3x+Ikmeiqf6L/PWrWrNRHmGY1s1SQuLk7eKv0e5V1r1gc/kW8b/i
xyuTijXhFklebc6iikdpZuceoG3xwoShm8pE4/5OLtHghsV3z9Ir57awooOxsze4khAeLHU6WKeX
vmmtLZ/G6TXaJEX3qtDejWrJ9S62osrxJB0fP5iYaI4EepNB6fQveOnVjib/78NA9oF6zqRG2k6U
5CpD54bTbsEkbvFEhmGVTw2PMWMFLl1dAAT3XtbKgIaSM5pn42AE3O2elk3C/J6GKEnZeDIg2HFf
2zDIp0WEolHZameCloX/fDArM+1E2KOX4rD2w6D1Ksb5CXpMqSDEYwbQ0p6hNcudTMqpJr72tXcl
5W/cXT7kic+3FaEbjzJyqWJ3xouhx8/rYYatCgVNvQFklFFQ4Di3qW9hLLALcxgYyXBYuNwX1beN
JxZYj6rTo8b+XvIlxMdRMnRrbMFC8zUUKIynI7/kmLU2dDoo30cPAT2q299/xwo/zw8dNRPjYwcN
AqmN6SeUGVIaRboNI3KrKp7M53CdS8AywxARROtX0/pyUcrMEtPBUII5gp8iDxmTvjH2lyVlo0kE
clcn+7gkM8Cw2lbuxJvH/ejmYrSpNlMUyUinnEcbbv+oavIekVhdEvCj6Ce3sZQcNhQcue2KroDZ
AjFoJ0U0Vg521RTPzVRjlyOYoa1ujVQREeBQvzaaO1PqABNO6/xwyoJvttlqoyqs5srQfn5smtXF
JUrR1fa3SE8drmHy9OPU9Mm9aMNY6m8wFK/Q1bCSqRHTh2uwKXSaWxOWt4vvfmOD6R1reXbhg1Hj
3Ayr6GuGvtGQBkATdP1Nuf2igIfy6z/hC9uOSn9JrtbE7ysLnxE1aPYHSmqQXtoMDguhn5EOnFgX
fgJApB3wucUKtDe9FSFyeOjL4DEnunMUy4aLLmFqSHkB6YdAFY0FiKXff8W4SB/EZLNQsYU1fPaD
9YsNcuz2wQgkFhZYTTLHvgSttaWGqvLOi/H23BaoCPhCGCVbGwoWleTi/97oau0yFUqItILXV/gK
4eog2kpBQWBhcpcvcEqcyerTfzHJzuyOghZCvD8mrAVmPm6UYnYI73FBoThKGWbAedKku5um41nE
otGCdX3VreUpwDvqb6PH5p72zY3pAqOnSgeGeAwZtQ2W6oBvL4isBS0pRiDLJswZmwFVljGDCwVh
WxsrKqFr7yNx1NnvingG1R0yP6NvpOKyXe8nN7nm+8LbrkZLADhsT3VxokhsOq8N3idF9EjK0gzT
ba5MgQK5dl+krbEgnrPCgs2iQQcdx+KenXsILSeug+EqpjUDVusEt2S3rvoULjCgNrb0HanvILp7
0SIvT1Ta/M6Ueiia92Nu/O3vUUFjm93b8uy6lABA/au2zONJSA4oQ0K1AgahnSX7UxRbqtZ6L5B4
A0a4MdBXENOsqEyXWk2C9zWO/gfIGuEs34LC+Le334EPvWzd3j/YHpkOhPWHaeXeNEhLlyfMO0Tq
aUiFi6JCTiC31zZgGJ+oU6BaTk0mnFyCa9AZ5rq8tsNQ1LKKiagJAlF6kcIf/o2is+2h97HdzoKE
jxnTE8blANGF1okLKvohL6zBJYes8ZfcM8B7A4ivG+5gD+pGwsVD8fU2Yiqi5r/5oY39w1rBJdXp
570KQPonSfHoBHlvtuXh7swHOA9y+0nMzPo6nDt5j3mjGq2NnXIdG3hJ/rsCkKllAbpjGLbznfcO
FTMVdzGSsbJOs9w06uoTDBrBciqBGFw6d/QbZYiMKLYenYTF/jkh03xjd6sOFfQHlhUdseEoOO5w
ekopWZRSU06fkzRTxVyv807d0ggw9eM7JWA+uDQpERJy3B9kj86QzURt+hmrx/qPq0tH4vOuzykM
epxZiol5N5vJFycDpdQG0OFDwlmn+mHRFs5eCjlcQongjYaJXwVwTJGRQImkpYhdrxYEP22/CRbS
K/wOGCLBnMRE/mOAOMnvVKe7+eMVcRVHFJeTvlVa7u/DsWDO2My4k9/PBcLAMTQXZWFQFnPwCHv7
tTIVWC4ys53ut4nLlWeZ1H72IJ2k11EkJ0yxuQo4SW/BgJvzw8EpPbLdUBAnKZqpNpMv+Lq7Trmu
YWI3MondnjaW4F/44RaFKSu1jTHb57mufotUWICyJFLdPaI/+lkbLSx1zEu4LzIoDY/pxUO3Zf6f
zc/uJvQEsio/oWDCwyCj/Zw4whLv8x62sCEC9EaXrUkILv+2NwRKtWzeBRXcEqUKp8QWvgOGYCmj
R+Cy+MLuMbNURR0GJ8JtVM3lhQ8c83b+GBFMwNZkcCa0E20TGrIB225mvzvBYAluoDDS0IEaf5ZN
jDchkwHNSMvapTqDPS08UILGAk2alToiLZhGMs4z1xD9bV+59qBFyMT+g/JNX6nrFJBun9Rz+3z3
+b3pF6lcbKS+4i0vo1fJshXgQoGl4zKXxC4esBuWlPP7VtHP8X/pSfcYkm3M14sclTMrw+xmJ7X+
s52dcXuQeiPNV4+bbeCfaHAkKVIOQk20QwS5FgZ3EDg2iJ6o9v8jXt4F8sAzG4hL1sQjNL4DDoV+
MdtOPxDVTViTM7EdgjVK75l9v8L6xO0Z9+jlp9mcM7V10hhjnLc1Y6tdcCIi1vQdga0Ra8teWCiI
BR9EU/5ScTuka+vqSP7njwIfX3nmq4ZVIgTLRBQj7yiz/AR1G21q/JHLNNNEx/+mXfmt6XZYZuUa
0sFbS7Ut4uNmUNjO6qA3UtEPkSNf1lrqqQKYDi6EXG68hA4GFqoguAWqY0UXziC+k9l6S8UGlYAD
TTmEKaHlG6eaAn5S+MLGCW4qwyJkfEu+hDvjKNdEPFXMq9KhKRRk+UD1VUwpQLbkUbg3zV1urw9k
pQi5Mc7zJkfw6jOZxvUcpN88uZt0aCf2lMQy4F35xD0XSez3Qr7+MUmAXXEJN4A3i4YNiLYoF2aW
yAPH4O9OCdsTFhXom0uTO3kJdXZeT2OyHJj2NALA2Ou89v/fkoaAYi7gRDUTz36PlQC4gYIxASEa
UxIhlnLHmWbyp/NWYBeFKCGn4I9G9iLHlzu+VOzgJNIAbh8k1xCCwWIeKUcMoE6u/B+Pmm6CdGnv
HxPfoS9RZ72iiTxGEPYEcovbZgkf6HwZScjrmYAOCDhoJjTFdTd5+sXruqNFPTqJvxUkPR5TeWim
m8lzyRhhfDGYpmvFW/2dNV2ZA4YU4PuhhPyB2O4QkUmvYibIhZpRJsiINQqiV4oWoi4J16v8Llbj
rhy4QyZ8dlT/0OPUxW6+Wk2/POKJVDZAAbGNuXHgceIRKBQparkm6EuC0Ke8Kwo540RbwCwgpPu5
4Z5Pv+BuJXGrkVgBgJqd921azPJQO8SxfQnHmgbiQbuffKh5evuYBMmV6Yse9cIM2TY4SMBzlMR/
GpnV4ukrJOr4z3Hm0ghUMt4uLGo+EK/zBZMly5x8ryb9vKTV1lNlXrzULqgndcASyC7dp0dUjab5
e/C8MYxMc0G2GBrMaxF8o5agxYGQw7PRp5U+cK3cwu5LPIRFSvpLh5m3PjOTPRccr/y8tGpbaIAL
MypdGJ7MBL7vGukSOa6DyB2Ca2e2lLb8bCWJsbtrjbOnNGptLqcshOgh22uZcuhsTlBSg0dMP8o0
Y/uLvi2kVePAi2cXQsHWYg8an6HMkdIfHHUhuTD/JQAEiOu8FbOkCPMpDLTaWcwbc8pO85wt4SkA
6aN7NQTePZlzLe6sg+BoE0FGjzGmi39iOAcKbHuBRdl2O5ih3oXUAdN7mXHtwiaflommAhWpMbBa
7c3KQUICj0o2c0Cp5YwD7prn9JpgNoT4c0pzViybtOu7hjccBnNlioAG7PMkwVOIcBSEMKv+UYd7
W8+BO2o6bW5/Po5ZemyPilTOhZLBIUMOxJgZfBBSO+3AhPjDxuktciCyYCeZ5Z4RNPui3ZhQuRa6
91PGH66Kh5/tbRBrF6RKzpm+6UTcs49SDY6Hu63/zGt6qKqjepwRYeppq/uDiwwqNJprMC2ISf4q
Rt1yGPu1U1Kk4dRhIaF+7lSQVE/hqcatIxHuqzivcrj+cYVakaHudeaPWT8riaTLEbGPTffSZKg+
kwsrHmWoOS6C0wKdmQ9uM8hwdjUhjb9oqHEU32bW/bzsHnoPzqoWenGUh0N4JOfyqRKm38ia8HE5
16p59gmFpylgMnrtm4UGJjsKlLFhSoSFmXwp2aDcH+8bmZf7WL0Zjj6O9Mgfm/Ip4zaqLSzSGkfd
sgw1Gr04d/w7NdGlV3kSJjUp3ulkaYyjRSjiJHmIQlAJk05lLnc66/MAtXWx4w8bIuM4yZOfnUJO
cwCl8MnAPkejlf981I4CwE8Q3c4io340k1pL7aeIBq92E79gRDZllJrT3fzVdqVs8VbRseNLRd42
UY5rgKWI6ow0AAeUUKn+YPYYM1B/eE0cG2F1uopV8MIXf6KsSTuHWDdXgb2hcrG1cAmdrpNZlyTV
zbAjtRd813DFw9aJNOM2jl9O7ZAxn82Q00BNfoCq1B6NMZMEZTo/o9QEHYxEhXhd9Sg7EEG8lJ6T
7Q9WEN6qWu5Ogowolpe4yM9xjWfrNZZwM3LMWsRlZyEaIbSUrXi3N+xxPElp2pajuDmcjRbsa8nc
R/MFTyHsa/BipE3lowU1xxRIMP0ItTSIy54k9Z7Iog/jndcebUcRLp3HGhRN9YdQxYVX/wxve25E
xPEKgx4VCVqRS01NLQqAeO5o59LNAEUQ61Hs6bWu/bdbzYEGTfC4TENlSIGx1Le0FrdIfR1EUovF
VO8J3cFmNid0YcIJFnBTYITLTQeTBOOftgHCLfmyejLsclppJo6enA6mSCxlUbJMn9oQ75cVwJO9
5uVym5txPz9qkUZXlyAXHE3QPnUl32/Ld87ypvDottoAGgRHM+rt5FfFMsksIZ3HqaGVt604Xo6o
8wLEm/Bakf/GAAO/oI4gmZv57QExjrn3uw8C6Bt3+JUysHZ6J3s9I+FbclZ6nSsn6TEdcU4diWKn
0SneZisMqmy75lFx4qjuUcarpmxcJTLanxGTFfebWWGg+h+axQVx9Qi3Phbqn3dJkLllJbW2wMA3
fE3u2heMNpJe2APB119E1O8Q8A2d+qY2W6Yrql6nocVc8V/1NRswxpsEuLV/FGmWAFYh3utB6bbS
IbX8x2T5t2WXqnZKSDMW6AaopVRV1IA09Uusv61F6/h+g6mTdZCcT2kJe9XTEJeUAK6Idrv3/2+G
gY073Y90xjwWPejQ3zKVZUCkAKPBQrNnXTLEgAcEpXVHUy+WIB1DBCVwTJBZsIzE9ACg2UzXtB/8
t6K99rZ6Ulj/ifpo6W74G4skCJoxaJtO74IRZl8E7zR/r1kyrfCQD8MnapBgcCrkwjP536rFV9mU
4n1/EXNFwL+UzrJUS4EWakE2ci24jgkBeLneQ6ye7X1ONhQzjo1RTFjjXSIu1GMuuiGgCDROP0tp
4jGS03WMcXDh6UNpJrmSuurO3pI7Cjz+DVYckhTZCH9YPHjjUF10kfe1A5dYL1sWFPJNwOvJK5Y6
oGrmXIpKkmSbRqWX80h9vfIzNZVOd237vcgwOc8WGx1tt0vLiT903MtLIhRNwzOIlE/XnYP7rdIy
5YO+EAJQwlMBWdNJhA+wqCwTB339vGtZmSHgj2djM7VnY77ZTBRr6Y1tLa+muov80SnHiviKdTM/
E2EBN0cX222xNsnmlcQwdkjCiMmPjuUT1B4vyJwQiRlc0ZIVA9BqidqORwtpOi+qc9Lfs/eKyU3X
Q96GazSRyZYvm3+WFbRipfiJKDggPrSKLSU2iQsJNuTgxVTeuguqdsKRG5dgTWTratF8ELijTNT+
HfGJ98Ij0SbPLjBjduniu0Zya24jnRekiPrNF396DG53B3IUtp/oJvT63At2QlobupU91Ek0F+Xy
3ZphK8N+cmrUYtxvmxNrO5sbCIyMv9ZvuvlSoO9X4feb2SFagbBgyCtqk9GOohogLHt3G0xQAC1v
3lLjCOCgx0QB56oJSvVKBjQgYTks3qP1VfIaX3EtqhhCfFtyxB9EQGpocSULKoic5hbCLoS64W0m
WkvBgmfr8o7Cm/4i4L3a/iZehxRFblgoXmQaMdgzSD+bkBgEYSaK10xF+8fhEXKWytPCN14ZoEuT
haI77NQsEwN3Y6c6zh0yrN5yp46zkOJIH76mHccQr/ClczaBfUJsG3shsVvYVT+zW3UBsUiF3AfG
M5jguyt/joxqX+miXEPYkmDoKeOeqXRkp2HKHFot9GvC3jZUFKCvhv3+1I26drw1mIr+fjTGI82H
QrnFpqxVf1PHmgPK4YhIUlxMRjo3YngzQ5pgLgfghCO4rmP1k1mNn1FJ47MJp3N88g27gkRIZpv/
UaTM/Zy/qWW/KpEfWejWgl29MAqokSdBlxpM7rk+3Qiv94+iFxWRu4VMTphniAzimjuwwYQ7usDB
jKX4w9iAeBn3EFxW4rn3EArkVb0BUvmtQBQCAWhVxfjrFW2fiRaW/fkTZDSP+ETOehda7Elyq05J
NUQT0yvKvLpZW1o7wlqe7GIeFyAzbsdzgiQZZdI97vd8WrXHSE9CPwfkt8Rf1+gM181+/Ev1vQUn
uh8+JtQPnpnLILxEw+rxxnNiNUuyvr+g6Moj1HUeu/J0iUfSkxC0ovoBvnr4FVWrWECF45W/Kv/C
eDG5UoAsoO8QOcM3zsCsexDAo5kVsd1IDbLCFzi4hOFks/K9pA99yNexQKt0uBf/o72057mRJ5yF
fnb5quhwEFQSUah+Z1sj0545rhjCjcSPNJRkWYkpHyrm8C1fOyQS7EBhKnm0jB1PZkyHGMs/Ew+8
gL3+FYx2gdakr4FI8TT76vHytCAaVUJW6v4+vZxIX66/pqrd9VmCWQMIE4dwv3dsSlP7uFHledvP
++g2WKymoJaXGHMfjYchjvJQlFRpCOhOf74hmA2TotHmZOou72bWgNz6jJIVQ1owsGOF8fqibAAB
A0r6Q7Z2mAZOBCK65lFtyisQswT/11A6qCHJblUk3XpJe/Lxy9v/363/4u56GV5dLz+Soip4kU8a
UcETfS8c6Yj1l3utk7dDmEawYR5d92sSZ3iG6k48RYoruTX5faVtJb3u6wEnG0jBr+YTeA6WaZEm
HPZ1JyDoyfNvkCIACWj/lIWjnC9Ck4jsHyQMXVUGn6JPr1e+7ai0NJaiX+I43PpRN8hkfb6dKmsQ
BpEZGv79uccufpes4o8NbvRPBaTvkmZYI0yZSuaFiCyv4JTm54v/RerEjq7FV7zfja/YSPKBRY/V
K8BuEsXnxmhItCwWZKw/1Z6b+NlfE+xSOeYlhUNceinO0qStEAdRcQR/cmUVoGDjfbvxtQfnT1qj
bfiZ14HeEj2tgeuTXjpYb5tgMych4PCftP6qAmaFsKPOf17yCfMUIjM4/0wMS9rA5v6ZRnd3woj7
RAVw6gjl9iOa+1L57VG8IEoTvbxBI2F94+AHBlpHBABt49B5oagniQ+H/aVNcYBM8EiLB4bO2thz
ZgxB1dTr5QVGINFqYhqy1M1PUsVnJ6dwdtoDDT1kK6dq1SPIelD042W4HyN2vHTCzJHXe0s0teGb
CKJkKNd2paEJ+eGQI+4pX3voDVXPWJ3ub+xUcOh4IlZkACRXopZGf06FjKHJ83+u0bGhFdLbKP2j
C1qqXXt3IDZt9C4Izm3JgFE4w6y+YNp/Ar4EDDVOY65jN557zs688OEVGhF/vOdaZglPmDPtRTY9
VTjBqgD0Wmry2RoJAI1cdXFKIowvFM0q8NGXDa9XW6vfY1cbQe66sNeXNAeP3rNNgJmnctBtzxHg
TEYdBDpwgf6P+oDyUIiMV0r7Y2XdEU1Uj52a8227pYDAodNbnHXoY15oxN3qcY7ZqEewmD7s5/6o
9vZYYkTxXeKV747PmXMkPYQgdz1xYdYC0aRSprCVGTLRZoNmrMaEeVP7CqTz2FUcqNBT0vyI42k8
ZjlizLjc/H8J2wb7t4XxoO2d3oA7xUtmJgNLnM4domrYUTa5f7aIE5EeaB5/BlItyiTVb9mS8lbK
2KbDMxySE410wEzXiY7ItGWp278AVYsvmIM3G3PMTTqGwnx+oHRWcBIsw/fzlcnzCQJEMAtyD5NZ
mOyXlLgzHmwbPrtjWGnWm2yU1E7HBKdZWOKv1Ab+iVbLcKRZeCIzNgYyXhVJRbaxfuBe9ILYVasf
Fqj3GWepAJT8rqjg1F0qJEkzGUDXmSRvcy4dOV9URJjIB7umi+V61Flud61pLOdhYeQrilcnJZQx
vq4CLL11RSQJjSi/l8i54fZr1KSFoFNo6cuzxLCjl9/vy9X2rHhRfk/QVQJCl6lNYML0WzWF+zjs
vVRb5Lr+i5VLHBU43mwM9G0SDiEQPaXGzMwbOTsRFg6NLcuqY73WFm2M/h3eFK+70k4rbVc0+cY5
N7wjYv+0UUE33mO4Xl/JP/IVo+yZNPjsCMQnvp0N93kOkk/5pRNJoAqZgBfbFnAyqO8U5hZAZAWy
hTGciFA7hYj3RaWD0UQSd2p6dw1551HreOdRi3eZOsejUg6BuYsCw58PSKw1tMRAUIelOyiKFkkm
NXBtFDZW3Os4QbI3stQq1QE1h/vtmFGzfUAuWHprg8QbpOe77b4Lgbp3eqngnOWX65klrObyEJa2
WRmAuQMWdzhp5U7MkD1i7Rz20j6kDBGeuwnRPbT2nuRSu+Pz/ftcNiCcmgj6EoTEBl4JZ6WmGe1a
jCi27HPA/O2Pt1amtjxhBpkdsMl8EEF35IoRT9RqLyUxBp3XRF1SAdoonaYTfidj5+1GSJvWYSNp
gybe//Rvo1GgEfHRi5XxcNICd/ywYxUEaDpJIU2IjVtxfYYfqgT8xyCuLmu6epx/4+dTlcW3xWZj
EbKhjHLME/+BT3vfYFTPFCQopomHXJc7YDQJP4NlOx0fhk/gBFBsGMerZD74CFiTa8cPRuGJVpXU
1zo63V2p7Nn1+zS+IE3V3ua3y5+BtpyciLSRitlzymE5rvIYuSH/5MJvyh7NI8IBolJ4QRg8B1+Y
wNniSDZydDO9+idA4mWXkJOH5SacZCpYAYNLM0W4pjQ2KVHe9ce/4LxPrrR6T1hqjML9X0vvWQpw
UAbFs9Cx7F55lFGZU66bSGtVjYcBk8qLVtTQgy9eica/xCeSudmFv6oqCnfTqu94RHFGjtYTklQV
wuyIY65E9mEJB9rXtzII0ECGUc2iK8dacYHzO1WAU3/T1hcr9GB6oGoUZasATM2NW0YS7zaYfxNB
CX4vn4nPUVxvpEXyJ8Vx8L9KdTYvtTR7zh3xVM8UI77RRTQhsGkqUc2RDqHDH/0UFqn0UUNHT3uf
E/zvy1XG2M/yzPVPRiF+iJQb6E1p7Yp77QBVD3C6cQchf28O9pAcFzQpvQFxDocjujKzP6JEtE/w
XI3IL7dRkPJovdcjIOBPuswmC5ETmyeZORiU/Uz2I6tjtZKTiBiaGgyKVPCCo2E3xlvZY5aFPqve
apj6ps9EOmyKfLs8rrjlSgJE6thMr5H7UaWNEhYTVI95PxVVgptMp8OrVnEArg35mo1g7X2xQDbe
gXHlBxdmN9f+en5SsXBNTI2zJz4sIVWNMikdEBjIQbiuUxF23AYq2LFvqTck9eqX0aEIzTll0piP
wbJoRcqOtTWiIJBSqHcOxR7EsGdWMBrq1k2z4HxylkZm0tCusklqEcWko5l59L8F6Hwgd5FaIKdm
FwyoEAlZyR8+fWWbZHaaixaTiPozR2s/dT7D3Un+xvvQmEjoONiBodtINDziD6/fDff+DfjiB5NO
g2+02voHwzRF/FwlWprPntVlE6v45H2aJksRgoT0OYozMq/QJn0WDu0IhqKy4jgjpH4uW0/emP/f
DVmqFrDCPLAekVgPTGz/LHCfNqSYyX5VnK/p6JG7hak9zFYRcDMM5AK0x4ByBjO3Mzr02tnZ7aYK
Zk+Hx5btbJoPrhNUfYlwIS0gQiU9T4zzkGLdMzRXF4AzFA1pbhmBCiFZIJGz61d3alCMllLKvoph
OMzh819+9y4NpMpXfkAuo4ShgFRV5z3vmGFKQ9ICZrHuk/M6Kh3gjIliOWNbVtBHhVRy6vAEqRvW
6+sxEc282JN94ek4KIe8aMFHay1+wQvcAN/mfQjMF4qWmtWTFoO+htoaWZ/Gip9b0VvUVFGDWWvd
KnPnIWSrd5y64AHUe7sQxruSMKxf0PJuk/+UxnMr/3oZJ9+aoQbGgKNEGIQqQSW67XoT4cidTqQc
qxt48DzKNCkElbaNdNlzn0ewB0TU36lze8FwIdmTsSreupV7vx4Pk5hVurShet4BsVuQDXPJR9dJ
Frto1gCsudqNLwzK0STEjyNldosI/8FnV2P1wiAc/YWjLFGx53mT3bMlRkLOO6S/eFDHBWUp+Ixm
Be7gFC/0b8QWmw9qQ7JRLuVySXZTCIftVtAHVTv+NNgM/Cyj8lMN/+7qtwclQJsXchxZU6J+E1IE
ryI5g/1Zq5pEb2n0fLJyKIYXG70MrbvZFyXqLl7KtgnFA7XYrM13ChTtvGRlhIf3OtgqpANCj5Vo
ba+ikMaLnr45ZpeniXMtOvM1YNgI/2hBlKSJyZ5kL2RVmBInfr1CgoVZo4X1WdD3h9ARHAQqqMHI
4qiiqw1zOvWnXglm4s4pJpiemvs00Ri8Mrtk+tJ6wkNedeDM/RiQ63XhLj02Nx+UYfgxb5QegenJ
PQPd3CjpMcpDEabzobWPE4nF6vzjhBdxrJYjX+GrdGO/AvmTZ6wT/V+LOB4njy7fq5G0LojSmJR8
Alxi2xMDALMKn0NHeuXB+eLOt2mTVx7RhmOT6Xahz13/6ZUhQdcKMhsoK7TNNzeStBecVAVTSVWJ
pvCX8Ytw3RlZdMglp1YpiO22kqsuWhXpdhoNgcHK3CWizcrfApG7kpP/JbpmOxEQN+dZFj7aYOjT
1LTy1UVhmQhuwxUcyUQtH+LAr6jzEHfSquzvbAz29vmtTlQ3c01GMaJrnU0/+BbrN4HsQasKFJkE
EXNi6boMOClbHpFyo6aWIfpQI8kifmq5BGNwrgxmWVnSSlMKLrvgp4nziIeUV5lfiJm8dBjouBtw
qWEQdh/9/ANb/cRroIBvPzAt9c/sXfC4JoK8l6lfsK8wc68RY1ylOO+qdFKg5quw6LX1gzMmFek0
yDe9XayXBGV+94yQBRVTHvNVKoV1W/TjoGpVupoxoa9AnFRIOOCJIsW9PtdLopfd9C+IN1X0+4dj
YzV0s7IABk2gXW7XXgi9esmvNM5X3m2XrxVgANPt5ozguOLnQiJcF8cYhMByV69lVuaHNhoWayJY
aTFlhXOdnN6bOuxAdjkYYMBHw9lHCgyz8tTjc/MlcTfPoN1NzO63Lg+fLwkFokAG4vZ18tI7ejD1
ePhtDwx31ap97uf1o+Z09tabQMGmg2p6b3HA5MLCMSGXBN/SQ1plc7HsgUwsVdwJte7ek+YgSAc0
LC6CrO2R211J26e9DGof5CusOfgCrvJWPEmaH2t5txzrQAXNGz5PZViU+2cpBC+Lh6r2j85J03yK
qeqFv00xfcSjyG09OpAVdfflzhAWays6j2I7A2Q/dUX+9bFjPtSi+2H5W5Ev/Ri8eQFyoJKs10uC
49xvyeCia9HrGR4vlKMbPFFUxhEH1+3pa2nJ4GwqqSKJFIiYMPhSqymS/Xn8JBWAQDYlv+4f/nbs
S6rnkCxZ2wWyX+BEUd/IgWmI8jDyZFzVYkyK4Y+KNB+Je+aZtZioD6APOF4XJ6odsbidGSZzp9VS
Os0Y20rSfRzIv5wy1+TFgQbzDO7RRgWIOhUWX52LRj/RjLwoCdL+lWl876ijMHCgDXAF1TUpGaLk
0hiv8tnYGbhZRSRkyAbBa7s89xfRrDQwjwgwv+RYlX5z1B3VHIsrvDFLJEct+pQaUbGVa0goajVE
ZCohxZrjJy5KrHb/dVzrEMVB1cogk3dpOuQcuoz0VjZPmcJUo+g4Q189ebAcOTcOUANyJD91H+y2
NgBIf6frDZCkFIpKKjzPCcVQMAS08FD/lm43gkLXXaixynyzdHde4H3djMBaV+KPKfMWSJ571rud
1NMpprpx+VLHI80v04OWeLjrVuZBGausdeA9M7PhOJkyDsH0pKFj9alV5enpcQfyoW44NkVXIL+P
IDx6n03KpLbzauC1jid3Tb14Zwt/jGSYb1+zV0O9PtXDHqepjEohCQVVhkbtTbc46A3rYJaBp+RT
A0UrsYX08hQzIEdX/9HptlDTBmPGF+Qw6iMjxPCLrzdLOMX1FBPkXLAp5WVIeUPLgqVH0kAfXJku
TNCLm40ZHhx6H+Gd+ynV43M46cdIfJWciF4s5iv5MwXELkmBy90yhPt0MAAxrmYyGt9VlTxou/R4
8jQgWPVnB68KIqaFNEiNF+Opti6uTBQQvWB6CM6yMwaYeVOYoqlxBbwN3OlEhc9wnSOlw37G7to1
J3OpU8kJksSxSFtKQZkgxfMcIQSJ+xXeMreakPi0ttkzQrkim2t1rsx7ydKIp3G67PZy+izqP+z2
iYJnyLQhqkkXMGOzIdXXYS8YT0q1JrUeUd9okirkhBBk5Mglv9rreGEhWGp3HFOvAp+rwrsvntML
rx4uTXvmV6LxjrTfd2Qu/V8rFUnxTlhd9Bv8DmV/zBEUCJ1wVPRilXGnLixFFwJWKR9KAyMQLVXV
ZWLLScTZ9kUBCCZTX27qY+O4WbR8Xqh+U5EsxD9E7jSFhDQAZuLlAkmmH2HdT7exy8JSFQtoAKBC
3PRdpysZb73Dx79N9GaSZV50i1isahLGKwL1CNb+lhy5cxq53+LkY16pddpNTeCQ2pe0y07r47ll
vKmHBw5GZ9fGEgzjcWHcIz87SOb/Y6jwqAz6KbW+xFYaowYqKnTgbWKj0zL6BqipFPgvAyw3CttI
GQo26pXC1eqOTVT87sgRzf+SDHbJce1Z4wrILVTiIADu9ORZ/kF16pQRLWz0ZjV0wwC0NvjE7/s1
sCtNEvUy1vwQFEp0LJGwgLDloZdiP7SY+EHC6uABOlqGpA3ZMt+nV8I3PX7WGjOIhG2DoIacenJ+
rFMB9WJKLL1OX5/E7Z4XuPWO6J1y3Y4nniDMerw7GfHw8lNQi0nQGrV5sCXLwhztIHTKpilDFmba
kl7B52F1s+X7OK5lkBFFB2CYjyD2G7fQl7E1LfhKlyq/cMl2zRukq95AfbAlXqBdkl2V6Oa3+1wh
FyTwksZYiQInnFShqoobKXJy39k7G4BPN2wQ6bbJY1GlFNZkfsMG6N39Uiszemv+iy3oj7nLfVkO
/QZzxuDOad10MSVu09sGT3COUhCLFOFiuJ9v5tPsU4ftCW+84MxPcmUp8bV0SW7dh+8wOHPjqZbf
zdXtmleT0uu3ADaDXm2LB2asQNRdQ4YZgXDDhw3WawrhxDIvxL+WYNU3TvjhFopKOgjC0n2thg1y
7K7tiiYDAIA3gqNM53UXPXJZdle9PBGWKlzj1g7abOYhSaX/PfJmApiUkaHm9391+uBotS0aYauj
yp/bcZW3oYmpShQ1YqEzmsaFhejWE7qTNp7doOFaPUyxE/E5W1YS5bOfnsYeN//E36cL2T+B3nKP
Q2e4myJJ0gZ2X4t34ZO9ZtSjC4a9LAmLz/XxiGo7ooBjp5yNryYnEZ9h6QHnmpb8dz17QalAyma+
4Qlz13H/nC6gfBVjvk6nK48bxY7m2RSSCCmROAx1x20bRJrx95FYSp8nxTPwhBoSqS39TBQI4+Ta
RgEBAGyDcAHSVzCQBGOL3yH6eSm8UxY+6Wp79RQTG9q54KEvqFUomAo38r5kD+LODrEGYaoN3Pp/
/3mRl89DhtoxP6nwzHrxhRKOQN7SwSa8fZzyAe5w4hAQ1K/bzTZeS/ZCn09soiccweTpVhcDaxbu
k07X06NXdvZFtvAlb9PI7LbS9JQjTN/EhMUt5FdhCziwt83dFKDgvUxZ3aBuNicrrvvzQPiUwYRV
RR+A3B/hdanhkDrBty1PUCcW5M0zJNrdZ4QiMlCsrZxffcYctDI7zTLOXl9Ie0dzElY9+d7+AlZ7
pMJZKLI21V7Ppuk181Np8lA98taIsuarczTRD8PApebGrAQRQ34wiGlVJS9/t0Vy6TL8ZtXiBQ4W
+z5yUmJZez60XyhV/lrk+rOkZ8Lp/gM5FCIXXCqtthxcOO1rp/D1mZnkRS9S70120dHnoBoBSpZf
UtECLRfaOK2lwWEH874YjNmsFpuc8rIVjJvIh0+KDgtWdNJfAmUIMtpFsgCEyLiEnXhBeKE9c4b1
sE5NWaFbl7Kz2lTtZj+lNJWi7rZkAgigo42YZbxRCDIXsUogu9aD+oVIY9gyJKn7zyZrB1E+qPa4
iua3ZPQJNDO2GSHim3G5UhwWi9bCOFnNseK2oh+IjMfH/XUUKJc8HQzd4WJ9eqm44pdflXaJkpgs
6ZZ514RudsoHgxIbFOMAMcp++7Ut9iMxQk+j8GgKFTe+PfUdprXahOLXZQ8QonMt8iKNBaGb0dYo
bec8pPeidI4erO8LhIRJo3U7ZneG8FYpVHCO+BiDi1auX+iVOZGIq0NxSYNBrOxT6wlHBaupuqsi
Z53Ha2bTLSvcp5RBXjFPFMxVMxKhwhdB9a+ZTSHSfuCH76LvBYFCeZe50ayZB7/x69T+rdfmTTpT
Be6aal9kqHKVkLEC+THHGTJ2kNv7ZTc+MC95olapQ5Jim1B4cn91xbY9JSxFjy0/c7w2VqlyHICn
g1VIRGi0SdfrVE+cOjN4IHndshmXM/dQQG0S/GBXIyCezNK1mU8F5EmCYM4OUi/xLOkmX96FCOtM
+hCjfQY5931585DImB6aje9Efp4dZEMCS0L1L+PUfO6XKz4cLoxtRMqFOd+O3SKrwuMwAOV5HiJ0
DtvD3JG6DdZ/oAxompLcpZSNB2unpLmYB4UzRMnVIGMC9TEJc+KhWFRxUXLg4WTQQgemYfT8mJ/Y
qqv4WMT6xM5NXvAlA/D1I4B1oklaIrZU267vhZlcDyulrPmQb1vITXtOk+e15hLcD7RfhWUc1SwE
Rt6umQa+Ft1GXKKfBYksyU6ZI41rDagZrBqXwJwhQc8O7xxnQZveW5NPWd/HP55p91GierrbU9uj
W2grvtXzKD8MAxIPQ5R6Yh2kcKOKhPpgmG9FnGnxDm+kfqtNUwOh/KcEQv0k2u4qTxJFfPvUpm7x
Q4d+EcsA+rLpC5Do4905daEIAv4/IOW8Iqgk1jcO0a9vZzZ5b5ZYVgkJrf1nI1dfEwqt8rgfPBtZ
pa5ejCpsCNfOJ3cMYRMqH9Cjmga4vbNP1XffPWGpQzI+dz3VA8oZtyIdott9lYtUZpLcNNfW3RK0
r3GAd37YBlskpmkq6Pq1iQm6h21apu4fanXiMiFyzxLcWzL8OWrkF6SIhXSUakDw8J8ROhZt4RNe
QCXSef2TW1G1If0DxgOWSg0am4dQwUxv7dfCH2pet0aB6GFUXbBGjlXbt+OC8z9C+nVDzUs7RVlc
LWwz9ccwPZ0IvawhjRSue34IRsx2kth5PRIP/zNZZX7XFOskoQuoSGhZ7/fqKVx7NLgI7lAbMTYk
oYvUakjCb4NPRDyDrVuCA2k6+GfYmvqDD1YHUNO0G7c8urcm7cVW4kVcmQqTvsz/vse8cwg45NvF
wgAysQedEhofTsRjVBsCNkeJnWVu5fIlvYu0tgjlNzzQX+ZD/sC1ZCXvEXv6CqYWSlp7q660dAk+
DkYiONmNtpe2WFfOgSE+YfwW252doX2hF4DMmq1UeqO3cBOT2zh3vYGaYNrOj7wj8bU9YnaJ5Skw
EjypSOVY6GrZ8PVsevtE04L8SAIIAPebMmwZE0XOVDBRfCyo9tsi29+DqZ1Jgxv0//YOrC8PN88z
tEOjEZWpMxYR2UsDIFypIj6TMGgchC553zBh/83J7cbS5Y3giJzrWzjR2gn6udmYXb6MRCq8UMTr
lppLt2UhGbupL77DK8Dw4MAQDMq2de4FqHphtrHumJcUxjLaIf0xzVhzVW9IZbRQLBHE6k8QY/D6
2P0Xr06VbXtLwsMlCcOfGqdkTO0HMfpcM3GRSRvtnfSYaSw0O54tSA4ZV/mHTraGsTtK6T5F3s9n
uyR8TCgJ9DHPQUwaW3Spzqd7wLzgPfsUqrm/pJEE7Ysvvm//4aHGepgPywW2R/eghUHK/I76GqEg
GyDS9HRmB4pRHCogpt55z+Fl+fiZdgyqVr6z/AHJtyQ4zMdpnu2838WuHd5E3MMXvQdR62YSSAGV
BN1T4HaiWBbLkdoIi9K1wCSBEOJzMCjX/RhyYNUn/Q8S8MCTrNllxCXCVCwHRSZyfE7anN2j5smR
Odt/Wgn4RRk4evd+qj7UVeGL80iQD2gHLKLHqSEojpKNV8A4rwA2kJqB3N161lB6X63hVGEIlMCc
Px3oAAE8jXIvqZrZ2neZ2HdsqewjlPvJ9Gz8s2d8g0ZgFufWa/9DJLD7SIngPU/BwZ/b7VpyHv4c
NM9lW1Vk4nu5ujhoGYCpDzGdNE5ZTOzZSjE93/BzwOajTc/iiG7i8UsU2OMOI4rvptsuvTy37QSo
PapyH6hFXT3hEIJZr4Du+LJkFrEE9YDf+JKM/DQdTogQGC1HiFCtaCzQUxIrNHskEDMkSZ3I7V1L
16MPt93+x3CNQptQuyF1R+HI5pmpgL7uueGk3L0JvBckXzfxsyX8MfFofCtwy8CCJTDMhB8nj1YE
mv0KzFmpLyq1oMEB86UfrY5M7go8M03HWL3EHqwLw+66/FeUsDehRG+vyx8gLuOBohmRDByJ2qzl
aMw9qIsV/M5HbsQMIeK9Z2WPWHNr+VDpyJjOFa44OguMe2a9PdySg7+7anut58H18vfZomSBOJ3c
uQnbizdCtw1SD6LtQ7pNrrn1XG/w6CjY8ao6pP4hdPpreSBpLihnmeB3VRfJadNuXil76TqSNvPL
MHayUeRXiYDMAMDbsTAiVLMMiRQ6VkJ+taQGGxw/fzyT/vD5ghJXXDxxqWNFbZ4XtklZErr7bcsS
20Av2FoyGmbjHF81xX7hhKBMP289lyszxDo4HTOlx0SD8qBwEcvSS7zx+87GRSBStEUZdUPCSm3M
K3XgTRDLtRlpeYIHSZeOCuDwGWHcAPNj7wVMw1rJMFp8GEWfwyRMxHS1BKGEX+w0KSCFmjGI/uV1
tfIOam+90gM0GYsFnjv2PD65ppYoQBlLYsTU80q8/DcQKvIZvwcdaa2sVmvMuUAkHPFDqjFV1hC8
z4leB8kbrbuJVH3a2L1MlgzNoxq8ptnZ1io+iuC7BfLbzTbCC0mib+nCuC6t+bOjoVqv7WUWEZDn
sreCHqFlyGKNXE7BeF933PDbkQf9n26ZU8LDLLNR5srOxx9CMEzXYOz2Ojgo0IV7mAsLWAv2hS61
jCh9CfXk3M6zyLFeZmMpkqNHZRNlP1wwXCIc4djJYk8Uz5s+oy706nQ14B/Aq9zW8fVDn/VC/+rh
Jr1/uEHtUH9jMjDHBmmEy2xFn/VIOK7Isy5WKkVttacpPgWoichje0beIF+xhifvHlejTdkrnuaG
I9XZYU1Bqz/mTVqG+WLjaCox/hYxhD8QaoZnYgPDaA4z/wwO6lDyKWO3HcKw+c47w0sEikQfpZY0
xoTI9nWJqkveUuAxYQ4nOp3B2ZrdpiwW7CGY+DtdstUt2uwGhEA8HTJ3RBXeWDmlwfUDMXuaNA77
6rHVaPoX/ppqLdZwgVpqK6dNpsvwH7LO5e0fvHsPbAQVfl+5CcEaBTopadqpjQfgFmZBg7PCcwn1
6n59jiJTJZa22W/tHt/7N+RsK3QkISypA2ZU6Gr39nw+RrHNHzXT+SoOuCz/AqE511b+h0vfoTMi
eIs+T3W6eIiRZ9JTc7UTL1onzZgMSX73GIvpXoir7/mIiNW4X83xZs1zdw9PWArVDT/UjZKlmwD8
EQlJ3W8Zc07CXLvo8xELz5kZD81DtNjqOLcpL8hzGN8Nqux1eHjwRHiSmhE9S6XglOXEB2o8u9+t
Aot0+77Nr7H0Obmv2Ij6/t8lRhYE6eY301WtGHaZZmvyG6lQYN31FJcRvm2MWR4nF673gLqlOmp1
2yWE7XxR+n0V48ECoRi0Is2FXpBOjyh/f//8BcSmwD8K+y2p2Ke8Nj1j8aSXLpYLGG9DZsAoslj0
axUKdh3mrHH2S8e0Vj0DHpGrPHRm5VGjK+NBrGjbkwJNA0VkKblAfJttehqW8RQ/EAuSdPdN09xj
OXuuw7r/o2bDMYWDqxDND7Lgbfp6zaTvbkuQvHglPWxRRw10EVSqSfotoxF16Sk3ecME72O1Bu83
tzhlj75kqaJ7AMSSrH/D8mQgMdhk1IwfghfyZu6jSYwlEiHXFh6xCs+JYqDJJ3W5L8cCcqgkui3j
w1kybms/2KufAysDaGnFgJU0+UrStVKmC6fmBs7Vnwg87cWiqirxxtXA/otq4aMqQMsNJnslhURo
enwcpai9L2dAFtVdpRrfIR0ZZ06tdLC1y9Ewx8QCF1TCkVVq3Hn7uAmxK+j2wcc9fbdY0itod5bU
oM1QNRCnMJ8WEOURo3dVKKjY0izOuyilys8p5iwXnIrge59eoUFaYjpUZGrv5cXRkHb7+s7COJ0/
C7rsGvdqziQYkl5ME+ZTcMM6W0ls/T48JzIVNrDtA7ZhlVAjL+zPf+xkbvPC2b1q02X0OTrTrPXT
KTXOhMc1H8zXSdbDt4gGrbKX7kLfzQtCsbzhgUPH66BbNuYK5QoGyRo62FvdQ8w4PErm+SjMjQiT
0PMnLZ/+PXPj30tvv1HqVK0TZjKYmku3GdIihrMp97CoFsxmroOoZtclTzsVN5LpOsYcDwbpBgjf
332PM75u2eQwnz7ueJztR1LrBCSeMKxsQPmkmvD0F7rIF/qetPkQQ5YiougsHG4XPzZmM6x7ua1F
0b+aj1awTS8Q8hnoLs+xzTCrecR1JuopOku7jGxOx3ZP604eiR24EW9cpxjG44hCuyHQslDmWM0t
/HgiEEIYR7Rt1MqHpVb8yFubrYUvcLLnmpJt+7yLksHCBiGJlQ79+wuuX71EZtRBFAOdMsAK+Vva
RMj+L2Xdj1ipGKCR3baTSZZrHigHzO95Bt3XNOMfymyzLwpwVYjthYMijbJdv+69iZJ00GySbk0+
bGJ4YmN+KfDxQVMV79udnr+VD3p4cF8hfMXK43WN0BGtiOGjlPLGw+mte0pYw9Eayg+NzJ3MV2cJ
XzQYov0XiT80PrvSdxtpQzdXsckXtwTFtJzGN0uSqt82xUCFKzfm1A8GnRWk/aY/42JkxYM1/Onc
SMQMjTJC2BMBBj1GbOpEh7C5kWsD2bw/NDsc3eRXCZQ3VpUStBACVDlUZHvnucfBW+RvmKtD2rqs
sH/LkAMzVbE0EEhDeEhkQif3cFOsfiGBpO3rXDIg29nZ4LTjXzqsCFSyicH1VKfp8nIiMWaHz1c8
xyy8obh+coXhS90j7mJDu5ZlVIQxY9ebYF/Apudj7CMTW5qNDX7BGTZokc6KOJ5UW3Nh3OVi1013
KHelS2MqvxwGdBUGsvnrp5Ji9jE66JREaRCZdYfyxojGlcjpQLdBR36/vr8rbji8cTFmUg1WLt5Z
VcPA7u4cjHUzXIZq6vsw982s+KqTm6U0Yv8624IbgsSY0q8GhTVFE5F+bba0iZnSrWrS0lo91S71
iyzZ4nAWZg6EtImCzfz4imPai90U4X0JbGqBlZbXauPDSg1R08iIwTZ6eDz0tUcRX3z86b28K0/u
CM39/C99vvadNWoEZOyS7ygTWf43qpaFaJbrVEsq/7Mksp5Us3Wq/EGic792HFCmjdZ4gWJ3wkAN
J8MZNS7NIvPzNqWLZpKAG7P/rv1EEGB/mKa+WdO6quM355SBVaoDRPIH9xSKaUUtmUmE/3GHlmRF
Drey/4V1KPGFLVGzAGjk/0VtBpwp9pxKkz6IH/PqsIsh6YjwyZC6RtAwEQ7LPbTI6klgBBvdziSR
1VjoUtzoqMl36tjp68unjK5kA1ZTsaG9hlwcMiPEnz44fxLZuU2YxbT+uV88IrBmuH2gBVyqUMAG
r1rV0lg8OXnk+eQuQMDgZU+q/jZF675qFg0urvPkqfQNcHEJVlhpqAo+ieogxjESuSsAasUY3iXw
HzmBEZMHaee2kWemDip9AP4Mzv64shQZvqiNgTDwpLNVmWmve4OY7oqUB+nKZbyPvhAbdC7467t5
7pD783E8qX1mq51nD+WYISF6V/MLTRh0pQwXESv/btQMDAezslTjM1RFUw/VM91ReqJU9olQ7YcS
pyRKUJ1WKR4vdisruOGq+Gazt7eMD/h+3k24jv2XdJO0R4D1N0OaBVD6NgSpBcrSyZ0f0sWxa3Y/
ZNyYIJJCA82aNL60lqkzUJ67qAK+8aAHhJ3ZvaFcqIWQYWRAsyqVdbfWHp/Qtpt7UhVxEH7vD3/7
I11a/AH0K64JcGOb4OHc0DGVQ0l2kGbgt4fd7XzD6cequ0t6syxTOLLkfZRzB3v7RlHhrMX78ooK
Psl9S9yOvK3HbUD9bMWGFh+TtoQy30bZbOGqRIWwHZ8qZsoVkarW8hFgp0zSI04t7x8gKsYnyhlO
5WkCrtkZAlWSFpwBzUE5qaQ6f++cTOITBM37iqrZK6yHuE63hxyRHP3B97nAC/RPauCppir3V34+
6IDMVQs3RgPzQjtm4Brjk66AyQZwm0E7/+B/mOhY/mveSneLGhk2IwQOHUTgXpSiYBFuzm3GXuaK
TtL3EwxeLyAmnr3NRkoG06em5QJLDEfTf2uFXRttApIBgrl5C8SPE32zyszhlVB9MQi4xZ7/JJne
xixvplxWgMw0g8V+cDDelKBTc5DL2LSjlOzRiYBOjLQYH+qkpTEAmDYK4tOR/VYjN55WBBQ9c73P
oOV5EsOMKcQmyBo3OCf+Z6DX8fbQThtMwDD9d3UI46t4G4imr4jHefSVA3ClhN0niZ7dsnZG/SLV
8PIXFD97u2SfXnX9zQNTiGepyKvDjUkY8nJGCjRgAgIg9K4uMCShfIJL+4pv8VofyueThtFTKjcz
eCD9HMRakSfVOMBVQRfnR1hhh9vmxpG4pA6B0qO273HJWBut10lC/JWGDK/qW3Ysx91jZkrc0rin
mSDsgBEsTTLLvKHCiiMCmmjX/AOTiyOQyEE7uDJdACqJO15UatveIYPCM/p90dhcfzQL6IKMff0h
T0U0JVTMVSh1z2038mO1DQQFvnEn5zcDwfbbKsQxivNj8gboMeHIX23cD9pGeM0TUo5MxbZSvPtA
XJf/nUrv7YfBX1G2B5rX02WIlFxvc0JVx9JiAUGOxlfFekaEvDc29iOvPmdWSo7taJjin8K7z6dd
c3h6FxbCINsw8JhMRA6HdevWitmcjPwA7DMG2wkNuDjKTmtKbemAxwbIxZsW6GkdrTeQDCIxj0C2
Y4HIfuTXU6uaeaTlEjIKW57mgnyB5wyBYH0gIP98T4zBxgYfq2Z6Qu4EK/soUw8revTDUtocO0mN
d6ItLP8TO+PtAQfvTIQm7Oc3DXsrIoB7hYpvQUavu1XNB3YU/GaZdFY0riiFUTZqt/NM8sSX2s+D
QkYnprO7imJewhM73BJJzCv7NgEs7fzqg8WMW3DpVabXaKM0kcz5C0WWPTrU9nQTpQEY0aOjnT5i
86Iyh833yPixUojhQHZiUWWzKOd8p4oapk2oEjs6nrA4cHrM2t8DS4ewhk0jdMvM4qFOwAdo2BJo
5EXSadIcus5jDO/maKjyT/3E5gUZCZqhMfblR/VTP0Lt4QlAuwuv6j32YR4OTGttPS/KF/e08IUP
6Q1UFOrwcUqwwhl7funQmfTTm5UPbVzzPY6KnXbGS8AUHLv508SyorWT63DuHp+7pqRLb+v/kBQ3
L/X6L/wgAitw51DNLGzeLJdf4sZxbJO2awjoglN9z+92UpTYM2kNnP46EtOp73DPmY1d6P1ylG3u
/sTrQrnqSXUJS1XSMSGFSuxF03klPPGsy7qO4+KmUECJyh1IlABp5kh7MFjHqVwWLnoiMJLCYPVf
QnNn4FQ6snYzVD5igjSqXw2oeMukESp396Xwv7wIFJ6LIJiL/BNNK03V25YItomQDGBr5WSJeiDZ
BhEsRZUSvFrk4p/BA/EqyGWymVyMvp1Sb1mfvFFb0MORfpA4rez/vZ4S/U3jNLjEKzj/qnEVVuVx
ClC11YIewE7FT4dlaLq2JZDm9K4vhSAxFSBY5wyqyyQFHe4qAMHtXJHeJcpkIcDymLIqROtiOJrP
XHGzE9IdMEfkTGs9OEjhL6uUlX0r2hqL4J/1sJs/b6Sujo0nHaztBWyczYelWuf4D3aE6LWOhAgc
+55wWBPPr1mobDsIoXC6Dr7p1lqJ95Ptar9kXziR6W+RASMrqOKB5m2pXv0cwmM7gp34RtvqvHDM
z1ANXjldgOVQzlBgOw3WEShsQIN5DxI5yFbW8Wg1XMIJN+eKSocDfc5dfxX+P3uu9JA7eGsHbD8i
mr+xOPoJzwv1yEr6hYgLXgF4NojHo2DndKdE+/Lxm0l1b9jhE70FFTWUXHbkZmOUKuWEWCYnWRt8
uZ92jFY2yUqSQSsRUWOst3Jsuaz8eJnFLpOpEcsCts4pxRfn6ykrer6/tvN9SmVedzFbcwJL6M3q
n2MQBEruuqUxKRobFBMG5Lxtai2uSOKizz71Sj//XGtfI0ah2G6Ff0mzfnGGbNBt9uwOXRGu88V8
Jl+3ZKuptzzZKYWFfVdjML6zZX6FTu2gUZU0cJKCH1p8gzGQUa/SL9dZbOvecOyJ57ZBd/16L39t
IsEVKHZX2/23VrVVlV0BlvyvHjP2it3MWN5zDHVMcxCX04qGY4zRIyzuVIEnUxhFZieD1eSXxjT6
DIv3KcI4VLLF+gyiWTV5+RixmNSWcS6xQWunl1YkbSRQ4X1QWAwFgvbqzzKQwzXGXavmVRHqFXK1
uAe78F0Wop6zWqJMkOWHVoqFJHxaNq8m7ogOEJJPxuSqXJ4yBhkC2Lj8coGUYIbM9iPlcirRqmr0
qMjYXZV6AZL2MRGtPN+62W//tdS5lSyS2hHkvZ6zqv6VGBq5WbBBxJrbbuGmFYlpjQ6vgic2hiGP
1jkpTszXNBRiEjrHliLwy4ie5TVPvStOtb1PyqAgeRAS9qys4Cj6eao41TILCKkt9M5IS1Hq2lXw
QjwvqcOOXBoOWW0x5Mh3kGzMrAeaiBLqPr9yrjQVdLJHcG5BlEMeYsa6lajntReso2T5Y6lYjfe8
lqmy1nj+xeyVwa1Ppi6uZzXEvoWM+mkw57/6ij5j7YipOqwPuqcvk5e+mtPSirYiYQR8QW2pg5o9
PbF7a2VrJqySF0refC6edxzYCcx6Uf6/tqfoF+zialoX8sc0LsA+nNZ8MA+LAYRbewegpkr8kwEz
ARaZOUida2cJ2sHWH6aME52zXcr0M46yL/hmHSi8Ta76n0zWCNeNyo5md+lQsrnc0FQ08LmseG7T
dHVv7pb5abCgSd5V0zr3Fy/O1/CQ4xuizfCcvLxVR3EQdBpt/SLk++hom9YyQvWIomvVwNhM8X4U
oqv4RmTuaExqgAUMzncegBG57EFI3081+8AM6BYQvxDH2CTA8TUqo8kb2ZpOTD0MR5Xuu/Qii347
ikYQiVbPVqsK0t7FH7n45dNKFohxACkoxRPHvCF4LkbNigqMaBQkN6591MPyBLR6iobemudKIFaB
u1J6t3pKK8KUPqW2SQWJPTT8Cb8Mwc09q6zWqEay9Z1Hx/rukMoe1Xjn6kR5+v91BiAaVjN+sKl7
o6r0Vmh738gRE847zNrhOWey6AlhToXMeptsyEswKIM1qA6UBXwiquI0HrmS00QrHvPioOWSw7Bz
mYyTwRtjTZ6gCSrxo2kUZFOXrPg+dRFF/9rYvDVvm8HSzoO6WOuBDnkV0O8jFjgaqcFC+KrK6oaN
nTeu7hhTQ3VB9Ich2DFmgLAXVijB4s8QDtGh4U0xP/g8x4VJxL6ILBHL3sMTBzGzcN2M9N9LP20H
wt3ArJP0+wz0phMFlpFgeUdacT4a7BVDuMVW1VaueAEC5+UoBB/XT3wB5BfY3Pk2o0fhP3SDfZmS
iwjJmFNKtVmgSWYcUCGJOuEv0fu2povLN/oY+sHorcnyoP2cerSu4YIOSTRhkZbdk7b30FFWeMQ8
tygyMkYQBlgP0rcAoVSk7RG6Vo14YxwRH/OGXDyCaduo8TMy5KVyPrmINMAIm5OicMpck7iH0pX6
fxpKm8xHpbFNC7xvc0l5MGi54DEaV+N26+8QEPhi9rTMzDmkrw1DUMWKPG8HPGAWlO0dbgrzZmIO
5f5v53UhAvRVW1K3PFlBg8yXV2gbgcKXNDK5KZ8GeRbT5QH9/Gx7XCWYAQItmPeAqvmkkFN7YutS
J1oBcLM2DGJY8AreE1oL9lnFIvr1JgUxYLYMvAzHrJtNub0mAoTUaQmbIuVI2uFbyFXxZXlMXtra
7NkHZ8e+numyzr2UVArobqiRRE31fn+Rj9FyXWlmUX25lXdQa/dZld8PfGGrog+ESpEKjDCZdmAG
0ZHiCzGNPnylQVVkgWXQg+44ek6ebQ8bJgHWDSRn3tulDu+9/d+1ToxbQ6+QRz4YW2Ha7OzW7WCO
GeLt9jw0mfzBXLuGJRLLvSj9eVwxMp/mOFWWKIqisdXCtn554xhLdu5UP3BO3pH1ATnFMvQM5uRr
CQGqyupYbOhzpcW2Gi1egxPbKFX/O437fm+OYy9GxsAuqoc8AI2RPvKF5jTyV598rxbtuLPyuGou
9NB9iLxIedPEKwiUq2HYX8UFEmk7peScTj2/lEoDOY1Jd70xx80H5cZhxqpAwQd8A/lz1QVqujrq
SQPZMQUS1Zed2vNSKd7iXtWpxJSaV2Fd8cdTsH82I7jbcVUVOSQkqHNBj65R0aHmlmZiuyOV0/bo
phEQB5XgEe8TY/wEVeGGQvEnV1MKKQuiunakv1aiWNQmFsg1Tc9byt0Jii+39BGpcZfp1fCXQsM2
RmZ542K9xgGf/eUO7cqIPk4oa6/JcPktbC7amcjEbY/ml8p85pEMYFTHPCezSUNHD/SaxXbGTPFv
COqj5pRZDsikBjMzmrD5K1DaDjWn9bxLK3BZY2shafTimYIbaxPooX/cZw6U0vilzCV/0m62EsKM
r+5/ywhNLnz5Qh/M1h4lRF0cZZ1c11Boh/qrBsoA/3/+yy1x6aqhk24TPE7rypq4BoGNqRHMJ2fe
BGEhlGMGmPhTUHQpTPqXWsn88+537rMfNDNFdlja55dSjMNtmC+RiOLVnzhFESw6qq2Gs3d/XNxp
b6Akl6ozf3p91XjK8n0/m8/u3JRd7ObhKY3DSDmRPfQpg7Zp9G9AL3+CULPRNZiztlVp0v/HV4iF
g8Y/bQjbDgnxPyMWgAvYd6u8TDDVfECFI/94hOM+7lvsfrAeqE9aI+lDrQHy96g4N0z5ByBZqaOI
mOaGv7Nu/KPF25dg5bztzUVytKRMXyqA8W746ZEArOZit2Sc7tlpRSTOuyD+i1oNjvIeXzaMJW7g
Ekw7YYqLU/QVIW8YRsU1etfqiApYt+QHOOGwom/Pz+VfX52uh8b/9g/3OqUdLH+/JPDFgzmNw6Gw
nySWzQm5oK1B6XVzmbLuFZJgtosCbDUbplYrWpmm5OY5YDyK9jZX0mZefZDr4eUYfKe5RmqgEZZt
VQagz7djMv5gR6ZQpmF14L3/C9jbjhRPj3yZBIUhnJJtCGYGohRN8Xbd8BfWXsjXfjzqfsO/XhdV
GR1H5Nk31XI1Ea3Tlfhat56OXwJ0TNV2P8Nxe18u/RH3ZzsEl6tvZfXHK4dSgKNENpwaCX1Y0OI0
MG+0Gjn4tD+8dEhbZb86by7i00/VF6riT8nSrK+59yMQzkt7ie5r8h0oz8gCxqv0BWBttJB0IxAq
36KtF4C+f5in9T4Chc/TII+0Svww5CTVNzm/9i8drxnzLCYzR7iS2ZkiuD0EC+SWDWWXWMd/z4Cr
q0wpsvCCkUcdq+vng9yNNLtFo44Jb76L0lwA4kdXJoLclZiPBxNIYq1tcxjBiUjggI5Q6Cx2A3RL
yui8akOHtbSiEsmQ0tl1xPAkxDgsazhlWLNeQr0VmlUBEXWN9JySZcAk+VZUHP+Xjcfzqr3cc8NL
hAMFV/VZcAJxb78Igo6zLBtQ0lv9ubTNjeHw2D1qGg0KDCm9aRTSS05Y+cIMNc2OmPHUjpjWUMOJ
DEz3zm8TW8hhrnR+Tp3JXtpMNQ2AHk/yahaMIctmGJ3fMQT2ZeTOxoLUjJ73NC4km1uRHSYZ0dTK
euXAxIETiQKQJxYu/1bVla8jsdMFH31W9taEJFmOf1BwTg7DVyfHVpKkSCgKQRCF0ILrIm5k4FxY
h1SGjuQ+cGIgo7mB373PEYRhu8pk7BKh8m+MD1swC0SG3OOaD/lmkOjeoB+Ia7rglNPjvJHMon+u
C4Auf0pUhF8rbc2QzpwU9gam7gu1esC7ulC4wb/2O2TbVcoUtAjpJNSx49Ou5RZlh3jw4/DQky+D
7zTL8Vis4UiuX4w0H0cBDtAV/BStdrKK/zld2ihKwY+gvILVkkQRNBr9Po4y1JfWFA6HB0D0YJ9X
dfYcPyY+4hLnPOy4P+XRIINEy+IsYsyybKzQKSZiKysnprpCFgrZGFdUmTOCZBMPTX50J9ugeka4
GFhVies+LbZnz6XvJZ1/zu00aeBYjWcjBBuTjZ5bo3y3si0Z7Hb9gtsj6+75SUbhcpomYUiLeKVR
VvLbYcDGQQhUJK9wP6fopNRovIxsF7nkDAPKvgMktWOxh2PPmE6eWez4ekxrKiV6zn2Kt/acPbWJ
lH+PZZwptTbqZsqkDfOLesAUymgzrAgzUlGxqbtb+KAkZCbalyQP1EE5JlVkqboXsA57/yYlF6tD
LVTSUBFJgaWxaofnTTTNDiplDVCQGveEJccZxWAc6v5PXShGdnjeTOOEBF1WCWxCzJN2nf31Tumi
PVceYYH72D9fowRw7NaNDX5DfgArTGsVC/ImNAuWN4KE2IxFjiVeKC0COvb+jqOKUwfjWY0qETUb
T6b37vTpOcB4OqxXBEShioCVNV0xLKht2PM6cc9HnYgllqeV0yPHdgupQWIKO50ubFGcWu+gAARx
HuhQwKRMaK7U9kLWH6ghVLe0d0XS0GYe0300oTIUzJk03Uo6/EsaN8U4/IGVONPsOUlxewWAxzea
yVhDabHpnkEU0e224b+mcMXfAZRfm+u+5sHoG2pa5RydGpR8FmII5JUMnkcXH/HFzQraiR+0OxVG
aK8BhIGAC+ecwIwawFmTS9Z1UBjF6KlQ7+SSuEKdO+k6gjm5S+Jta2+QCcHHALRiDz9YMyjFqmEz
UHrHQx0s9MawfGVmO/lEppvg+7UZIVzrFfW4AXiymScP7PIHUGy1R/aKuYrPi0fphfhc9dQ3hBOv
B6VlfRdrA8yxh1NBGvsBShKuo7KKbiZqO5+34Z/nMe5TGJaDIl7W8HB2Q1byU1xyTT49y+T6iYZX
3NB+3LblmWBmEtBxp4B2iiL9nb+Fh0O9btNz+OiLqxVHvKFTIJ6D2U+Rjo7+rR+V5qcgvFI3/6bM
1KEagtyiNcj5qFkAWvZzdinXrzM/4fwoMLFXHv2UBM06tFqlVZFZbw2mhRYcDdgFu+xvhCItkEAK
6UjWeG5xXSxN2XnIxjiYj1WUsY6RkJaZs88nwcu44EZyGapvRi1qrs/5YRMQ3gEezNX8qn915Uu5
FAIsLOnb1CUqYNgXXTcNu3CMO7WH9NXe+dD2pMQ0YLaAVYzwbN62NNqldtBFQTq7ibx9tH8ZWqxE
W+6mo0A4ypDCg/d3VUI1QvAtLcGFUfzfN6BAbO49+t/eWwCDUnJTeSttsv8UjiDPr9KCrkXDOBz9
utEyIndaGWuL6VbsTsiB0I7HFMQwZc8bbmdtFpfOmTGiS6k8iAgh74xysmd7ncNmVIAzWhd6Ppmf
x2OT2ypX7MHPViCUyoMkfXqP8pfU3w5yw+SPAJv6V9jigP2kaiCKM5da9nJbbyGxNXmSUCbO7mSJ
qHo0L+6Kor8z8JjpvlL08RRXEppVtifS4RC5Hn73ws6DJfTZm6pXdN0R5m98f8wvCb/jzi1W6B4Y
M3AFs2JTxJkaM9kiIYOgTQqipHYD+Yupv2ex0ac6cN/etAlKZ2BI4ZvCP2WGxYBcRPZ7ABMkwzLC
cZlCfaCLby/WgKMtbMtWrlVvIO8zi1alRSgmzIEnOdNBYwgoW07KF7MZNjWknIvys0NV/e3PWiF+
C/OuxC7CBIUmbPpYMIToML0HKRwwA2BZMwDRkgJ1sYBRbBhEiuOQbIP9ja3OBLkSK9mvnH+aMhfW
CpcETyz1aMqWcvjYLAw0whmOc0Tv+EmF5tc531ZNlKBn3Au4xnLPyjXCVFntzgsPOhrsKxvut3Ld
17pdXOgGL5OHZywW9OtqZcyxjmSOlhi6TfWjvVl8WEO+dagU8CNpPZlrh/ZUIX/gIMmASZfP9Jwe
05t9NdXETknHsv/91XYOvbDAieBzR31oDf4Rh7GqZ84dTVguesW1NvXrjdM0LmYU9K+ra2Ul0fqn
5zZiws8R65jPwK+LNmZA24kfB0KzKeNbwlFv3CXlkGMaWI9kaHJfZU+q7OdcBf0EskPAN+FQVe/t
xGjxtUfbmUZbKesPc7GfG4gmejYNzmF8wu1y1/c/YIoDg0Bc1+1XVi6++DrM1yD328k/H567afgw
x9CibmP84Cb5yqM+L6+f4+X2dlpBzPfOAaRvK0ybvsiZqjAAiVACoiadLwZS3KzztMG5LL2wHhVG
kYTZM0jOD+JXvCOvo+J86lEFzMk4PMcSUmns5Ib9Pg8rWpFT7APbdzxCB3bfU12sX3rl1obiKZIu
I6qrjajy3MlZqnxU+TSVotqbXPFA3SWYcRCqgz4suF2LEbLgSLwQpJ2exT6mY610c/yCrubQ8knt
8HPvOMjUMtztmfmbtlZnyAtv2Zi38pRZlY3MsBCFp3Jul80KFQnXWchQawNyf0mOqSAQ9ryp3XGa
mMa8Gbuh/unKtgN1FZDQketL8WIW51LQLmgHihsBZ+k2lChAWhtTydrFLS38a3QkA1zbKBbcpHrK
fVK6KPEisMyiTHuYJJc/HnRJFE44hboS9RmBIt69cvTqIQ8+WA3KqUN0Pz0SyvwcqsQPcQ/4PPBJ
2K/W8LZ6t/TpVJMTQ+dSM/gr9L2BHY7tIUddUk5OvQQywu2Y8wNvb9pGAB6+dtvCAxDZeXPTpFoq
pph87PfkwhVkqg0Su1+l7i3ocx5Tsuo/jrqvg89Z9+uIwUElu4ZvuVFU6EWus+ddaJlR5WXK0p6k
CchePz3Makp3pb5gL07cF5FGahPz/2BgqQN3eVCooeANPWs4FpHr1Qd95dwZl/NUj9hDWofIn19Y
dLRos3qZjXwkcNPaIfrEkqLZpXo/hgxacKnzb4Yb/r1EgMd5BAB6CcDEKUVXhPVll/kfEGRG/9gv
wpN4Osg2Dxx/Le8afKJtW3fdmGR5GG5/uqTIoWqloqzrGNWY4ad1izDwN7rEjar4V+zfk9+ZPBCw
ZNeSuCn7R0Vu/YNp6z4lbr/gFiPZWtLXNffi4bBSrgFNthskDX3tubnVRkdGsP0yKn88B3PBFnwN
4ymq8aFRxL2SBjya0SKhqQZiJEFW3YQz7MBOA7z9w22zbXX/oLaFUcnA1nYYSoRPS4XvNWnYYgxP
csVRDlqLJtMeaoBoqaH7qMvjjpTzdGfmJLTR7HWCYHPgZLclu9Ei9U4uVEw3b+flGc0d4ekGlC2S
Pp3Ry07n2JEV6KU4F97LMyocTshDMQeq+HNVVfkTE0vXMOFFYbfVFvSb5V+gZ4JPIVBIJpAG/DM/
G8YcOVV93k9bSgaeS5LWEs/FtuP0ugYtaf0RqjodfVmxN+6sQI+pSNESJmHOkf2AuezlyEqlSnoD
xyLAbXCRtune/9ZPwZS5ywqoKKFLzbCw0y6ixUjYwMly26QtUmLLDkx5YIXRXgkin2gdcCgeWVnI
uUEfAwIdNZTvjZOJaiJviJ7Vzly1l0GfdW9O1SaOnYpnS8pLB7ZEt9USQNkEUt6CaWSH2G/t6soQ
1Pkvd8s6AydFwA6NGid2e6SOJjCzL7foZEtQK6Sdvx4ME58D7Sm8bd7svVEPr3EnymxuBd17EYWS
U5hfnnZ0JFTE6jvwY8Im9wuVBpeOXfX7gJjmegoip4Slrc7kVD0Zj/vrNJlr6IhwD9BFT0hxrk/H
WtSpzk87ZhpPBpnfhm6zjrMcpbFis8yC5J8dc5IY8ULNUYZEMsIEMTXGAULgAADyEBTXYflCqBNA
iPKOTLGdKa2C00v3UEo6JRzoLc4Qr78P8UhgQq4OgA3pAv85k+SoVROqj4ytdyMIy+r3R/X3aBHW
iITaGMMG8IUqBJ6X7vAomgyqIy/WMm6XkfR9pnCmsgZK7jylvXM7WbPnolXFeavhoEpMbQA9HFE0
bl98xm/IoSr0ClBwrN8pDnnR2BKf+FfrNhyPkaJ53Jl3l0NzkF2G1izB06QWRJdwbKznzHVEjZK1
/NHiSk+AEswLxApzSzscWWyO4gozohEIBwYB0+GxbGfCBhMMgi+dTG96eTjIM8GquMKcDhpSAPJi
Kc4KDcztPC6xJt+gpqfPZIbtvrkFrZkqh0fL/yXrxlRW88qCtuZbIb2nq2Xq7H4eGGNvL8d8cSTG
Y5A5SYnso7nvCny+nB/d7RCfHPhh+oe9J4/eHfSWZsblwYOJTCGvUIlCvyoWTEwJK3k84IIv0hyV
QiSFnBk512Vb70QU6oOjShDKvALqSuPSQuelpqqdTyu3Sgs4xbwrQv3XqrmqL1xpDgZZazcKTpNx
VdVGj85XpJYjb0Ur7D+kx1KECAkw71jdY3ZIX+9HXJagTZrulxhYBG+JlBg+KSzngvrgtTh15tS3
i6xtmzS1iBu3BtNm7rmpk8rZco1jPnlg1s1HagONyWNgb5+K9G3JEUVQjsc6N23pQPNfFNAR6Klv
r5tQq/AaPuBQXZU/jLFOPSC58Mn5QTDtXR+c2HLkA5lxI0j8+RvlaVmDz4I8g6VpIto6tUXSJJV5
5ynlNzxXptCfViz/lbjPGe+P7uxhYBj+8qUjQRrbc7SuzseDzVp2QY5yifSF5VA07q3Ryv3+mW2X
X1Z+xyMMFiImcKBvfvEo/kkO86HXXx0Pm6s3yq1wOVsBjKe1BuU00y+jwJGG5W+zQdpEtKSE9sDX
0CiEAwLQZadXKkXa0yv1UPlouE8YaQnrGulAZbUHHJYhbpO2/PP6vuk2ReeQwFRI0iD2JZZC+R45
AaR5RFkZ4mKEL+KrxFytDx9Yod9saeVFpxHHDcJDJR0nJWELFx9N1AuwKAuxHtpoi5sYVfE1IkWS
TavyUgoA6ASWVQpKYUGU9RDdwuP706RXF8fZBexi8BlH/OTEgkG7vjqBF4st94apSGQRFu4TxjW1
a3n0qIdf0XC14viiyfRjv/HxgGtbXRewar7zG0D3jt8s+OaRcg3E5CAnVQWG+GhtImG/GpFjeY35
dCchuzqzQlyLUirFa4R8JcghYAmcH+7f2d6cDvarQo4HGqFKkxw35fPqVNy9F2BLF4Jbpf5kRWY6
rHXXF017ycb1py7Xc/2Mr2HGmlNBx3+dA1rIwAPE8WB4kGgJ0lQcnekEOnXSzPxkBUKuPsT1QxdI
R2r4mxkHdpnJEloAxQGFuUQGrm3P+5reyrHzfse4MWM9NZI6TQA3wc6hOSpaxeOe1PStTviqK8KS
1xDiNVbx5i3cGhTBJui+TLFw0nWN7bm+CtSZMMAbLf65PG8NgkabMsjyL49gBZWPlkuZ1AonTTwm
yDAvqehJFwhtVTx9PIqj0IMtQ3lv6wXhC7cmAUVvws784ytALsCsH93dEJuZnvGVcAwnVAW+/ZhN
ozuFfxb+bqtU1i+K2xHjL9IPHWe07wsYgqSmtLeie8JlIriAypdGH3p3URlGW+d7rJPKEFXbgOXm
841S9xoJJrBsDr8Rc/3l4NWYNTKTcY9smo/+FzenUcm9kBteB0MHeTvsI38IlN+zWfuycV4llqV8
i1xMllo3JZw7k2aSqs/xkjR4FQ5PhYiKL1i8t+se73LxyAhPtMOvoAlOyDSRfnHLsBKXkohRbodl
cqB1LZec3hBNV4ZQXrOlnuJRvcuRfaxKKsVAIzyV3bhFgIzPIvoFb0FLjloWdSIO5Xu+qLhA1hXW
o4fRK4USDLDdY3ycK8YLaY03DZQK5P/0A1POgCAaNiDjR5UqG3PnUH0Nj+drzdDDiIn0NEWUAa9C
9U0NOyAXzkZu+jr6lC9yHQrw+YVv7xIZY0ezEqxyHXa1HolIuErEtBvk6yf9C92ErAa2NKJOgLG9
dYafPoq/S8jupp6BsXL6FmflIAxum6f7RvErZlB6KWVS9BzJXFHZd09dEUtg1FEdnnmcvsV7LIc1
McgUmLlw9d9PMLNRrz7VAuZsr0crD47o1r24nNk35GmUW85vyafAcYgJh4I+fWeqBAAAcfaCsZT/
Xl2i4R7YR9S9eQfv+58+AQcDd+kHpq3r6MbGI8+T4cSwxpX7INbI1uX9Fzx0srKyoZhXmdXHiOT2
HZYw1HXXbAgmvyH9h3AQCRH4sMCvWxtdgVofUA0kqa6zZblxRNAYDXiBduyUjApUZjEarIOg0E8U
scH9ZN7fHRIZis6wspbHnJEH3BghsQn+uMKg36lfa3Gt80mOLCH1u4M+0DZwPzG8TN5V5bHdoxpZ
53dITT9g1dr2KojpETfAzIRdZNn5yGH+Ml50vtbdUTwolRWc0NqbPENiRN41jobBrJYVKfSj2M6Q
dXGyehwghbuBevFwD2pvvD+NKNV1ntlGvtPyivtRBiJ8r/FU582A9rVkoqbEKXphzGm8E03O44d+
VzRQTVzXapR9Zru5ePDG0u9ZegLNVSLnELizoon/l7ZzebQ5hkXzqMPMexcvox4BCQi9H2TrQsYn
YzOQBPoLKNvnM3365tovyz3MUoEPOEtMKvOS8ss2I/5ARhymyJcgl76zMARWEZabIufVItJWIpzu
ZlR0rT9/CO6XM+O3QT63R2+WVIv8HpA+oS1gIpsct9uVF9t2AK6VU8mAOitaaesygNeb1JASnflQ
ZVwHE5TNuaMSoFiEnfAt3d0SNACoPhk43pUGLm8lU+y6wefZPaKHMFVBvz2ZSCPtCIfPrtqHxuKr
4jToneaQgjH+DhOBDxmVoWajHI3wPrWcFr7e4LOb1jYrK14GZpNv6x8vVQMUGgPWWpBqOEnRlK76
nqU6E33MOlYZr0HRIL2zi3P2l1pkomWFTzb+0aWDuaTlRUYTuWHUEVoQ7rcdQDSGmdyKLVRGFcMz
MitQabNdvzCrJtaJFY+3HOrguFwRysodA/AupZpuYZLjCtooRd5yFwqYScHFjzVLcHXnKoJClrbT
RyY+nTUHkoucEIuuM7aOLK6htzrcaidWasCDb3UvoUKhfFYNCeTGQNId7pexAo3LWtuJvalLU4A0
+KFsYMwN7iRv2IRgETu7BoK4JNYXaVV/OfwMLFND24LMXhMyniiLDAw/Vl79GjtV5vn535Uk7IXU
c32ylKLe65HL535BEnCRoJ+KsHYwY7ZvQ1yM4B3/Vfc9aQ9gEgvRqWqQcUFAkxgYGITJqsjpFG2T
il9VaLyhs7wTFEBeS+Dt7UHF90HzZ6gmLIsunNocI/C+kG90jKxzlxMeavlqBuhS8VKmlbFhW9LZ
ccPsDpm0DoiZ/RPkHIeQrnN4wiKk90L20K0vZoithiqZfZByafH/epk2iAfZlfJaW3Ik9J+vMPpq
dqMXIV0hNvBPtMd6EtSFzqWqKu4oygLeB7OvWLhJE1nAdh0u6GihXDoGn+HE0zr79nWvhdUCwPUP
VP0kpsKH2qfHlk1cTEcJLIohQPbUCjZE7BvhbrTd08b94Y3slqC46Je72a//ArAH/k8L7x9D2w/V
2X7SWfyC6cp+b0SIMddI4KARc35GlaXDohMFkkJp7sBa0CuZthxZD9Kc4yii+wAtXQ/kq0hGTkhY
9e+De0RE9HYQKt7zpDLEv/jxwOxwaJGAUdcSSIeH+0glhvOneb9Nvrz7BT2VBTNb+4DeZgBuQoi0
YlAilpXGPwb1BnDX5eD1wH/y4RkvVxuh8D0klOZDEsWBAJPBdsLAszNWRFjY1OnXIhMj010xmMFv
gNN9EC7fK9ED3o6aKG+M6hrs4NrCVzvMPboox4XxHF+wre3tci6uL3c1G0ZM6uE12Z9tPFARLf30
BwVw/0nw77w20S/uK2eBKJgMmg29AilP+3Yn3Tr8guvCua9XVe8LZPYjZ2mkEcs4iO657MX8yQnl
HqpfdYohhZaxdaYykrpyAYAIr8ye6KwTQhHTJZ1scMQn7LBSlIPx/5mcYcJo3O3mHlbZpe8Wxlrb
/vPbvGVKvozzBXbonb0a+3YPVGMb0x5ru2+bAD2aJZOyPGW5wkuoSbC5G2S/UPWvoqUHIJmzX/eP
QG5YdmA21CxZrh6bsBo+oZUBW50DEiscW0oh52Y8mSvjYLAYKD+rBZIcaR8Y9tlKTdss4eDAQt2l
fkcFsaWNd936w94lSRZ2GI5WRES9q1C+CQNsvultKrOB3MiUvFz5CaS2Pnw+4l1O7aLp/74/pjsG
dCHmnVpW3QyroXTpkHxYklhbYzfcYvnwJEuBxO7EnoxdVcDmBET9GImP4+b9ksT373qPesOK5LpV
kNeBV3McfCCAWlULeuwZM4isJhCRVBi0+oTE0URSD4UZOwrDX23/YtXVGSaL9tRtj4KktRrseS8D
gS/fHvANyqJopeLi+HXNItaskBzRegdBjw21BH/bBHATvdIADtnhGg7NbwAoDrwBBZ3pachWP34X
ZTzluUF75Utvds0jNqq5g/H7M6Zrwi1mZmrIpq5P66v1TksC7oJ6rtlbKqJ3InqFSZYLoJd4upX6
AgsgoaOXQoiiFd+bWyepyLq4azEPuQw1z1K3b9Kh/up51Tcruk8dbO3dKYAwHdF04CBRVnm64eM8
Kt0K7uM9oxB7l+9TWhEtI6eJDrr6jAJ0+BaNfZ2h1/uNcSDxiww64q7+OSML+TZE86KeZdemLZN1
MfAIZH7MRArE7ClCWR+9XZrpeObqWBw2LVXxFztGX9MemBm7NQPURtiOzpkpddyXdYfof/4w62iK
9B0v3k4+JY/mCy0Ky4gxJFHdJKOEgYvyIQ2scrIm+ACuH98mGZxywq6MitoUlU6HSb+AFUYC2SjA
dQBDty9mNtqDTIXVcjotjR809B7y/aG1xJB6Vyf6tpuGDAfEd7lSSCBhhDvCjErfcUbifC+WKbzR
GCDd2UcjoEFKvNlJaEoyH/cSbIpr9wot9VqDacCA2vIEmzkFTUcyAQ39mIKBEMHiFqqRk4A5QKGS
qm7eF4LY4Mo/yGhmR5SoKPfQmFLxY4ipXtO8GXqP/606nLUrdSfqup7ucoPse7r8EiRsOZgzRjkC
U+kAhEroy8v9/mw+6nq3IagMcR7rjeSqSsyj3t+huI0wddGQKPwqSlLxtvkmn7orHzJSGsmckG+k
AK7c4stZPcFga2nSIoPi0ie/n7885tAszgFjKyCQB0E8CYn8l4i+hfvubfEjEK6PkCr8gfOlV4Os
w94kLcJxHqQP6bmgWxRJwFsdR3ca4fxqG0Jgb38jB42QLP/P0EjjCFhtFdImPodvzXNlP8Jd2BsP
KSOE7X75FsCjfqvp5oxzWd2ivlWh70mnloU4YXnAAq1xslIThStlwC2aalccT0MXIk4uMStDisDg
vNZ52Z87iYy3g+jsgf624uFIpqLa4xACehRzirYwQVJD+8cjC4vmTqqvH9Itstj/lD6ZFOp+R+Ex
+PaOuRYXDR0F4ZRXO6g+glP1xXNc5b+DLlxHbiVU27FTergBeJYwOJVCixKFdDjpQQc6QHrk4oxC
w6a8dL0pLXOpk5Ip0/h/L33pyfuEw4hEuTDAY0fcGoEGCFxhuSZmhQDvz4dMkFHdzW4tjDVP5pTJ
8Wnai9XfzuE2pB9pPfWhUSFmruG0ZWDuYQpfHRmXmQnlxjGO6hh5G0rtbWGDJK8oy+Iz5ZavtHRb
w0VhRqcY2qnRulV9ueGESWdIFrNPTqgi1zUgJSiy+cStaWDsJCThRl1BdWqivUqqyjfNnFqW5I1l
yHW+zMmpkR9/zg0xM1UcgeeKR2zWABG2x+8aN6O0eBGdJZ6cVBafiYL7jaV3qfX9c1WvseOs5bQR
T2v5Hb4tI0cAghrKoEFUymnS5HBKH6YhoMtHIp/sZqdEbBxfPbKXVtPvQioDHU/r4NMheKhg9kYr
Z3AZFVo2f9SaBW9XNPpIZgeNfRhehAiGPWQ9QvCgdinyYhY1xRFpcpbL0KggSwggaWD78vgnrMi4
EdQq4rr1nOrbzf4ibJUh/GE/7Ojin2X7HhnnVkgjX+mmro9KiPq74A/wbg8Vof/NAywL4nM9jB/m
C+gdz2t9qA5Bs59wYafQgs/MZegH84hD1wDehqEZ2mMwE6YhN7zWtnOD0s3hYJ0/bX2FzSeF9D+j
y7leNbVdRn03xChAJHqmg0+ybxEKcIx7ag0mbuHsU/iz1FZgZ/SHSfcjGT0YQhOkUqXhrodPOs0V
ZueCE9f4BQ39ev1SJnQrugbEMXSDLYDy3EZcnX6xyTbSO0Wa/Ybqnm+GUJTFY5PeGSTookXAncG+
Who0bwgQag1bnBBuIVqmg+VC7YFRUfgnVCp1obLX9aMfexClIDxJqpiGp3jIspbFilXbzv+6hpz7
VaqfQ38Qmas4Qb/hQKL2dFmw5hm6Hzw6qJ/5vE0hf5BmDC5i8mN76mGn9p4wo4oIAuXt+u8OJScu
6Ei7V92yYLERhCsARQbGICUJ7ih0bFm7//Y4mKT0n25FP5wSOaFmyNH6AgpmBbhmb3Nshc5PzQM8
KR+DIcjS7TG1FytC+bYZhCA+qvUQ4t/vlq8yZYsla7ClVHKeoghCMeJQr5pRo5jyPyfbKT36Evz2
E4TDMOmSbmrmJ6xsaE4o6S+79jNimcz4yeWrzbXU/vsMXDtd4c6IT+DZ5FhemLhVN6hPEU26qg1I
y1m0s1wiYNI67lSK5YYCCxCdaUjeiGYVgl8GaeybXYEn+KLHL7BgHYgJjG/T6JdMd8EzqWlzUnoN
pAiGeJ1nM3+TPgOHrRFZ/CeSqLa3wBC3J1XuK2bwAhs3LS/xQpXDvL2wpP6OySA3P8hqjOAIKJ40
DoQHZc7d/TKnoEwb/bib5jcwPr2SSd/hHe3yv6hi+FYMISE9Pv3EPs4vuGBglKkMK90D7qqFAHns
FbWLC6/1yl6mubsH03QvIPZbsDlpD3aXeFXyFukjbAc4VMWLxZGDLmINfCdFKCZzO+dGtjOXFaGy
kgszlun7WMqpRJVaBXuP75B28MI8FM9jMotYYtVq1tOOHVY44ldF9/WP65tMXpNXDxHoanJLkw4T
XnBiTkht1vf0Vm5/shW+X2kTWvnP2xgHaPN4+4AJ8pw0ob9fNY+JpiXKCK3L+4cHpx7dft6EYr20
i5qBFdamSPEvTZnh5icsmJBABCrkkJsXlbjD1IPHlXoOUg+1r0pnGTyrqQhfUDr9BxC7qrzgQCBn
0F4Vt236gHoKw5yptKTWOQ1etYNRRUgPMpvU+5d6TSEaV2r7jrKd6RoiqMOR/nrIESLxz0HIVwZF
SV9h5vX1jUIFD+PN78ixMUKpLAoypigOkCpSvOC9M8pmEg2DFa0WrRU2450kPrpVnRM+/CB+5Dqx
peMy6GVX6U8hVF2Mi8EmKkdzevW/MWNQ9pzl8CyW0NjkEc/henZZIYSF/SoLz4Cfmp2XRPoCcs/r
HyBeMSdJRwcRUFWTMZhbXE4PdvWGGr3bT3oDKQs4p+cIA97MH106FhgfsaP0xi4z2niuC2/1eEj+
LJz/iNShEyBCt5sx2xlpTbN1pXN6UCE3QtPTQ5Aj1jtp+g7IANFra3lFjX3dbBQmihOnl4CaPHqG
haE7DvNDPZsxweBWHjGzkEPs+5Wbbrbc4YwHdreuaf3PpT6mt1llEAfaEGje5qZSVblRuFg5e2OL
GWH3MhpqoW6UeSt656A5zS2EtvERzEYZS90bxDQ4AOzSNX5NdPrkbEEo96h+Vg3ZBJbjYoeCFBOV
mcbDid3C0gwIMLcch0dkstOMA5nzO9f8Ppqi95x00VuAUZ9NRTd/Zg1l8s5xAnx86Ts/JFIuzmsk
7kgL/7gktgMnYPVOW9s4TOQGbvIzljSrqzGmYXfFoHrWKZE5J8IhNwuCnBVOdxOaFi7TrZUyxTp3
qLR54zQ+1hQxtaMsSlTOCV9xoHKSySOlomp6vDiw7egYyaH0Mlw4Ha5nQYMdrt9QSsXvyffgeGyf
wj/Nfs5CGeLScUR114zcVwLKNFtSQQ5GTkp+40B5xDU4VUjqS9gkQtBiyfQrnOGcJS740M+mC1xB
to5LSahd2HwJdaFicR67gfFpSX0Ynkq88A+jYwZ8fcbg5jQBQkt8xsk3dnvz8hmNsXtbUGgrqmjp
eKKjLerx+rNch1Cybgtj6d06aZQopC1jxfCP78kNB69wgrHOYOr5AH+xohDA6Yn4YRzNkbX1l0KX
bQv7HdIE+9WiNGTlGoakdYEjECR5ac+cpv2OHPWrtLdYBX61vCQ1bjpoOgeqInQNiskTcAornQSL
YkE6kWI7QRV5lpUpJWAWno7zseAVIAO3toeJ748CJHp37FYYMrBHvRjqCoSCYnh43bYd2186kFun
SjN0rwor2sUThW2NCIKo1JalAP/pElcPGloYdDZg4UtP78nk9O7owv4R1Jliw30EhSNaTx+tY+wI
h3LlVgwWFEWV7PUbmR8+4WMVP33bPN27ea6O7qoehUiXc8+qRSQ9FsA2gC9gy0ofuQM7t/TQ4acp
FZS/yPE8UHkW0tVD1EY42VfMuHHE+pa8Usc6rYlM/XAuxoFHVsZAqTpqCmj5uVu5y8FFA8Paecad
BWy19ZOhOQCLILxzjWPhX91rP3zWdQOmbMrO8nl9vDEH96c3xgsQNG026sbxrxP4rCnUdRHc1TS7
nWe3GA9d6VO+i2teMRPQhMNmRrj3Zy+cO4SEMhsZ6jmUREG1To1dUiwGYSvWhuf4sB/dxXuQuVAU
6Y1OgoxLlpFgxz1PGiscoWJzCHso8+TQIg6A20vn6Fznd0YXZvWUI8/VxlN7z9f973YsWz1ytlhH
qk+QuVpNFyP8x/2waliA1TFxYm9jUsQctxboFLlxiTuY+QRPb69H87tbNLNQTK1CJkwLT55Tt5Ss
SHUEaFiF19Ue7saatVIqr29f6rZ/c/ZsiI8Pi5JVDwf+QznoGszoV90Wvb8BIVFAqcJycxhvkYPl
siv+nmSAvkaYXOlLbWyIh752Qf1DRJALXIXrbr3b+Pzcus+YmyfJGiIYBfeeH6fpQcYZyYyNMLg/
v6hVkdq7Y3ezoqjgZOS/lNjvBvRGonuhwu2UfbvJzq0wRoks/dFYNqurzAtNXU+JlG3cd2cfS5sm
bih1ibthgyX16EZ2eQ3Q89dZJWXUkEzpHjiitNKlZ69H0ak6hoIsP9J09b0K4xHO5oYXsiZ+7bXT
79UbZpbQNOwMK/Odma/u+FgCxfzDpE34bJrhO3haKpYAYq4L6PODZlwaNxeK413JEdWqnytIFk+B
ifdm06gHpncwGhyc6a+IQIngFisi6IgbjjfZ0xQ1N1IINT5QIrkdCBY+M6iERg4v0VVp7ljak6X+
2wAkcJVmwdVunHT/Zra/wLFCRD8E8JcJuUmvbSPGlhyGo2svi0GbmRIbdnpzGwqXE+fupW3xJQo4
5vtZNfYfukfjOIf2SeNWae6hxYY4iHNSPV52LprvFiBS4hl5lsaq4u7dkE4TSrvQCyQJIlBRLO6c
RljMAQOadSN2V1TN09uvaxxlmdAm+RYf1Ibe+rryYAIuLe/OVSUI1rjVyaQ4JZsF17KmQQK1VC35
Ci9JdURTddkpFbn9M2qucGi/hAP3jskW2boeVhYKxl1FRt9GlnSFq7V4PYj10UdzUlxWrUW6Ltt5
T4i1QfojKwKJOXfX/l+HKenzrm4ZybLBCE4oGv7SENlAROtL8HOsUG4nKOYom8MtMMDWonQSK86O
9xgAiIACiMwlykbHnWVustXAcGeIPnYnJkPiKOpYMU2RWY6MU1BZEkJ1HYpoFQX8+ZULuV3LiXfz
zllDaemk7Wj6whq0Pd2IPrPxrNYqrDduV9fXPK9gHRqpdAHmFAnE1Tmk0mdN/vcOhO3hSL1Nvcw/
YgcxEiVCM2iFhw7SjPdOcnldXaghsWsqpqzXidleKOIGQAPjIJ/W6gJrDxJ5yAKfN9rq1Cvs5Gte
5DWAh9/a8HMM7TWdoFKfvAhbf1tL8tNkNtSgQUwR9hRrdA7BwosGc40cI+RgWqD+Wcknb2UGF0M4
tTwRQxdDgm7iUStXPMoogOEO/SBxToT1VBgGjNXLOp5CZf4tfJu8MfY+VTwH0fXD/27Y2cMp4w6G
IFI6ZefYgjxyh3YaZ9E/Kiw2idFA3p1ie7tcBj/IxPElVS3mceIut5lw6oW6szdFZ42PWPO2OEiP
BQHuwMq9oVtUn3bN7ZnHrb7HDHElfIqx7KQKNnZd8nlFAT6IlspAQ3HoSvbM3F2XlnwNs2wmaoKP
hJF8TI+aFEoR3EiA0TmlvaGo7AYR70U5L0xsnM7OUJq17CZdHHduRp1wTpxsK7/h0lh1yZgoMwnR
1lFkTM999BRLsu/Hriful4CSj9iER1Is/nPeUYnCq3lde2dAqydyZXucsUL2Yn5I8SrSEJw1l8W8
Pg/kcYaQCnQKnlUpXsrhPeq236nd3oiMxbYWGPE3Xmp27jENpUVMvOuCtGRAkc36YVez1Y1zVyvI
pdnIjnEvrZ1uBj93eEb4kjn2jJKH3v9USjM7R9kksrtpkUdNVUWI9ZVvNy36JLDyWcYsF/scHsay
y4Wdr/o3gpN7XxiOcgMN+/gVMwLctHyvg8X5JIO/PkgxEdSHnOZSLCWkW6XOybPW1bpmsNaQJNgt
be2zgKYhuq3kbAuD45ONnb+XTp8XT0NLtQJeRKKkVEembhwNoAwpBuBtglO96Hb2h/P28vLwaulu
u3Y3G2NV1wtRwlsa2uEfAfBPtH2v4MaSkmUZwJctcld543VGlCDgha9y0Ku0G0EIyebyNesP5sh3
bKOqO7pw9U9EDvDqP+tS2WSTkuIXqRhnZhnYbY54Lf/GDa6mlKJRmAVfRJPz3ammNY5Bb91afq4X
V9bBwxO1AdiqzgNFgvlxUvUWbr/u3qliklIq2mdKulLJIJ/+GAkKfzzRXss8V3HeD9EDKQwU1UWT
j7qn0LHpyBEkzqLd3DqCLf6dw3J1wxOPb/7PtdDQQV2aKDT/qpklPNubfBKHz+0NkbmfG8I+zo/n
c858Lns/WqUq244sZXnmuQEL57sD4uow9HfZmXydS5VZnHt8lyn76jw5BwvQT+OxPNVN7CAZhnZD
x91lKVSoUClH4+1hNVe+XNdG6eNjlLBrMB86ixkzjeTEb4XwI8XkXrBOIwyTHBXNuzZcSbrklD7N
HkRHpoPVoPG6yLU5P0zhZqYNkdcD4nzLdr76a1YoMAuC4s7Db8xKa3gLfBUVKCp54DkK9NCOR3Ti
ijD/QQD+pd+zelzfQ8hk/iMLxC4MBB7IfKl0Qu2EV1mZbbpo42kFBHshAmH6q1zU4keHX/u6qLWy
I8CXRH6rPgyX5mzuHxnW83EZ5201KK+dj7wh+dBgHE2EAWyTT4KiOLr2J6FpRhJnD/de+IzmnAKK
LzB1bPJblaF6LVLfIMp7ORrB5Gj03zU5eOu+J5u+n4/huaXpYVq3PRc1aqW01CZmsqGfxjH1ZS1J
pxY6iH4rW2MrgbvSPd99/ZLlD9Cg28W7w3Qe2/ZcBp0yWMOAPeRShPjVIPV80ku9wJDQvcI2DZ29
Tsf4pKgoh703dQ8UbzZFwYxxNiYoatVKAPTx53S7AAhp7He+nM0U4jlqOKDFxAMSh1uxIhY9M1zz
g7xLpkanfFtOrutvLBw9C1DziiLjEuHt74PCv3x/IPg20LTQdTGkwHQAADVLGRyrVPS0MXLY90k2
Jp7TeHd/oaSHb005mcD79wZcGcRChDqQDwj+92M0qDhfFqneNSFqCe2IFVTBNIwMW8opEVA/PWI8
11xX9eoX2N7mb8dvoFd5nNAuuQ6IDNkCmGXCCypL+ST4FW6Jbi5bINW5xjXkfpLpVo9W/okh6A2t
R0WXA2v7KJxi7S/IZ+vQYRb/NaF/Szbemfjhrtje9Xf05+0Od1VIFxe0EFvadOBAEHlNEDBbFwy9
wu9TmSNzzlRetP6XIxzv4RM0Gu3tAgEhT5WTGIS0+tlydLMVnghZhagm5yiA6G7a06ZWPkZc0bCj
Im3vQdKFyFeR/aN/hCjGp4M2bM9dZvNoVFWuC15S4t8ek2pKdpHqi7JJ2fQueN5fAC2KMSi4UB7I
B2RMAAtNrNmFqKvqfzW/F3Yay01cpQMxyzrl8MuC5TvWodDaG08Is+XB8s/x0C93QT/rKEdUO8N+
B5nocxGr54yLbWISmtEydq2bDaBVxYe4wG4d1u0aYP7xg4MKnaSAvCtaHPM9RLilJr4Vn+C4S22D
/B4FrSwDjTHs0oMB8tK+TiaS5j1AFiXoE3aEtUJ2QHXnUJEJebY43kzAjx4JmW/G5M1k3aHoltNc
dVWGeNpsecti8Z/b5DvZWFUwmHxqVdBMywfnnraxJXfnhCi2YRCn6LcryYNNIlsMBSfNp4isDTzy
XKjjaMFSCJuEAaObBeB5airmzfFC/Y/kYITHANbI/xOAqgKyjiJphErNjvduW47pFHG6GnjPOzEJ
BBlUnAd8WeQZ3iEkMqolyfVywUqmLX4OPpkxLXPA6UYobEHmrmqNQgascXTklegqIMDFYPHKjAY2
bHfLTKxkRz6NpEPpoB7obadcBukKbfB81mmySvkMsbp8Td8F+lupr5N5dRnfoEZwsV8jaxe3HeIN
y6CoGUYEWsfrQJeUzQaEFlJG3DwPzMilHH4bneAnLepMdxlv0njT3gX8RPRfuo09Wu0CuciGuruC
QcGjxBqa0ZuTpyvJU1XTcUYPTitH3mbrwQRcQHsp+XjY9QMgzX4ZqKKIjGppmsDuKX3DUt8kzPgx
DycNgBWFYy+RpLR99YPe/8fd503dPNxdtUkZVdU6eZuc/TFJoTAf850gBjSCRpGm4U5pdMpGIsF8
xgKyRkI7bw/0Ndsc9OWquPXX/nK6To9m/STser396sMfJR5cCjGUtMxJeW+ZrmJ+L3P4NVo2YRMg
JF1Y/ULEv9NOTekSeTj2LhrZRlsmslfUvzUihE/QvtCbtddaDlHB+fuKt/Fuf41RZ3Ygv/lM5Jy/
XI66j4w0aZEj7Ak7uvPW7aHIXAS7setiVEJJRI0iXnddI0X+GfKmdmFHWN8b6pMbX19hvUrveM97
nkBIXVR8tMmpMLlB3BFPSiJLh05fBFpBZLjJtjvB4PjqApFu381jrDAg6AqKSwsz1BdCSFwLSN9T
uTJYMS+EljY29axy6Zth/d/Y5d4fDor+G+RO1fX3xfSie9oKjVH0rkr1ygx0I7exLqzdLekU1sBi
MpnMzibXwDV51JOHzH36Uva4h/ImlKJi1Ik0vb5Yu9yrv2DxWav3MQho2oORNF7xaP04b+L5bKfD
vw5xlFjbnGb6EuIgXUfeXffpo6Ce8JC485yeWy/cT+hC1TPOHLkAWY/TzMU4C9Cpo86FvMayYsgy
Uh2Iv0JYe9CnvsLN5AxSiMzwjjwC+oTXSpszRDLn+nnBjQJWRfBVfl6KdwTVJkVqPrz8m9nqiy4i
h3T7JdPuTfBWtDfj6UM8O4Zox00DgxdFAQhhWpax9rXPwRpYinO9JQX32tcqhn8jR40uppijirEy
JQ7wJ1QpsYlgP5NgQYzutW5Pq3NF3wC15CWkbyFI3eS7EFDEdV9mgDRUDlLpSIEUG/CxXfs0RsuJ
2WGscUzQmzsOKa80y6trYqTejHtUTYzAYSr1eOhqrMFOn2Fw2ko9XpHd9xFEtqTcjucGK//EdXNF
ee4rQ7Vx/80ETWQoJaOjYkU3V+4kLFtMmfzhHeNXrORh8msEb+kwCSe1akrTHZmhzT1W2BvL5KQ/
qlgHbz2Bu+4GuIhggGo1OBB1Z6VohAasDQVDzBkCcSdBi9SvDSwN9IElbsMmRFcp8fsl/wwoFWNH
hvp6m2Bi0NZa+hwkpKOZ6GLGguK9tbvy32XopVOxQb8N2JjfrtEuPL3x0NjGs/9r7lU5AJlRhqsG
v0zCSGmZtSKfHkvTmfxscf8FNWRUSkzWtbifN5+OFC9OiHBVEiPAT7PLSCJgXfCZfVYsec8bN1oK
XHm2PReRu3rZMrDU4HfkpCrp0rY4Ddg1IPLkpt6xF0qnwSUgGL3jX1AIkCrtN3V892nsNbr7fNXp
zQMywEBxNd5OCFWTjyfn4n6uyOHUmdZ6hr4eFcv2Djs++wU2Jw8WTBvermgdIW9g6oD3/ZhR2SYb
g1DclrmmdmJyMyDt8u4sL/CUmw3rwL2OVbt9m+wO90XjJBfkQOwHeRrBaCyZ0QZSXzzBlVoYWgJP
i0D+E+gGE1ZHcBYlNkfb0ChnzyiGtIrA8O8ScyGyoUP/A8GIH4+ZXZUvMa3LQDaR+/kg6/rJR2S8
dU3bVgu45HFgJODmSA2ybr1fdYGlfIDeSv2H1yjOvzZJDsKam8k4C2k0c8gFqqzvChSiS2/hMMbR
ECL1TxdpADwNfElzeTFvsH8GDGp4LQAdAA9R7K008EnHWzNhffZvAo3DA6RkwBPlhHxEw5VEfwen
vCOrQGZItcikcuNeVQjOUEcODjxzFR+ryj0jec7rg/j2XyzMO9BBv+//fensjj9UTCOhnSW2RmRY
H0fhNjmctauP+5zc2bN7fga6gftKH7i35tF08QnA4bli3T4jyNOetHU8nHTqMLgfMHfFdMBWZd16
n58uAxPYGMFdbn3aUU7GrpPFPcNOym+yaaNp4vIta1vMaGLk8O2o+rs5QkP59BS9L9c7i8BvnRHb
AtGT+0bS7F4/HSYDMLNrmljF3z/6vRHraD01/9VmFCHZynGSAhnZGiu+kz59rVoB2mMRQybRv3o3
t2zNO7tglyvHlA82al+ZNmjrjMOplAJFwronZrtOkY4/kbbggK4nSwSMt8wmxIJP9pSJx+ZH/xwd
UMquLDzKVflM1cUNd6dF08sMpXArxK8ED5PoMSk7En+OsUBamioqu6wmuFJBCx+IpRUrXg+raIiU
mSQZC64Qxggog8TTLLcYTIuJA0yqVRvxlBcWfnoMhkld8VzsQ3x3RApFscBlb/SawIog3R4Gqp+y
Vrb/6YiXTu5X8einuE35s9x/R2B5vE2h65jgmFfNuDG2cp/vFUM3TTDcgSeSsEhR0j06xQeSvBPC
gWOKVidqQW+d0TvfwrZkh3LBrayQrj7ktQNIHHOP+XuH39CClx+NxcgWQvdvoQyRlf9hlVnCU94S
ww6MM5in2n9UKyfbZn+K6kDl97gIX+3CuuAGpoCwlk3s9JNoSZaKoFjwoi6DGiDUdi5jPOgnbwAR
omSVHmwLTChPfU7xYg2nqhE99HQEYLBBVlvL2k3Fae8Ths3zfgyxnhbMVCsEp5yrWUYF9I2ON6o+
tPHhUNlRY/RfP6ci0PEfRCgrQRJwQ3nTcZRJtL01JKRsqg/pn5f1IP+ulT6I0AhnvgklJTLfM7yX
Clyd6Jtdxxyou2dBQrT19Q9g2FXGPgNjSFkmKaH4kxgitXBYKbglFFb1swCsl2ai++UQW7ogeSOW
9ibofrZTeNWx6tCYP2y7Vq2SSwi8UNDzw1CfqBk1i+gsxXp1lhrbUU2FeuW85bXCGhmkA+Qj3ALT
bGPPum2Meyg5DkThjh9HtNJ9RsJ5gb5aOpxtS1GJBzV10WsUpfAJG1gocXURRKtWc8GVom9846M+
avrQzXck+I3vIgFSRacv46ZrKZw1PudEwcehMiPdUB0MgQQnA8/nJIoMahJ4kfLxV9fMSD6un6r2
tZ5FxG+PjQWCoibUZWJfkv9vNS4qjzAqtr8Fzv7ffKRgyeRx/TPqaB/8R3s8klx9YOteAcyYGwCj
LMuLZlWvt6QJcyoOlXrhFuCmtmlfC3KqO8KK+6GNi6q/3n2+49AeeGm3tlxReFHBQvwU0nFzJP5T
sdiQlEPS7sBqtPkhzqD4Ay5jp/dz/DTAa2Yt4nGgn8kkzarhcmV3ThLz14scqcxVdelKO6gPWdqv
Cvqc24BPyKfoFvIHRC5aTAfBY21MwcIT8hgIe+dUgVF6MAnPk9ePbWCl4QI60L+MRxnuT/C7nBPt
craluqjkS222jX1Cftf/Jb5gnvhY/S9wf9oUdxiyi5ISHCaqpkFkfERoNsiV5tLh6gtHyv03/lRL
h4gX8Sb3x8vtGM0IKdDcyBtN6JtQHf1/ceM+g77Zmq9xKnIFR7WKE3ulsVJENnmZjEFliShkZ5Ry
d9NwD97aoDGhW++z4bBoTPwvG+XEWG5xQu7Bn9Vy7VSZRp0+I7lcPi9joOEiaeQ+qwqWvWTP/bNR
BF4Dt3I8VzaQHzlbuKBc21c6YI3mXO1Wvth8WZsjumhP+P/Q9SQ7GEeewqIcpQkJb0kh58B5C04V
IhSmozC6MRoZFggCzXwyANFqhrES3uGQ9sX712bWr1E2P0AF4bm601nhmbhek6UJL+prdacGg51h
uCbhKEcqxEOh0gW9akpIG9qKAEQuzzK/kkIa21hPK92cVhm+I//ZqL/e9oc6o62RpBJCa9/t0gc+
nz3B7yvc/9KY/MvbLyoUnjhQnmrYV32xtnsqqitFA9pJP+pKjSMT4PpXHQi3cfFXP59oZovlhBAD
sTlhgF4zwfT3ZyQfbkddC/G1BQHDj+WViFgfTXScdCajSLhnsd/Hmeccrww2aKnQ5ueBaRvHfpcU
qacB2BR3jzY76n0dmC0nnp5JEtZ4tURTnHN5MBXoLnf2EGjcjnw4J1smmivcPQZmA+hXvhQD2UqO
urNSxMBiKIArctB78aCdExVpwbf6wvZkUTq131qCmqVfj81e9xkZj9LU2y2CG8sH0lB6kX3PDqlh
hx+1za4MYmfzP618Bz/F1390XkYwCujAEAgp7D7fKyZE+FIOmFA2HZ6uNVVKWpD9eq4OIcO5hYqT
lb/EEpsj7fDUgZ3B2/cUFAJU/mUFd4tA1umEwoR+lFoljs2X0VHq3a2Xy+A2LNTyxuwOi62UDEd5
rmCBxmGoRwuGKzbgt0sjQrtCi5e9bqmCdI8mzgt/PmjZhRocO0fnf6IVeYwWQ9RdoljElPKrOfGo
In+2BPzYro0NrPy1TidvFBbe5gRyIeMtnnyJdKheiAZ7c+6ESddWi7BpbgON9xM7+e0yktYc4V9+
FLE43T3a7g2xBOWGY6CcskhByeuRfYwIFbWpyiv6h4YKvF4HNXLdi1W47kcToKyUvc1mWqBleUhW
WIlOjgkTKuRFEogmC7fbKvP8aRueelnfaBCpnILdASkmxNT4zvfCIFVjt5PyF2pEh07vfW8vgQsw
1Ekv8mZIINMBQkiLvWDHwjgsj/HvoeX/38aLsvgl8uWCoIORsqzXIloyXFjYmS3C5t6HO56BTXCP
vvHhpaCkPrwZcY8XwVygmSjghYvrnidMPKQ8AXYpP4MkSXTaDAPTAuexRUjdl3z8QqrCgh8MsQCi
sbIxkyUGRV8xVDPrDQEjdM5dzheGOrpsJx8pq8SGAjL/sdag/y4xYyBopvRP4OySZVUxI922um7B
NI8slRVYhMG7cyHC1smtR5+VEAGSZhFxGFPCUVO53eiaajS8xj7JsyxrZj9KURbHVwDCy3d6LyPO
RN0R8WquRcw0+kw8LOhBFrzfYETF/Tl1f1gdaZMIBiKYqORV0D3iE++jd3rvz7VGlOQRsVA3U898
4W1xCjw08w3N1ERNkyyjoN8MU5hbQlguddEzGJUvpyi8PDKEIKuIQMtJVg/6NRWtnVE9fJJuWpfF
Xrw02lpK8OoEhVZOdcwBDwK3kyRxLbjlm1j0MS7nyQmit2nmKH+Nzc60JAImXwEjjjBflWf8ebKo
Lx9bBkZ7HLXQsM1RWOSwDc6T3StSp4FNfhNQNifIywfqxImifj3ZrGr4g9M6qzsSPBtAtP7q+RF7
INaY09j8KHSGuD2RanZrPb8K9gnUXoOkCI5Z9rDvQD8XbLN/JcJPVVD7rZn4xez+8AJNIaO2f6mU
F6gTcBXd4NWQA24XV8lSbDjCYMv6l3YqPnCL5iKABDmEbBKGV+UtfgYPLSP7XYj1ubEak8YfoGYq
RaQX3yStnei8ngKwJtD07kmcpg9s66uJhach6wk0HMgHIO7mRmLi1V0URklW/aHdoCz0xYzJGwLO
3Xt/Qp4IGrwBRXDQuK587tnDtiwXu/yo5RWSzPdUk0w7wlThJQvx8TjfF4yp8UHl9II3ar9ISVXt
L5qMWSIS8/h14Y2s3Um82tC0SKO68K8Wj/p8HJfevuv4jZfwHCf4TSDZK6Kk34/LO6+oBTiZFjl8
79rI7mG/Y5jnOzkyK2d/opoVrnom3EC8rDLmffDia3nB20L1RLgbeiGGDTJG94ATareBGZergXOM
x2tQT7A94AmtF8yr58YXnjKpttbJpEtEGZNBf4bYTjHV7P+QvmoWemonVDrls0rsuIm1h7fR7YTO
TaeqwEU0PXVM77KXG4krX8LI+32CR8nbNBbeQgllqCoHq+jh6Ur6wzPU0uIug8PW/ndjXBGdeb2s
gV2U2PYejloJ6tLQTv/cyYq/N3wuUC3XHuRH5xc2g337h0BSOBLNzQFP4mPazDyo5nvPM0JgUyF0
cAXZ3ARWbpK2xOZFXJjrDrRgv1a0ENhXJOwO4jre6gIaI549r4ig7WviuCiLu+wxlSlk+RxlGKuc
oSygq9ruKRgnz3oegiCa0h/XWIZGtSq8q1t/XIxC4+Sd6K6ctOzp3Lm1q85EpEOeRX3gwoNXhP/U
NN6GxkSPYdX5EjKeCtykvLBOvJHB5CxGONs7fp/lu6PkulIkRCglPiOdQ5fuJdu9dmQ/9c93AQc4
NXTX4fYKv4P7DTg0CJWfmKvUNVbBMl3Ki8k/FXTVRRfNeWOW4kY6c/9TYAuyfP34k++9AqV354IM
tbd4XzOXAeJaMpxTf678sT7Hb5rzNXdPAu71edSRbUXXmuTC7unm3JO+u6j3oaDwWJiFJQLMZAwc
4J6ozrvnp0/ZU6w1Quyx5U6idOA/oQOmoU8RnG87lOIlsjIJyqc81ZrpbiciHe53LyEMtsJ1QdSD
B/GnU5QdT1JNDR84vaWyHhnj2Rscf+l+rkNFr63iKnz8F91Qvkl2ZBejBrONUrum1brIhxrglH2u
ziEQxPHG2gg9Tutyc8xmaX7xM1TY083WjK/NZOSt+hC3wsYnaAQwbAwY9nI/GfSm0JzCy0HcTBOA
r8zrBSU/5xpF4HJxwrW5r5Zl1e29rWROD3paN7/PwAfyXulHoEqDmTQDgtQy3xj5ZWJT8T0Kd0k+
8Cq6KGMQ1SiJp8OaIRfw/lFH8IKxG6lIorx5FpBPXXCcRHhpxiUCR/6WAcctmql6TxuOcKTQn+uK
tWCvSOtIu+UyX1JNCOpgag84lcwiYsgckkyFkx59AN8Sfuo71K9M4Jkj/A4pEDh0zt212KycRKKQ
xVMNe4ypGorhWPPPcSFmrBtEg3vV0HFPO5TMPXz81c/x5acdgaeauwkgEa5fnTc/KkZ0LKRNJfTy
ZQgvPRTUcAhSUOcrb68Ul6HMm9KnyPEPLD23Gk7xPLbZYdnaKLo1eauca9tjAP1hoh1/tlEHVGOf
uY0yff9y4F0be9W054/FKBSb7cGh9XseoCBYsjTYksas94VDXffGVLNnoqjl5PI7pL+GiJuQgu6r
UCRJJXXbHZZp1ogavOmQSmK4PNOl5L/K9fW7iA7fQky+fACk3PhnC9ceiAG3CeOdIsY7bB0ZGDYB
785m0yY/jwCiloRS3T+xlcoeYZFfeXNiewVJGDtj6Y3JCWfjwrLa4nkRrlKmPnMVpkhEWCV+QMxi
NXWQX3QyPEZNu4X8SspQ/ygOqFIlzekDGReKm/T9mVBwmPTAvQPhLg6rtTdmizXkTzJLIGlq72dz
Bw7XfsaHcxWxxKnRAang1BZWUdP84xWycOkaCMM3AWEMPk//OFfZyKDwpZC08amqMuFLxBx4jWD/
TMSS7ZFJk4sJ6ghElD+LrYuTQlWjRWOl51oeBLvE4xdiLGN53nihWUAKNujpawNNXNbGNsNO6BUH
bguDWVpx/xPFL8yKypf+Urlhaxk82Id8XHF7LC2eREZxr0r4uPSVqziuF2EHc6Rknjj61NDijcmo
cG2iPGVo9tjkfmKoeEwQX9qI/6HtuAZ2Fe6/I2iZcYK3XFHEjN9xusPNmHGxjK30ShEWepBZWIQa
xBC5CrPL2yFu0JOnpxTGeCPsVV/D6lmtBWlrdRsRTaJ/mtVd2WCwYtG6xLvmTk78TiVAwuR/4rVl
BFg5q0mFH0hQkOTzbx0upyHv7ANAFWEOFi9/A84zJoa1hjqhRCUVVhNl+jzNWMtkE8leJq7OvXcm
BSaQ4elRQ1UuHoC9ZzD8L8/U1HAXQei6WnQ9GetEbw8MFOorGbFdJh7Ab41Dnu2VlyMujtvQc2uZ
W76i9SCi8e+F0AW4qZvkHnpBSlfL66qpDWrm4J+UHPmGrvDQ66KF5QlEhz0parPyRmPqkgnvp0Ha
2+xsR9P3xyeOa58MZ8uKt2RNDCf2Kb5QeqUP4BGHJg9KB4epjecGBwsjiXtw+sAC1rztjU4+FGvG
ig+C5Odh6u8tJfg98uCXaurvXSyfrxjIEjaSX7qmlX4QiSmZtwqTFw+ogu6kbnLKYjFrmEW9/gmy
whV2RMX1Xc4SCKnM3RwuBmT6j9NiF4IHJRX7yj/IovL2haIS7yrsokqmp2QoXROn9kd7VWbCqKDb
AormSox5c1I6fXdeao8TGIcfYGTt+r0DxRWNyGyQjZj6NtOqkSMcGr7xmo80z3kCCSOh4f0R9nMf
Q25sdQQPm06eORb04jud/DdlbmcKxLw8YcJwRFiv6tyRVbW9h9wOrtFXfJGt6d8Yj5V5sywAORYO
mO6xBiCS4rs+ERh90FzRMeijGEIFeRFSC9dpoMSK2KgNJULg1pLm7RjiTddmcE6DXZqImP0E2RT+
IG9qGKgtUKy0J8BN1Q56ZmofnrlBL6hHKss6fxW6VkrRvelmATLSera4MWiTXkajtMOeA0Lm9mvw
Jpl+4DvuiF+gM1sNGAcN+viDlWdZvw14T+4BOFw0FfP4aA3f33eNn9LFPBMs3b1JztYpmiJBbRVS
PcWqOOwjfgcYnorvUR5v9KTUrz/6+LXk5hxYejU9XkkGrIfQn2FKmAtsNxBGZJQMLo6ooq/QKXC7
AqPdtUfjdLW9mic7VaExnDWOCY/+/G22rvGN/CNA8DPO0QTtGyhla/xPDaRVrNC9Zq5atssHa9td
02frhAlo2uBCULRxe+2Py0S7G+MpdR3jNcN+dGPcCgEHnPUfFJ8jiSoUrGv2aUK90zpI4TMRdLMT
CZmqr7EcrqgM9lTeqzKME5QSStDjLBlhJoNu/mC6K2ExWgtrhBYyZhzbE+DqGxYMpudUWlLz1a9L
qlUqFR71xic0TQKvxdAAUdUpWVPrkMXqviA/KfDlCFdmdI9RobcEZblo7FtSiiL7hX7DeBVGvdGw
6MWDp3Gv0mTjSWW7X1kmCJ7NuEgIuY2akJtx3FUGHRqMEUFlu0SLSLHTbdiE5BzERwbBzfwSmlFR
1MtcCGtGrnEZ0KnIJvpYxbhkJTn/QJuggUxfVwt2yMzUFWbBmpfUWsMHZ4DDFcHMJMEWrxAk/ZXu
U4+E9xj+MJ49pUE4mSrR1hIuiO/SW9cQxeTTCp+FVerVv6DR4aD3xqkdJ50CJYn+tUb3pceeUOcY
2gAeRcYXstsLYtRmpWuEA+i8s2u6DZbbQomem2b/c0RH9NcrTZpY+ysPsA2mSY36HL9+84nSDZH2
rmWaCAQEAQbpZPc2XAO5Al2z4UXNGYHeFw1s0dtGDYIzFtt8fTHedI9yj8uv89qnq+QzQCh8nAsy
tqjgvJ6t2s6OyZjO3Hl077kT7bAcAv11Db7tz9LpO5Fy0Cjv/Wyc3iAkFcCqA0cmc1OPYUV2+qQR
gbqs/KTYY7p9JKxBRqXUcXIfRDB/JVJMrNOZLTpHY9wb7qW1ViY4jG10SKlQmLXFJjPNKgNMh4gI
odhMtnBdPNMJhxJzGNpxkcNh7CCqetRS469rAv4KMVoHmklkp/Qp9WvTipqX4r4VfFHNGtgrPxiu
L2GoryIRLAeD8qghMBtMSkqEtxpWqfqrIev7G6WQBoHKVHc6k+KbmmlX/FqzAdPswmUVzId5JjSd
IOSumYg2Pxc6ONOgOtlhLCA0bZlpz0eh1zqSSKku13bf4l0BXaFFzlP9ZdWfDjYTGQpe8TemvBLG
pVc4zutzqoc04yoXI6y5p4fqXZ0kelSocCaE6hMuNgm+yH8pdr4MbwqfQM+wUkPupcjYbs0BJgRP
wlB/6voiHE93ORbtAyZkpQD2BBvI6wZwOHGyinpyYsezrHvVDAIl2qigCRSDMS04/C/AvVTcZbAS
pKxAUSU2FQ5ORDctiLrZhVy+UG/OW5sO9/TG7Sn5W9c+m1BlGLhSRv5YeSqG4B0PpdKyBFQnDQnK
fHzONfGPNQgCTxg4QrkvOWP1dxppy+b0Vvtv1OFRKCN2BA5wOi7cbDURKV6+qD+CDfyhS8HYCuvz
VEmLkIGS7GxIi/kV21lvhukeddZmJPjJ1rWsPuOFtsdhrjx/fKGOeIPPxxgMJoaQjgiWKkMC7wo/
pGKtMBqnaUBIxIIWTpXYPgMdEY4hlcR1kwm0UgyuVleUG5nQ+mZthrNIFAHlOAC6FWwpxTE3wHXm
SIiN2hRYN1NyndCi9ym3UP7GbyoVke30cfQA57xE77qAVV7LQyd8IbhVbWD7AJcfOlcpnuD9BWQL
UVfgf1aqizwIUOyEIj7sqU7gAFG7a1bJLv2eNj+QhoaoTDyVQa+G+KYo1Ke+6NjOHkjAQXvPz8Z8
IWT3n46O86r5MuS6uapzm9tVpn3GVssK4Nv0M3emx7LyUjbVufDKDWMMswEoRBpv2VDPJy9zedDc
bzDFS+6e4XovKTRztmJh4AzI1tbI8X/YzThtEwvLuLK3J6NQPxzAfcfHuPab+fwc4Rw7uyt5djgb
u8EQA77Qzgf7KWfMZJ+hE/Fdzz7hg3A1CZ7DY4Z5uG7VdI3mSFIDZjJWjYwQeXAVeKjBd1aa/H7y
DWDvoe1316GTqn0oVSGubxUGEhOuASLOc7yrsQw6abWTl2DbkWKIiT9FZ92EOleccyxE06ekhVlv
45hLnH8y9TfRgC6aQDdDxcMlSuxAsAex2OSzdCH29h/Zqcv7fs8BeqJR9qhpGuPlIKRIoRlPZMou
A8i3n9P5iKdm2SGi9i+qgSkdE1+grsIiaU/0xJ5XzxoxXDNdOoJsLzkfpwN1YKRpVODl9O8MGovr
lFJE4EVHcUCUzNxNMJ9SNR4sHV2m1B7S04ySmb+DKgLgjR2PCGs+dTSgQPvDeO62INqLDci+gfGa
bMDNj4GAHlWTGm3dYmYMHQ4+LrYnUVz0oaakFCP0lNZPxpkciIPrDAa5bU6ex2F0ktFa5N3k7rIq
m2Q3x33DdcOYOg9yl4t7xRrTX0/CVW7GWW7aqufHR3Yph3Dm9Bzl9OWfEs6qBiiP+gKD6pQwZgym
l0txfh0MneZu8ILqgSegjMin93BW7Ftt+S6whnA0/Hv+OfI1CAdqtugFFo2fUPBvKqdMOSE2ULj+
b/B+TVT10zqLfoVM6PvJipWHbGaXmCRnN9ToAcKfuWmnWlIBcBaD7y9a5VE9sixaPbzZMjBmx4vE
uDzaTldD0Qx3Ms0qtv3250QmACgukECaM3Lfnuql+yB4eiwoM1auIhIo5QuBGA+MbccP99E1AfzE
6513ne/6xBB0PzhhpZ7BbBN18QADS9HYZCZkQv4esPkBYiyRzNZo0fKMuDq27KIcZAwo2BC8Qjmx
8+Egi0i8950PV2PgCJ+nOo+YKXC5ZADrsVX+urPh4GUvKZYOMxbmvGCGcKItGtFS5ynsQPgkqyoz
PaNG/3gsQ10D9wPMSVlUBvOHFWhOEPvZ7u06DEX31crYWJslyW8QiQ5EaqCRAy0QsZwqKfyX4SeJ
ROALEihmsCZ1jXxGbLdbXhy+urIa87gG2IRANnzfdmX42tp0OPTiuzQhx6Izq232Bz3z3sAll05M
AMwsUHtVvHwDVDTQV1jS2rm9G1f8WBpev1DwULpJDeJQk6iUnpKb7LEz4ieglhZn5sZ03H6osHI6
81d3nQIjL2ZCp1EWD3EuCHitZbLgRQ7a+NbgvzQVXGQUZRS94YzrVx4/fbFLH0e2AN+HixYNTxft
bkFrLI6X55+KJ7zEkHi6UlTmbC9VI80glPlWGc+Q2VRqIMQszFSoWB/NQeDFr1QgNYHg6Z4ovwry
3A6EZ0NUF5Cqj2YvbEiqh5d4GO4ZbYXLMMdPMMuBAPn78Tz/9MgfA+eYGnvsUIekgth6meWY5yb3
F5BDZZ9ySj/ameGl8MLfrHqAznhY12ZS2NTxK+8ceAK2+zDVm1+WXtXU9l/jsNMz3KrmL3Mjt4KV
+3fg5RtQKdu+XUXve7T4IJfkUhMPhmMxlZiS0RAM7G3DvUpVd/d2ulfwiQEW7NJ3/7CgGcdtAoXP
j4SRc46kZxbtSUtTyCDhbjqHA1A4dMTBslRL8C9sIz6IQ53vBgJG+3KOZf941xuOP7N6qJjguHJT
moF93dzTKdUXuC9PIjEx+TeCZnj8oyhDV2++mw2glIPXdMVpUc1uygiRHARFye2C/lpwZxJmNrgv
XEjrWhxSoIzqCkefoSXPaVn0/gZjwHlDcB2biphruzK09E1+G5/jMwk0pCE1w4IDW/kbxVFeuH9X
jWEI5d351keYePcOxsWTJxMUiMtb+45DjkQNcrBrsvjG2wZ4ov/M6huaIhPX4aqzCScqHhqhKb29
MzlBtu5oaxbCFmymtPpWCY1QfV4Ewu5o39Y0oXC5fllUsRABKfj6BoZ9UUDDP7ftVoQ3FHTUnCS+
LXKep/xIxgafMoWTAz9EgEx0vHQ79ae0RjtvpoC8gABQssqLb7kzmfCsNcB+AOabu4zKD+iyb3/Q
AuqMPuUtMdBPdzDFwVhLZGGr1XOSdovavNlxp5NCBWgCzt6z/lHNH6IxcMHm1A3t0NmhL4i9auxt
lRjWnee/BCxE4tyNkOegmKj3gQqdb8TbjmVvTS82/b0Q7gd//JDmyodBRv0dC0ZsJEbcvJP+CHX7
l3jKXXpy8fchw9QSMwmU2SGb/MYAa0fLE9+RaEdbtXAaN0vuWhAb8TmPsJwpttNdCn+GQE8Oku1K
sCZZbIhPhF+qvizbSHarQxEhTWBALg+JIP0l69bf9tuTWygTTnGCj+aksTjaKA7WG628xAJA2mbu
ZADEJGizPPOYutDYOG5D9hvkIfVYBxOTSSJU9HIDkWwh1E6DUdAeFLloFRR6fSWdRmwhTRSuBJ2Z
Xwi609Xiez2Zkq9WTnINTzMeqQK0CcvBM1OOpkmGp4SFBGWwTLasCFW/miKUNz4Luq6O2QKzNult
XizEaZsR5XIT/mj+t19/d+hY6763W0nF32Dw87Um6u9SkjJUl6BGIYSR9Szb1rlXKlCJVSHY6b8j
NRVZ4tU+EtT5NTU88A0z6Ry0i2/cu3/n+52ntw76GOR8EZ5PM07FO33YzdxpEKOlEg8I2CmdsMV7
vhECGg0dtSUg5vsNwExaOw7HBJgXOBBFgi9IGGYSkkruH7ZZLq+b6+LnllQTL5HBMKWcNa0EPflt
SiMb5/UOqweSKU70hALEBqtWYW2vLsg7Hz/kls5ubz8jciupVr3C9N+rdtJK0TmM4Y+wJ8Ma3hex
NhDD/uzdwlKe3LC2/bwm70gn0++sz6Qn08WkwcKkY7QsReuykhgoZ526gXQfgyhzJeDY0RSxvUuh
uWFFavCcH9BYfrnadvDnWVwkRYQBTcAb/MfWRAuNYbpC3Io+BuYNHQ3qgaFOdqB1sh5l+uz+mPkf
ivOSGX872pOh/1q8Y1D2JrFLpI1CfNQLqdplqJeWIuN8zZYii/+EZs+6fKylp22OhtW/HPjicCDE
T3uITviZoIJMM7mWiEoso/M81SRj9Uc2PRc//r0B5XaH/ciS+aatp30nZMlyLjFA0oE/Vn5lwxFG
lB4m+c4MmT3iYLXEzedsyDDnazC2IrNcmYK30rpqRelsxf/aBdULcHu4EXCou8gcoMmUcoy/niYP
b/RhwbtEut+p50/ooAtvCiN0qN42DvZhpl10avSbiF3mgqG8xHgo/jgjq/IGU4yoHtslsQL6GM5p
C5wTN2oKbZxXMb6x5DJmaXU07YzamMd6EAXygOylWwH1aVPgXnNQLAEqeAkk31ObfZkt290r8Qjp
mHX3gydtWuXkNG2cW4HvsglD7yf/akvGfrTnH+R/IM90T5hh46HjVvTQ1JQIlwRnawcEZhcHABtU
v0e9jLc0VMP1qratCsZ7g+kkxkS6RuWNRBMMjRgP6cp9xMq3QLmH6jd4Zo76bstOrUnc2BREsF4o
g3EL77WQU5u1/pdUZF34zHzQqvVu5kZzyyXT85dFcmmI7sGNtbgB2cxQvx1f4fVRPNYx8tRkSRko
tsZ0lXn2ivPrZyXMLXFivXN93GT8Opo+xqehU3+RLbmBraN8sqrB6XnJVDksWfOB52R+4+LuraVn
cUdFQTpK87SSzQKkCgFKhhmIbezuE0mZ3HLP/JSH/3SiWDov5i+sFIJiinuF/pXl0qkOHXn30dvF
aJ26PzQ+wR+xEfOvBglFmrHlypy+/4VqWwqaRLvLDyAqVYnyAW8rLB//8TbnOLLSxcstDIllpUNX
3krSJzk0iTJIZlR4GWud/JgjvSgt8EkaEOAS7mBkjx/6bkQjTGgDSaVJjUaUjuTULJ6nIM/o21qg
H9CGw/gD/dSdCTgBzBs0Yk2P2QfAo3pAnXdCrbSjJlARAvBTMxwLQs2k9/WIRYwDIh0QS0c7TDH5
EYMeaUD0nXJ4JdBkRqQs9eEZ/CC2jqYREVQ4aiXk1WfPZ47Bu4IgjCpb2Ro5x3ORs7vbmZj+IpRJ
AlejdEHtkufFAG9DEV/W3D+OvdKAeifsp/jEefKoWxJorm3o/Phl35neEOPNN7Mko+b/F+qhLRhS
EdU8CfqBFW0QDlONwryiGQgeOFQ1CuXASW1/Y3yTZ4hx4hSpxRrOp1P/lcLHsoUG5trUOOfjCFBs
zcP1+JMy4F6KIYjPOJH2lDU1VHzBmF/wFuBfDo/tGQ89ByBrC3tFvplRrri7u4y7pHqoOvFvmAwt
agoWjPxsiLy99g6A2SAHWQFYQKieQSC6gN77h52iy4Av+84Is5dRGVbqfcVDjH9u4v3fyCStH287
Mst+1edR65G5Rp1EdrktQN7jh3Lnc7NLZLeeeMQKzvtdz4vOvgbJ74a2JXmKGhn4XlZRYczgt/XK
2aiCE/A5W4INK1ASB0M7hGlWH+5T3WUqhjhUNY/q1qqQFg09cCaUUxUesYiEQu0685GpydwBjFjm
tiTzw5HTueV5g43F/XqsP4OR8IgkRbfznxSwGYMzWeZP5mlbAaRh0HdEVNN2w6yH+Nl6GJjiuZty
UUFlX+NF2olJb+ulVdHyGGmOoUsWb2Vn6mg58HdjKeUdq0EXa22KJGhsGOmB3OEW4vo5kRdWUnh/
XOtp9zzfi7nz7ZG4DdbjZoOc16NkUP7ECRCAzdHF4ISP3a120hWF5u42lzXuyVf+F6vmHiJ6IwG9
OrJsYMsqX3loRxvF4ttGMp6TzfxMUHmxxSfMkUGywlhAYoLEiDIdsuCCqzVnGzsMtxGrDMGx1rqb
a4Gv/Z31hwNCzyQVIJvxu57pcqd6NOPP+x2VWI7oW3TCs4roanFuYnmiKsJyOqa9F1UCEj0EC5ef
s5kUBaDTNkbsB0N6p8hUDvqAfe+d/VCT3MSi6WsyMRlp+gVZ31xjKNwGGknXMeEFsJdcZCspkliT
NCgYF6W//1hjhoKmOr0Ckndq2F+xnCNct9tSPL4Vyj9kIQl+bpv3QhFWjMIA7nFrDUfh9AOHJiVg
SY0IYHoeVxRjvOMkswxF3eFwYTVSbbRdTxGXhe8bbQQndNmBjGkkO0eeeobYBDd79PM8jydjksA+
MPuIVU95s9fjbQTasukBoNwEHu7ZOATYZIMQezC9ApZyt4X1yOFgqo67VGaF7xGlECoPryG6UTQA
wi+aT697FJXBVrZD7p3YK5W8F6TbDB4eRECZ1UD/xE//7pmS/p5ziAYboe5f0RsuojhghokoOQAS
lymjmwXGwwfKka6xPjDVLPZ+IQhg1OQFfVHicHoLIpD5UQXJz0IR9pORcXxIPSqxvH6HAr7ArDUC
e58iitSLO6/hxt77iQ6BsEPggRnAKRSM/KmNFaBMwc91e/7OI8+FSUkiRMNk7npJk3YQHbtOBh2n
NCfdA4e2VTsqkLSMt7tyTikR+qUL+U+cWVFNWKdRo2hahSDMls8Fp8oHogcDCd5bWrIv3BOlMUS1
sO8KIV221DbQNPYMVi5rx1GbG1tjACmnygMyubKjcE3h5MgzP0fQeN/2ClLkCcHpOBT7mqpb2cGm
4Br8fqBvjkuoH40B+GAk/NI7vc5EjlhS0/o8wJlZqUDw+BWBqsavmV1mNtrlCn2KOmNP/Z4lX39P
mFgqihr7NrkifC9aCExqq2tEZOrbaDyvgX5NbAIMhQmCNI/7HnDqjweXdRqZJG5+6B/mnnzZoKCB
FAUqxy55HOCKbHQSOWH2TOeAiZ035/mCphhWMZNx9FRYPRJaZKSrrtcpF+HhAEpficRWavhz8Zf8
SemKBz4zWg7YtZMfMmG4aY3turbpnmjoLhTkAaFuL6OQlMwbLhahhgm22gMizMOZ72enUwjwjW8t
er/7MHqxTKC3rFRtkeaSd56ERtL2POBF8VUUr3vaNk5r3g4DXpS2uLdlDSrMZm3rKgLn9ZkGCsw5
NnrN709KT/pmtKIAkA1Heb7Hw4AaIaTmUx/rmxNn22HHIylFPtpT8Z8k7HRNlRTMXGk0bRBsNuEn
BRI1Kjt6aefdCOakuOcb1MO+tbvYEsp8fKzxSWyrB/fGb8QgxcPXEukML41QmqVhQ4Qiv2sgyz9Q
mFxGig37d4nivzVhWusIEIjdgaf4PJj/m6PgSuEcj58CA9NTenkI7cjRLd2uYcEF9i2EgxGySskv
i7/YFajyoVjeebJQ7FgTMIYY8RcRibN9Kybp03SYGgP7XPTPyYMVzOQHGYjNKPcWYLUxauJFKzy3
rZJSj/c7Fa2X5SaJANggcPT3q4aRn5h1XXNa+dhZq/6HdiUW+BgxKqh3QEfiOpi1BR53K8Knx1D0
Llcp1yYKc6xJkJAHXoUD3lIrHIFpFsZVQgjrx5XgPt6nDdpGpv0jnoT4L3cp9Kgl8Eqnim00gZbK
byYveQ4sZgKfpM2SozqJurfqzcScw5HdkrjCOlk6DfYmR0ZbOeP13VRWQVRUTqRLUv8FIqWCIvYm
nznUU+3zpjL2Vh1+SShMHRfrg+rOBFxmsd3fNQjSm53sOvkhq79lBpMkTq/0NWVTQKtLzW1fqb00
xmgtd4E+EMBmO7/IG2bzLXO+ROBgb8H5gr4T9RrElvXjDuDimyUqUMArO+2iv2kqtfNHTzN1jEJ2
7AehBGHZAHJamD1yNrWDmve024aaHc5Q1BESJWQm9bkRiGh/Yo4k32cCxoQ3BOUwO19QTJ1Qy663
5j+2G66+vMDi8yQZAFrBPBMLmLTD7b6noxbh4EOqU9y/lqQAMcOrekTxwkRo60yDf+vJfgHvzhCy
SjRaG8A2OcXqYOICktN+euOXBnMxvdshxB36tfY4OPEVrO2aXN4gxs9Ozi6JRy7s9KckdthnFVuQ
ZdkLArGA7QOFpBmgIUVJPY2nM3nStPpNXQhG8ECR1Xe9WQh7UfzHE2afSL7jJ9nJRvUo5bAHsvgm
APMLt9TYyA/WhQEVKBD9jttr+Y4fh7VTn++eqWP9tqk98hju0ruEfqi5IqbrIxmcdktvriEvUnOe
xCsGQL9p9P7LRIZZsRVsm3NMeCfjKWYtWgwcZ5YyOzIz3OkaCYPYSNMc6RDE+OBLnhVci3tfcm3V
NVF7j3e+S5o3hsObJGN/wbYB9Bjo/lM8neqvjrmPfGDKIjj0P5HbspAWSS5DTF4E/ms9KRYYHNbR
4vY5AUq9uV9YfycYvVWYAn4mPCKjUxPO+Uttv5ZfIaqeNIa33OWkFKlo9r+ZW3s3GUirIvVEspTx
o47HmwZHLZxerHqQlJr6qLoKfSNnp96wotC6l0ng5igfmTKUMvkT4qnu2UJVGQNjgg1uMWy2bmkC
woWHF1E6kPG46zPvLkJTrwJfySiAEAcDq3bsy9eFgVneo1Qe+I+oEQUSTUuk3Mhv+maKO8IEJ0Kq
XdJM9q3oddSq3VdBAOz7MCIFsApf3gBT8t3U+ZZl0LtaMHK8z5jawAinJ0Yw4hPjKzzAm74SLu4i
szLXjQOcBHjIT3fA28vKi/WAlEtApFbS2WFeXZt0tbEhBT1g9Nuz2cwBrYkY7Feg42vFnoDt1nNx
tkMOEiojMpkbEd0+dtfdJ/vB3bAZ9tyWavNFrs6+RgRFvoT3l+yHHBl560klFBWtmWb1h9KXkobq
bpnChTsoFQRT1axc8HywDVrqCdE1itW0sNvFwiaDK0SQkakkgDMctm53YahJhKigXp1bAo9i2ev9
7thkLCuC25faycARhK9j/I+aIoOxfC1k+rPz360+p2koKU2z3hEspx4k4yta/e8uAPK8HoY1Odvs
dbULmFmtjT4OKFJyH+fMuRdzxowGXTxe3LR3eNNDvSzN52tfBarQ7iIm8BNLQy6vQMSqD9kk7t7U
Lw36qMlSBtO0RZYP8sbK3WU5R2A9hCnC47kbmNI0Rs0LkzdoEauIC/8QS7o6P2u456QKezsN/xZ0
5eic8JlPwpfeM97hu9y9fQyjLthpuzpQyOwCXCO2SPNbph5PnhcUmNqo7UoMevNDn6NJZo7+NhjB
jE70k201fxL13JHfLyedYeMJTdJvjBSxW64h82NjRjKgeueipqHxhnniclpUEa2XkKPA2gtUba8E
ZdYrVbf3fo9dms8VPtw6Bu7a4A6NgRzOZMkgHi8UjXk8cW2ieBPlIAeXVaD1u9RNcuIedwhejgqM
wCVEAATd4xRPkWZNzcokYmimP6LZQhdxwkjfLpa2AeIFldj8hPaluTlqRC4IvQk/YcaCjVZLGgzi
VaLER3DPlQHxK3/XNFViOBQnuQbEjHZFGJTT8NUlZlm5JlkDuzLL8KWZdlmEkPRkFZsamSop8wkA
OKBEuBu0rTwfUoYNnBrwkkEirhcW67g/eqlC8N7nlsfsXq/+tf0iQqnFhkQF5Ajw0y69RWAT7kBi
mKnZO46EoIFOneT7u9P6w1A76MJWZNp1Vkzge5nJJPtv+3zKOuydlQloj5pnXPg8IlKzCCipM3fu
3mTwA5zqsEXBAxYQUCtcOxzUBqHaMw0azquYyvfHGzTEJeR5jQ6MI5u74/Tn4DJ8Rb/vojzM1Cid
jyRID4Vp1uyECZKtX+C/SUpPKCS9qR/UqFWtrRlx/rwsY0Jqu+d1AqyuGTYmNyTCWo3synYUzMWf
b8RRC9/k0K35LYzGtFdCXHfpcpOwhC5XwfZSgO4h3YtWb1IZyGO6rNn/YzXYl9IL9thmRLO/ozdp
dVVXQFCSScbsTK9CUHlOcK/TqpGcZFtMvKjCDKPabwXtzE99CmUI/QQcjIag8qwSUrYWzOMFjapy
H5nhBqtVT6FwqajeRHZob2YQ3QhhzjZ2F1ULSkk3wO01E5sRqLOFYEWHn5D2p/X+M5eUvwUYnj9f
pn6BhblEKuE6faqbWoqI496jThuSy8Qi0s3GWChiVbIJHylqcJKJu0ikoeYK9YSwgKG5lSvb4aqW
41lLXRgBbYunOgbvKHx3igL2nCGwuwVY7knguPnNuwljiu00L0mEkKj7r4M8am8/VZHkAHRCYmdI
IQW/Zfrqyg47sxpz0RunW0GZy2GNyyKEORITEbfO2yWj/KX5gD4raTx6Pd6Oum6v++jENRoQYo9k
ALmfAcSCBlyvDBQ+RN4ey3qRAnY/2HramhRUSiOlDE8n6WY30rf4uunEHWOuzk4xR9+FPbpXCSzb
zoMEAhJCXbwE1TbTj4Os42S2qPKYu6bE0Xut+9RqW2ghc5UXximgNvWmBQAV5vsycT5qq5bdWT4G
wzgA2OGqheP0KwjA4XHVFn/cJQ0L9TgredPr1kO+JgJyto28SSBP6lOPqV/axr4R/1d0SK6n1MYB
wh17LkCM/TfwTLHCYR06Q3L0IsT7wnuICTVDMlhMBFjKYwiCfW8R75Uq+2LvuXLdVDJwxyRNR+T/
Kl4JSQQsBeptTwSCQzOSq3+a425D+RMZI9lJBZFvPog7n5OwzliTTfgn9xUiQUKF3kJyc2YXniGm
6HvOEK61CYYUf2YP++NTuH6ntnc1oa7T1B8RV20DCYNc/2Tdleh4d31pWfmqDdi7HWoYYWy8C4IS
Y7wSuI00of1mfbnReoYajhotGlt4SHX4p0N5JkAKyoR8otZWCWv5WxXKH36zy2uEZYlc8WR1d+BQ
rAaBOBQWP4j/CLBQln4/94IEPCkgVogEnNKP1WmkyHf+/UAsCQaah2cnxrQ++AVqrnPQeOGChfm/
G2+hKpBURNco86aWW9Lz125ekpLlyvQmcfVyJv1ClxwaJ0utCVgu9ncxyHy70GIPYHxLN3kEmAxB
Lij0bd9QBNj0ZJOJk3XcxKn40k+3C0lvrSu1nv7sDgFVf8grBMKFXIhtI3jq+l3HkUQC10asn+fG
Czrj8MGOZl3xG3E/+wcwMhBC978Q0Y10cjGC6iaNNcEFtrUw+MAgtE/h26Nk7Jv0/0OiwGGWL2aC
I7AOeU/s4DvsTvSNY2LFfNObU9QDQPSZ9hALLL2whI+/3oXw4JHRYQtK1lUOQhMju7hGvIsWSrZ/
wkJjNBBpyV9YmqjTAc2Kdyxrs2iymoiyFs3tNrjqy1Sdqj3/hRdss08ofmIl5/oqGvHJ0sPEQK8e
YLc45BOxGCqJD077Bn/eMuwS2DBPjwxjza0/92isJMtcreWIipfW0cUs/KevEEjnjMOvJRFb6tqb
m6h7pimWUf7/0VL56nepN2iDvyNbK9ZYz8xJaVZJORO23YGpBnIG0MKYXvWb+d24ljD2egpWv32J
fmtBaBqBcHjsb3hFbzNLktrjfzh5LHpyOapUFiXVI6S+exohGXusxig/eNVu1i5wcRmQcUlhXHJs
BT2SJa+XEY+qDIQkIsnHY5EqgczEcUTJaNj7olzJKUThvdNfeyo1drXt57ppzzH9pLF4IxpGOTy3
SvA1lP/Q4oCbCpi1n4lt/U2gY2XnnX6th8vpmmGAb64eO02UWh0152Zi0Fqw7nefWLuLBeca4k+w
Z4neH+hHlWwbuKpjptpiptdSo1syyxlnJA4tzLmNoDRPjzRhbFVSGYwIij4awfV1NK4vxP3IzO+u
4N+f12VduI2EETDcqtUsE7UTeACr46CKHVIP3/vlJXS7X+5aNrFjhFTx3WUyXfSx2wGV5rYhZi/+
8ZohlzD+gg0F4O5C5wVVkwq8zsMO6BlElG1I/8PRVDI3+tuOeLvCjJhw9kmo+lLcyFmpiyPC+Qn1
OxHeTSGnPS8pg0XNbE53gyf7FbtpM87ZBKohqrPtkApiyI1jtpBCZSGUyTZtcDMRevycYweVIWe4
cUCL9/VxyApQJ2LL3LqYgCmwSjjTLvd8jrpyOwDYYux+etwBqEVdPlkvapAROYxIIgEVSGY3vhOe
1Qc3QLfpxIsAQ5MjZoanqwiKW8Dkr9t0UOcT50tY00cu1ZcOV/b4kFuQiOyzmimuefGb+6iPB+Ur
4K4MRNKht2evE1HtKbC3Y0btYMybT7xLNfE7K1kZ0f/+QYKuEkmwlow02wiIkpJmj0NayUcIneKS
O9ebkgSDKBPZcOE2svgSoVclgZtlA1wbYaivA4UASplGQGooVpPK6+lXupYiRRdTWoq80EsFw/er
ovYfkOknc/611HR+AOjIRbjnSFNOPtprG+JiSJqo5CyA4TlxIN4drGCF3/EaPIimsc+/uuEQZwPh
5XQceqPDEQu32cUcDe/EDrzYm3DjSmsA4vHoKBdpPzS4PSOZjEuu9deRBQmXbotYvJOFMsE4VJMY
voH+WbDTxbM19gnCTNvw8TLNIf6Fs69LZXNkKCaF+iurIJZ3y869Aa4V32VAkPoz5FQn4hodsCgt
Z8AtJaml+3Mhx2onQsWTSC9L0+/ogq/+Z2cvjn2fOtCplkYvF535VJAb+bDQx3fGHsNAQX/+WEeH
q0UCoXMonnh3neMb8ZF5iIOvoPQcyEXrJBJyhZf3UNTbuSjiWfDxN0BU2mlC97UP/rxYYxmXo1GZ
m6ozOxwGpdaJmgZRngb2gKYjAGX1CgQGcpx36B3eU4/prJ06PutijXA0pCR+GIi3VOO2V3saUhV7
PCJhR8c1Jsn/56ZyVSaRYfNFqZ7Dt2YkAk/ZlaJo9xIwTGbRE32nwk2JPVtHM08qnoQt2a3UPws9
AMcKHAEIXjCXvhU27VDtjlxVtXQiqWhcoI76NhqjBoquTSbPfzQexVsGLMQgA1G8jxajEi68Ev/6
8rRXLX2BxGRiswVUIODYCkLRmwewk7xI3gXnQWAmO7MJwBdPkL11VPRrZcESydZ+0mHMYOonTN2v
dDgYRYlbgtYA+0PMZgU9/FYUnSa33x2rYS6ZDETsat16+Bv5RP9wiqkbf2ep9W+ipKwDrMw1L0K8
4trvckXm0N6jDDZ4MD7P+4oRmKjLdULHi75DcLsLjPc0/m5VlVL/9j3fMB8EnM6i8Y/xhU8e4s+Z
xWSEXNjFAebOU5vtBPDgn++jooIo1MnlVmw688CZFWGBmPm7yxaxXHNQ4gE0zG5SZFt367mSL+Pv
4wNI++mjZWj6QT29EZxz31b02BBYEjy0pa8GVKKtbq9kGMfA0/xrr1rQZhSPS496+qmzPIzMo4fX
CIOrA8tMe2kPqJXhn4a9Z/bCP4bUMocm7EyoaZJBLMw1IGokzCdw/v4JQj/K8vEZ7tKVlP3I0/LW
YD1uhRczyYhlIQhwH0mtV4PCUEz3BSr1HwG62n67a5ojJkNgc5N5U6YO2Ab3anObrLEs3ttJxcR6
DlNl7Pq18aPAJ0CyvmEvgNIcKgxWp0qsvekXP9uCk1fVPw+D3ZqagN87LZl5lPexAiKeaCR5Acqv
+WT6fQfkW9oZgyTZKbEMnrOnJe/yQFG0vax1ytjpKh7chbv5hf9s/6wWWNCzfGxtdhjLQNV/myKP
wpROsokXgJa4iPeWHpBqSbw1Qxd+M6GCCREZr24d42ErOzzT33u7Xja4XAFp25xxc+YDfsF+Udsh
Qzo917j1NMJ7l20ti/rSgaASyNox04B2oyZjFkC7MkfCiRqnHBlBRDpNemqZ+XzXY64AkQvC/RrV
tApXkd8aw1z3Nl+OLl2N92E8ArWPzjg1YF/fm/l+gCU79yuhHCWR/pZDHZQ1hxrdsaxe4IwGsKh9
cqAZVmIIUby/ND5CjPcv5pjwHjb5YxdV1oqespDxdPx/UwBaKOX+EoFUfHwrUcPONPT1yzdbOtfa
A0mOh57s8rsmKYq7RXj8CM7I+8YguuOvhagVV5exKnRGwa+bmNWpqojGzY/lYa55m1g0kvQLObUX
ghVUKFRMVFZ8nFUnUmH6Jofwc7T2EfcBg+086W7ExLTj7VQkpDNYCAGi510P3+9Lp+C51iChExKR
QLW2HurxRYLcaaZeGUAyA7nSHDkTHoP6uRvCYLwxDtJDhGLaORkUyY8fRV44n4x3a4CMGSyygumR
0lyR9QoytqoDZeiVx3DnVlst4W3wJg6bwUNwMJNJ2RWtv84JwVPQpWVStHrjSd0TviRIY5Tb9vjc
J/xG2xi+3TBX5OX/h9rTasS8xit/lxcHrpEvAem+FgNIuKiqYXTgUd60eQqbO9lX9FxVV1hvdSQb
4wh6BRLTUVt6kjbJFIkRRuVY4ZZdsFBNyrF50UV3Q1Teon23Z9UgYLLoF65sP50E3DA3npMDZ7/H
7WSABsAsSyzu3HTYsTtkRlZM6qjLpWa1FAaosygXheIICANO+AcxKCdLkYHW3h+D0roGe+428jmt
vn1jEFnAnCsucZ1OQ5dFIsfKJ8b3jbO7B8vidsQ1XZXtu1CYc2pjoh+MP+g0tqpPJhU6ZMMCmMe3
r7i6+4NHqnGTjGGP84LsOT7KDCrufCIp5lDyRdJBjkw++hYYeVy7UsBEoYVdaRsHJLCrCvKDQ97W
T2WFa+SpMOqmFzYeBiE6V9vmL6nIICuly8Hpi8wckI8gZdabo8gGoTaa1mk2pu/r9CevxCqcvbv9
66rFwlJWBrippIK1DNeFK+0XQKJ8cRof2G+jCC+YjtaBQDsQ66saxSB3+z5eWwqobKJynxFr1DLd
15O7ciXDHys7ahgfWrbB2Nq/YBJjNyOQd8w1EgM7l2sjCExSnp0cpMca3VYmjMhHW7zo5MfkGdKg
fDfyzW3GK7BjAP+g7aourqoNaMJiIxJmPqOpPjMUNGq8do+XrEOClnOFSz6Hr5edXw917k6v2TV1
cpU/6N9sYWid5tXtyK/+QTptz3ajPLjvVpMb7sZ30g3ngeFT6mM49Se1XpxuJsOOpzJOvgCN9jG3
j5tk6kSp/M10eERAwUdKCgIJnHT4UwOTH5+KUMcDMFWebxD0cKrR41jLXBnZas+vFP05RKuYzWD0
Tmmat9JG6zqyLj33ll2HjoVysccSWkfMO6J4cfqnSbBX626UR1RNTM+G7MmTB/nuLw9h1CT2gVkV
2mCN29BJKQCcwRtf9m4QaDUO14dqWbyoc8mwDs6oOZo5DMUqB6xf6xcQMaCKV/hE79P1jU4BDGeA
s+c2ixALnQJ7YMnjxPjKP1LV+DLu6hr9xHsPei5EBtqaNhkgcJ8SQ4Rz5TkWbsRwUG6wG/jrx6hQ
r3sGUm6YFwFF4LhwevNkWmbqurrQw4D9BmxzHas+FeIE+JRIByizpxofbwmog0gnG1EoiBkgrMUX
413GClixydoEnnZKb4XtfJ+9stw7n8hHptAIEi0oVIEabV8SKHse88cxbs+dQdqdRh1goojmzmRf
YRTI5oy1SUDY+TXgiiggmKNR1oE8QN0Aln8/7ErRwNtRIdsYnIsXh08m4A5L/5hCcYB6jqf+9TkF
7+Mx5ZWmvKB66fCGgwM8o6Heb9QrSW320S+9G0YIeNwd/1wmx8UEBAnldbD+x50Has+Vc55Xa0gN
h9PkNcQEiesjZnYa9HHhl8ooBnNpbL59iLuOGuE+smz8+J0ty3ZJ6/adR20zrkKfn1mYmhNCeK6c
nkqS0Wltq9necavwOVZQV1UrVykpvGEJ/4FlVScmqkqphaL2nprYxiCba8DnFqSE+F8lAEE6X2ZH
VmIQhCYY9hoOI50dqr4kLSc9xAEQDwaqPLx6odyOrNc3IVywQDnZVeuxisQCl8InJhf5SAWxjxdJ
tjv0cFbENc3jUbKMfi4O5rgqr4XVxxNYmzJMLsNbWYbbkP2ohfgGT1v+wNxxeoA1ZWgf//2QFjCt
R86M/3trfgZ32Q==
`protect end_protected
